magic
tech gf180mcuD
magscale 1 10
timestamp 1702351822
<< metal1 >>
rect 12562 56814 12574 56866
rect 12626 56863 12638 56866
rect 13346 56863 13358 56866
rect 12626 56817 13358 56863
rect 12626 56814 12638 56817
rect 13346 56814 13358 56817
rect 13410 56814 13422 56866
rect 54226 56814 54238 56866
rect 54290 56863 54302 56866
rect 55010 56863 55022 56866
rect 54290 56817 55022 56863
rect 54290 56814 54302 56817
rect 55010 56814 55022 56817
rect 55074 56814 55086 56866
rect 13458 56590 13470 56642
rect 13522 56639 13534 56642
rect 14802 56639 14814 56642
rect 13522 56593 14814 56639
rect 13522 56590 13534 56593
rect 14802 56590 14814 56593
rect 14866 56590 14878 56642
rect 20178 56590 20190 56642
rect 20242 56639 20254 56642
rect 20738 56639 20750 56642
rect 20242 56593 20750 56639
rect 20242 56590 20254 56593
rect 20738 56590 20750 56593
rect 20802 56590 20814 56642
rect 23650 56590 23662 56642
rect 23714 56639 23726 56642
rect 24658 56639 24670 56642
rect 23714 56593 24670 56639
rect 23714 56590 23726 56593
rect 24658 56590 24670 56593
rect 24722 56590 24734 56642
rect 28690 56590 28702 56642
rect 28754 56639 28766 56642
rect 29362 56639 29374 56642
rect 28754 56593 29374 56639
rect 28754 56590 28766 56593
rect 29362 56590 29374 56593
rect 29426 56590 29438 56642
rect 35410 56590 35422 56642
rect 35474 56639 35486 56642
rect 36754 56639 36766 56642
rect 35474 56593 36766 56639
rect 35474 56590 35486 56593
rect 36754 56590 36766 56593
rect 36818 56590 36830 56642
rect 43026 56590 43038 56642
rect 43090 56639 43102 56642
rect 43586 56639 43598 56642
rect 43090 56593 43598 56639
rect 43090 56590 43102 56593
rect 43586 56590 43598 56593
rect 43650 56590 43662 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 4622 56306 4674 56318
rect 4622 56242 4674 56254
rect 5518 56306 5570 56318
rect 5518 56242 5570 56254
rect 6190 56306 6242 56318
rect 6190 56242 6242 56254
rect 7422 56306 7474 56318
rect 7422 56242 7474 56254
rect 8654 56306 8706 56318
rect 8654 56242 8706 56254
rect 10110 56306 10162 56318
rect 10110 56242 10162 56254
rect 11230 56306 11282 56318
rect 11230 56242 11282 56254
rect 12126 56306 12178 56318
rect 12126 56242 12178 56254
rect 14366 56306 14418 56318
rect 14366 56242 14418 56254
rect 18734 56306 18786 56318
rect 18734 56242 18786 56254
rect 31054 56306 31106 56318
rect 31054 56242 31106 56254
rect 35310 56306 35362 56318
rect 35310 56242 35362 56254
rect 36766 56306 36818 56318
rect 36766 56242 36818 56254
rect 39118 56306 39170 56318
rect 39118 56242 39170 56254
rect 40574 56306 40626 56318
rect 40574 56242 40626 56254
rect 41134 56306 41186 56318
rect 41134 56242 41186 56254
rect 44046 56306 44098 56318
rect 44046 56242 44098 56254
rect 45054 56306 45106 56318
rect 45054 56242 45106 56254
rect 46398 56306 46450 56318
rect 46398 56242 46450 56254
rect 47854 56306 47906 56318
rect 47854 56242 47906 56254
rect 49086 56306 49138 56318
rect 49086 56242 49138 56254
rect 50430 56306 50482 56318
rect 50430 56242 50482 56254
rect 51774 56306 51826 56318
rect 51774 56242 51826 56254
rect 53118 56306 53170 56318
rect 53118 56242 53170 56254
rect 55022 56306 55074 56318
rect 55022 56242 55074 56254
rect 55918 56306 55970 56318
rect 55918 56242 55970 56254
rect 15038 56194 15090 56206
rect 5842 56142 5854 56194
rect 5906 56142 5918 56194
rect 15038 56130 15090 56142
rect 17838 56194 17890 56206
rect 41358 56194 41410 56206
rect 23650 56142 23662 56194
rect 23714 56142 23726 56194
rect 17838 56130 17890 56142
rect 41358 56130 41410 56142
rect 41694 56194 41746 56206
rect 41694 56130 41746 56142
rect 42366 56194 42418 56206
rect 42366 56130 42418 56142
rect 15934 56082 15986 56094
rect 14802 56030 14814 56082
rect 14866 56030 14878 56082
rect 15474 56030 15486 56082
rect 15538 56030 15550 56082
rect 15934 56018 15986 56030
rect 18734 56082 18786 56094
rect 30270 56082 30322 56094
rect 37550 56082 37602 56094
rect 21186 56030 21198 56082
rect 21250 56030 21262 56082
rect 22754 56030 22766 56082
rect 22818 56030 22830 56082
rect 24658 56030 24670 56082
rect 24722 56030 24734 56082
rect 28690 56030 28702 56082
rect 28754 56030 28766 56082
rect 32274 56030 32286 56082
rect 32338 56030 32350 56082
rect 34290 56030 34302 56082
rect 34354 56030 34366 56082
rect 36082 56030 36094 56082
rect 36146 56030 36158 56082
rect 18734 56018 18786 56030
rect 30270 56018 30322 56030
rect 37550 56018 37602 56030
rect 39790 56082 39842 56094
rect 39790 56018 39842 56030
rect 42030 56082 42082 56094
rect 42030 56018 42082 56030
rect 4958 55970 5010 55982
rect 4958 55906 5010 55918
rect 6974 55970 7026 55982
rect 6974 55906 7026 55918
rect 8206 55970 8258 55982
rect 8206 55906 8258 55918
rect 9662 55970 9714 55982
rect 9662 55906 9714 55918
rect 10782 55970 10834 55982
rect 10782 55906 10834 55918
rect 11678 55970 11730 55982
rect 11678 55906 11730 55918
rect 12574 55970 12626 55982
rect 12574 55906 12626 55918
rect 13470 55970 13522 55982
rect 13470 55906 13522 55918
rect 13918 55970 13970 55982
rect 13918 55906 13970 55918
rect 16494 55970 16546 55982
rect 16494 55906 16546 55918
rect 19070 55970 19122 55982
rect 19070 55906 19122 55918
rect 20750 55970 20802 55982
rect 42702 55970 42754 55982
rect 21970 55918 21982 55970
rect 22034 55918 22046 55970
rect 25330 55918 25342 55970
rect 25394 55918 25406 55970
rect 27458 55918 27470 55970
rect 27522 55918 27534 55970
rect 29362 55918 29374 55970
rect 29426 55918 29438 55970
rect 32610 55918 32622 55970
rect 32674 55918 32686 55970
rect 34626 55918 34638 55970
rect 34690 55918 34702 55970
rect 37986 55918 37998 55970
rect 38050 55918 38062 55970
rect 20750 55906 20802 55918
rect 42702 55906 42754 55918
rect 43598 55970 43650 55982
rect 43598 55906 43650 55918
rect 44606 55970 44658 55982
rect 44606 55906 44658 55918
rect 45950 55970 46002 55982
rect 45950 55906 46002 55918
rect 47406 55970 47458 55982
rect 47406 55906 47458 55918
rect 48638 55970 48690 55982
rect 48638 55906 48690 55918
rect 49982 55970 50034 55982
rect 49982 55906 50034 55918
rect 51326 55970 51378 55982
rect 51326 55906 51378 55918
rect 52670 55970 52722 55982
rect 52670 55906 52722 55918
rect 54014 55970 54066 55982
rect 54014 55906 54066 55918
rect 55470 55970 55522 55982
rect 55470 55906 55522 55918
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 42254 55522 42306 55534
rect 17042 55470 17054 55522
rect 17106 55470 17118 55522
rect 17602 55470 17614 55522
rect 17666 55470 17678 55522
rect 19618 55470 19630 55522
rect 19682 55470 19694 55522
rect 42254 55458 42306 55470
rect 14702 55410 14754 55422
rect 5058 55358 5070 55410
rect 5122 55358 5134 55410
rect 11666 55358 11678 55410
rect 11730 55358 11742 55410
rect 14702 55346 14754 55358
rect 16494 55410 16546 55422
rect 16494 55346 16546 55358
rect 16718 55410 16770 55422
rect 41582 55410 41634 55422
rect 24210 55358 24222 55410
rect 24274 55358 24286 55410
rect 28578 55358 28590 55410
rect 28642 55358 28654 55410
rect 29586 55358 29598 55410
rect 29650 55358 29662 55410
rect 34290 55358 34302 55410
rect 34354 55358 34366 55410
rect 35074 55358 35086 55410
rect 35138 55358 35150 55410
rect 39890 55358 39902 55410
rect 39954 55358 39966 55410
rect 40674 55358 40686 55410
rect 40738 55358 40750 55410
rect 16718 55346 16770 55358
rect 41582 55346 41634 55358
rect 15374 55298 15426 55310
rect 2146 55246 2158 55298
rect 2210 55246 2222 55298
rect 8754 55246 8766 55298
rect 8818 55246 8830 55298
rect 15374 55234 15426 55246
rect 15598 55298 15650 55310
rect 15598 55234 15650 55246
rect 15934 55298 15986 55310
rect 18958 55298 19010 55310
rect 18386 55246 18398 55298
rect 18450 55246 18462 55298
rect 15934 55234 15986 55246
rect 18958 55234 19010 55246
rect 19854 55298 19906 55310
rect 19854 55234 19906 55246
rect 20302 55298 20354 55310
rect 40238 55298 40290 55310
rect 21410 55246 21422 55298
rect 21474 55246 21486 55298
rect 25666 55246 25678 55298
rect 25730 55246 25742 55298
rect 31490 55246 31502 55298
rect 31554 55246 31566 55298
rect 34738 55246 34750 55298
rect 34802 55246 34814 55298
rect 37090 55246 37102 55298
rect 37154 55246 37166 55298
rect 20302 55234 20354 55246
rect 40238 55234 40290 55246
rect 13694 55186 13746 55198
rect 2930 55134 2942 55186
rect 2994 55134 3006 55186
rect 9538 55134 9550 55186
rect 9602 55134 9614 55186
rect 13694 55122 13746 55134
rect 15038 55186 15090 55198
rect 18846 55186 18898 55198
rect 17490 55134 17502 55186
rect 17554 55134 17566 55186
rect 15038 55122 15090 55134
rect 18846 55122 18898 55134
rect 20638 55186 20690 55198
rect 24558 55186 24610 55198
rect 22082 55134 22094 55186
rect 22146 55134 22158 55186
rect 20638 55122 20690 55134
rect 24558 55122 24610 55134
rect 25342 55186 25394 55198
rect 30942 55186 30994 55198
rect 36206 55186 36258 55198
rect 41806 55186 41858 55198
rect 26450 55134 26462 55186
rect 26514 55134 26526 55186
rect 32162 55134 32174 55186
rect 32226 55134 32238 55186
rect 37762 55134 37774 55186
rect 37826 55134 37838 55186
rect 25342 55122 25394 55134
rect 30942 55122 30994 55134
rect 36206 55122 36258 55134
rect 41806 55122 41858 55134
rect 42702 55186 42754 55198
rect 42702 55122 42754 55134
rect 5966 55074 6018 55086
rect 30382 55074 30434 55086
rect 6290 55022 6302 55074
rect 6354 55022 6366 55074
rect 5966 55010 6018 55022
rect 30382 55010 30434 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 7310 54738 7362 54750
rect 7310 54674 7362 54686
rect 15486 54738 15538 54750
rect 15486 54674 15538 54686
rect 16718 54738 16770 54750
rect 21534 54738 21586 54750
rect 17602 54686 17614 54738
rect 17666 54686 17678 54738
rect 16718 54674 16770 54686
rect 21534 54674 21586 54686
rect 21982 54738 22034 54750
rect 21982 54674 22034 54686
rect 22654 54738 22706 54750
rect 22654 54674 22706 54686
rect 22990 54738 23042 54750
rect 22990 54674 23042 54686
rect 23438 54738 23490 54750
rect 23438 54674 23490 54686
rect 24670 54738 24722 54750
rect 24670 54674 24722 54686
rect 25230 54738 25282 54750
rect 25230 54674 25282 54686
rect 27806 54738 27858 54750
rect 27806 54674 27858 54686
rect 28590 54738 28642 54750
rect 28590 54674 28642 54686
rect 32174 54738 32226 54750
rect 32174 54674 32226 54686
rect 33070 54738 33122 54750
rect 33070 54674 33122 54686
rect 38894 54738 38946 54750
rect 38894 54674 38946 54686
rect 39342 54738 39394 54750
rect 39342 54674 39394 54686
rect 9886 54626 9938 54638
rect 9886 54562 9938 54574
rect 10670 54626 10722 54638
rect 10670 54562 10722 54574
rect 16606 54626 16658 54638
rect 16606 54562 16658 54574
rect 16942 54626 16994 54638
rect 20750 54626 20802 54638
rect 17826 54574 17838 54626
rect 17890 54574 17902 54626
rect 18386 54574 18398 54626
rect 18450 54574 18462 54626
rect 16942 54562 16994 54574
rect 20750 54562 20802 54574
rect 21086 54626 21138 54638
rect 21086 54562 21138 54574
rect 10446 54514 10498 54526
rect 1810 54462 1822 54514
rect 1874 54462 1886 54514
rect 6290 54462 6302 54514
rect 6354 54462 6366 54514
rect 10446 54450 10498 54462
rect 10782 54514 10834 54526
rect 10782 54450 10834 54462
rect 16382 54514 16434 54526
rect 16382 54450 16434 54462
rect 17390 54514 17442 54526
rect 19294 54514 19346 54526
rect 18946 54462 18958 54514
rect 19010 54462 19022 54514
rect 17390 54450 17442 54462
rect 19294 54450 19346 54462
rect 19518 54514 19570 54526
rect 19518 54450 19570 54462
rect 19854 54514 19906 54526
rect 19854 54450 19906 54462
rect 24222 54514 24274 54526
rect 24222 54450 24274 54462
rect 25566 54514 25618 54526
rect 28142 54514 28194 54526
rect 26338 54462 26350 54514
rect 26402 54462 26414 54514
rect 31826 54462 31838 54514
rect 31890 54462 31902 54514
rect 32386 54462 32398 54514
rect 32450 54462 32462 54514
rect 35746 54462 35758 54514
rect 35810 54462 35822 54514
rect 40898 54462 40910 54514
rect 40962 54462 40974 54514
rect 47058 54462 47070 54514
rect 47122 54462 47134 54514
rect 25566 54450 25618 54462
rect 28142 54450 28194 54462
rect 15822 54402 15874 54414
rect 2482 54350 2494 54402
rect 2546 54350 2558 54402
rect 4610 54350 4622 54402
rect 4674 54350 4686 54402
rect 6178 54350 6190 54402
rect 6242 54350 6254 54402
rect 9762 54350 9774 54402
rect 9826 54350 9838 54402
rect 15822 54338 15874 54350
rect 19406 54402 19458 54414
rect 20290 54350 20302 54402
rect 20354 54350 20366 54402
rect 26674 54350 26686 54402
rect 26738 54350 26750 54402
rect 28914 54350 28926 54402
rect 28978 54350 28990 54402
rect 31042 54350 31054 54402
rect 31106 54350 31118 54402
rect 36418 54350 36430 54402
rect 36482 54350 36494 54402
rect 38546 54350 38558 54402
rect 38610 54350 38622 54402
rect 41682 54350 41694 54402
rect 41746 54350 41758 54402
rect 43810 54350 43822 54402
rect 43874 54350 43886 54402
rect 44146 54350 44158 54402
rect 44210 54350 44222 54402
rect 46274 54350 46286 54402
rect 46338 54350 46350 54402
rect 19406 54338 19458 54350
rect 6974 54290 7026 54302
rect 5506 54238 5518 54290
rect 5570 54238 5582 54290
rect 6974 54226 7026 54238
rect 7198 54290 7250 54302
rect 7198 54226 7250 54238
rect 7310 54290 7362 54302
rect 7310 54226 7362 54238
rect 10110 54290 10162 54302
rect 10110 54226 10162 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 17726 53954 17778 53966
rect 17726 53890 17778 53902
rect 19070 53954 19122 53966
rect 19070 53890 19122 53902
rect 21870 53954 21922 53966
rect 21870 53890 21922 53902
rect 2494 53842 2546 53854
rect 18846 53842 18898 53854
rect 3714 53790 3726 53842
rect 3778 53790 3790 53842
rect 5954 53790 5966 53842
rect 6018 53790 6030 53842
rect 8082 53790 8094 53842
rect 8146 53790 8158 53842
rect 9986 53790 9998 53842
rect 10050 53790 10062 53842
rect 16370 53790 16382 53842
rect 16434 53790 16446 53842
rect 2494 53778 2546 53790
rect 18846 53778 18898 53790
rect 20526 53842 20578 53854
rect 20526 53778 20578 53790
rect 23662 53842 23714 53854
rect 37102 53842 37154 53854
rect 42478 53842 42530 53854
rect 34738 53790 34750 53842
rect 34802 53790 34814 53842
rect 41682 53790 41694 53842
rect 41746 53790 41758 53842
rect 44818 53790 44830 53842
rect 44882 53790 44894 53842
rect 50978 53790 50990 53842
rect 51042 53790 51054 53842
rect 23662 53778 23714 53790
rect 37102 53778 37154 53790
rect 42478 53778 42530 53790
rect 23438 53730 23490 53742
rect 3826 53678 3838 53730
rect 3890 53678 3902 53730
rect 8754 53678 8766 53730
rect 8818 53678 8830 53730
rect 12786 53678 12798 53730
rect 12850 53678 12862 53730
rect 13570 53678 13582 53730
rect 13634 53678 13646 53730
rect 21858 53678 21870 53730
rect 21922 53678 21934 53730
rect 22866 53678 22878 53730
rect 22930 53678 22942 53730
rect 23438 53666 23490 53678
rect 24334 53730 24386 53742
rect 24334 53666 24386 53678
rect 24894 53730 24946 53742
rect 24894 53666 24946 53678
rect 29710 53730 29762 53742
rect 36990 53730 37042 53742
rect 42366 53730 42418 53742
rect 30370 53678 30382 53730
rect 30434 53678 30446 53730
rect 31938 53678 31950 53730
rect 32002 53678 32014 53730
rect 38770 53678 38782 53730
rect 38834 53678 38846 53730
rect 29710 53666 29762 53678
rect 36990 53666 37042 53678
rect 42366 53666 42418 53678
rect 43038 53730 43090 53742
rect 43038 53666 43090 53678
rect 43486 53730 43538 53742
rect 47730 53678 47742 53730
rect 47794 53678 47806 53730
rect 48178 53678 48190 53730
rect 48242 53678 48254 53730
rect 43486 53666 43538 53678
rect 2606 53618 2658 53630
rect 2606 53554 2658 53566
rect 2942 53618 2994 53630
rect 18174 53618 18226 53630
rect 12114 53566 12126 53618
rect 12178 53566 12190 53618
rect 14242 53566 14254 53618
rect 14306 53566 14318 53618
rect 2942 53554 2994 53566
rect 18174 53554 18226 53566
rect 19854 53618 19906 53630
rect 19854 53554 19906 53566
rect 21534 53618 21586 53630
rect 21534 53554 21586 53566
rect 27134 53618 27186 53630
rect 27134 53554 27186 53566
rect 28478 53618 28530 53630
rect 28478 53554 28530 53566
rect 29934 53618 29986 53630
rect 29934 53554 29986 53566
rect 30606 53618 30658 53630
rect 35646 53618 35698 53630
rect 32610 53566 32622 53618
rect 32674 53566 32686 53618
rect 30606 53554 30658 53566
rect 35646 53554 35698 53566
rect 35982 53618 36034 53630
rect 39554 53566 39566 53618
rect 39618 53566 39630 53618
rect 46946 53566 46958 53618
rect 47010 53566 47022 53618
rect 48850 53566 48862 53618
rect 48914 53566 48926 53618
rect 35982 53554 36034 53566
rect 2382 53506 2434 53518
rect 17054 53506 17106 53518
rect 42590 53506 42642 53518
rect 16706 53454 16718 53506
rect 16770 53454 16782 53506
rect 23090 53454 23102 53506
rect 23154 53454 23166 53506
rect 23986 53454 23998 53506
rect 24050 53454 24062 53506
rect 29362 53454 29374 53506
rect 29426 53454 29438 53506
rect 2382 53442 2434 53454
rect 17054 53442 17106 53454
rect 42590 53442 42642 53454
rect 43934 53506 43986 53518
rect 43934 53442 43986 53454
rect 51550 53506 51602 53518
rect 51550 53442 51602 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 3278 53170 3330 53182
rect 7198 53170 7250 53182
rect 6626 53118 6638 53170
rect 6690 53118 6702 53170
rect 3278 53106 3330 53118
rect 7198 53106 7250 53118
rect 11678 53170 11730 53182
rect 22430 53170 22482 53182
rect 30494 53170 30546 53182
rect 41470 53170 41522 53182
rect 16034 53118 16046 53170
rect 16098 53118 16110 53170
rect 28354 53118 28366 53170
rect 28418 53118 28430 53170
rect 31266 53118 31278 53170
rect 31330 53118 31342 53170
rect 11678 53106 11730 53118
rect 22430 53106 22482 53118
rect 30494 53106 30546 53118
rect 41470 53106 41522 53118
rect 44158 53170 44210 53182
rect 44158 53106 44210 53118
rect 47070 53170 47122 53182
rect 47070 53106 47122 53118
rect 47518 53170 47570 53182
rect 47518 53106 47570 53118
rect 48078 53170 48130 53182
rect 48078 53106 48130 53118
rect 3502 53058 3554 53070
rect 3502 52994 3554 53006
rect 6078 53058 6130 53070
rect 6078 52994 6130 53006
rect 6190 53058 6242 53070
rect 6190 52994 6242 53006
rect 10110 53058 10162 53070
rect 30718 53058 30770 53070
rect 23650 53006 23662 53058
rect 23714 53006 23726 53058
rect 23874 53006 23886 53058
rect 23938 53006 23950 53058
rect 10110 52994 10162 53006
rect 30718 52994 30770 53006
rect 41358 53058 41410 53070
rect 41358 52994 41410 53006
rect 41582 53058 41634 53070
rect 41582 52994 41634 53006
rect 42030 53058 42082 53070
rect 42030 52994 42082 53006
rect 44382 53058 44434 53070
rect 44382 52994 44434 53006
rect 44494 53058 44546 53070
rect 44494 52994 44546 53006
rect 44830 53058 44882 53070
rect 44830 52994 44882 53006
rect 47966 53058 48018 53070
rect 47966 52994 48018 53006
rect 48750 53058 48802 53070
rect 49858 53006 49870 53058
rect 49922 53006 49934 53058
rect 48750 52994 48802 53006
rect 6862 52946 6914 52958
rect 5842 52894 5854 52946
rect 5906 52894 5918 52946
rect 6862 52882 6914 52894
rect 7310 52946 7362 52958
rect 7310 52882 7362 52894
rect 7422 52946 7474 52958
rect 11454 52946 11506 52958
rect 10546 52894 10558 52946
rect 10610 52894 10622 52946
rect 7422 52882 7474 52894
rect 11454 52882 11506 52894
rect 11678 52946 11730 52958
rect 11678 52882 11730 52894
rect 11902 52946 11954 52958
rect 11902 52882 11954 52894
rect 15822 52946 15874 52958
rect 15822 52882 15874 52894
rect 16158 52946 16210 52958
rect 22878 52946 22930 52958
rect 16594 52894 16606 52946
rect 16658 52894 16670 52946
rect 18274 52894 18286 52946
rect 18338 52894 18350 52946
rect 19170 52894 19182 52946
rect 19234 52894 19246 52946
rect 16158 52882 16210 52894
rect 22878 52882 22930 52894
rect 28030 52946 28082 52958
rect 28030 52882 28082 52894
rect 28590 52946 28642 52958
rect 28590 52882 28642 52894
rect 28926 52946 28978 52958
rect 28926 52882 28978 52894
rect 29150 52946 29202 52958
rect 29150 52882 29202 52894
rect 29598 52946 29650 52958
rect 42142 52946 42194 52958
rect 33170 52894 33182 52946
rect 33234 52894 33246 52946
rect 38994 52894 39006 52946
rect 39058 52894 39070 52946
rect 29598 52882 29650 52894
rect 42142 52882 42194 52894
rect 48974 52946 49026 52958
rect 48974 52882 49026 52894
rect 49422 52946 49474 52958
rect 49422 52882 49474 52894
rect 50206 52946 50258 52958
rect 53778 52894 53790 52946
rect 53842 52894 53854 52946
rect 50206 52882 50258 52894
rect 5182 52834 5234 52846
rect 13134 52834 13186 52846
rect 18734 52834 18786 52846
rect 27806 52834 27858 52846
rect 3154 52782 3166 52834
rect 3218 52782 3230 52834
rect 10434 52782 10446 52834
rect 10498 52782 10510 52834
rect 17938 52782 17950 52834
rect 18002 52782 18014 52834
rect 19842 52782 19854 52834
rect 19906 52782 19918 52834
rect 21970 52782 21982 52834
rect 22034 52782 22046 52834
rect 5182 52770 5234 52782
rect 13134 52770 13186 52782
rect 18734 52770 18786 52782
rect 27806 52770 27858 52782
rect 28814 52834 28866 52846
rect 39454 52834 39506 52846
rect 33842 52782 33854 52834
rect 33906 52782 33918 52834
rect 35970 52782 35982 52834
rect 36034 52782 36046 52834
rect 28814 52770 28866 52782
rect 39454 52770 39506 52782
rect 40462 52834 40514 52846
rect 40462 52770 40514 52782
rect 48190 52834 48242 52846
rect 48190 52770 48242 52782
rect 48862 52834 48914 52846
rect 50866 52782 50878 52834
rect 50930 52782 50942 52834
rect 52994 52782 53006 52834
rect 53058 52782 53070 52834
rect 48862 52770 48914 52782
rect 5070 52722 5122 52734
rect 5070 52658 5122 52670
rect 5406 52722 5458 52734
rect 5406 52658 5458 52670
rect 5518 52722 5570 52734
rect 5518 52658 5570 52670
rect 16270 52722 16322 52734
rect 16270 52658 16322 52670
rect 22990 52722 23042 52734
rect 22990 52658 23042 52670
rect 24222 52722 24274 52734
rect 24222 52658 24274 52670
rect 24558 52722 24610 52734
rect 24558 52658 24610 52670
rect 29822 52722 29874 52734
rect 29822 52658 29874 52670
rect 30046 52722 30098 52734
rect 30046 52658 30098 52670
rect 30942 52722 30994 52734
rect 30942 52658 30994 52670
rect 42030 52722 42082 52734
rect 42030 52658 42082 52670
rect 44942 52722 44994 52734
rect 44942 52658 44994 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 6974 52386 7026 52398
rect 6402 52334 6414 52386
rect 6466 52334 6478 52386
rect 6974 52322 7026 52334
rect 7086 52386 7138 52398
rect 7086 52322 7138 52334
rect 7422 52386 7474 52398
rect 7422 52322 7474 52334
rect 17950 52386 18002 52398
rect 17950 52322 18002 52334
rect 19406 52386 19458 52398
rect 19406 52322 19458 52334
rect 19742 52386 19794 52398
rect 30046 52386 30098 52398
rect 27906 52334 27918 52386
rect 27970 52334 27982 52386
rect 19742 52322 19794 52334
rect 30046 52322 30098 52334
rect 30382 52386 30434 52398
rect 30382 52322 30434 52334
rect 11790 52274 11842 52286
rect 2482 52222 2494 52274
rect 2546 52222 2558 52274
rect 4610 52222 4622 52274
rect 4674 52222 4686 52274
rect 11330 52222 11342 52274
rect 11394 52222 11406 52274
rect 11790 52210 11842 52222
rect 16158 52274 16210 52286
rect 16158 52210 16210 52222
rect 18510 52274 18562 52286
rect 30270 52274 30322 52286
rect 34974 52274 35026 52286
rect 40798 52274 40850 52286
rect 50766 52274 50818 52286
rect 24882 52222 24894 52274
rect 24946 52222 24958 52274
rect 26898 52222 26910 52274
rect 26962 52222 26974 52274
rect 31042 52222 31054 52274
rect 31106 52222 31118 52274
rect 34066 52222 34078 52274
rect 34130 52222 34142 52274
rect 38994 52222 39006 52274
rect 39058 52222 39070 52274
rect 46722 52222 46734 52274
rect 46786 52222 46798 52274
rect 18510 52210 18562 52222
rect 30270 52210 30322 52222
rect 34974 52210 35026 52222
rect 40798 52210 40850 52222
rect 50766 52210 50818 52222
rect 52782 52274 52834 52286
rect 52782 52210 52834 52222
rect 5854 52162 5906 52174
rect 1810 52110 1822 52162
rect 1874 52110 1886 52162
rect 5618 52110 5630 52162
rect 5682 52110 5694 52162
rect 5854 52098 5906 52110
rect 7310 52162 7362 52174
rect 7310 52098 7362 52110
rect 7758 52162 7810 52174
rect 7758 52098 7810 52110
rect 7870 52162 7922 52174
rect 15710 52162 15762 52174
rect 8418 52110 8430 52162
rect 8482 52110 8494 52162
rect 7870 52098 7922 52110
rect 15710 52098 15762 52110
rect 16270 52162 16322 52174
rect 16270 52098 16322 52110
rect 16606 52162 16658 52174
rect 17838 52162 17890 52174
rect 26462 52162 26514 52174
rect 29150 52162 29202 52174
rect 17042 52110 17054 52162
rect 17106 52110 17118 52162
rect 19730 52110 19742 52162
rect 19794 52110 19806 52162
rect 21858 52110 21870 52162
rect 21922 52110 21934 52162
rect 22754 52110 22766 52162
rect 22818 52110 22830 52162
rect 23986 52110 23998 52162
rect 24050 52110 24062 52162
rect 24434 52110 24446 52162
rect 24498 52110 24510 52162
rect 27122 52110 27134 52162
rect 27186 52110 27198 52162
rect 27346 52110 27358 52162
rect 27410 52110 27422 52162
rect 16606 52098 16658 52110
rect 17838 52098 17890 52110
rect 26462 52098 26514 52110
rect 29150 52098 29202 52110
rect 29374 52162 29426 52174
rect 29374 52098 29426 52110
rect 29598 52162 29650 52174
rect 40126 52162 40178 52174
rect 31266 52110 31278 52162
rect 31330 52110 31342 52162
rect 31490 52110 31502 52162
rect 31554 52110 31566 52162
rect 34290 52110 34302 52162
rect 34354 52110 34366 52162
rect 38882 52110 38894 52162
rect 38946 52110 38958 52162
rect 29598 52098 29650 52110
rect 40126 52098 40178 52110
rect 40910 52162 40962 52174
rect 40910 52098 40962 52110
rect 41358 52162 41410 52174
rect 41358 52098 41410 52110
rect 41582 52162 41634 52174
rect 42142 52162 42194 52174
rect 44942 52162 44994 52174
rect 48078 52162 48130 52174
rect 49310 52162 49362 52174
rect 41794 52110 41806 52162
rect 41858 52110 41870 52162
rect 44034 52110 44046 52162
rect 44098 52110 44110 52162
rect 45154 52110 45166 52162
rect 45218 52110 45230 52162
rect 46610 52110 46622 52162
rect 46674 52110 46686 52162
rect 47730 52110 47742 52162
rect 47794 52110 47806 52162
rect 48514 52110 48526 52162
rect 48578 52110 48590 52162
rect 41582 52098 41634 52110
rect 42142 52098 42194 52110
rect 44942 52098 44994 52110
rect 48078 52098 48130 52110
rect 49310 52098 49362 52110
rect 49646 52162 49698 52174
rect 50878 52162 50930 52174
rect 50530 52110 50542 52162
rect 50594 52110 50606 52162
rect 49646 52098 49698 52110
rect 50878 52098 50930 52110
rect 51326 52162 51378 52174
rect 51326 52098 51378 52110
rect 51886 52162 51938 52174
rect 51886 52098 51938 52110
rect 5966 52050 6018 52062
rect 11902 52050 11954 52062
rect 9202 51998 9214 52050
rect 9266 51998 9278 52050
rect 5966 51986 6018 51998
rect 11902 51986 11954 51998
rect 15486 52050 15538 52062
rect 15486 51986 15538 51998
rect 16046 52050 16098 52062
rect 16046 51986 16098 51998
rect 17950 52050 18002 52062
rect 39454 52050 39506 52062
rect 21970 51998 21982 52050
rect 22034 51998 22046 52050
rect 24658 51998 24670 52050
rect 24722 51998 24734 52050
rect 33282 51998 33294 52050
rect 33346 51998 33358 52050
rect 17950 51986 18002 51998
rect 39454 51986 39506 51998
rect 40350 52050 40402 52062
rect 40350 51986 40402 51998
rect 42702 52050 42754 52062
rect 42702 51986 42754 51998
rect 45838 52050 45890 52062
rect 48974 52050 49026 52062
rect 46386 51998 46398 52050
rect 46450 51998 46462 52050
rect 45838 51986 45890 51998
rect 48974 51986 49026 51998
rect 49870 52050 49922 52062
rect 49870 51986 49922 51998
rect 51438 52050 51490 52062
rect 51438 51986 51490 51998
rect 11678 51938 11730 51950
rect 11678 51874 11730 51886
rect 12126 51938 12178 51950
rect 12126 51874 12178 51886
rect 15598 51938 15650 51950
rect 15598 51874 15650 51886
rect 17278 51938 17330 51950
rect 17278 51874 17330 51886
rect 17502 51938 17554 51950
rect 17502 51874 17554 51886
rect 17614 51938 17666 51950
rect 17614 51874 17666 51886
rect 18398 51938 18450 51950
rect 25902 51938 25954 51950
rect 22642 51886 22654 51938
rect 22706 51886 22718 51938
rect 18398 51874 18450 51886
rect 25902 51874 25954 51886
rect 32286 51938 32338 51950
rect 32286 51874 32338 51886
rect 33630 51938 33682 51950
rect 41694 51938 41746 51950
rect 39778 51886 39790 51938
rect 39842 51886 39854 51938
rect 33630 51874 33682 51886
rect 41694 51874 41746 51886
rect 43262 51938 43314 51950
rect 49534 51938 49586 51950
rect 44258 51886 44270 51938
rect 44322 51886 44334 51938
rect 43262 51874 43314 51886
rect 49534 51874 49586 51886
rect 51214 51938 51266 51950
rect 51214 51874 51266 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 5070 51602 5122 51614
rect 5070 51538 5122 51550
rect 6974 51602 7026 51614
rect 6974 51538 7026 51550
rect 7198 51602 7250 51614
rect 7198 51538 7250 51550
rect 9998 51602 10050 51614
rect 16494 51602 16546 51614
rect 10994 51550 11006 51602
rect 11058 51550 11070 51602
rect 9998 51538 10050 51550
rect 16494 51538 16546 51550
rect 22542 51602 22594 51614
rect 22542 51538 22594 51550
rect 27246 51602 27298 51614
rect 27246 51538 27298 51550
rect 28926 51602 28978 51614
rect 28926 51538 28978 51550
rect 32174 51602 32226 51614
rect 32174 51538 32226 51550
rect 33182 51602 33234 51614
rect 33182 51538 33234 51550
rect 33406 51602 33458 51614
rect 34190 51602 34242 51614
rect 33842 51550 33854 51602
rect 33906 51550 33918 51602
rect 33406 51538 33458 51550
rect 34190 51538 34242 51550
rect 39902 51602 39954 51614
rect 39902 51538 39954 51550
rect 41694 51602 41746 51614
rect 41694 51538 41746 51550
rect 43150 51602 43202 51614
rect 43150 51538 43202 51550
rect 46846 51602 46898 51614
rect 46846 51538 46898 51550
rect 48750 51602 48802 51614
rect 48750 51538 48802 51550
rect 4622 51490 4674 51502
rect 4622 51426 4674 51438
rect 5182 51490 5234 51502
rect 5182 51426 5234 51438
rect 6750 51490 6802 51502
rect 16718 51490 16770 51502
rect 10770 51438 10782 51490
rect 10834 51438 10846 51490
rect 12338 51438 12350 51490
rect 12402 51438 12414 51490
rect 6750 51426 6802 51438
rect 16718 51426 16770 51438
rect 16830 51490 16882 51502
rect 16830 51426 16882 51438
rect 23214 51490 23266 51502
rect 23214 51426 23266 51438
rect 23326 51490 23378 51502
rect 23326 51426 23378 51438
rect 23886 51490 23938 51502
rect 23886 51426 23938 51438
rect 25454 51490 25506 51502
rect 25454 51426 25506 51438
rect 25566 51490 25618 51502
rect 25566 51426 25618 51438
rect 26462 51490 26514 51502
rect 26462 51426 26514 51438
rect 27134 51490 27186 51502
rect 27134 51426 27186 51438
rect 27694 51490 27746 51502
rect 27694 51426 27746 51438
rect 28702 51490 28754 51502
rect 28702 51426 28754 51438
rect 31838 51490 31890 51502
rect 31838 51426 31890 51438
rect 32398 51490 32450 51502
rect 37102 51490 37154 51502
rect 40350 51490 40402 51502
rect 36194 51438 36206 51490
rect 36258 51438 36270 51490
rect 39666 51438 39678 51490
rect 39730 51438 39742 51490
rect 32398 51426 32450 51438
rect 37102 51426 37154 51438
rect 40350 51426 40402 51438
rect 40910 51490 40962 51502
rect 40910 51426 40962 51438
rect 41022 51490 41074 51502
rect 51662 51490 51714 51502
rect 43698 51438 43710 51490
rect 43762 51438 43774 51490
rect 47282 51438 47294 51490
rect 47346 51438 47358 51490
rect 51986 51438 51998 51490
rect 52050 51438 52062 51490
rect 41022 51426 41074 51438
rect 51662 51426 51714 51438
rect 4846 51378 4898 51390
rect 5854 51378 5906 51390
rect 5618 51326 5630 51378
rect 5682 51326 5694 51378
rect 4846 51314 4898 51326
rect 5854 51314 5906 51326
rect 6078 51378 6130 51390
rect 6078 51314 6130 51326
rect 9886 51378 9938 51390
rect 9886 51314 9938 51326
rect 10222 51378 10274 51390
rect 10222 51314 10274 51326
rect 10446 51378 10498 51390
rect 23550 51378 23602 51390
rect 11442 51326 11454 51378
rect 11506 51326 11518 51378
rect 12450 51326 12462 51378
rect 12514 51326 12526 51378
rect 13122 51326 13134 51378
rect 13186 51326 13198 51378
rect 17602 51326 17614 51378
rect 17666 51326 17678 51378
rect 18050 51326 18062 51378
rect 18114 51326 18126 51378
rect 19282 51326 19294 51378
rect 19346 51326 19358 51378
rect 10446 51314 10498 51326
rect 23550 51314 23602 51326
rect 23774 51378 23826 51390
rect 31726 51378 31778 51390
rect 28242 51326 28254 51378
rect 28306 51326 28318 51378
rect 23774 51314 23826 51326
rect 31726 51314 31778 51326
rect 32510 51378 32562 51390
rect 32510 51314 32562 51326
rect 33070 51378 33122 51390
rect 33070 51314 33122 51326
rect 35870 51378 35922 51390
rect 35870 51314 35922 51326
rect 36542 51378 36594 51390
rect 36542 51314 36594 51326
rect 37438 51378 37490 51390
rect 37438 51314 37490 51326
rect 37886 51378 37938 51390
rect 37886 51314 37938 51326
rect 38110 51378 38162 51390
rect 40126 51378 40178 51390
rect 39442 51326 39454 51378
rect 39506 51326 39518 51378
rect 38110 51314 38162 51326
rect 40126 51314 40178 51326
rect 41246 51378 41298 51390
rect 41246 51314 41298 51326
rect 41918 51378 41970 51390
rect 41918 51314 41970 51326
rect 42142 51378 42194 51390
rect 42142 51314 42194 51326
rect 42366 51378 42418 51390
rect 43262 51378 43314 51390
rect 42914 51326 42926 51378
rect 42978 51326 42990 51378
rect 42366 51314 42418 51326
rect 43262 51314 43314 51326
rect 45278 51378 45330 51390
rect 45278 51314 45330 51326
rect 45726 51378 45778 51390
rect 49198 51378 49250 51390
rect 48850 51326 48862 51378
rect 48914 51326 48926 51378
rect 45726 51314 45778 51326
rect 49198 51314 49250 51326
rect 49534 51378 49586 51390
rect 53902 51378 53954 51390
rect 50754 51326 50766 51378
rect 50818 51326 50830 51378
rect 51874 51326 51886 51378
rect 51938 51326 51950 51378
rect 49534 51314 49586 51326
rect 53902 51314 53954 51326
rect 17390 51266 17442 51278
rect 27806 51266 27858 51278
rect 39230 51266 39282 51278
rect 13906 51214 13918 51266
rect 13970 51214 13982 51266
rect 16034 51214 16046 51266
rect 16098 51214 16110 51266
rect 19954 51214 19966 51266
rect 20018 51214 20030 51266
rect 22082 51214 22094 51266
rect 22146 51214 22158 51266
rect 26338 51214 26350 51266
rect 26402 51214 26414 51266
rect 29026 51214 29038 51266
rect 29090 51214 29102 51266
rect 17390 51202 17442 51214
rect 27806 51202 27858 51214
rect 39230 51202 39282 51214
rect 41806 51266 41858 51278
rect 41806 51202 41858 51214
rect 47966 51266 48018 51278
rect 47966 51202 48018 51214
rect 50094 51266 50146 51278
rect 53342 51266 53394 51278
rect 50866 51214 50878 51266
rect 50930 51214 50942 51266
rect 52546 51214 52558 51266
rect 52610 51214 52622 51266
rect 50094 51202 50146 51214
rect 53342 51202 53394 51214
rect 6190 51154 6242 51166
rect 6190 51090 6242 51102
rect 7310 51154 7362 51166
rect 7310 51090 7362 51102
rect 23886 51154 23938 51166
rect 23886 51090 23938 51102
rect 25566 51154 25618 51166
rect 25566 51090 25618 51102
rect 26686 51154 26738 51166
rect 26686 51090 26738 51102
rect 27358 51154 27410 51166
rect 27358 51090 27410 51102
rect 28030 51154 28082 51166
rect 28030 51090 28082 51102
rect 31838 51154 31890 51166
rect 31838 51090 31890 51102
rect 37662 51154 37714 51166
rect 37662 51090 37714 51102
rect 38558 51154 38610 51166
rect 38558 51090 38610 51102
rect 39902 51154 39954 51166
rect 39902 51090 39954 51102
rect 49086 51154 49138 51166
rect 49086 51090 49138 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 25566 50818 25618 50830
rect 15586 50766 15598 50818
rect 15650 50815 15662 50818
rect 16034 50815 16046 50818
rect 15650 50769 16046 50815
rect 15650 50766 15662 50769
rect 16034 50766 16046 50769
rect 16098 50766 16110 50818
rect 16818 50766 16830 50818
rect 16882 50766 16894 50818
rect 25566 50754 25618 50766
rect 25902 50818 25954 50830
rect 25902 50754 25954 50766
rect 27134 50818 27186 50830
rect 27134 50754 27186 50766
rect 27470 50818 27522 50830
rect 27470 50754 27522 50766
rect 28142 50818 28194 50830
rect 28142 50754 28194 50766
rect 28590 50818 28642 50830
rect 28590 50754 28642 50766
rect 30382 50818 30434 50830
rect 30382 50754 30434 50766
rect 38670 50818 38722 50830
rect 38670 50754 38722 50766
rect 39006 50818 39058 50830
rect 39006 50754 39058 50766
rect 50766 50818 50818 50830
rect 50766 50754 50818 50766
rect 11342 50706 11394 50718
rect 4610 50654 4622 50706
rect 4674 50654 4686 50706
rect 6402 50654 6414 50706
rect 6466 50654 6478 50706
rect 11342 50642 11394 50654
rect 15934 50706 15986 50718
rect 15934 50642 15986 50654
rect 18174 50706 18226 50718
rect 22766 50706 22818 50718
rect 20066 50654 20078 50706
rect 20130 50654 20142 50706
rect 18174 50642 18226 50654
rect 22766 50642 22818 50654
rect 28478 50706 28530 50718
rect 40238 50706 40290 50718
rect 49422 50706 49474 50718
rect 31826 50654 31838 50706
rect 31890 50654 31902 50706
rect 32498 50654 32510 50706
rect 32562 50654 32574 50706
rect 36418 50654 36430 50706
rect 36482 50654 36494 50706
rect 37986 50654 37998 50706
rect 38050 50654 38062 50706
rect 46722 50654 46734 50706
rect 46786 50654 46798 50706
rect 54450 50654 54462 50706
rect 54514 50654 54526 50706
rect 28478 50642 28530 50654
rect 40238 50642 40290 50654
rect 49422 50642 49474 50654
rect 10894 50594 10946 50606
rect 1810 50542 1822 50594
rect 1874 50542 1886 50594
rect 5730 50542 5742 50594
rect 5794 50542 5806 50594
rect 10894 50530 10946 50542
rect 11230 50594 11282 50606
rect 11230 50530 11282 50542
rect 11454 50594 11506 50606
rect 11454 50530 11506 50542
rect 11902 50594 11954 50606
rect 16270 50594 16322 50606
rect 12226 50542 12238 50594
rect 12290 50542 12302 50594
rect 11902 50530 11954 50542
rect 16270 50530 16322 50542
rect 16606 50594 16658 50606
rect 17726 50594 17778 50606
rect 17042 50542 17054 50594
rect 17106 50542 17118 50594
rect 16606 50530 16658 50542
rect 17726 50530 17778 50542
rect 18958 50594 19010 50606
rect 22654 50594 22706 50606
rect 23998 50594 24050 50606
rect 19954 50542 19966 50594
rect 20018 50542 20030 50594
rect 21522 50542 21534 50594
rect 21586 50542 21598 50594
rect 23762 50542 23774 50594
rect 23826 50542 23838 50594
rect 18958 50530 19010 50542
rect 22654 50530 22706 50542
rect 23998 50530 24050 50542
rect 24110 50594 24162 50606
rect 24110 50530 24162 50542
rect 26798 50594 26850 50606
rect 28254 50594 28306 50606
rect 30270 50594 30322 50606
rect 32174 50594 32226 50606
rect 40014 50594 40066 50606
rect 44158 50594 44210 50606
rect 27122 50542 27134 50594
rect 27186 50542 27198 50594
rect 29698 50542 29710 50594
rect 29762 50542 29774 50594
rect 31266 50542 31278 50594
rect 31330 50542 31342 50594
rect 33618 50542 33630 50594
rect 33682 50542 33694 50594
rect 40674 50542 40686 50594
rect 40738 50542 40750 50594
rect 41682 50542 41694 50594
rect 41746 50542 41758 50594
rect 42466 50542 42478 50594
rect 42530 50542 42542 50594
rect 26798 50530 26850 50542
rect 28254 50530 28306 50542
rect 30270 50530 30322 50542
rect 32174 50530 32226 50542
rect 40014 50530 40066 50542
rect 44158 50530 44210 50542
rect 46510 50594 46562 50606
rect 50878 50594 50930 50606
rect 46834 50542 46846 50594
rect 46898 50542 46910 50594
rect 46510 50530 46562 50542
rect 50878 50530 50930 50542
rect 51102 50594 51154 50606
rect 53006 50594 53058 50606
rect 51314 50542 51326 50594
rect 51378 50542 51390 50594
rect 52770 50542 52782 50594
rect 52834 50542 52846 50594
rect 54562 50542 54574 50594
rect 54626 50542 54638 50594
rect 54898 50542 54910 50594
rect 54962 50542 54974 50594
rect 51102 50530 51154 50542
rect 53006 50530 53058 50542
rect 10110 50482 10162 50494
rect 2482 50430 2494 50482
rect 2546 50430 2558 50482
rect 9762 50430 9774 50482
rect 9826 50430 9838 50482
rect 10110 50418 10162 50430
rect 10782 50482 10834 50494
rect 10782 50418 10834 50430
rect 12462 50482 12514 50494
rect 18846 50482 18898 50494
rect 17378 50430 17390 50482
rect 17442 50430 17454 50482
rect 12462 50418 12514 50430
rect 18846 50418 18898 50430
rect 19294 50482 19346 50494
rect 19294 50418 19346 50430
rect 22430 50482 22482 50494
rect 25342 50482 25394 50494
rect 24546 50430 24558 50482
rect 24610 50430 24622 50482
rect 22430 50418 22482 50430
rect 25342 50418 25394 50430
rect 26238 50482 26290 50494
rect 26238 50418 26290 50430
rect 29150 50482 29202 50494
rect 30494 50482 30546 50494
rect 29922 50430 29934 50482
rect 29986 50430 29998 50482
rect 29150 50418 29202 50430
rect 30494 50418 30546 50430
rect 30942 50482 30994 50494
rect 30942 50418 30994 50430
rect 31502 50482 31554 50494
rect 31502 50418 31554 50430
rect 33182 50482 33234 50494
rect 37550 50482 37602 50494
rect 34290 50430 34302 50482
rect 34354 50430 34366 50482
rect 33182 50418 33234 50430
rect 37550 50418 37602 50430
rect 38446 50482 38498 50494
rect 38446 50418 38498 50430
rect 39566 50482 39618 50494
rect 39566 50418 39618 50430
rect 39790 50482 39842 50494
rect 39790 50418 39842 50430
rect 40350 50482 40402 50494
rect 43822 50482 43874 50494
rect 41906 50430 41918 50482
rect 41970 50430 41982 50482
rect 42690 50430 42702 50482
rect 42754 50430 42766 50482
rect 43250 50430 43262 50482
rect 43314 50430 43326 50482
rect 40350 50418 40402 50430
rect 43822 50418 43874 50430
rect 44046 50482 44098 50494
rect 44046 50418 44098 50430
rect 45390 50482 45442 50494
rect 45390 50418 45442 50430
rect 47406 50482 47458 50494
rect 47406 50418 47458 50430
rect 49534 50482 49586 50494
rect 49534 50418 49586 50430
rect 49870 50482 49922 50494
rect 49870 50418 49922 50430
rect 50318 50482 50370 50494
rect 50318 50418 50370 50430
rect 51774 50482 51826 50494
rect 51774 50418 51826 50430
rect 16382 50370 16434 50382
rect 8642 50318 8654 50370
rect 8706 50318 8718 50370
rect 16382 50306 16434 50318
rect 21310 50370 21362 50382
rect 21310 50306 21362 50318
rect 22878 50370 22930 50382
rect 22878 50306 22930 50318
rect 29262 50370 29314 50382
rect 29262 50306 29314 50318
rect 30718 50370 30770 50382
rect 30718 50306 30770 50318
rect 31726 50370 31778 50382
rect 31726 50306 31778 50318
rect 31838 50370 31890 50382
rect 31838 50306 31890 50318
rect 32510 50370 32562 50382
rect 32510 50306 32562 50318
rect 32734 50370 32786 50382
rect 32734 50306 32786 50318
rect 33070 50370 33122 50382
rect 43598 50370 43650 50382
rect 41794 50318 41806 50370
rect 41858 50318 41870 50370
rect 33070 50306 33122 50318
rect 43598 50306 43650 50318
rect 49086 50370 49138 50382
rect 49086 50306 49138 50318
rect 49310 50370 49362 50382
rect 49310 50306 49362 50318
rect 49982 50370 50034 50382
rect 49982 50306 50034 50318
rect 50094 50370 50146 50382
rect 50094 50306 50146 50318
rect 53342 50370 53394 50382
rect 55010 50318 55022 50370
rect 55074 50318 55086 50370
rect 53342 50306 53394 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 2046 50034 2098 50046
rect 2046 49970 2098 49982
rect 2158 50034 2210 50046
rect 9662 50034 9714 50046
rect 19070 50034 19122 50046
rect 6290 49982 6302 50034
rect 6354 49982 6366 50034
rect 7634 49982 7646 50034
rect 7698 49982 7710 50034
rect 17378 49982 17390 50034
rect 17442 49982 17454 50034
rect 2158 49970 2210 49982
rect 9662 49970 9714 49982
rect 19070 49970 19122 49982
rect 22430 50034 22482 50046
rect 28814 50034 28866 50046
rect 26562 49982 26574 50034
rect 26626 49982 26638 50034
rect 22430 49970 22482 49982
rect 28814 49970 28866 49982
rect 29486 50034 29538 50046
rect 29486 49970 29538 49982
rect 32622 50034 32674 50046
rect 32622 49970 32674 49982
rect 33070 50034 33122 50046
rect 33070 49970 33122 49982
rect 33182 50034 33234 50046
rect 33182 49970 33234 49982
rect 40238 50034 40290 50046
rect 40238 49970 40290 49982
rect 40798 50034 40850 50046
rect 40798 49970 40850 49982
rect 42702 50034 42754 50046
rect 42702 49970 42754 49982
rect 46286 50034 46338 50046
rect 46286 49970 46338 49982
rect 9550 49922 9602 49934
rect 4946 49870 4958 49922
rect 5010 49870 5022 49922
rect 6402 49870 6414 49922
rect 6466 49870 6478 49922
rect 9550 49858 9602 49870
rect 10670 49922 10722 49934
rect 10670 49858 10722 49870
rect 16606 49922 16658 49934
rect 16606 49858 16658 49870
rect 19518 49922 19570 49934
rect 19518 49858 19570 49870
rect 22542 49922 22594 49934
rect 24782 49922 24834 49934
rect 23874 49870 23886 49922
rect 23938 49870 23950 49922
rect 24434 49870 24446 49922
rect 24498 49870 24510 49922
rect 22542 49858 22594 49870
rect 24782 49858 24834 49870
rect 27358 49922 27410 49934
rect 27358 49858 27410 49870
rect 27582 49922 27634 49934
rect 33294 49922 33346 49934
rect 28018 49870 28030 49922
rect 28082 49870 28094 49922
rect 30370 49870 30382 49922
rect 30434 49870 30446 49922
rect 31266 49870 31278 49922
rect 31330 49870 31342 49922
rect 27582 49858 27634 49870
rect 33294 49858 33346 49870
rect 33406 49922 33458 49934
rect 36542 49922 36594 49934
rect 40126 49922 40178 49934
rect 33618 49870 33630 49922
rect 33682 49870 33694 49922
rect 37314 49870 37326 49922
rect 37378 49870 37390 49922
rect 33406 49858 33458 49870
rect 36542 49858 36594 49870
rect 40126 49858 40178 49870
rect 42590 49922 42642 49934
rect 45614 49922 45666 49934
rect 43138 49870 43150 49922
rect 43202 49870 43214 49922
rect 44594 49870 44606 49922
rect 44658 49870 44670 49922
rect 45266 49870 45278 49922
rect 45330 49870 45342 49922
rect 42590 49858 42642 49870
rect 45614 49858 45666 49870
rect 47966 49922 48018 49934
rect 47966 49858 48018 49870
rect 50206 49922 50258 49934
rect 50206 49858 50258 49870
rect 56702 49922 56754 49934
rect 56702 49858 56754 49870
rect 2270 49810 2322 49822
rect 2270 49746 2322 49758
rect 2606 49810 2658 49822
rect 6974 49810 7026 49822
rect 3490 49758 3502 49810
rect 3554 49758 3566 49810
rect 4834 49758 4846 49810
rect 4898 49758 4910 49810
rect 5842 49758 5854 49810
rect 5906 49758 5918 49810
rect 2606 49746 2658 49758
rect 6974 49746 7026 49758
rect 7086 49810 7138 49822
rect 7086 49746 7138 49758
rect 7198 49810 7250 49822
rect 7198 49746 7250 49758
rect 11006 49810 11058 49822
rect 11006 49746 11058 49758
rect 11566 49810 11618 49822
rect 11566 49746 11618 49758
rect 11902 49810 11954 49822
rect 11902 49746 11954 49758
rect 12350 49810 12402 49822
rect 12350 49746 12402 49758
rect 12462 49810 12514 49822
rect 12462 49746 12514 49758
rect 12574 49810 12626 49822
rect 12574 49746 12626 49758
rect 12798 49810 12850 49822
rect 12798 49746 12850 49758
rect 16830 49810 16882 49822
rect 16830 49746 16882 49758
rect 17726 49810 17778 49822
rect 17726 49746 17778 49758
rect 18734 49810 18786 49822
rect 18734 49746 18786 49758
rect 18958 49810 19010 49822
rect 19742 49810 19794 49822
rect 19170 49758 19182 49810
rect 19234 49758 19246 49810
rect 18958 49746 19010 49758
rect 19742 49746 19794 49758
rect 20078 49810 20130 49822
rect 20078 49746 20130 49758
rect 20638 49810 20690 49822
rect 22206 49810 22258 49822
rect 26126 49810 26178 49822
rect 27470 49810 27522 49822
rect 21298 49758 21310 49810
rect 21362 49758 21374 49810
rect 21634 49758 21646 49810
rect 21698 49758 21710 49810
rect 21858 49758 21870 49810
rect 21922 49758 21934 49810
rect 23650 49758 23662 49810
rect 23714 49758 23726 49810
rect 26226 49758 26238 49810
rect 26290 49758 26302 49810
rect 20638 49746 20690 49758
rect 22206 49746 22258 49758
rect 26126 49746 26178 49758
rect 27470 49746 27522 49758
rect 28254 49810 28306 49822
rect 28254 49746 28306 49758
rect 28702 49810 28754 49822
rect 28702 49746 28754 49758
rect 28926 49810 28978 49822
rect 28926 49746 28978 49758
rect 29374 49810 29426 49822
rect 29374 49746 29426 49758
rect 29598 49810 29650 49822
rect 29598 49746 29650 49758
rect 30046 49810 30098 49822
rect 45950 49810 46002 49822
rect 30594 49758 30606 49810
rect 30658 49758 30670 49810
rect 31154 49758 31166 49810
rect 31218 49758 31230 49810
rect 32050 49758 32062 49810
rect 32114 49758 32126 49810
rect 34402 49758 34414 49810
rect 34466 49758 34478 49810
rect 37874 49758 37886 49810
rect 37938 49758 37950 49810
rect 38658 49758 38670 49810
rect 38722 49758 38734 49810
rect 41458 49758 41470 49810
rect 41522 49758 41534 49810
rect 41794 49758 41806 49810
rect 41858 49758 41870 49810
rect 43586 49758 43598 49810
rect 43650 49758 43662 49810
rect 44034 49758 44046 49810
rect 44098 49758 44110 49810
rect 30046 49746 30098 49758
rect 45950 49746 46002 49758
rect 46286 49810 46338 49822
rect 46286 49746 46338 49758
rect 46622 49810 46674 49822
rect 46622 49746 46674 49758
rect 46846 49810 46898 49822
rect 46846 49746 46898 49758
rect 46958 49810 47010 49822
rect 46958 49746 47010 49758
rect 47070 49810 47122 49822
rect 47070 49746 47122 49758
rect 47518 49810 47570 49822
rect 47518 49746 47570 49758
rect 48750 49810 48802 49822
rect 51774 49810 51826 49822
rect 49298 49758 49310 49810
rect 49362 49758 49374 49810
rect 49634 49758 49646 49810
rect 49698 49758 49710 49810
rect 51538 49758 51550 49810
rect 51602 49758 51614 49810
rect 48750 49746 48802 49758
rect 51774 49746 51826 49758
rect 52670 49810 52722 49822
rect 52670 49746 52722 49758
rect 53118 49810 53170 49822
rect 54574 49810 54626 49822
rect 56478 49810 56530 49822
rect 53778 49758 53790 49810
rect 53842 49758 53854 49810
rect 54674 49758 54686 49810
rect 54738 49758 54750 49810
rect 55234 49758 55246 49810
rect 55298 49758 55310 49810
rect 53118 49746 53170 49758
rect 54574 49746 54626 49758
rect 56478 49746 56530 49758
rect 56814 49810 56866 49822
rect 56814 49746 56866 49758
rect 17950 49698 18002 49710
rect 3378 49646 3390 49698
rect 3442 49646 3454 49698
rect 17950 49634 18002 49646
rect 19966 49698 20018 49710
rect 39230 49698 39282 49710
rect 48078 49698 48130 49710
rect 26674 49646 26686 49698
rect 26738 49646 26750 49698
rect 34178 49646 34190 49698
rect 34242 49646 34254 49698
rect 36642 49646 36654 49698
rect 36706 49646 36718 49698
rect 41906 49646 41918 49698
rect 41970 49646 41982 49698
rect 44146 49646 44158 49698
rect 44210 49646 44222 49698
rect 19966 49634 20018 49646
rect 39230 49634 39282 49646
rect 48078 49634 48130 49646
rect 50094 49698 50146 49710
rect 50094 49634 50146 49646
rect 50878 49698 50930 49710
rect 50878 49634 50930 49646
rect 52782 49698 52834 49710
rect 54462 49698 54514 49710
rect 54114 49646 54126 49698
rect 54178 49646 54190 49698
rect 52782 49634 52834 49646
rect 54462 49634 54514 49646
rect 9662 49586 9714 49598
rect 9662 49522 9714 49534
rect 11454 49586 11506 49598
rect 11454 49522 11506 49534
rect 11790 49586 11842 49598
rect 11790 49522 11842 49534
rect 16494 49586 16546 49598
rect 16494 49522 16546 49534
rect 36318 49586 36370 49598
rect 36318 49522 36370 49534
rect 40350 49586 40402 49598
rect 40350 49522 40402 49534
rect 48190 49586 48242 49598
rect 48190 49522 48242 49534
rect 48862 49586 48914 49598
rect 48862 49522 48914 49534
rect 49086 49586 49138 49598
rect 49086 49522 49138 49534
rect 49870 49586 49922 49598
rect 49870 49522 49922 49534
rect 53006 49586 53058 49598
rect 53006 49522 53058 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 2718 49250 2770 49262
rect 2718 49186 2770 49198
rect 18846 49250 18898 49262
rect 23662 49250 23714 49262
rect 20178 49198 20190 49250
rect 20242 49198 20254 49250
rect 18846 49186 18898 49198
rect 23662 49186 23714 49198
rect 26574 49250 26626 49262
rect 26574 49186 26626 49198
rect 27806 49250 27858 49262
rect 27806 49186 27858 49198
rect 29262 49250 29314 49262
rect 47294 49250 47346 49262
rect 45490 49198 45502 49250
rect 45554 49198 45566 49250
rect 52882 49198 52894 49250
rect 52946 49198 52958 49250
rect 29262 49186 29314 49198
rect 47294 49186 47346 49198
rect 5742 49138 5794 49150
rect 28590 49138 28642 49150
rect 10322 49086 10334 49138
rect 10386 49086 10398 49138
rect 17154 49086 17166 49138
rect 17218 49086 17230 49138
rect 26786 49086 26798 49138
rect 26850 49086 26862 49138
rect 5742 49074 5794 49086
rect 28590 49074 28642 49086
rect 29822 49138 29874 49150
rect 32174 49138 32226 49150
rect 42590 49138 42642 49150
rect 30818 49086 30830 49138
rect 30882 49086 30894 49138
rect 37202 49086 37214 49138
rect 37266 49086 37278 49138
rect 40226 49086 40238 49138
rect 40290 49086 40302 49138
rect 29822 49074 29874 49086
rect 32174 49074 32226 49086
rect 42590 49074 42642 49086
rect 47182 49138 47234 49150
rect 51662 49138 51714 49150
rect 48738 49086 48750 49138
rect 48802 49086 48814 49138
rect 51090 49086 51102 49138
rect 51154 49086 51166 49138
rect 47182 49074 47234 49086
rect 51662 49074 51714 49086
rect 51998 49138 52050 49150
rect 56690 49086 56702 49138
rect 56754 49086 56766 49138
rect 57474 49086 57486 49138
rect 57538 49086 57550 49138
rect 51998 49074 52050 49086
rect 4734 49026 4786 49038
rect 4734 48962 4786 48974
rect 5966 49026 6018 49038
rect 5966 48962 6018 48974
rect 6190 49026 6242 49038
rect 6190 48962 6242 48974
rect 9774 49026 9826 49038
rect 9774 48962 9826 48974
rect 9998 49026 10050 49038
rect 9998 48962 10050 48974
rect 12014 49026 12066 49038
rect 18622 49026 18674 49038
rect 19518 49026 19570 49038
rect 12226 48974 12238 49026
rect 12290 48974 12302 49026
rect 12786 48974 12798 49026
rect 12850 48974 12862 49026
rect 14354 48974 14366 49026
rect 14418 48974 14430 49026
rect 19058 48974 19070 49026
rect 19122 48974 19134 49026
rect 12014 48962 12066 48974
rect 18622 48962 18674 48974
rect 19518 48962 19570 48974
rect 19630 49026 19682 49038
rect 19630 48962 19682 48974
rect 19742 49026 19794 49038
rect 19742 48962 19794 48974
rect 21310 49026 21362 49038
rect 21310 48962 21362 48974
rect 21534 49026 21586 49038
rect 21534 48962 21586 48974
rect 21870 49026 21922 49038
rect 21870 48962 21922 48974
rect 22094 49026 22146 49038
rect 25678 49026 25730 49038
rect 22978 48974 22990 49026
rect 23042 48974 23054 49026
rect 22094 48962 22146 48974
rect 25678 48962 25730 48974
rect 26238 49026 26290 49038
rect 27134 49026 27186 49038
rect 29934 49026 29986 49038
rect 31726 49026 31778 49038
rect 26898 48974 26910 49026
rect 26962 48974 26974 49026
rect 28242 48974 28254 49026
rect 28306 48974 28318 49026
rect 31378 48974 31390 49026
rect 31442 48974 31454 49026
rect 26238 48962 26290 48974
rect 27134 48962 27186 48974
rect 29934 48962 29986 48974
rect 31726 48962 31778 48974
rect 31950 49026 32002 49038
rect 31950 48962 32002 48974
rect 32286 49026 32338 49038
rect 36542 49026 36594 49038
rect 40014 49026 40066 49038
rect 42142 49026 42194 49038
rect 32722 48974 32734 49026
rect 32786 48974 32798 49026
rect 38994 48974 39006 49026
rect 39058 48974 39070 49026
rect 40338 48974 40350 49026
rect 40402 48974 40414 49026
rect 32286 48962 32338 48974
rect 36542 48962 36594 48974
rect 40014 48962 40066 48974
rect 42142 48962 42194 48974
rect 42478 49026 42530 49038
rect 42478 48962 42530 48974
rect 43822 49026 43874 49038
rect 43822 48962 43874 48974
rect 43934 49026 43986 49038
rect 43934 48962 43986 48974
rect 44382 49026 44434 49038
rect 44382 48962 44434 48974
rect 44942 49026 44994 49038
rect 46286 49026 46338 49038
rect 48414 49026 48466 49038
rect 52110 49026 52162 49038
rect 53118 49026 53170 49038
rect 45602 48974 45614 49026
rect 45666 48974 45678 49026
rect 46610 48974 46622 49026
rect 46674 48974 46686 49026
rect 47954 48974 47966 49026
rect 48018 48974 48030 49026
rect 50530 48974 50542 49026
rect 50594 48974 50606 49026
rect 52658 48974 52670 49026
rect 52722 48974 52734 49026
rect 44942 48962 44994 48974
rect 46286 48962 46338 48974
rect 48414 48962 48466 48974
rect 52110 48962 52162 48974
rect 53118 48962 53170 48974
rect 53454 49026 53506 49038
rect 57038 49026 57090 49038
rect 53890 48974 53902 49026
rect 53954 48974 53966 49026
rect 53454 48962 53506 48974
rect 57038 48962 57090 48974
rect 2942 48914 2994 48926
rect 5630 48914 5682 48926
rect 3490 48862 3502 48914
rect 3554 48862 3566 48914
rect 4386 48862 4398 48914
rect 4450 48862 4462 48914
rect 2942 48850 2994 48862
rect 5630 48850 5682 48862
rect 10670 48914 10722 48926
rect 10670 48850 10722 48862
rect 10894 48914 10946 48926
rect 10894 48850 10946 48862
rect 11902 48914 11954 48926
rect 18510 48914 18562 48926
rect 15026 48862 15038 48914
rect 15090 48862 15102 48914
rect 11902 48850 11954 48862
rect 18510 48850 18562 48862
rect 22430 48914 22482 48926
rect 23998 48914 24050 48926
rect 22866 48862 22878 48914
rect 22930 48862 22942 48914
rect 22430 48850 22482 48862
rect 23998 48850 24050 48862
rect 28030 48914 28082 48926
rect 28030 48850 28082 48862
rect 29374 48914 29426 48926
rect 29374 48850 29426 48862
rect 30158 48914 30210 48926
rect 30158 48850 30210 48862
rect 30942 48914 30994 48926
rect 30942 48850 30994 48862
rect 36206 48914 36258 48926
rect 36206 48850 36258 48862
rect 36318 48914 36370 48926
rect 36318 48850 36370 48862
rect 41246 48914 41298 48926
rect 46174 48914 46226 48926
rect 45154 48862 45166 48914
rect 45218 48862 45230 48914
rect 41246 48850 41298 48862
rect 46174 48850 46226 48862
rect 53342 48914 53394 48926
rect 54562 48862 54574 48914
rect 54626 48862 54638 48914
rect 53342 48850 53394 48862
rect 2830 48802 2882 48814
rect 2830 48738 2882 48750
rect 3838 48802 3890 48814
rect 3838 48738 3890 48750
rect 10782 48802 10834 48814
rect 17502 48802 17554 48814
rect 20750 48802 20802 48814
rect 11442 48750 11454 48802
rect 11506 48750 11518 48802
rect 12562 48750 12574 48802
rect 12626 48750 12638 48802
rect 17826 48750 17838 48802
rect 17890 48750 17902 48802
rect 10782 48738 10834 48750
rect 17502 48738 17554 48750
rect 20750 48738 20802 48750
rect 21422 48802 21474 48814
rect 21422 48738 21474 48750
rect 22318 48802 22370 48814
rect 22318 48738 22370 48750
rect 27470 48802 27522 48814
rect 27470 48738 27522 48750
rect 27694 48802 27746 48814
rect 27694 48738 27746 48750
rect 28478 48802 28530 48814
rect 28478 48738 28530 48750
rect 29262 48802 29314 48814
rect 29262 48738 29314 48750
rect 29710 48802 29762 48814
rect 29710 48738 29762 48750
rect 30606 48802 30658 48814
rect 30606 48738 30658 48750
rect 30830 48802 30882 48814
rect 35870 48802 35922 48814
rect 32946 48750 32958 48802
rect 33010 48750 33022 48802
rect 30830 48738 30882 48750
rect 35870 48738 35922 48750
rect 44158 48802 44210 48814
rect 44158 48738 44210 48750
rect 45726 48802 45778 48814
rect 45726 48738 45778 48750
rect 46062 48802 46114 48814
rect 46062 48738 46114 48750
rect 47070 48802 47122 48814
rect 47070 48738 47122 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 6974 48466 7026 48478
rect 26238 48466 26290 48478
rect 32062 48466 32114 48478
rect 45166 48466 45218 48478
rect 11106 48414 11118 48466
rect 11170 48414 11182 48466
rect 20962 48414 20974 48466
rect 21026 48414 21038 48466
rect 26562 48414 26574 48466
rect 26626 48414 26638 48466
rect 39666 48414 39678 48466
rect 39730 48414 39742 48466
rect 44370 48414 44382 48466
rect 44434 48414 44446 48466
rect 6974 48402 7026 48414
rect 26238 48402 26290 48414
rect 32062 48402 32114 48414
rect 45166 48402 45218 48414
rect 45726 48466 45778 48478
rect 45726 48402 45778 48414
rect 46062 48466 46114 48478
rect 46062 48402 46114 48414
rect 46174 48466 46226 48478
rect 46174 48402 46226 48414
rect 48862 48466 48914 48478
rect 48862 48402 48914 48414
rect 49310 48466 49362 48478
rect 49310 48402 49362 48414
rect 49870 48466 49922 48478
rect 49870 48402 49922 48414
rect 50542 48466 50594 48478
rect 50542 48402 50594 48414
rect 7982 48354 8034 48366
rect 2482 48302 2494 48354
rect 2546 48302 2558 48354
rect 6626 48302 6638 48354
rect 6690 48302 6702 48354
rect 7982 48290 8034 48302
rect 8094 48354 8146 48366
rect 8094 48290 8146 48302
rect 8766 48354 8818 48366
rect 16046 48354 16098 48366
rect 13570 48302 13582 48354
rect 13634 48302 13646 48354
rect 8766 48290 8818 48302
rect 16046 48290 16098 48302
rect 20526 48354 20578 48366
rect 27022 48354 27074 48366
rect 31950 48354 32002 48366
rect 22530 48302 22542 48354
rect 22594 48302 22606 48354
rect 28242 48302 28254 48354
rect 28306 48302 28318 48354
rect 20526 48290 20578 48302
rect 27022 48290 27074 48302
rect 31950 48290 32002 48302
rect 39230 48354 39282 48366
rect 45054 48354 45106 48366
rect 40338 48302 40350 48354
rect 40402 48302 40414 48354
rect 42466 48302 42478 48354
rect 42530 48302 42542 48354
rect 39230 48290 39282 48302
rect 45054 48290 45106 48302
rect 49646 48354 49698 48366
rect 49646 48290 49698 48302
rect 54014 48354 54066 48366
rect 54014 48290 54066 48302
rect 5630 48242 5682 48254
rect 1810 48190 1822 48242
rect 1874 48190 1886 48242
rect 5630 48178 5682 48190
rect 5854 48242 5906 48254
rect 5854 48178 5906 48190
rect 8318 48242 8370 48254
rect 8318 48178 8370 48190
rect 9998 48242 10050 48254
rect 14814 48242 14866 48254
rect 14354 48190 14366 48242
rect 14418 48190 14430 48242
rect 9998 48178 10050 48190
rect 14814 48178 14866 48190
rect 16158 48242 16210 48254
rect 16158 48178 16210 48190
rect 16382 48242 16434 48254
rect 20862 48242 20914 48254
rect 39006 48242 39058 48254
rect 16594 48190 16606 48242
rect 16658 48190 16670 48242
rect 17938 48190 17950 48242
rect 18002 48190 18014 48242
rect 21074 48190 21086 48242
rect 21138 48190 21150 48242
rect 21858 48190 21870 48242
rect 21922 48190 21934 48242
rect 27346 48190 27358 48242
rect 27410 48190 27422 48242
rect 28130 48190 28142 48242
rect 28194 48190 28206 48242
rect 31042 48190 31054 48242
rect 31106 48190 31118 48242
rect 31602 48190 31614 48242
rect 31666 48190 31678 48242
rect 37986 48190 37998 48242
rect 38050 48190 38062 48242
rect 16382 48178 16434 48190
rect 20862 48178 20914 48190
rect 39006 48178 39058 48190
rect 39118 48242 39170 48254
rect 44158 48242 44210 48254
rect 44606 48242 44658 48254
rect 40114 48190 40126 48242
rect 40178 48190 40190 48242
rect 40898 48190 40910 48242
rect 40962 48190 40974 48242
rect 42130 48190 42142 48242
rect 42194 48190 42206 48242
rect 42690 48190 42702 48242
rect 42754 48190 42766 48242
rect 43810 48190 43822 48242
rect 43874 48190 43886 48242
rect 44370 48190 44382 48242
rect 44434 48190 44446 48242
rect 39118 48178 39170 48190
rect 44158 48178 44210 48190
rect 44606 48178 44658 48190
rect 45950 48242 46002 48254
rect 50990 48242 51042 48254
rect 52334 48242 52386 48254
rect 53566 48242 53618 48254
rect 46610 48190 46622 48242
rect 46674 48190 46686 48242
rect 47170 48190 47182 48242
rect 47234 48190 47246 48242
rect 51314 48190 51326 48242
rect 51378 48190 51390 48242
rect 52770 48190 52782 48242
rect 52834 48190 52846 48242
rect 45950 48178 46002 48190
rect 50990 48178 51042 48190
rect 52334 48178 52386 48190
rect 53566 48178 53618 48190
rect 53790 48242 53842 48254
rect 57026 48190 57038 48242
rect 57090 48190 57102 48242
rect 53790 48178 53842 48190
rect 8878 48130 8930 48142
rect 4610 48078 4622 48130
rect 4674 48078 4686 48130
rect 8878 48066 8930 48078
rect 9886 48130 9938 48142
rect 9886 48066 9938 48078
rect 10558 48130 10610 48142
rect 35646 48130 35698 48142
rect 45278 48130 45330 48142
rect 51886 48130 51938 48142
rect 11442 48078 11454 48130
rect 11506 48078 11518 48130
rect 19730 48078 19742 48130
rect 19794 48078 19806 48130
rect 24658 48078 24670 48130
rect 24722 48078 24734 48130
rect 27234 48078 27246 48130
rect 27298 48078 27310 48130
rect 29026 48078 29038 48130
rect 29090 48078 29102 48130
rect 36194 48078 36206 48130
rect 36258 48078 36270 48130
rect 48066 48078 48078 48130
rect 48130 48078 48142 48130
rect 10558 48066 10610 48078
rect 35646 48066 35698 48078
rect 45278 48066 45330 48078
rect 51886 48066 51938 48078
rect 53230 48130 53282 48142
rect 53230 48066 53282 48078
rect 53678 48130 53730 48142
rect 53678 48066 53730 48078
rect 54574 48130 54626 48142
rect 54574 48066 54626 48078
rect 56590 48130 56642 48142
rect 56590 48066 56642 48078
rect 8990 48018 9042 48030
rect 6178 47966 6190 48018
rect 6242 47966 6254 48018
rect 8990 47954 9042 47966
rect 9550 48018 9602 48030
rect 9550 47954 9602 47966
rect 9662 48018 9714 48030
rect 9662 47954 9714 47966
rect 10782 48018 10834 48030
rect 32062 48018 32114 48030
rect 21074 47966 21086 48018
rect 21138 47966 21150 48018
rect 10782 47954 10834 47966
rect 32062 47954 32114 47966
rect 49982 48018 50034 48030
rect 49982 47954 50034 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 5070 47682 5122 47694
rect 5070 47618 5122 47630
rect 10894 47682 10946 47694
rect 20526 47682 20578 47694
rect 20178 47630 20190 47682
rect 20242 47630 20254 47682
rect 10894 47618 10946 47630
rect 20526 47618 20578 47630
rect 21646 47682 21698 47694
rect 21646 47618 21698 47630
rect 22206 47682 22258 47694
rect 22206 47618 22258 47630
rect 22542 47682 22594 47694
rect 22542 47618 22594 47630
rect 28254 47682 28306 47694
rect 31278 47682 31330 47694
rect 28578 47630 28590 47682
rect 28642 47630 28654 47682
rect 28254 47618 28306 47630
rect 31278 47618 31330 47630
rect 49534 47682 49586 47694
rect 49534 47618 49586 47630
rect 50206 47682 50258 47694
rect 50206 47618 50258 47630
rect 50318 47682 50370 47694
rect 50318 47618 50370 47630
rect 50542 47682 50594 47694
rect 50542 47618 50594 47630
rect 50654 47682 50706 47694
rect 50654 47618 50706 47630
rect 51102 47682 51154 47694
rect 51102 47618 51154 47630
rect 51438 47682 51490 47694
rect 51438 47618 51490 47630
rect 51774 47682 51826 47694
rect 51774 47618 51826 47630
rect 5742 47570 5794 47582
rect 9886 47570 9938 47582
rect 7746 47518 7758 47570
rect 7810 47518 7822 47570
rect 5742 47506 5794 47518
rect 9886 47506 9938 47518
rect 11230 47570 11282 47582
rect 11230 47506 11282 47518
rect 11790 47570 11842 47582
rect 19854 47570 19906 47582
rect 31166 47570 31218 47582
rect 42142 47570 42194 47582
rect 43374 47570 43426 47582
rect 17266 47518 17278 47570
rect 17330 47518 17342 47570
rect 19394 47518 19406 47570
rect 19458 47518 19470 47570
rect 30818 47518 30830 47570
rect 30882 47518 30894 47570
rect 36306 47518 36318 47570
rect 36370 47518 36382 47570
rect 38546 47518 38558 47570
rect 38610 47518 38622 47570
rect 39554 47518 39566 47570
rect 39618 47518 39630 47570
rect 43026 47518 43038 47570
rect 43090 47518 43102 47570
rect 11790 47506 11842 47518
rect 19854 47506 19906 47518
rect 31166 47506 31218 47518
rect 42142 47506 42194 47518
rect 43374 47506 43426 47518
rect 43822 47570 43874 47582
rect 43822 47506 43874 47518
rect 44158 47570 44210 47582
rect 44158 47506 44210 47518
rect 45502 47570 45554 47582
rect 47954 47518 47966 47570
rect 48018 47518 48030 47570
rect 51986 47518 51998 47570
rect 52050 47518 52062 47570
rect 57586 47518 57598 47570
rect 57650 47518 57662 47570
rect 45502 47506 45554 47518
rect 4958 47458 5010 47470
rect 4958 47394 5010 47406
rect 5966 47458 6018 47470
rect 5966 47394 6018 47406
rect 6078 47458 6130 47470
rect 11006 47458 11058 47470
rect 6962 47406 6974 47458
rect 7026 47406 7038 47458
rect 6078 47394 6130 47406
rect 11006 47394 11058 47406
rect 12014 47458 12066 47470
rect 12574 47458 12626 47470
rect 20750 47458 20802 47470
rect 12226 47406 12238 47458
rect 12290 47406 12302 47458
rect 15922 47406 15934 47458
rect 15986 47406 15998 47458
rect 16594 47406 16606 47458
rect 16658 47406 16670 47458
rect 12014 47394 12066 47406
rect 12574 47394 12626 47406
rect 20750 47394 20802 47406
rect 21422 47458 21474 47470
rect 21422 47394 21474 47406
rect 21758 47458 21810 47470
rect 21758 47394 21810 47406
rect 28030 47458 28082 47470
rect 44270 47458 44322 47470
rect 46174 47458 46226 47470
rect 29250 47406 29262 47458
rect 29314 47406 29326 47458
rect 29810 47406 29822 47458
rect 29874 47406 29886 47458
rect 33506 47406 33518 47458
rect 33570 47406 33582 47458
rect 37090 47406 37102 47458
rect 37154 47406 37166 47458
rect 37426 47406 37438 47458
rect 37490 47406 37502 47458
rect 38882 47406 38894 47458
rect 38946 47406 38958 47458
rect 40002 47406 40014 47458
rect 40066 47406 40078 47458
rect 41010 47406 41022 47458
rect 41074 47406 41086 47458
rect 42914 47406 42926 47458
rect 42978 47406 42990 47458
rect 45826 47406 45838 47458
rect 45890 47406 45902 47458
rect 28030 47394 28082 47406
rect 44270 47394 44322 47406
rect 46174 47394 46226 47406
rect 46286 47458 46338 47470
rect 48750 47458 48802 47470
rect 47058 47406 47070 47458
rect 47122 47406 47134 47458
rect 48066 47406 48078 47458
rect 48130 47406 48142 47458
rect 46286 47394 46338 47406
rect 48750 47394 48802 47406
rect 48974 47458 49026 47470
rect 49758 47458 49810 47470
rect 52670 47458 52722 47470
rect 49298 47406 49310 47458
rect 49362 47406 49374 47458
rect 52098 47406 52110 47458
rect 52162 47406 52174 47458
rect 48974 47394 49026 47406
rect 49758 47394 49810 47406
rect 52670 47394 52722 47406
rect 53006 47458 53058 47470
rect 53006 47394 53058 47406
rect 53230 47458 53282 47470
rect 54786 47406 54798 47458
rect 54850 47406 54862 47458
rect 53230 47394 53282 47406
rect 4846 47346 4898 47358
rect 4846 47282 4898 47294
rect 5630 47346 5682 47358
rect 5630 47282 5682 47294
rect 11342 47346 11394 47358
rect 11342 47282 11394 47294
rect 11678 47346 11730 47358
rect 22318 47346 22370 47358
rect 53790 47346 53842 47358
rect 16146 47294 16158 47346
rect 16210 47294 16222 47346
rect 34178 47294 34190 47346
rect 34242 47294 34254 47346
rect 40338 47294 40350 47346
rect 40402 47294 40414 47346
rect 41234 47294 41246 47346
rect 41298 47294 41310 47346
rect 41794 47294 41806 47346
rect 41858 47294 41870 47346
rect 47730 47294 47742 47346
rect 47794 47294 47806 47346
rect 55458 47294 55470 47346
rect 55522 47294 55534 47346
rect 11678 47282 11730 47294
rect 22318 47282 22370 47294
rect 53790 47282 53842 47294
rect 12686 47234 12738 47246
rect 12686 47170 12738 47182
rect 12798 47234 12850 47246
rect 12798 47170 12850 47182
rect 21758 47234 21810 47246
rect 21758 47170 21810 47182
rect 22990 47234 23042 47246
rect 22990 47170 23042 47182
rect 44942 47234 44994 47246
rect 44942 47170 44994 47182
rect 46398 47234 46450 47246
rect 46398 47170 46450 47182
rect 48526 47234 48578 47246
rect 48526 47170 48578 47182
rect 48862 47234 48914 47246
rect 48862 47170 48914 47182
rect 49422 47234 49474 47246
rect 49422 47170 49474 47182
rect 51326 47234 51378 47246
rect 51326 47170 51378 47182
rect 52894 47234 52946 47246
rect 52894 47170 52946 47182
rect 53454 47234 53506 47246
rect 53454 47170 53506 47182
rect 53678 47234 53730 47246
rect 53678 47170 53730 47182
rect 54238 47234 54290 47246
rect 54238 47170 54290 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 15262 46898 15314 46910
rect 8978 46846 8990 46898
rect 9042 46846 9054 46898
rect 15262 46834 15314 46846
rect 20302 46898 20354 46910
rect 37102 46898 37154 46910
rect 20626 46846 20638 46898
rect 20690 46846 20702 46898
rect 20302 46834 20354 46846
rect 37102 46834 37154 46846
rect 37550 46898 37602 46910
rect 37550 46834 37602 46846
rect 39678 46898 39730 46910
rect 39678 46834 39730 46846
rect 39790 46898 39842 46910
rect 42478 46898 42530 46910
rect 41906 46846 41918 46898
rect 41970 46846 41982 46898
rect 39790 46834 39842 46846
rect 42478 46834 42530 46846
rect 44382 46898 44434 46910
rect 44382 46834 44434 46846
rect 45054 46898 45106 46910
rect 45054 46834 45106 46846
rect 45278 46898 45330 46910
rect 45278 46834 45330 46846
rect 52110 46898 52162 46910
rect 52110 46834 52162 46846
rect 7310 46786 7362 46798
rect 38334 46786 38386 46798
rect 2930 46734 2942 46786
rect 2994 46734 3006 46786
rect 6850 46734 6862 46786
rect 6914 46734 6926 46786
rect 14018 46734 14030 46786
rect 14082 46734 14094 46786
rect 23650 46734 23662 46786
rect 23714 46734 23726 46786
rect 31714 46734 31726 46786
rect 31778 46734 31790 46786
rect 36754 46734 36766 46786
rect 36818 46734 36830 46786
rect 7310 46722 7362 46734
rect 38334 46722 38386 46734
rect 38670 46786 38722 46798
rect 38670 46722 38722 46734
rect 39006 46786 39058 46798
rect 39006 46722 39058 46734
rect 39230 46786 39282 46798
rect 51662 46786 51714 46798
rect 41234 46734 41246 46786
rect 41298 46734 41310 46786
rect 39230 46722 39282 46734
rect 51662 46722 51714 46734
rect 5518 46674 5570 46686
rect 6302 46674 6354 46686
rect 8430 46674 8482 46686
rect 2258 46622 2270 46674
rect 2322 46622 2334 46674
rect 5954 46622 5966 46674
rect 6018 46622 6030 46674
rect 7634 46622 7646 46674
rect 7698 46622 7710 46674
rect 5518 46610 5570 46622
rect 6302 46610 6354 46622
rect 8430 46610 8482 46622
rect 8654 46674 8706 46686
rect 10558 46674 10610 46686
rect 31390 46674 31442 46686
rect 35870 46674 35922 46686
rect 10210 46622 10222 46674
rect 10274 46622 10286 46674
rect 14802 46622 14814 46674
rect 14866 46622 14878 46674
rect 17938 46622 17950 46674
rect 18002 46622 18014 46674
rect 24322 46622 24334 46674
rect 24386 46622 24398 46674
rect 28130 46622 28142 46674
rect 28194 46622 28206 46674
rect 32050 46622 32062 46674
rect 32114 46622 32126 46674
rect 8654 46610 8706 46622
rect 10558 46610 10610 46622
rect 31390 46610 31442 46622
rect 35870 46610 35922 46622
rect 36318 46674 36370 46686
rect 37998 46674 38050 46686
rect 37538 46622 37550 46674
rect 37602 46622 37614 46674
rect 36318 46610 36370 46622
rect 37998 46610 38050 46622
rect 39566 46674 39618 46686
rect 39566 46610 39618 46622
rect 40238 46674 40290 46686
rect 42702 46674 42754 46686
rect 40898 46622 40910 46674
rect 40962 46622 40974 46674
rect 41794 46622 41806 46674
rect 41858 46622 41870 46674
rect 40238 46610 40290 46622
rect 42702 46610 42754 46622
rect 42926 46674 42978 46686
rect 42926 46610 42978 46622
rect 43262 46674 43314 46686
rect 43262 46610 43314 46622
rect 44606 46674 44658 46686
rect 50206 46674 50258 46686
rect 51886 46674 51938 46686
rect 45602 46622 45614 46674
rect 45666 46622 45678 46674
rect 49634 46622 49646 46674
rect 49698 46622 49710 46674
rect 51090 46622 51102 46674
rect 51154 46622 51166 46674
rect 44606 46610 44658 46622
rect 50206 46610 50258 46622
rect 51886 46610 51938 46622
rect 52222 46674 52274 46686
rect 52222 46610 52274 46622
rect 52558 46674 52610 46686
rect 52558 46610 52610 46622
rect 52894 46674 52946 46686
rect 52894 46610 52946 46622
rect 53230 46674 53282 46686
rect 53230 46610 53282 46622
rect 53454 46674 53506 46686
rect 53454 46610 53506 46622
rect 53678 46674 53730 46686
rect 53678 46610 53730 46622
rect 54126 46674 54178 46686
rect 54126 46610 54178 46622
rect 55358 46674 55410 46686
rect 55358 46610 55410 46622
rect 57710 46674 57762 46686
rect 57710 46610 57762 46622
rect 8094 46562 8146 46574
rect 11902 46562 11954 46574
rect 21310 46562 21362 46574
rect 28590 46562 28642 46574
rect 5058 46510 5070 46562
rect 5122 46510 5134 46562
rect 9762 46510 9774 46562
rect 9826 46510 9838 46562
rect 19618 46510 19630 46562
rect 19682 46510 19694 46562
rect 21522 46510 21534 46562
rect 21586 46510 21598 46562
rect 25218 46510 25230 46562
rect 25282 46510 25294 46562
rect 27346 46510 27358 46562
rect 27410 46510 27422 46562
rect 8094 46498 8146 46510
rect 11902 46498 11954 46510
rect 21310 46498 21362 46510
rect 28590 46498 28642 46510
rect 31054 46562 31106 46574
rect 31054 46498 31106 46510
rect 32286 46562 32338 46574
rect 32286 46498 32338 46510
rect 35534 46562 35586 46574
rect 35534 46498 35586 46510
rect 37886 46562 37938 46574
rect 37886 46498 37938 46510
rect 38782 46562 38834 46574
rect 38782 46498 38834 46510
rect 42814 46562 42866 46574
rect 45166 46562 45218 46574
rect 50766 46562 50818 46574
rect 43698 46510 43710 46562
rect 43762 46510 43774 46562
rect 47954 46510 47966 46562
rect 48018 46510 48030 46562
rect 49858 46510 49870 46562
rect 49922 46510 49934 46562
rect 42814 46498 42866 46510
rect 45166 46498 45218 46510
rect 50766 46498 50818 46510
rect 53006 46562 53058 46574
rect 53006 46498 53058 46510
rect 53902 46562 53954 46574
rect 53902 46498 53954 46510
rect 54462 46562 54514 46574
rect 54462 46498 54514 46510
rect 54910 46562 54962 46574
rect 54910 46498 54962 46510
rect 57150 46562 57202 46574
rect 57150 46498 57202 46510
rect 5406 46450 5458 46462
rect 5406 46386 5458 46398
rect 5742 46450 5794 46462
rect 5742 46386 5794 46398
rect 6526 46450 6578 46462
rect 6526 46386 6578 46398
rect 7646 46450 7698 46462
rect 32398 46450 32450 46462
rect 10322 46398 10334 46450
rect 10386 46398 10398 46450
rect 7646 46386 7698 46398
rect 32398 46386 32450 46398
rect 35982 46450 36034 46462
rect 35982 46386 36034 46398
rect 36430 46450 36482 46462
rect 54350 46450 54402 46462
rect 50642 46398 50654 46450
rect 50706 46398 50718 46450
rect 36430 46386 36482 46398
rect 54350 46386 54402 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 5070 46114 5122 46126
rect 5070 46050 5122 46062
rect 17278 46114 17330 46126
rect 17278 46050 17330 46062
rect 25790 46114 25842 46126
rect 25790 46050 25842 46062
rect 38446 46114 38498 46126
rect 38446 46050 38498 46062
rect 39566 46114 39618 46126
rect 39566 46050 39618 46062
rect 4958 46002 5010 46014
rect 17614 46002 17666 46014
rect 6962 45950 6974 46002
rect 7026 45950 7038 46002
rect 10098 45950 10110 46002
rect 10162 45950 10174 46002
rect 16930 45950 16942 46002
rect 16994 45950 17006 46002
rect 4958 45938 5010 45950
rect 17614 45938 17666 45950
rect 17838 46002 17890 46014
rect 17838 45938 17890 45950
rect 18622 46002 18674 46014
rect 18622 45938 18674 45950
rect 20414 46002 20466 46014
rect 35198 46002 35250 46014
rect 32610 45950 32622 46002
rect 32674 45950 32686 46002
rect 34738 45950 34750 46002
rect 34802 45950 34814 46002
rect 20414 45938 20466 45950
rect 35198 45938 35250 45950
rect 36542 46002 36594 46014
rect 36542 45938 36594 45950
rect 37214 46002 37266 46014
rect 37214 45938 37266 45950
rect 40014 46002 40066 46014
rect 40014 45938 40066 45950
rect 43934 46002 43986 46014
rect 50206 46002 50258 46014
rect 48626 45950 48638 46002
rect 48690 45950 48702 46002
rect 52658 45950 52670 46002
rect 52722 45950 52734 46002
rect 57810 45950 57822 46002
rect 57874 45950 57886 46002
rect 43934 45938 43986 45950
rect 50206 45938 50258 45950
rect 12238 45890 12290 45902
rect 18958 45890 19010 45902
rect 29822 45890 29874 45902
rect 37326 45890 37378 45902
rect 8754 45838 8766 45890
rect 8818 45838 8830 45890
rect 9762 45838 9774 45890
rect 9826 45838 9838 45890
rect 14130 45838 14142 45890
rect 14194 45838 14206 45890
rect 19506 45838 19518 45890
rect 19570 45838 19582 45890
rect 25778 45838 25790 45890
rect 25842 45838 25854 45890
rect 31938 45838 31950 45890
rect 32002 45838 32014 45890
rect 12238 45826 12290 45838
rect 18958 45826 19010 45838
rect 29822 45826 29874 45838
rect 37326 45826 37378 45838
rect 37550 45890 37602 45902
rect 37550 45826 37602 45838
rect 37774 45890 37826 45902
rect 37774 45826 37826 45838
rect 38670 45890 38722 45902
rect 38670 45826 38722 45838
rect 39230 45890 39282 45902
rect 39230 45826 39282 45838
rect 41806 45890 41858 45902
rect 41806 45826 41858 45838
rect 42142 45890 42194 45902
rect 42142 45826 42194 45838
rect 42478 45890 42530 45902
rect 45614 45890 45666 45902
rect 43026 45838 43038 45890
rect 43090 45838 43102 45890
rect 42478 45826 42530 45838
rect 45614 45826 45666 45838
rect 45726 45890 45778 45902
rect 50094 45890 50146 45902
rect 50878 45890 50930 45902
rect 51326 45890 51378 45902
rect 53902 45890 53954 45902
rect 46274 45838 46286 45890
rect 46338 45838 46350 45890
rect 49522 45838 49534 45890
rect 49586 45838 49598 45890
rect 50754 45838 50766 45890
rect 50818 45838 50830 45890
rect 51090 45838 51102 45890
rect 51154 45838 51166 45890
rect 53442 45838 53454 45890
rect 53506 45838 53518 45890
rect 45726 45826 45778 45838
rect 50094 45826 50146 45838
rect 50878 45826 50930 45838
rect 51326 45826 51378 45838
rect 53902 45826 53954 45838
rect 54126 45890 54178 45902
rect 54126 45826 54178 45838
rect 54350 45890 54402 45902
rect 54898 45838 54910 45890
rect 54962 45838 54974 45890
rect 54350 45826 54402 45838
rect 4846 45778 4898 45790
rect 25454 45778 25506 45790
rect 9650 45726 9662 45778
rect 9714 45726 9726 45778
rect 10658 45726 10670 45778
rect 10722 45726 10734 45778
rect 14802 45726 14814 45778
rect 14866 45726 14878 45778
rect 4846 45714 4898 45726
rect 25454 45714 25506 45726
rect 30158 45778 30210 45790
rect 39006 45778 39058 45790
rect 45838 45778 45890 45790
rect 38098 45726 38110 45778
rect 38162 45726 38174 45778
rect 41570 45726 41582 45778
rect 41634 45726 41646 45778
rect 30158 45714 30210 45726
rect 39006 45714 39058 45726
rect 45838 45714 45890 45726
rect 53006 45778 53058 45790
rect 53666 45726 53678 45778
rect 53730 45726 53742 45778
rect 55682 45726 55694 45778
rect 55746 45726 55758 45778
rect 53006 45714 53058 45726
rect 19070 45666 19122 45678
rect 19070 45602 19122 45614
rect 19182 45666 19234 45678
rect 19182 45602 19234 45614
rect 20078 45666 20130 45678
rect 20078 45602 20130 45614
rect 21422 45666 21474 45678
rect 21422 45602 21474 45614
rect 21870 45666 21922 45678
rect 21870 45602 21922 45614
rect 25118 45666 25170 45678
rect 25118 45602 25170 45614
rect 26238 45666 26290 45678
rect 26238 45602 26290 45614
rect 26686 45666 26738 45678
rect 26686 45602 26738 45614
rect 37102 45666 37154 45678
rect 37102 45602 37154 45614
rect 40462 45666 40514 45678
rect 40462 45602 40514 45614
rect 41246 45666 41298 45678
rect 41246 45602 41298 45614
rect 42142 45666 42194 45678
rect 44270 45666 44322 45678
rect 50542 45666 50594 45678
rect 42802 45614 42814 45666
rect 42866 45614 42878 45666
rect 45154 45614 45166 45666
rect 45218 45614 45230 45666
rect 42142 45602 42194 45614
rect 44270 45602 44322 45614
rect 50542 45602 50594 45614
rect 51774 45666 51826 45678
rect 51774 45602 51826 45614
rect 52782 45666 52834 45678
rect 52782 45602 52834 45614
rect 54462 45666 54514 45678
rect 54462 45602 54514 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 8878 45330 8930 45342
rect 8878 45266 8930 45278
rect 9662 45330 9714 45342
rect 25902 45330 25954 45342
rect 11106 45278 11118 45330
rect 11170 45278 11182 45330
rect 9662 45266 9714 45278
rect 25902 45266 25954 45278
rect 33182 45330 33234 45342
rect 33182 45266 33234 45278
rect 34638 45330 34690 45342
rect 34638 45266 34690 45278
rect 37886 45330 37938 45342
rect 37886 45266 37938 45278
rect 37998 45330 38050 45342
rect 37998 45266 38050 45278
rect 38782 45330 38834 45342
rect 42142 45330 42194 45342
rect 41234 45278 41246 45330
rect 41298 45278 41310 45330
rect 38782 45266 38834 45278
rect 42142 45266 42194 45278
rect 42366 45330 42418 45342
rect 42366 45266 42418 45278
rect 43150 45330 43202 45342
rect 43150 45266 43202 45278
rect 43486 45330 43538 45342
rect 43486 45266 43538 45278
rect 44270 45330 44322 45342
rect 44270 45266 44322 45278
rect 45950 45330 46002 45342
rect 45950 45266 46002 45278
rect 48862 45330 48914 45342
rect 48862 45266 48914 45278
rect 49758 45330 49810 45342
rect 49758 45266 49810 45278
rect 10222 45218 10274 45230
rect 34862 45218 34914 45230
rect 5058 45166 5070 45218
rect 5122 45166 5134 45218
rect 13346 45166 13358 45218
rect 13410 45166 13422 45218
rect 18722 45166 18734 45218
rect 18786 45166 18798 45218
rect 10222 45154 10274 45166
rect 34862 45154 34914 45166
rect 38670 45218 38722 45230
rect 38670 45154 38722 45166
rect 49982 45218 50034 45230
rect 55582 45218 55634 45230
rect 50754 45166 50766 45218
rect 50818 45166 50830 45218
rect 49982 45154 50034 45166
rect 55582 45154 55634 45166
rect 56590 45218 56642 45230
rect 56590 45154 56642 45166
rect 14590 45106 14642 45118
rect 34414 45106 34466 45118
rect 4386 45054 4398 45106
rect 4450 45054 4462 45106
rect 8082 45054 8094 45106
rect 8146 45054 8158 45106
rect 8418 45054 8430 45106
rect 8482 45054 8494 45106
rect 14130 45054 14142 45106
rect 14194 45054 14206 45106
rect 18050 45054 18062 45106
rect 18114 45054 18126 45106
rect 21186 45054 21198 45106
rect 21250 45054 21262 45106
rect 26338 45054 26350 45106
rect 26402 45054 26414 45106
rect 29586 45054 29598 45106
rect 29650 45054 29662 45106
rect 14590 45042 14642 45054
rect 34414 45042 34466 45054
rect 34526 45106 34578 45118
rect 34526 45042 34578 45054
rect 35310 45106 35362 45118
rect 35310 45042 35362 45054
rect 37774 45106 37826 45118
rect 37774 45042 37826 45054
rect 38446 45106 38498 45118
rect 42254 45106 42306 45118
rect 38994 45054 39006 45106
rect 39058 45054 39070 45106
rect 41010 45054 41022 45106
rect 41074 45054 41086 45106
rect 38446 45042 38498 45054
rect 42254 45042 42306 45054
rect 42814 45106 42866 45118
rect 42814 45042 42866 45054
rect 43038 45106 43090 45118
rect 43038 45042 43090 45054
rect 43262 45106 43314 45118
rect 43262 45042 43314 45054
rect 44158 45106 44210 45118
rect 44158 45042 44210 45054
rect 44494 45106 44546 45118
rect 44942 45106 44994 45118
rect 44706 45054 44718 45106
rect 44770 45054 44782 45106
rect 44494 45042 44546 45054
rect 44942 45042 44994 45054
rect 45166 45106 45218 45118
rect 53566 45106 53618 45118
rect 45378 45054 45390 45106
rect 45442 45054 45454 45106
rect 51090 45054 51102 45106
rect 51154 45054 51166 45106
rect 52658 45054 52670 45106
rect 52722 45054 52734 45106
rect 45166 45042 45218 45054
rect 53566 45042 53618 45054
rect 53790 45106 53842 45118
rect 53790 45042 53842 45054
rect 54126 45106 54178 45118
rect 54126 45042 54178 45054
rect 55358 45106 55410 45118
rect 57138 45054 57150 45106
rect 57202 45054 57214 45106
rect 55358 45042 55410 45054
rect 17502 44994 17554 45006
rect 25342 44994 25394 45006
rect 36878 44994 36930 45006
rect 7186 44942 7198 44994
rect 7250 44942 7262 44994
rect 8530 44942 8542 44994
rect 8594 44942 8606 44994
rect 20850 44942 20862 44994
rect 20914 44942 20926 44994
rect 21970 44942 21982 44994
rect 22034 44942 22046 44994
rect 24098 44942 24110 44994
rect 24162 44942 24174 44994
rect 27122 44942 27134 44994
rect 27186 44942 27198 44994
rect 29250 44942 29262 44994
rect 29314 44942 29326 44994
rect 30370 44942 30382 44994
rect 30434 44942 30446 44994
rect 32498 44942 32510 44994
rect 32562 44942 32574 44994
rect 17502 44930 17554 44942
rect 25342 44930 25394 44942
rect 36878 44930 36930 44942
rect 39454 44994 39506 45006
rect 46398 44994 46450 45006
rect 54686 44994 54738 45006
rect 45266 44942 45278 44994
rect 45330 44942 45342 44994
rect 48738 44942 48750 44994
rect 48802 44942 48814 44994
rect 49634 44942 49646 44994
rect 49698 44942 49710 44994
rect 51202 44942 51214 44994
rect 51266 44942 51278 44994
rect 39454 44930 39506 44942
rect 46398 44930 46450 44942
rect 54686 44930 54738 44942
rect 55022 44994 55074 45006
rect 57362 44942 57374 44994
rect 57426 44942 57438 44994
rect 55022 44930 55074 44942
rect 25678 44882 25730 44894
rect 25678 44818 25730 44830
rect 26014 44882 26066 44894
rect 26014 44818 26066 44830
rect 35422 44882 35474 44894
rect 35422 44818 35474 44830
rect 49086 44882 49138 44894
rect 49086 44818 49138 44830
rect 52894 44882 52946 44894
rect 52894 44818 52946 44830
rect 53342 44882 53394 44894
rect 53342 44818 53394 44830
rect 54350 44882 54402 44894
rect 54350 44818 54402 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 11790 44546 11842 44558
rect 55582 44546 55634 44558
rect 53330 44494 53342 44546
rect 53394 44494 53406 44546
rect 11790 44482 11842 44494
rect 55582 44482 55634 44494
rect 12126 44434 12178 44446
rect 7410 44382 7422 44434
rect 7474 44382 7486 44434
rect 9538 44382 9550 44434
rect 9602 44382 9614 44434
rect 12126 44370 12178 44382
rect 12798 44434 12850 44446
rect 12798 44370 12850 44382
rect 14814 44434 14866 44446
rect 21422 44434 21474 44446
rect 19506 44382 19518 44434
rect 19570 44382 19582 44434
rect 14814 44370 14866 44382
rect 21422 44370 21474 44382
rect 22206 44434 22258 44446
rect 38222 44434 38274 44446
rect 25442 44382 25454 44434
rect 25506 44382 25518 44434
rect 27570 44382 27582 44434
rect 27634 44382 27646 44434
rect 31042 44382 31054 44434
rect 31106 44382 31118 44434
rect 32498 44382 32510 44434
rect 32562 44382 32574 44434
rect 22206 44370 22258 44382
rect 38222 44370 38274 44382
rect 43038 44434 43090 44446
rect 43038 44370 43090 44382
rect 43374 44434 43426 44446
rect 43374 44370 43426 44382
rect 57262 44434 57314 44446
rect 57262 44370 57314 44382
rect 8318 44322 8370 44334
rect 15150 44322 15202 44334
rect 20414 44322 20466 44334
rect 34862 44322 34914 44334
rect 37102 44322 37154 44334
rect 7298 44270 7310 44322
rect 7362 44270 7374 44322
rect 7858 44270 7870 44322
rect 7922 44270 7934 44322
rect 10322 44270 10334 44322
rect 10386 44270 10398 44322
rect 16034 44270 16046 44322
rect 16098 44270 16110 44322
rect 16706 44270 16718 44322
rect 16770 44270 16782 44322
rect 22418 44270 22430 44322
rect 22482 44270 22494 44322
rect 23314 44270 23326 44322
rect 23378 44270 23390 44322
rect 28354 44270 28366 44322
rect 28418 44270 28430 44322
rect 31378 44270 31390 44322
rect 31442 44270 31454 44322
rect 32162 44270 32174 44322
rect 32226 44270 32238 44322
rect 33282 44270 33294 44322
rect 33346 44270 33358 44322
rect 34290 44270 34302 44322
rect 34354 44270 34366 44322
rect 35186 44270 35198 44322
rect 35250 44270 35262 44322
rect 35970 44270 35982 44322
rect 36034 44270 36046 44322
rect 8318 44258 8370 44270
rect 15150 44258 15202 44270
rect 20414 44258 20466 44270
rect 34862 44258 34914 44270
rect 37102 44258 37154 44270
rect 37662 44322 37714 44334
rect 37662 44258 37714 44270
rect 37774 44322 37826 44334
rect 37774 44258 37826 44270
rect 38670 44322 38722 44334
rect 42478 44322 42530 44334
rect 50430 44322 50482 44334
rect 53902 44322 53954 44334
rect 55358 44322 55410 44334
rect 40786 44270 40798 44322
rect 40850 44270 40862 44322
rect 43922 44270 43934 44322
rect 43986 44270 43998 44322
rect 46050 44270 46062 44322
rect 46114 44270 46126 44322
rect 48066 44270 48078 44322
rect 48130 44270 48142 44322
rect 49298 44270 49310 44322
rect 49362 44270 49374 44322
rect 53106 44270 53118 44322
rect 53170 44270 53182 44322
rect 53666 44270 53678 44322
rect 53730 44270 53742 44322
rect 54786 44270 54798 44322
rect 54850 44270 54862 44322
rect 38670 44258 38722 44270
rect 42478 44258 42530 44270
rect 50430 44258 50482 44270
rect 53902 44258 53954 44270
rect 55358 44258 55410 44270
rect 56366 44322 56418 44334
rect 56366 44258 56418 44270
rect 56814 44322 56866 44334
rect 56814 44258 56866 44270
rect 57486 44322 57538 44334
rect 57486 44258 57538 44270
rect 57598 44322 57650 44334
rect 57598 44258 57650 44270
rect 12350 44210 12402 44222
rect 19854 44210 19906 44222
rect 7186 44158 7198 44210
rect 7250 44158 7262 44210
rect 9874 44158 9886 44210
rect 9938 44158 9950 44210
rect 10546 44158 10558 44210
rect 10610 44158 10622 44210
rect 16258 44158 16270 44210
rect 16322 44158 16334 44210
rect 17378 44158 17390 44210
rect 17442 44158 17454 44210
rect 12350 44146 12402 44158
rect 19854 44146 19906 44158
rect 20190 44210 20242 44222
rect 20190 44146 20242 44158
rect 22094 44210 22146 44222
rect 22094 44146 22146 44158
rect 22990 44210 23042 44222
rect 22990 44146 23042 44158
rect 32846 44210 32898 44222
rect 38110 44210 38162 44222
rect 34626 44158 34638 44210
rect 34690 44158 34702 44210
rect 35298 44158 35310 44210
rect 35362 44158 35374 44210
rect 32846 44146 32898 44158
rect 38110 44146 38162 44158
rect 38446 44210 38498 44222
rect 50318 44210 50370 44222
rect 43474 44158 43486 44210
rect 43538 44158 43550 44210
rect 43810 44158 43822 44210
rect 43874 44158 43886 44210
rect 45714 44158 45726 44210
rect 45778 44158 45790 44210
rect 48962 44158 48974 44210
rect 49026 44158 49038 44210
rect 38446 44146 38498 44158
rect 50318 44146 50370 44158
rect 50766 44210 50818 44222
rect 50766 44146 50818 44158
rect 50878 44210 50930 44222
rect 50878 44146 50930 44158
rect 51102 44210 51154 44222
rect 56254 44210 56306 44222
rect 55010 44158 55022 44210
rect 55074 44158 55086 44210
rect 51102 44146 51154 44158
rect 56254 44146 56306 44158
rect 56590 44210 56642 44222
rect 56590 44146 56642 44158
rect 57150 44210 57202 44222
rect 57150 44146 57202 44158
rect 15486 44098 15538 44110
rect 15486 44034 15538 44046
rect 20078 44098 20130 44110
rect 20078 44034 20130 44046
rect 23102 44098 23154 44110
rect 23102 44034 23154 44046
rect 29262 44098 29314 44110
rect 37550 44098 37602 44110
rect 33506 44046 33518 44098
rect 33570 44046 33582 44098
rect 29262 44034 29314 44046
rect 37550 44034 37602 44046
rect 39118 44098 39170 44110
rect 44382 44098 44434 44110
rect 50094 44098 50146 44110
rect 41010 44046 41022 44098
rect 41074 44046 41086 44098
rect 46162 44046 46174 44098
rect 46226 44046 46238 44098
rect 39118 44034 39170 44046
rect 44382 44034 44434 44046
rect 50094 44034 50146 44046
rect 51438 44098 51490 44110
rect 51438 44034 51490 44046
rect 52222 44098 52274 44110
rect 52222 44034 52274 44046
rect 52894 44098 52946 44110
rect 54350 44098 54402 44110
rect 53554 44046 53566 44098
rect 53618 44046 53630 44098
rect 55906 44046 55918 44098
rect 55970 44046 55982 44098
rect 52894 44034 52946 44046
rect 54350 44034 54402 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 37998 43762 38050 43774
rect 10098 43710 10110 43762
rect 10162 43710 10174 43762
rect 37998 43698 38050 43710
rect 40014 43762 40066 43774
rect 40014 43698 40066 43710
rect 45502 43762 45554 43774
rect 45502 43698 45554 43710
rect 48638 43762 48690 43774
rect 48638 43698 48690 43710
rect 18510 43650 18562 43662
rect 9762 43598 9774 43650
rect 9826 43598 9838 43650
rect 11442 43598 11454 43650
rect 11506 43598 11518 43650
rect 18050 43598 18062 43650
rect 18114 43598 18126 43650
rect 18510 43586 18562 43598
rect 18958 43650 19010 43662
rect 18958 43586 19010 43598
rect 21310 43650 21362 43662
rect 27918 43650 27970 43662
rect 28702 43650 28754 43662
rect 27234 43598 27246 43650
rect 27298 43598 27310 43650
rect 28242 43598 28254 43650
rect 28306 43598 28318 43650
rect 21310 43586 21362 43598
rect 27918 43586 27970 43598
rect 28702 43586 28754 43598
rect 30158 43650 30210 43662
rect 30158 43586 30210 43598
rect 30494 43650 30546 43662
rect 35646 43650 35698 43662
rect 33954 43598 33966 43650
rect 34018 43598 34030 43650
rect 30494 43586 30546 43598
rect 35646 43586 35698 43598
rect 36654 43650 36706 43662
rect 36654 43586 36706 43598
rect 39790 43650 39842 43662
rect 39790 43586 39842 43598
rect 43038 43650 43090 43662
rect 52782 43650 52834 43662
rect 52434 43598 52446 43650
rect 52498 43598 52510 43650
rect 43038 43586 43090 43598
rect 52782 43586 52834 43598
rect 53006 43650 53058 43662
rect 53006 43586 53058 43598
rect 53790 43650 53842 43662
rect 53790 43586 53842 43598
rect 56030 43650 56082 43662
rect 56030 43586 56082 43598
rect 57038 43650 57090 43662
rect 57038 43586 57090 43598
rect 20862 43538 20914 43550
rect 6962 43486 6974 43538
rect 7026 43486 7038 43538
rect 9538 43486 9550 43538
rect 9602 43486 9614 43538
rect 10546 43486 10558 43538
rect 10610 43486 10622 43538
rect 10994 43486 11006 43538
rect 11058 43486 11070 43538
rect 11666 43486 11678 43538
rect 11730 43486 11742 43538
rect 12226 43486 12238 43538
rect 12290 43486 12302 43538
rect 17826 43486 17838 43538
rect 17890 43486 17902 43538
rect 20862 43474 20914 43486
rect 21198 43538 21250 43550
rect 21198 43474 21250 43486
rect 21422 43538 21474 43550
rect 27582 43538 27634 43550
rect 24546 43486 24558 43538
rect 24610 43486 24622 43538
rect 21422 43474 21474 43486
rect 27582 43474 27634 43486
rect 33630 43538 33682 43550
rect 33630 43474 33682 43486
rect 34414 43538 34466 43550
rect 35870 43538 35922 43550
rect 34850 43486 34862 43538
rect 34914 43486 34926 43538
rect 34414 43474 34466 43486
rect 35870 43474 35922 43486
rect 36094 43538 36146 43550
rect 36094 43474 36146 43486
rect 36206 43538 36258 43550
rect 36206 43474 36258 43486
rect 36542 43538 36594 43550
rect 36542 43474 36594 43486
rect 36878 43538 36930 43550
rect 36878 43474 36930 43486
rect 38782 43538 38834 43550
rect 38782 43474 38834 43486
rect 39230 43538 39282 43550
rect 39230 43474 39282 43486
rect 42478 43538 42530 43550
rect 42478 43474 42530 43486
rect 42814 43538 42866 43550
rect 47294 43538 47346 43550
rect 46162 43486 46174 43538
rect 46226 43486 46238 43538
rect 46498 43486 46510 43538
rect 46562 43486 46574 43538
rect 42814 43474 42866 43486
rect 47294 43474 47346 43486
rect 47630 43538 47682 43550
rect 47630 43474 47682 43486
rect 48190 43538 48242 43550
rect 50318 43538 50370 43550
rect 49410 43486 49422 43538
rect 49474 43486 49486 43538
rect 49634 43486 49646 43538
rect 49698 43486 49710 43538
rect 48190 43474 48242 43486
rect 50318 43474 50370 43486
rect 51774 43538 51826 43550
rect 51774 43474 51826 43486
rect 52110 43538 52162 43550
rect 52110 43474 52162 43486
rect 55470 43538 55522 43550
rect 55470 43474 55522 43486
rect 55806 43538 55858 43550
rect 55806 43474 55858 43486
rect 56590 43538 56642 43550
rect 56590 43474 56642 43486
rect 56814 43538 56866 43550
rect 56814 43474 56866 43486
rect 19742 43426 19794 43438
rect 33406 43426 33458 43438
rect 7522 43374 7534 43426
rect 7586 43374 7598 43426
rect 12898 43374 12910 43426
rect 12962 43374 12974 43426
rect 15026 43374 15038 43426
rect 15090 43374 15102 43426
rect 21746 43374 21758 43426
rect 21810 43374 21822 43426
rect 23874 43374 23886 43426
rect 23938 43374 23950 43426
rect 28578 43374 28590 43426
rect 28642 43374 28654 43426
rect 19742 43362 19794 43374
rect 33406 43362 33458 43374
rect 35310 43426 35362 43438
rect 39342 43426 39394 43438
rect 38994 43374 39006 43426
rect 39058 43374 39070 43426
rect 35310 43362 35362 43374
rect 39342 43362 39394 43374
rect 42926 43426 42978 43438
rect 55918 43426 55970 43438
rect 45826 43374 45838 43426
rect 45890 43374 45902 43426
rect 49522 43374 49534 43426
rect 49586 43374 49598 43426
rect 51314 43374 51326 43426
rect 51378 43374 51390 43426
rect 53106 43374 53118 43426
rect 53170 43374 53182 43426
rect 42926 43362 42978 43374
rect 55918 43362 55970 43374
rect 18846 43314 18898 43326
rect 18846 43250 18898 43262
rect 28926 43314 28978 43326
rect 28926 43250 28978 43262
rect 38558 43314 38610 43326
rect 38558 43250 38610 43262
rect 40126 43314 40178 43326
rect 40126 43250 40178 43262
rect 47406 43314 47458 43326
rect 47406 43250 47458 43262
rect 50542 43314 50594 43326
rect 53566 43314 53618 43326
rect 50866 43262 50878 43314
rect 50930 43262 50942 43314
rect 50542 43250 50594 43262
rect 53566 43250 53618 43262
rect 53902 43314 53954 43326
rect 57362 43262 57374 43314
rect 57426 43262 57438 43314
rect 53902 43250 53954 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 22654 42978 22706 42990
rect 22654 42914 22706 42926
rect 37550 42978 37602 42990
rect 43822 42978 43874 42990
rect 40450 42926 40462 42978
rect 40514 42926 40526 42978
rect 37550 42914 37602 42926
rect 43822 42914 43874 42926
rect 17054 42866 17106 42878
rect 9538 42814 9550 42866
rect 9602 42814 9614 42866
rect 17054 42802 17106 42814
rect 17838 42866 17890 42878
rect 22318 42866 22370 42878
rect 33742 42866 33794 42878
rect 36318 42866 36370 42878
rect 21746 42814 21758 42866
rect 21810 42814 21822 42866
rect 24322 42814 24334 42866
rect 24386 42814 24398 42866
rect 26450 42814 26462 42866
rect 26514 42814 26526 42866
rect 34626 42814 34638 42866
rect 34690 42814 34702 42866
rect 17838 42802 17890 42814
rect 22318 42802 22370 42814
rect 33742 42802 33794 42814
rect 36318 42802 36370 42814
rect 38670 42866 38722 42878
rect 38670 42802 38722 42814
rect 38782 42866 38834 42878
rect 42478 42866 42530 42878
rect 48974 42866 49026 42878
rect 40562 42814 40574 42866
rect 40626 42814 40638 42866
rect 45826 42814 45838 42866
rect 45890 42814 45902 42866
rect 38782 42802 38834 42814
rect 42478 42802 42530 42814
rect 48974 42802 49026 42814
rect 53118 42866 53170 42878
rect 55682 42814 55694 42866
rect 55746 42814 55758 42866
rect 57810 42814 57822 42866
rect 57874 42814 57886 42866
rect 53118 42802 53170 42814
rect 14926 42754 14978 42766
rect 6738 42702 6750 42754
rect 6802 42702 6814 42754
rect 14926 42690 14978 42702
rect 16270 42754 16322 42766
rect 16270 42690 16322 42702
rect 18062 42754 18114 42766
rect 18062 42690 18114 42702
rect 18286 42754 18338 42766
rect 31278 42754 31330 42766
rect 18834 42702 18846 42754
rect 18898 42702 18910 42754
rect 23538 42702 23550 42754
rect 23602 42702 23614 42754
rect 18286 42690 18338 42702
rect 31278 42690 31330 42702
rect 31950 42754 32002 42766
rect 31950 42690 32002 42702
rect 32510 42754 32562 42766
rect 36206 42754 36258 42766
rect 34290 42702 34302 42754
rect 34354 42702 34366 42754
rect 35858 42702 35870 42754
rect 35922 42702 35934 42754
rect 32510 42690 32562 42702
rect 36206 42690 36258 42702
rect 37662 42754 37714 42766
rect 42814 42754 42866 42766
rect 38098 42702 38110 42754
rect 38162 42702 38174 42754
rect 39218 42702 39230 42754
rect 39282 42702 39294 42754
rect 40114 42702 40126 42754
rect 40178 42702 40190 42754
rect 37662 42690 37714 42702
rect 42814 42690 42866 42702
rect 43150 42754 43202 42766
rect 43150 42690 43202 42702
rect 43598 42754 43650 42766
rect 43598 42690 43650 42702
rect 43934 42754 43986 42766
rect 43934 42690 43986 42702
rect 44270 42754 44322 42766
rect 51662 42754 51714 42766
rect 44930 42702 44942 42754
rect 44994 42702 45006 42754
rect 46274 42702 46286 42754
rect 46338 42702 46350 42754
rect 47170 42702 47182 42754
rect 47234 42702 47246 42754
rect 50978 42702 50990 42754
rect 51042 42702 51054 42754
rect 44270 42690 44322 42702
rect 51662 42690 51714 42702
rect 52558 42754 52610 42766
rect 52558 42690 52610 42702
rect 53006 42754 53058 42766
rect 54898 42702 54910 42754
rect 54962 42702 54974 42754
rect 53006 42690 53058 42702
rect 17390 42642 17442 42654
rect 21310 42642 21362 42654
rect 7410 42590 7422 42642
rect 7474 42590 7486 42642
rect 17602 42590 17614 42642
rect 17666 42590 17678 42642
rect 17390 42578 17442 42590
rect 21310 42578 21362 42590
rect 22542 42642 22594 42654
rect 22542 42578 22594 42590
rect 30606 42642 30658 42654
rect 30606 42578 30658 42590
rect 30830 42642 30882 42654
rect 42366 42642 42418 42654
rect 46734 42642 46786 42654
rect 53230 42642 53282 42654
rect 38434 42590 38446 42642
rect 38498 42590 38510 42642
rect 42914 42590 42926 42642
rect 42978 42590 42990 42642
rect 45154 42590 45166 42642
rect 45218 42590 45230 42642
rect 47282 42590 47294 42642
rect 47346 42590 47358 42642
rect 50866 42590 50878 42642
rect 50930 42590 50942 42642
rect 30830 42578 30882 42590
rect 42366 42578 42418 42590
rect 46734 42578 46786 42590
rect 53230 42578 53282 42590
rect 9998 42530 10050 42542
rect 9998 42466 10050 42478
rect 10782 42530 10834 42542
rect 10782 42466 10834 42478
rect 11790 42530 11842 42542
rect 11790 42466 11842 42478
rect 14590 42530 14642 42542
rect 14590 42466 14642 42478
rect 16382 42530 16434 42542
rect 18622 42530 18674 42542
rect 17714 42478 17726 42530
rect 17778 42478 17790 42530
rect 16382 42466 16434 42478
rect 18622 42466 18674 42478
rect 21534 42530 21586 42542
rect 21534 42466 21586 42478
rect 21758 42530 21810 42542
rect 21758 42466 21810 42478
rect 21870 42530 21922 42542
rect 21870 42466 21922 42478
rect 23214 42530 23266 42542
rect 23214 42466 23266 42478
rect 27806 42530 27858 42542
rect 27806 42466 27858 42478
rect 31054 42530 31106 42542
rect 31054 42466 31106 42478
rect 37550 42530 37602 42542
rect 37550 42466 37602 42478
rect 41470 42530 41522 42542
rect 41470 42466 41522 42478
rect 44158 42530 44210 42542
rect 44158 42466 44210 42478
rect 51438 42530 51490 42542
rect 51438 42466 51490 42478
rect 51774 42530 51826 42542
rect 51774 42466 51826 42478
rect 51886 42530 51938 42542
rect 51886 42466 51938 42478
rect 53678 42530 53730 42542
rect 53678 42466 53730 42478
rect 54126 42530 54178 42542
rect 54126 42466 54178 42478
rect 54574 42530 54626 42542
rect 54574 42466 54626 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 9886 42194 9938 42206
rect 9886 42130 9938 42142
rect 10670 42194 10722 42206
rect 10670 42130 10722 42142
rect 10894 42194 10946 42206
rect 10894 42130 10946 42142
rect 21422 42194 21474 42206
rect 21422 42130 21474 42142
rect 22094 42194 22146 42206
rect 22094 42130 22146 42142
rect 37998 42194 38050 42206
rect 37998 42130 38050 42142
rect 40126 42194 40178 42206
rect 40126 42130 40178 42142
rect 43710 42194 43762 42206
rect 47854 42194 47906 42206
rect 47282 42142 47294 42194
rect 47346 42142 47358 42194
rect 43710 42130 43762 42142
rect 47854 42130 47906 42142
rect 48750 42194 48802 42206
rect 48750 42130 48802 42142
rect 55806 42194 55858 42206
rect 55806 42130 55858 42142
rect 14478 42082 14530 42094
rect 15822 42082 15874 42094
rect 10210 42030 10222 42082
rect 10274 42030 10286 42082
rect 14802 42030 14814 42082
rect 14866 42030 14878 42082
rect 14478 42018 14530 42030
rect 15822 42018 15874 42030
rect 19630 42082 19682 42094
rect 37886 42082 37938 42094
rect 19954 42030 19966 42082
rect 20018 42030 20030 42082
rect 31266 42030 31278 42082
rect 31330 42030 31342 42082
rect 19630 42018 19682 42030
rect 37886 42018 37938 42030
rect 39454 42082 39506 42094
rect 39454 42018 39506 42030
rect 39566 42082 39618 42094
rect 39566 42018 39618 42030
rect 40238 42082 40290 42094
rect 49534 42082 49586 42094
rect 45826 42030 45838 42082
rect 45890 42030 45902 42082
rect 56690 42030 56702 42082
rect 56754 42030 56766 42082
rect 40238 42018 40290 42030
rect 49534 42018 49586 42030
rect 10558 41970 10610 41982
rect 14366 41970 14418 41982
rect 17726 41970 17778 41982
rect 6066 41918 6078 41970
rect 6130 41918 6142 41970
rect 11106 41918 11118 41970
rect 11170 41918 11182 41970
rect 15250 41918 15262 41970
rect 15314 41918 15326 41970
rect 16034 41918 16046 41970
rect 16098 41918 16110 41970
rect 10558 41906 10610 41918
rect 14366 41906 14418 41918
rect 17726 41906 17778 41918
rect 17950 41970 18002 41982
rect 17950 41906 18002 41918
rect 18174 41970 18226 41982
rect 18174 41906 18226 41918
rect 18398 41970 18450 41982
rect 18398 41906 18450 41918
rect 18734 41970 18786 41982
rect 18734 41906 18786 41918
rect 18846 41970 18898 41982
rect 18846 41906 18898 41918
rect 19070 41970 19122 41982
rect 19070 41906 19122 41918
rect 19294 41970 19346 41982
rect 21198 41970 21250 41982
rect 20962 41918 20974 41970
rect 21026 41918 21038 41970
rect 19294 41906 19346 41918
rect 21198 41906 21250 41918
rect 21310 41970 21362 41982
rect 21310 41906 21362 41918
rect 21534 41970 21586 41982
rect 21534 41906 21586 41918
rect 25566 41970 25618 41982
rect 32510 41970 32562 41982
rect 25890 41918 25902 41970
rect 25954 41918 25966 41970
rect 31938 41918 31950 41970
rect 32002 41918 32014 41970
rect 25566 41906 25618 41918
rect 32510 41906 32562 41918
rect 34526 41970 34578 41982
rect 38222 41970 38274 41982
rect 39790 41970 39842 41982
rect 34850 41918 34862 41970
rect 34914 41918 34926 41970
rect 38994 41918 39006 41970
rect 39058 41918 39070 41970
rect 34526 41906 34578 41918
rect 38222 41906 38274 41918
rect 39790 41906 39842 41918
rect 41022 41970 41074 41982
rect 41022 41906 41074 41918
rect 41582 41970 41634 41982
rect 41582 41906 41634 41918
rect 41806 41970 41858 41982
rect 41806 41906 41858 41918
rect 42030 41970 42082 41982
rect 42030 41906 42082 41918
rect 42142 41970 42194 41982
rect 42142 41906 42194 41918
rect 42366 41970 42418 41982
rect 42366 41906 42418 41918
rect 43038 41970 43090 41982
rect 43038 41906 43090 41918
rect 43598 41970 43650 41982
rect 43598 41906 43650 41918
rect 45278 41970 45330 41982
rect 45278 41906 45330 41918
rect 45502 41970 45554 41982
rect 45502 41906 45554 41918
rect 46958 41970 47010 41982
rect 46958 41906 47010 41918
rect 47630 41970 47682 41982
rect 47630 41906 47682 41918
rect 48302 41970 48354 41982
rect 49198 41970 49250 41982
rect 53118 41970 53170 41982
rect 48962 41918 48974 41970
rect 49026 41918 49038 41970
rect 51314 41918 51326 41970
rect 51378 41918 51390 41970
rect 52210 41918 52222 41970
rect 52274 41918 52286 41970
rect 52434 41918 52446 41970
rect 52498 41918 52510 41970
rect 48302 41906 48354 41918
rect 49198 41906 49250 41918
rect 53118 41906 53170 41918
rect 53454 41970 53506 41982
rect 53454 41906 53506 41918
rect 56030 41970 56082 41982
rect 57026 41918 57038 41970
rect 57090 41918 57102 41970
rect 56030 41906 56082 41918
rect 34302 41858 34354 41870
rect 6850 41806 6862 41858
rect 6914 41806 6926 41858
rect 8978 41806 8990 41858
rect 9042 41806 9054 41858
rect 11890 41806 11902 41858
rect 11954 41806 11966 41858
rect 14018 41806 14030 41858
rect 14082 41806 14094 41858
rect 15474 41806 15486 41858
rect 15538 41806 15550 41858
rect 26674 41806 26686 41858
rect 26738 41806 26750 41858
rect 28802 41806 28814 41858
rect 28866 41806 28878 41858
rect 29138 41806 29150 41858
rect 29202 41806 29214 41858
rect 34302 41794 34354 41806
rect 38446 41858 38498 41870
rect 38446 41794 38498 41806
rect 43262 41858 43314 41870
rect 43262 41794 43314 41806
rect 46622 41858 46674 41870
rect 46622 41794 46674 41806
rect 47742 41858 47794 41870
rect 52894 41858 52946 41870
rect 50194 41806 50206 41858
rect 50258 41806 50270 41858
rect 51090 41806 51102 41858
rect 51154 41806 51166 41858
rect 47742 41794 47794 41806
rect 52894 41794 52946 41806
rect 53006 41858 53058 41870
rect 53006 41794 53058 41806
rect 53566 41858 53618 41870
rect 53566 41794 53618 41806
rect 54014 41858 54066 41870
rect 54014 41794 54066 41806
rect 54462 41858 54514 41870
rect 54462 41794 54514 41806
rect 54910 41858 54962 41870
rect 55682 41806 55694 41858
rect 55746 41806 55758 41858
rect 57250 41806 57262 41858
rect 57314 41806 57326 41858
rect 54910 41794 54962 41806
rect 38670 41746 38722 41758
rect 38670 41682 38722 41694
rect 40126 41746 40178 41758
rect 40126 41682 40178 41694
rect 40910 41746 40962 41758
rect 40910 41682 40962 41694
rect 42814 41746 42866 41758
rect 42814 41682 42866 41694
rect 49086 41746 49138 41758
rect 49086 41682 49138 41694
rect 52670 41746 52722 41758
rect 54002 41694 54014 41746
rect 54066 41743 54078 41746
rect 54226 41743 54238 41746
rect 54066 41697 54238 41743
rect 54066 41694 54078 41697
rect 54226 41694 54238 41697
rect 54290 41694 54302 41746
rect 52670 41682 52722 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 17278 41410 17330 41422
rect 17278 41346 17330 41358
rect 18062 41410 18114 41422
rect 18062 41346 18114 41358
rect 19518 41410 19570 41422
rect 19518 41346 19570 41358
rect 51662 41410 51714 41422
rect 51662 41346 51714 41358
rect 9886 41298 9938 41310
rect 9886 41234 9938 41246
rect 14254 41298 14306 41310
rect 14254 41234 14306 41246
rect 16718 41298 16770 41310
rect 16718 41234 16770 41246
rect 19854 41298 19906 41310
rect 19854 41234 19906 41246
rect 21422 41298 21474 41310
rect 40126 41298 40178 41310
rect 22418 41246 22430 41298
rect 22482 41246 22494 41298
rect 25666 41246 25678 41298
rect 25730 41246 25742 41298
rect 30594 41246 30606 41298
rect 30658 41246 30670 41298
rect 34626 41246 34638 41298
rect 34690 41246 34702 41298
rect 21422 41234 21474 41246
rect 40126 41234 40178 41246
rect 41918 41298 41970 41310
rect 50654 41298 50706 41310
rect 46162 41246 46174 41298
rect 46226 41246 46238 41298
rect 41918 41234 41970 41246
rect 50654 41234 50706 41246
rect 51550 41298 51602 41310
rect 53442 41246 53454 41298
rect 53506 41246 53518 41298
rect 55570 41246 55582 41298
rect 55634 41246 55646 41298
rect 57250 41246 57262 41298
rect 57314 41246 57326 41298
rect 51550 41234 51602 41246
rect 10110 41186 10162 41198
rect 14366 41186 14418 41198
rect 13570 41134 13582 41186
rect 13634 41134 13646 41186
rect 10110 41122 10162 41134
rect 14366 41122 14418 41134
rect 14814 41186 14866 41198
rect 14814 41122 14866 41134
rect 15038 41186 15090 41198
rect 15038 41122 15090 41134
rect 15262 41186 15314 41198
rect 15262 41122 15314 41134
rect 16270 41186 16322 41198
rect 16270 41122 16322 41134
rect 16942 41186 16994 41198
rect 16942 41122 16994 41134
rect 18286 41186 18338 41198
rect 19742 41186 19794 41198
rect 29262 41186 29314 41198
rect 19282 41134 19294 41186
rect 19346 41134 19358 41186
rect 25330 41134 25342 41186
rect 25394 41134 25406 41186
rect 28578 41134 28590 41186
rect 28642 41134 28654 41186
rect 18286 41122 18338 41134
rect 19742 41122 19794 41134
rect 29262 41122 29314 41134
rect 31390 41186 31442 41198
rect 39230 41186 39282 41198
rect 31714 41134 31726 41186
rect 31778 41134 31790 41186
rect 31390 41122 31442 41134
rect 39230 41122 39282 41134
rect 39790 41186 39842 41198
rect 39790 41122 39842 41134
rect 39902 41186 39954 41198
rect 39902 41122 39954 41134
rect 40350 41186 40402 41198
rect 49982 41186 50034 41198
rect 44930 41134 44942 41186
rect 44994 41134 45006 41186
rect 48962 41134 48974 41186
rect 49026 41134 49038 41186
rect 40350 41122 40402 41134
rect 49982 41122 50034 41134
rect 50094 41186 50146 41198
rect 50094 41122 50146 41134
rect 50542 41186 50594 41198
rect 50542 41122 50594 41134
rect 50990 41186 51042 41198
rect 50990 41122 51042 41134
rect 51886 41186 51938 41198
rect 52658 41134 52670 41186
rect 52722 41134 52734 41186
rect 57586 41134 57598 41186
rect 57650 41134 57662 41186
rect 51886 41122 51938 41134
rect 15934 41074 15986 41086
rect 15934 41010 15986 41022
rect 17614 41074 17666 41086
rect 18510 41074 18562 41086
rect 17826 41022 17838 41074
rect 17890 41022 17902 41074
rect 17614 41010 17666 41022
rect 18510 41010 18562 41022
rect 19070 41074 19122 41086
rect 19070 41010 19122 41022
rect 19966 41074 20018 41086
rect 19966 41010 20018 41022
rect 20638 41074 20690 41086
rect 31054 41074 31106 41086
rect 24546 41022 24558 41074
rect 24610 41022 24622 41074
rect 27794 41022 27806 41074
rect 27858 41022 27870 41074
rect 30818 41022 30830 41074
rect 30882 41022 30894 41074
rect 20638 41010 20690 41022
rect 31054 41010 31106 41022
rect 31166 41074 31218 41086
rect 35086 41074 35138 41086
rect 32498 41022 32510 41074
rect 32562 41022 32574 41074
rect 31166 41010 31218 41022
rect 35086 41010 35138 41022
rect 35198 41074 35250 41086
rect 35198 41010 35250 41022
rect 39454 41074 39506 41086
rect 39454 41010 39506 41022
rect 40910 41074 40962 41086
rect 40910 41010 40962 41022
rect 41358 41074 41410 41086
rect 41358 41010 41410 41022
rect 41470 41074 41522 41086
rect 50206 41074 50258 41086
rect 43026 41022 43038 41074
rect 43090 41022 43102 41074
rect 45154 41022 45166 41074
rect 45218 41022 45230 41074
rect 48290 41022 48302 41074
rect 48354 41022 48366 41074
rect 41470 41010 41522 41022
rect 50206 41010 50258 41022
rect 50878 41074 50930 41086
rect 50878 41010 50930 41022
rect 51998 41074 52050 41086
rect 51998 41010 52050 41022
rect 56702 41074 56754 41086
rect 56702 41010 56754 41022
rect 5070 40962 5122 40974
rect 5070 40898 5122 40910
rect 9214 40962 9266 40974
rect 14142 40962 14194 40974
rect 10434 40910 10446 40962
rect 10498 40910 10510 40962
rect 13794 40910 13806 40962
rect 13858 40910 13870 40962
rect 9214 40898 9266 40910
rect 14142 40898 14194 40910
rect 15150 40962 15202 40974
rect 15150 40898 15202 40910
rect 15486 40962 15538 40974
rect 15486 40898 15538 40910
rect 16046 40962 16098 40974
rect 20302 40962 20354 40974
rect 17938 40910 17950 40962
rect 18002 40910 18014 40962
rect 16046 40898 16098 40910
rect 20302 40898 20354 40910
rect 21310 40962 21362 40974
rect 21310 40898 21362 40910
rect 21534 40962 21586 40974
rect 21534 40898 21586 40910
rect 21758 40962 21810 40974
rect 21758 40898 21810 40910
rect 34862 40962 34914 40974
rect 34862 40898 34914 40910
rect 35646 40962 35698 40974
rect 35646 40898 35698 40910
rect 36094 40962 36146 40974
rect 36094 40898 36146 40910
rect 37550 40962 37602 40974
rect 40574 40962 40626 40974
rect 39778 40910 39790 40962
rect 39842 40910 39854 40962
rect 37550 40898 37602 40910
rect 40574 40898 40626 40910
rect 40798 40962 40850 40974
rect 40798 40898 40850 40910
rect 41134 40962 41186 40974
rect 41134 40898 41186 40910
rect 42702 40962 42754 40974
rect 42702 40898 42754 40910
rect 43374 40962 43426 40974
rect 43374 40898 43426 40910
rect 43822 40962 43874 40974
rect 43822 40898 43874 40910
rect 49758 40962 49810 40974
rect 49758 40898 49810 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 8094 40626 8146 40638
rect 8094 40562 8146 40574
rect 8878 40626 8930 40638
rect 12014 40626 12066 40638
rect 8878 40562 8930 40574
rect 11230 40570 11282 40582
rect 9886 40514 9938 40526
rect 7634 40462 7646 40514
rect 7698 40462 7710 40514
rect 9886 40450 9938 40462
rect 10110 40514 10162 40526
rect 10110 40450 10162 40462
rect 10558 40514 10610 40526
rect 12014 40562 12066 40574
rect 13470 40626 13522 40638
rect 16382 40626 16434 40638
rect 20638 40626 20690 40638
rect 23214 40626 23266 40638
rect 14802 40574 14814 40626
rect 14866 40574 14878 40626
rect 19282 40574 19294 40626
rect 19346 40574 19358 40626
rect 22306 40574 22318 40626
rect 22370 40574 22382 40626
rect 13470 40562 13522 40574
rect 16382 40562 16434 40574
rect 20638 40562 20690 40574
rect 23214 40562 23266 40574
rect 26462 40626 26514 40638
rect 26462 40562 26514 40574
rect 27918 40626 27970 40638
rect 27918 40562 27970 40574
rect 33518 40626 33570 40638
rect 33518 40562 33570 40574
rect 39678 40626 39730 40638
rect 39678 40562 39730 40574
rect 41022 40626 41074 40638
rect 41022 40562 41074 40574
rect 41806 40626 41858 40638
rect 41806 40562 41858 40574
rect 42030 40626 42082 40638
rect 42030 40562 42082 40574
rect 43038 40626 43090 40638
rect 43038 40562 43090 40574
rect 43598 40626 43650 40638
rect 43598 40562 43650 40574
rect 47294 40626 47346 40638
rect 47294 40562 47346 40574
rect 47854 40626 47906 40638
rect 47854 40562 47906 40574
rect 48750 40626 48802 40638
rect 48750 40562 48802 40574
rect 49534 40626 49586 40638
rect 56914 40574 56926 40626
rect 56978 40574 56990 40626
rect 49534 40562 49586 40574
rect 10882 40462 10894 40514
rect 10946 40462 10958 40514
rect 11230 40506 11282 40518
rect 11342 40514 11394 40526
rect 16270 40514 16322 40526
rect 24222 40514 24274 40526
rect 15922 40462 15934 40514
rect 15986 40462 15998 40514
rect 18498 40462 18510 40514
rect 18562 40462 18574 40514
rect 10558 40450 10610 40462
rect 11342 40450 11394 40462
rect 16270 40450 16322 40462
rect 24222 40450 24274 40462
rect 24558 40514 24610 40526
rect 39902 40514 39954 40526
rect 27570 40462 27582 40514
rect 27634 40462 27646 40514
rect 31154 40462 31166 40514
rect 31218 40462 31230 40514
rect 36530 40462 36542 40514
rect 36594 40462 36606 40514
rect 24558 40450 24610 40462
rect 39902 40450 39954 40462
rect 40126 40514 40178 40526
rect 40126 40450 40178 40462
rect 44046 40514 44098 40526
rect 44046 40450 44098 40462
rect 47630 40514 47682 40526
rect 47630 40450 47682 40462
rect 49086 40514 49138 40526
rect 54686 40514 54738 40526
rect 50866 40462 50878 40514
rect 50930 40462 50942 40514
rect 49086 40450 49138 40462
rect 54686 40450 54738 40462
rect 55022 40514 55074 40526
rect 57026 40462 57038 40514
rect 57090 40462 57102 40514
rect 57362 40462 57374 40514
rect 57426 40462 57438 40514
rect 55022 40450 55074 40462
rect 7310 40402 7362 40414
rect 4050 40350 4062 40402
rect 4114 40350 4126 40402
rect 4834 40350 4846 40402
rect 4898 40350 4910 40402
rect 7310 40338 7362 40350
rect 8542 40402 8594 40414
rect 8542 40338 8594 40350
rect 10222 40402 10274 40414
rect 12462 40402 12514 40414
rect 12002 40350 12014 40402
rect 12066 40350 12078 40402
rect 10222 40338 10274 40350
rect 12462 40338 12514 40350
rect 12798 40402 12850 40414
rect 12798 40338 12850 40350
rect 13582 40402 13634 40414
rect 13582 40338 13634 40350
rect 13806 40402 13858 40414
rect 13806 40338 13858 40350
rect 14254 40402 14306 40414
rect 14254 40338 14306 40350
rect 14478 40402 14530 40414
rect 20862 40402 20914 40414
rect 15698 40350 15710 40402
rect 15762 40350 15774 40402
rect 18834 40350 18846 40402
rect 18898 40350 18910 40402
rect 19506 40350 19518 40402
rect 19570 40350 19582 40402
rect 14478 40338 14530 40350
rect 20862 40338 20914 40350
rect 21086 40402 21138 40414
rect 26350 40402 26402 40414
rect 22530 40350 22542 40402
rect 22594 40350 22606 40402
rect 21086 40338 21138 40350
rect 26350 40338 26402 40350
rect 26574 40402 26626 40414
rect 32062 40402 32114 40414
rect 26898 40350 26910 40402
rect 26962 40350 26974 40402
rect 30930 40350 30942 40402
rect 30994 40350 31006 40402
rect 26574 40338 26626 40350
rect 32062 40338 32114 40350
rect 32510 40402 32562 40414
rect 32510 40338 32562 40350
rect 33070 40402 33122 40414
rect 33070 40338 33122 40350
rect 33406 40402 33458 40414
rect 33406 40338 33458 40350
rect 33742 40402 33794 40414
rect 38782 40402 38834 40414
rect 37202 40350 37214 40402
rect 37266 40350 37278 40402
rect 37874 40350 37886 40402
rect 37938 40350 37950 40402
rect 33742 40338 33794 40350
rect 38782 40338 38834 40350
rect 39454 40402 39506 40414
rect 39454 40338 39506 40350
rect 42254 40402 42306 40414
rect 42254 40338 42306 40350
rect 42926 40402 42978 40414
rect 42926 40338 42978 40350
rect 43262 40402 43314 40414
rect 43262 40338 43314 40350
rect 43374 40402 43426 40414
rect 43374 40338 43426 40350
rect 43822 40402 43874 40414
rect 43822 40338 43874 40350
rect 44382 40402 44434 40414
rect 44382 40338 44434 40350
rect 44718 40402 44770 40414
rect 46062 40402 46114 40414
rect 51662 40402 51714 40414
rect 54350 40402 54402 40414
rect 55918 40402 55970 40414
rect 44930 40350 44942 40402
rect 44994 40350 45006 40402
rect 45490 40350 45502 40402
rect 45554 40350 45566 40402
rect 50194 40350 50206 40402
rect 50258 40350 50270 40402
rect 51874 40350 51886 40402
rect 51938 40350 51950 40402
rect 54002 40350 54014 40402
rect 54066 40350 54078 40402
rect 55682 40350 55694 40402
rect 55746 40350 55758 40402
rect 44718 40338 44770 40350
rect 46062 40338 46114 40350
rect 51662 40338 51714 40350
rect 54350 40338 54402 40350
rect 55918 40338 55970 40350
rect 56590 40402 56642 40414
rect 56590 40338 56642 40350
rect 3278 40290 3330 40302
rect 9774 40290 9826 40302
rect 6962 40238 6974 40290
rect 7026 40238 7038 40290
rect 3278 40226 3330 40238
rect 9774 40226 9826 40238
rect 20974 40290 21026 40302
rect 31614 40290 31666 40302
rect 42142 40290 42194 40302
rect 23202 40238 23214 40290
rect 23266 40238 23278 40290
rect 34402 40238 34414 40290
rect 34466 40238 34478 40290
rect 38098 40238 38110 40290
rect 38162 40238 38174 40290
rect 20974 40226 21026 40238
rect 31614 40226 31666 40238
rect 42142 40226 42194 40238
rect 44494 40290 44546 40302
rect 53678 40290 53730 40302
rect 47954 40238 47966 40290
rect 48018 40238 48030 40290
rect 53890 40238 53902 40290
rect 53954 40238 53966 40290
rect 44494 40226 44546 40238
rect 53678 40226 53730 40238
rect 2942 40178 2994 40190
rect 2942 40114 2994 40126
rect 3054 40178 3106 40190
rect 3054 40114 3106 40126
rect 3390 40178 3442 40190
rect 3390 40114 3442 40126
rect 8766 40178 8818 40190
rect 8766 40114 8818 40126
rect 8878 40178 8930 40190
rect 8878 40114 8930 40126
rect 11342 40178 11394 40190
rect 11342 40114 11394 40126
rect 12350 40178 12402 40190
rect 12350 40114 12402 40126
rect 13470 40178 13522 40190
rect 13470 40114 13522 40126
rect 22990 40178 23042 40190
rect 22990 40114 23042 40126
rect 44830 40178 44882 40190
rect 44830 40114 44882 40126
rect 45838 40178 45890 40190
rect 50978 40126 50990 40178
rect 51042 40126 51054 40178
rect 45838 40114 45890 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 10110 39842 10162 39854
rect 41010 39790 41022 39842
rect 41074 39790 41086 39842
rect 50866 39790 50878 39842
rect 50930 39790 50942 39842
rect 10110 39778 10162 39790
rect 5742 39730 5794 39742
rect 11118 39730 11170 39742
rect 2482 39678 2494 39730
rect 2546 39678 2558 39730
rect 7970 39678 7982 39730
rect 8034 39678 8046 39730
rect 9314 39678 9326 39730
rect 9378 39678 9390 39730
rect 5742 39666 5794 39678
rect 11118 39666 11170 39678
rect 13582 39730 13634 39742
rect 17166 39730 17218 39742
rect 16146 39678 16158 39730
rect 16210 39678 16222 39730
rect 13582 39666 13634 39678
rect 17166 39666 17218 39678
rect 17502 39730 17554 39742
rect 17502 39666 17554 39678
rect 18846 39730 18898 39742
rect 18846 39666 18898 39678
rect 19294 39730 19346 39742
rect 19294 39666 19346 39678
rect 26350 39730 26402 39742
rect 26350 39666 26402 39678
rect 26910 39730 26962 39742
rect 26910 39666 26962 39678
rect 27582 39730 27634 39742
rect 27582 39666 27634 39678
rect 30494 39730 30546 39742
rect 30494 39666 30546 39678
rect 38222 39730 38274 39742
rect 43486 39730 43538 39742
rect 41234 39678 41246 39730
rect 41298 39678 41310 39730
rect 38222 39666 38274 39678
rect 43486 39666 43538 39678
rect 44942 39730 44994 39742
rect 54126 39730 54178 39742
rect 51314 39678 51326 39730
rect 51378 39678 51390 39730
rect 55794 39678 55806 39730
rect 55858 39678 55870 39730
rect 57922 39678 57934 39730
rect 57986 39678 57998 39730
rect 44942 39666 44994 39678
rect 54126 39666 54178 39678
rect 6078 39618 6130 39630
rect 7422 39618 7474 39630
rect 9662 39618 9714 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 6402 39566 6414 39618
rect 6466 39566 6478 39618
rect 8306 39566 8318 39618
rect 8370 39566 8382 39618
rect 6078 39554 6130 39566
rect 7422 39554 7474 39566
rect 9662 39554 9714 39566
rect 9886 39618 9938 39630
rect 9886 39554 9938 39566
rect 11006 39618 11058 39630
rect 11006 39554 11058 39566
rect 13470 39618 13522 39630
rect 13470 39554 13522 39566
rect 13694 39618 13746 39630
rect 13694 39554 13746 39566
rect 14030 39618 14082 39630
rect 14030 39554 14082 39566
rect 15486 39618 15538 39630
rect 16606 39618 16658 39630
rect 15810 39566 15822 39618
rect 15874 39566 15886 39618
rect 15486 39554 15538 39566
rect 16606 39554 16658 39566
rect 17838 39618 17890 39630
rect 17838 39554 17890 39566
rect 18286 39618 18338 39630
rect 18286 39554 18338 39566
rect 18510 39618 18562 39630
rect 18510 39554 18562 39566
rect 22094 39618 22146 39630
rect 30718 39618 30770 39630
rect 23426 39566 23438 39618
rect 23490 39566 23502 39618
rect 26562 39566 26574 39618
rect 26626 39566 26638 39618
rect 27794 39566 27806 39618
rect 27858 39566 27870 39618
rect 28018 39566 28030 39618
rect 28082 39566 28094 39618
rect 22094 39554 22146 39566
rect 30718 39554 30770 39566
rect 36094 39618 36146 39630
rect 38110 39618 38162 39630
rect 42926 39618 42978 39630
rect 37762 39566 37774 39618
rect 37826 39566 37838 39618
rect 40002 39566 40014 39618
rect 40066 39566 40078 39618
rect 41122 39566 41134 39618
rect 41186 39566 41198 39618
rect 36094 39554 36146 39566
rect 38110 39554 38162 39566
rect 42926 39554 42978 39566
rect 45166 39618 45218 39630
rect 45166 39554 45218 39566
rect 45390 39618 45442 39630
rect 51090 39566 51102 39618
rect 51154 39566 51166 39618
rect 51426 39566 51438 39618
rect 51490 39566 51502 39618
rect 55010 39566 55022 39618
rect 55074 39566 55086 39618
rect 45390 39554 45442 39566
rect 5630 39506 5682 39518
rect 8766 39506 8818 39518
rect 5842 39454 5854 39506
rect 5906 39454 5918 39506
rect 7074 39454 7086 39506
rect 7138 39454 7150 39506
rect 5630 39442 5682 39454
rect 8766 39442 8818 39454
rect 10446 39506 10498 39518
rect 10446 39442 10498 39454
rect 12910 39506 12962 39518
rect 12910 39442 12962 39454
rect 17726 39506 17778 39518
rect 17726 39442 17778 39454
rect 20078 39506 20130 39518
rect 20078 39442 20130 39454
rect 21534 39506 21586 39518
rect 21534 39442 21586 39454
rect 23774 39506 23826 39518
rect 44830 39506 44882 39518
rect 40114 39454 40126 39506
rect 40178 39454 40190 39506
rect 23774 39442 23826 39454
rect 44830 39442 44882 39454
rect 52894 39506 52946 39518
rect 52894 39442 52946 39454
rect 53006 39506 53058 39518
rect 54350 39506 54402 39518
rect 53106 39454 53118 39506
rect 53170 39454 53182 39506
rect 53006 39442 53058 39454
rect 54350 39442 54402 39454
rect 9214 39394 9266 39406
rect 4722 39342 4734 39394
rect 4786 39342 4798 39394
rect 9214 39330 9266 39342
rect 9438 39394 9490 39406
rect 9438 39330 9490 39342
rect 10558 39394 10610 39406
rect 10558 39330 10610 39342
rect 10782 39394 10834 39406
rect 10782 39330 10834 39342
rect 11566 39394 11618 39406
rect 11566 39330 11618 39342
rect 12798 39394 12850 39406
rect 12798 39330 12850 39342
rect 20190 39394 20242 39406
rect 20190 39330 20242 39342
rect 23662 39394 23714 39406
rect 23662 39330 23714 39342
rect 26238 39394 26290 39406
rect 26238 39330 26290 39342
rect 26462 39394 26514 39406
rect 36430 39394 36482 39406
rect 31042 39342 31054 39394
rect 31106 39342 31118 39394
rect 26462 39330 26514 39342
rect 36430 39330 36482 39342
rect 44046 39394 44098 39406
rect 44046 39330 44098 39342
rect 48414 39394 48466 39406
rect 48414 39330 48466 39342
rect 50430 39394 50482 39406
rect 50430 39330 50482 39342
rect 52670 39394 52722 39406
rect 52670 39330 52722 39342
rect 52782 39394 52834 39406
rect 53778 39342 53790 39394
rect 53842 39342 53854 39394
rect 52782 39330 52834 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 3950 39058 4002 39070
rect 10334 39058 10386 39070
rect 3490 39006 3502 39058
rect 3554 39006 3566 39058
rect 7186 39006 7198 39058
rect 7250 39006 7262 39058
rect 8530 39006 8542 39058
rect 8594 39006 8606 39058
rect 3950 38994 4002 39006
rect 10334 38994 10386 39006
rect 11566 39058 11618 39070
rect 11566 38994 11618 39006
rect 11902 39058 11954 39070
rect 11902 38994 11954 39006
rect 13470 39058 13522 39070
rect 13470 38994 13522 39006
rect 15934 39058 15986 39070
rect 24446 39058 24498 39070
rect 15934 38994 15986 39006
rect 17726 39002 17778 39014
rect 19730 39006 19742 39058
rect 19794 39006 19806 39058
rect 2942 38946 2994 38958
rect 2942 38882 2994 38894
rect 10222 38946 10274 38958
rect 12798 38946 12850 38958
rect 10658 38894 10670 38946
rect 10722 38894 10734 38946
rect 10222 38882 10274 38894
rect 12798 38882 12850 38894
rect 13582 38946 13634 38958
rect 13582 38882 13634 38894
rect 14926 38946 14978 38958
rect 14926 38882 14978 38894
rect 15374 38946 15426 38958
rect 15374 38882 15426 38894
rect 17614 38946 17666 38958
rect 24446 38994 24498 39006
rect 24558 39058 24610 39070
rect 27806 39058 27858 39070
rect 27010 39006 27022 39058
rect 27074 39006 27086 39058
rect 24558 38994 24610 39006
rect 27806 38994 27858 39006
rect 28030 39058 28082 39070
rect 28030 38994 28082 39006
rect 30046 39058 30098 39070
rect 30046 38994 30098 39006
rect 30942 39058 30994 39070
rect 30942 38994 30994 39006
rect 34302 39058 34354 39070
rect 34302 38994 34354 39006
rect 34638 39058 34690 39070
rect 34638 38994 34690 39006
rect 36990 39058 37042 39070
rect 36990 38994 37042 39006
rect 37214 39058 37266 39070
rect 37214 38994 37266 39006
rect 37774 39058 37826 39070
rect 37774 38994 37826 39006
rect 40238 39058 40290 39070
rect 40238 38994 40290 39006
rect 40462 39058 40514 39070
rect 40462 38994 40514 39006
rect 41022 39058 41074 39070
rect 41022 38994 41074 39006
rect 44382 39058 44434 39070
rect 44382 38994 44434 39006
rect 48078 39058 48130 39070
rect 48078 38994 48130 39006
rect 50990 39058 51042 39070
rect 50990 38994 51042 39006
rect 51438 39058 51490 39070
rect 55022 39058 55074 39070
rect 53666 39006 53678 39058
rect 53730 39006 53742 39058
rect 51438 38994 51490 39006
rect 55022 38994 55074 39006
rect 55470 39058 55522 39070
rect 57486 39058 57538 39070
rect 57138 39006 57150 39058
rect 57202 39006 57214 39058
rect 55470 38994 55522 39006
rect 57486 38994 57538 39006
rect 17726 38938 17778 38950
rect 19182 38946 19234 38958
rect 18274 38894 18286 38946
rect 18338 38894 18350 38946
rect 17614 38882 17666 38894
rect 19182 38882 19234 38894
rect 21534 38946 21586 38958
rect 25230 38946 25282 38958
rect 21746 38894 21758 38946
rect 21810 38894 21822 38946
rect 23538 38894 23550 38946
rect 23602 38894 23614 38946
rect 21534 38882 21586 38894
rect 25230 38882 25282 38894
rect 27582 38946 27634 38958
rect 36654 38946 36706 38958
rect 40126 38946 40178 38958
rect 28354 38894 28366 38946
rect 28418 38894 28430 38946
rect 28914 38894 28926 38946
rect 28978 38894 28990 38946
rect 29698 38894 29710 38946
rect 29762 38894 29774 38946
rect 39554 38894 39566 38946
rect 39618 38894 39630 38946
rect 27582 38882 27634 38894
rect 36654 38882 36706 38894
rect 40126 38882 40178 38894
rect 41358 38946 41410 38958
rect 41358 38882 41410 38894
rect 43598 38946 43650 38958
rect 51326 38946 51378 38958
rect 43810 38894 43822 38946
rect 43874 38894 43886 38946
rect 46834 38894 46846 38946
rect 46898 38894 46910 38946
rect 50642 38894 50654 38946
rect 50706 38894 50718 38946
rect 43598 38882 43650 38894
rect 51326 38882 51378 38894
rect 53118 38946 53170 38958
rect 53118 38882 53170 38894
rect 53230 38946 53282 38958
rect 53230 38882 53282 38894
rect 55918 38946 55970 38958
rect 55918 38882 55970 38894
rect 3054 38834 3106 38846
rect 2706 38782 2718 38834
rect 2770 38782 2782 38834
rect 3054 38770 3106 38782
rect 3726 38834 3778 38846
rect 3726 38770 3778 38782
rect 4174 38834 4226 38846
rect 4174 38770 4226 38782
rect 4286 38834 4338 38846
rect 4286 38770 4338 38782
rect 4734 38834 4786 38846
rect 4734 38770 4786 38782
rect 5182 38834 5234 38846
rect 6302 38834 6354 38846
rect 6066 38782 6078 38834
rect 6130 38782 6142 38834
rect 5182 38770 5234 38782
rect 6302 38770 6354 38782
rect 6414 38834 6466 38846
rect 6414 38770 6466 38782
rect 7534 38834 7586 38846
rect 8542 38834 8594 38846
rect 8990 38834 9042 38846
rect 8306 38782 8318 38834
rect 8370 38782 8382 38834
rect 8754 38782 8766 38834
rect 8818 38782 8830 38834
rect 7534 38770 7586 38782
rect 8542 38770 8594 38782
rect 8990 38770 9042 38782
rect 9662 38834 9714 38846
rect 10894 38834 10946 38846
rect 9986 38782 9998 38834
rect 10050 38782 10062 38834
rect 9662 38770 9714 38782
rect 10894 38770 10946 38782
rect 11342 38834 11394 38846
rect 11342 38770 11394 38782
rect 12350 38834 12402 38846
rect 12350 38770 12402 38782
rect 13022 38834 13074 38846
rect 13022 38770 13074 38782
rect 13694 38834 13746 38846
rect 13694 38770 13746 38782
rect 14142 38834 14194 38846
rect 14142 38770 14194 38782
rect 14254 38834 14306 38846
rect 14254 38770 14306 38782
rect 14590 38834 14642 38846
rect 14590 38770 14642 38782
rect 15486 38834 15538 38846
rect 16830 38834 16882 38846
rect 16370 38782 16382 38834
rect 16434 38782 16446 38834
rect 15486 38770 15538 38782
rect 16830 38770 16882 38782
rect 18510 38834 18562 38846
rect 19406 38834 19458 38846
rect 18722 38782 18734 38834
rect 18786 38782 18798 38834
rect 18510 38770 18562 38782
rect 19406 38770 19458 38782
rect 20302 38834 20354 38846
rect 20302 38770 20354 38782
rect 20862 38834 20914 38846
rect 20862 38770 20914 38782
rect 21086 38834 21138 38846
rect 21086 38770 21138 38782
rect 21870 38834 21922 38846
rect 24110 38834 24162 38846
rect 22082 38782 22094 38834
rect 22146 38782 22158 38834
rect 22866 38782 22878 38834
rect 22930 38782 22942 38834
rect 21870 38770 21922 38782
rect 24110 38770 24162 38782
rect 24334 38834 24386 38846
rect 24334 38770 24386 38782
rect 25342 38834 25394 38846
rect 25342 38770 25394 38782
rect 26686 38834 26738 38846
rect 26686 38770 26738 38782
rect 27470 38834 27522 38846
rect 27470 38770 27522 38782
rect 29262 38834 29314 38846
rect 31838 38834 31890 38846
rect 31378 38782 31390 38834
rect 31442 38782 31454 38834
rect 29262 38770 29314 38782
rect 31838 38770 31890 38782
rect 35198 38834 35250 38846
rect 37326 38834 37378 38846
rect 35746 38782 35758 38834
rect 35810 38782 35822 38834
rect 35198 38770 35250 38782
rect 37326 38770 37378 38782
rect 37662 38834 37714 38846
rect 37662 38770 37714 38782
rect 37998 38834 38050 38846
rect 41694 38834 41746 38846
rect 42366 38834 42418 38846
rect 38546 38782 38558 38834
rect 38610 38782 38622 38834
rect 39218 38782 39230 38834
rect 39282 38782 39294 38834
rect 39442 38782 39454 38834
rect 39506 38782 39518 38834
rect 41906 38782 41918 38834
rect 41970 38782 41982 38834
rect 37998 38770 38050 38782
rect 41694 38770 41746 38782
rect 42366 38770 42418 38782
rect 42702 38834 42754 38846
rect 42702 38770 42754 38782
rect 42926 38834 42978 38846
rect 50430 38834 50482 38846
rect 44146 38782 44158 38834
rect 44210 38782 44222 38834
rect 47618 38782 47630 38834
rect 47682 38782 47694 38834
rect 48850 38782 48862 38834
rect 48914 38782 48926 38834
rect 42926 38770 42978 38782
rect 50430 38770 50482 38782
rect 52222 38834 52274 38846
rect 56702 38834 56754 38846
rect 52882 38782 52894 38834
rect 52946 38782 52958 38834
rect 52222 38770 52274 38782
rect 56702 38770 56754 38782
rect 4846 38722 4898 38734
rect 10558 38722 10610 38734
rect 6850 38670 6862 38722
rect 6914 38670 6926 38722
rect 4846 38658 4898 38670
rect 10558 38658 10610 38670
rect 13134 38722 13186 38734
rect 13134 38658 13186 38670
rect 14478 38722 14530 38734
rect 14478 38658 14530 38670
rect 18174 38722 18226 38734
rect 18174 38658 18226 38670
rect 20078 38722 20130 38734
rect 26462 38722 26514 38734
rect 22754 38670 22766 38722
rect 22818 38670 22830 38722
rect 20078 38658 20130 38670
rect 26462 38658 26514 38670
rect 30382 38722 30434 38734
rect 41470 38722 41522 38734
rect 36082 38670 36094 38722
rect 36146 38670 36158 38722
rect 30382 38658 30434 38670
rect 41470 38658 41522 38670
rect 42590 38722 42642 38734
rect 52334 38722 52386 38734
rect 44706 38670 44718 38722
rect 44770 38670 44782 38722
rect 49186 38670 49198 38722
rect 49250 38670 49262 38722
rect 42590 38658 42642 38670
rect 52334 38658 52386 38670
rect 54126 38722 54178 38734
rect 54126 38658 54178 38670
rect 54574 38722 54626 38734
rect 54574 38658 54626 38670
rect 56590 38722 56642 38734
rect 56590 38658 56642 38670
rect 5406 38610 5458 38622
rect 12574 38610 12626 38622
rect 5730 38558 5742 38610
rect 5794 38558 5806 38610
rect 5406 38546 5458 38558
rect 12574 38546 12626 38558
rect 15374 38610 15426 38622
rect 15374 38546 15426 38558
rect 17614 38610 17666 38622
rect 23886 38610 23938 38622
rect 20626 38558 20638 38610
rect 20690 38558 20702 38610
rect 17614 38546 17666 38558
rect 23886 38546 23938 38558
rect 41806 38610 41858 38622
rect 44146 38558 44158 38610
rect 44210 38558 44222 38610
rect 52434 38558 52446 38610
rect 52498 38558 52510 38610
rect 54002 38558 54014 38610
rect 54066 38607 54078 38610
rect 54450 38607 54462 38610
rect 54066 38561 54462 38607
rect 54066 38558 54078 38561
rect 54450 38558 54462 38561
rect 54514 38607 54526 38610
rect 55010 38607 55022 38610
rect 54514 38561 55022 38607
rect 54514 38558 54526 38561
rect 55010 38558 55022 38561
rect 55074 38558 55086 38610
rect 41806 38546 41858 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 4062 38274 4114 38286
rect 4062 38210 4114 38222
rect 20526 38274 20578 38286
rect 20526 38210 20578 38222
rect 20638 38274 20690 38286
rect 20638 38210 20690 38222
rect 36318 38274 36370 38286
rect 36318 38210 36370 38222
rect 37326 38274 37378 38286
rect 37326 38210 37378 38222
rect 37662 38274 37714 38286
rect 37662 38210 37714 38222
rect 38110 38274 38162 38286
rect 39554 38222 39566 38274
rect 39618 38222 39630 38274
rect 38110 38210 38162 38222
rect 14142 38162 14194 38174
rect 28478 38162 28530 38174
rect 43934 38162 43986 38174
rect 48414 38162 48466 38174
rect 53342 38162 53394 38174
rect 15698 38110 15710 38162
rect 15762 38110 15774 38162
rect 19618 38110 19630 38162
rect 19682 38110 19694 38162
rect 34738 38110 34750 38162
rect 34802 38110 34814 38162
rect 40562 38110 40574 38162
rect 40626 38110 40638 38162
rect 42690 38110 42702 38162
rect 42754 38110 42766 38162
rect 45938 38110 45950 38162
rect 46002 38110 46014 38162
rect 51314 38110 51326 38162
rect 51378 38110 51390 38162
rect 56802 38110 56814 38162
rect 56866 38110 56878 38162
rect 14142 38098 14194 38110
rect 28478 38098 28530 38110
rect 43934 38098 43986 38110
rect 48414 38098 48466 38110
rect 53342 38098 53394 38110
rect 7646 38050 7698 38062
rect 4834 37998 4846 38050
rect 4898 37998 4910 38050
rect 5842 37998 5854 38050
rect 5906 37998 5918 38050
rect 7646 37986 7698 37998
rect 10222 38050 10274 38062
rect 10222 37986 10274 37998
rect 10558 38050 10610 38062
rect 12686 38050 12738 38062
rect 14030 38050 14082 38062
rect 11106 37998 11118 38050
rect 11170 37998 11182 38050
rect 11554 37998 11566 38050
rect 11618 37998 11630 38050
rect 13794 37998 13806 38050
rect 13858 37998 13870 38050
rect 10558 37986 10610 37998
rect 12686 37986 12738 37998
rect 14030 37986 14082 37998
rect 14366 38050 14418 38062
rect 19742 38050 19794 38062
rect 15810 37998 15822 38050
rect 15874 37998 15886 38050
rect 17490 37998 17502 38050
rect 17554 37998 17566 38050
rect 18834 37998 18846 38050
rect 18898 37998 18910 38050
rect 14366 37986 14418 37998
rect 19742 37986 19794 37998
rect 24558 38050 24610 38062
rect 24558 37986 24610 37998
rect 24894 38050 24946 38062
rect 24894 37986 24946 37998
rect 25230 38050 25282 38062
rect 26238 38050 26290 38062
rect 35422 38050 35474 38062
rect 25666 37998 25678 38050
rect 25730 37998 25742 38050
rect 29138 37998 29150 38050
rect 29202 37998 29214 38050
rect 30034 37998 30046 38050
rect 30098 37998 30110 38050
rect 31266 37998 31278 38050
rect 31330 37998 31342 38050
rect 31938 37998 31950 38050
rect 32002 37998 32014 38050
rect 25230 37986 25282 37998
rect 26238 37986 26290 37998
rect 35422 37986 35474 37998
rect 36206 38050 36258 38062
rect 37886 38050 37938 38062
rect 45502 38050 45554 38062
rect 37650 37998 37662 38050
rect 37714 37998 37726 38050
rect 38770 37998 38782 38050
rect 38834 37998 38846 38050
rect 43474 37998 43486 38050
rect 43538 37998 43550 38050
rect 45042 37998 45054 38050
rect 45106 37998 45118 38050
rect 36206 37986 36258 37998
rect 37886 37986 37938 37998
rect 45502 37986 45554 37998
rect 49870 38050 49922 38062
rect 53118 38050 53170 38062
rect 51426 37998 51438 38050
rect 51490 37998 51502 38050
rect 51650 37998 51662 38050
rect 51714 37998 51726 38050
rect 49870 37986 49922 37998
rect 53118 37986 53170 37998
rect 53566 38050 53618 38062
rect 57374 38050 57426 38062
rect 54002 37998 54014 38050
rect 54066 37998 54078 38050
rect 53566 37986 53618 37998
rect 57374 37986 57426 37998
rect 3502 37938 3554 37950
rect 3502 37874 3554 37886
rect 3950 37938 4002 37950
rect 3950 37874 4002 37886
rect 6862 37938 6914 37950
rect 6862 37874 6914 37886
rect 10446 37938 10498 37950
rect 10446 37874 10498 37886
rect 11678 37938 11730 37950
rect 11678 37874 11730 37886
rect 12798 37938 12850 37950
rect 22206 37938 22258 37950
rect 23662 37938 23714 37950
rect 16034 37886 16046 37938
rect 16098 37886 16110 37938
rect 19954 37886 19966 37938
rect 20018 37886 20030 37938
rect 22530 37886 22542 37938
rect 22594 37886 22606 37938
rect 12798 37874 12850 37886
rect 22206 37874 22258 37886
rect 23662 37874 23714 37886
rect 23998 37938 24050 37950
rect 23998 37874 24050 37886
rect 24222 37938 24274 37950
rect 24222 37874 24274 37886
rect 27694 37938 27746 37950
rect 27694 37874 27746 37886
rect 27806 37938 27858 37950
rect 27806 37874 27858 37886
rect 28366 37938 28418 37950
rect 39790 37938 39842 37950
rect 50206 37938 50258 37950
rect 29250 37886 29262 37938
rect 29314 37886 29326 37938
rect 31490 37886 31502 37938
rect 31554 37886 31566 37938
rect 32610 37886 32622 37938
rect 32674 37886 32686 37938
rect 44818 37886 44830 37938
rect 44882 37886 44894 37938
rect 46722 37886 46734 37938
rect 46786 37886 46798 37938
rect 28366 37874 28418 37886
rect 39790 37874 39842 37886
rect 50206 37874 50258 37886
rect 50318 37938 50370 37950
rect 50318 37874 50370 37886
rect 50542 37938 50594 37950
rect 50542 37874 50594 37886
rect 52670 37938 52722 37950
rect 52882 37886 52894 37938
rect 52946 37886 52958 37938
rect 54674 37886 54686 37938
rect 54738 37886 54750 37938
rect 52670 37874 52722 37886
rect 3726 37826 3778 37838
rect 3726 37762 3778 37774
rect 4510 37826 4562 37838
rect 4510 37762 4562 37774
rect 5070 37826 5122 37838
rect 5070 37762 5122 37774
rect 8206 37826 8258 37838
rect 8206 37762 8258 37774
rect 9214 37826 9266 37838
rect 9214 37762 9266 37774
rect 13022 37826 13074 37838
rect 13022 37762 13074 37774
rect 14254 37826 14306 37838
rect 14254 37762 14306 37774
rect 14926 37826 14978 37838
rect 20190 37826 20242 37838
rect 15250 37774 15262 37826
rect 15314 37774 15326 37826
rect 14926 37762 14978 37774
rect 20190 37762 20242 37774
rect 21310 37826 21362 37838
rect 23886 37826 23938 37838
rect 21634 37774 21646 37826
rect 21698 37774 21710 37826
rect 21310 37762 21362 37774
rect 23886 37762 23938 37774
rect 24894 37826 24946 37838
rect 26350 37826 26402 37838
rect 25890 37774 25902 37826
rect 25954 37774 25966 37826
rect 24894 37762 24946 37774
rect 26350 37762 26402 37774
rect 26574 37826 26626 37838
rect 26574 37762 26626 37774
rect 27470 37826 27522 37838
rect 35870 37826 35922 37838
rect 30034 37774 30046 37826
rect 30098 37774 30110 37826
rect 35074 37774 35086 37826
rect 35138 37774 35150 37826
rect 27470 37762 27522 37774
rect 35870 37762 35922 37774
rect 36318 37826 36370 37838
rect 36318 37762 36370 37774
rect 43822 37826 43874 37838
rect 43822 37762 43874 37774
rect 46398 37826 46450 37838
rect 53678 37826 53730 37838
rect 51986 37774 51998 37826
rect 52050 37774 52062 37826
rect 46398 37762 46450 37774
rect 53678 37762 53730 37774
rect 57038 37826 57090 37838
rect 57038 37762 57090 37774
rect 57262 37826 57314 37838
rect 57262 37762 57314 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 2382 37490 2434 37502
rect 2382 37426 2434 37438
rect 9550 37490 9602 37502
rect 17726 37490 17778 37502
rect 17378 37438 17390 37490
rect 17442 37438 17454 37490
rect 9550 37426 9602 37438
rect 17726 37426 17778 37438
rect 23102 37490 23154 37502
rect 23102 37426 23154 37438
rect 28254 37490 28306 37502
rect 28254 37426 28306 37438
rect 35982 37490 36034 37502
rect 35982 37426 36034 37438
rect 40126 37490 40178 37502
rect 40126 37426 40178 37438
rect 44606 37490 44658 37502
rect 44606 37426 44658 37438
rect 45502 37490 45554 37502
rect 45502 37426 45554 37438
rect 48862 37490 48914 37502
rect 55694 37490 55746 37502
rect 51090 37438 51102 37490
rect 51154 37438 51166 37490
rect 48862 37426 48914 37438
rect 55694 37426 55746 37438
rect 55806 37490 55858 37502
rect 55806 37426 55858 37438
rect 4510 37378 4562 37390
rect 7758 37378 7810 37390
rect 22542 37378 22594 37390
rect 2706 37326 2718 37378
rect 2770 37326 2782 37378
rect 5282 37326 5294 37378
rect 5346 37326 5358 37378
rect 12338 37326 12350 37378
rect 12402 37326 12414 37378
rect 13570 37326 13582 37378
rect 13634 37326 13646 37378
rect 18274 37326 18286 37378
rect 18338 37326 18350 37378
rect 20514 37326 20526 37378
rect 20578 37326 20590 37378
rect 4510 37314 4562 37326
rect 7758 37314 7810 37326
rect 22542 37314 22594 37326
rect 23326 37378 23378 37390
rect 23326 37314 23378 37326
rect 27582 37378 27634 37390
rect 27582 37314 27634 37326
rect 34750 37378 34802 37390
rect 34750 37314 34802 37326
rect 34974 37378 35026 37390
rect 34974 37314 35026 37326
rect 36430 37378 36482 37390
rect 36430 37314 36482 37326
rect 42702 37378 42754 37390
rect 52222 37378 52274 37390
rect 46386 37326 46398 37378
rect 46450 37326 46462 37378
rect 49746 37326 49758 37378
rect 49810 37326 49822 37378
rect 42702 37314 42754 37326
rect 52222 37314 52274 37326
rect 54126 37378 54178 37390
rect 54126 37314 54178 37326
rect 54910 37378 54962 37390
rect 54910 37314 54962 37326
rect 55582 37378 55634 37390
rect 55582 37314 55634 37326
rect 3054 37266 3106 37278
rect 2146 37214 2158 37266
rect 2210 37214 2222 37266
rect 3054 37202 3106 37214
rect 3502 37266 3554 37278
rect 3502 37202 3554 37214
rect 4622 37266 4674 37278
rect 8878 37266 8930 37278
rect 11230 37266 11282 37278
rect 14926 37266 14978 37278
rect 19854 37266 19906 37278
rect 21982 37266 22034 37278
rect 5170 37214 5182 37266
rect 5234 37214 5246 37266
rect 10882 37214 10894 37266
rect 10946 37214 10958 37266
rect 11778 37214 11790 37266
rect 11842 37214 11854 37266
rect 15922 37214 15934 37266
rect 15986 37214 15998 37266
rect 16706 37214 16718 37266
rect 16770 37214 16782 37266
rect 18498 37214 18510 37266
rect 18562 37214 18574 37266
rect 20290 37214 20302 37266
rect 20354 37214 20366 37266
rect 21298 37214 21310 37266
rect 21362 37214 21374 37266
rect 21522 37214 21534 37266
rect 21586 37214 21598 37266
rect 4622 37202 4674 37214
rect 8878 37202 8930 37214
rect 11230 37202 11282 37214
rect 14926 37202 14978 37214
rect 19854 37202 19906 37214
rect 21982 37202 22034 37214
rect 22206 37266 22258 37278
rect 22206 37202 22258 37214
rect 22766 37266 22818 37278
rect 27358 37266 27410 37278
rect 25778 37214 25790 37266
rect 25842 37214 25854 37266
rect 26450 37214 26462 37266
rect 26514 37214 26526 37266
rect 22766 37202 22818 37214
rect 27358 37202 27410 37214
rect 27694 37266 27746 37278
rect 27694 37202 27746 37214
rect 28478 37266 28530 37278
rect 28478 37202 28530 37214
rect 28926 37266 28978 37278
rect 35534 37266 35586 37278
rect 31826 37214 31838 37266
rect 31890 37214 31902 37266
rect 28926 37202 28978 37214
rect 35534 37202 35586 37214
rect 36654 37266 36706 37278
rect 36654 37202 36706 37214
rect 37438 37266 37490 37278
rect 38782 37266 38834 37278
rect 37762 37214 37774 37266
rect 37826 37214 37838 37266
rect 37438 37202 37490 37214
rect 38782 37202 38834 37214
rect 39454 37266 39506 37278
rect 39454 37202 39506 37214
rect 42366 37266 42418 37278
rect 42366 37202 42418 37214
rect 42590 37266 42642 37278
rect 42590 37202 42642 37214
rect 45166 37266 45218 37278
rect 45166 37202 45218 37214
rect 46062 37266 46114 37278
rect 46062 37202 46114 37214
rect 46734 37266 46786 37278
rect 46734 37202 46786 37214
rect 51326 37266 51378 37278
rect 54238 37266 54290 37278
rect 53442 37214 53454 37266
rect 53506 37214 53518 37266
rect 53778 37214 53790 37266
rect 53842 37214 53854 37266
rect 51326 37202 51378 37214
rect 54238 37202 54290 37214
rect 54350 37266 54402 37278
rect 54350 37202 54402 37214
rect 54686 37266 54738 37278
rect 54686 37202 54738 37214
rect 55246 37266 55298 37278
rect 55246 37202 55298 37214
rect 57262 37266 57314 37278
rect 57262 37202 57314 37214
rect 3614 37154 3666 37166
rect 9662 37154 9714 37166
rect 15710 37154 15762 37166
rect 8306 37102 8318 37154
rect 8370 37102 8382 37154
rect 10322 37102 10334 37154
rect 10386 37102 10398 37154
rect 15026 37102 15038 37154
rect 15090 37102 15102 37154
rect 3614 37090 3666 37102
rect 9662 37090 9714 37102
rect 15710 37090 15762 37102
rect 16270 37154 16322 37166
rect 22430 37154 22482 37166
rect 28366 37154 28418 37166
rect 39230 37154 39282 37166
rect 20178 37102 20190 37154
rect 20242 37102 20254 37154
rect 26338 37102 26350 37154
rect 26402 37102 26414 37154
rect 31490 37102 31502 37154
rect 31554 37102 31566 37154
rect 16270 37090 16322 37102
rect 22430 37090 22482 37102
rect 28366 37090 28418 37102
rect 39230 37090 39282 37102
rect 43710 37154 43762 37166
rect 43710 37090 43762 37102
rect 47406 37154 47458 37166
rect 47406 37090 47458 37102
rect 55134 37154 55186 37166
rect 57598 37154 57650 37166
rect 57138 37102 57150 37154
rect 57202 37102 57214 37154
rect 55134 37090 55186 37102
rect 57598 37090 57650 37102
rect 3838 37042 3890 37054
rect 3838 36978 3890 36990
rect 3950 37042 4002 37054
rect 3950 36978 4002 36990
rect 4734 37042 4786 37054
rect 15598 37042 15650 37054
rect 11330 36990 11342 37042
rect 11394 36990 11406 37042
rect 4734 36978 4786 36990
rect 15598 36978 15650 36990
rect 22990 37042 23042 37054
rect 35086 37042 35138 37054
rect 26786 36990 26798 37042
rect 26850 36990 26862 37042
rect 22990 36978 23042 36990
rect 35086 36978 35138 36990
rect 36990 37042 37042 37054
rect 36990 36978 37042 36990
rect 39678 37042 39730 37054
rect 39678 36978 39730 36990
rect 42030 37042 42082 37054
rect 42030 36978 42082 36990
rect 42142 37042 42194 37054
rect 42142 36978 42194 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 5070 36706 5122 36718
rect 5070 36642 5122 36654
rect 7646 36706 7698 36718
rect 7646 36642 7698 36654
rect 7982 36706 8034 36718
rect 7982 36642 8034 36654
rect 8318 36706 8370 36718
rect 8318 36642 8370 36654
rect 10222 36706 10274 36718
rect 10222 36642 10274 36654
rect 14478 36706 14530 36718
rect 14478 36642 14530 36654
rect 15486 36706 15538 36718
rect 15486 36642 15538 36654
rect 36318 36706 36370 36718
rect 51314 36654 51326 36706
rect 51378 36654 51390 36706
rect 36318 36642 36370 36654
rect 21422 36594 21474 36606
rect 29262 36594 29314 36606
rect 2482 36542 2494 36594
rect 2546 36542 2558 36594
rect 4610 36542 4622 36594
rect 4674 36542 4686 36594
rect 11554 36542 11566 36594
rect 11618 36542 11630 36594
rect 28578 36542 28590 36594
rect 28642 36542 28654 36594
rect 21422 36530 21474 36542
rect 29262 36530 29314 36542
rect 30158 36594 30210 36606
rect 44158 36594 44210 36606
rect 34514 36542 34526 36594
rect 34578 36542 34590 36594
rect 49522 36542 49534 36594
rect 49586 36542 49598 36594
rect 56130 36542 56142 36594
rect 56194 36542 56206 36594
rect 30158 36530 30210 36542
rect 44158 36530 44210 36542
rect 6190 36482 6242 36494
rect 10110 36482 10162 36494
rect 14030 36482 14082 36494
rect 1810 36430 1822 36482
rect 1874 36430 1886 36482
rect 8642 36430 8654 36482
rect 8706 36430 8718 36482
rect 9426 36430 9438 36482
rect 9490 36430 9502 36482
rect 10658 36430 10670 36482
rect 10722 36430 10734 36482
rect 6190 36418 6242 36430
rect 10110 36418 10162 36430
rect 14030 36418 14082 36430
rect 14142 36482 14194 36494
rect 15374 36482 15426 36494
rect 20414 36482 20466 36494
rect 14802 36430 14814 36482
rect 14866 36430 14878 36482
rect 16034 36430 16046 36482
rect 16098 36430 16110 36482
rect 17602 36430 17614 36482
rect 17666 36430 17678 36482
rect 19618 36430 19630 36482
rect 19682 36430 19694 36482
rect 14142 36418 14194 36430
rect 15374 36418 15426 36430
rect 20414 36418 20466 36430
rect 20750 36482 20802 36494
rect 20750 36418 20802 36430
rect 21534 36482 21586 36494
rect 21534 36418 21586 36430
rect 21982 36482 22034 36494
rect 21982 36418 22034 36430
rect 22990 36482 23042 36494
rect 22990 36418 23042 36430
rect 23438 36482 23490 36494
rect 23438 36418 23490 36430
rect 24110 36482 24162 36494
rect 24110 36418 24162 36430
rect 24334 36482 24386 36494
rect 26910 36482 26962 36494
rect 29598 36482 29650 36494
rect 26226 36430 26238 36482
rect 26290 36430 26302 36482
rect 26450 36430 26462 36482
rect 26514 36430 26526 36482
rect 28466 36430 28478 36482
rect 28530 36430 28542 36482
rect 24334 36418 24386 36430
rect 26910 36418 26962 36430
rect 29598 36418 29650 36430
rect 29822 36482 29874 36494
rect 29822 36418 29874 36430
rect 30046 36482 30098 36494
rect 35534 36482 35586 36494
rect 37998 36482 38050 36494
rect 31714 36430 31726 36482
rect 31778 36430 31790 36482
rect 35970 36430 35982 36482
rect 36034 36430 36046 36482
rect 30046 36418 30098 36430
rect 35534 36418 35586 36430
rect 37998 36418 38050 36430
rect 38446 36482 38498 36494
rect 38446 36418 38498 36430
rect 39566 36482 39618 36494
rect 39566 36418 39618 36430
rect 43374 36482 43426 36494
rect 43374 36418 43426 36430
rect 43822 36482 43874 36494
rect 46846 36482 46898 36494
rect 44930 36430 44942 36482
rect 44994 36430 45006 36482
rect 46274 36430 46286 36482
rect 46338 36430 46350 36482
rect 43822 36418 43874 36430
rect 46846 36418 46898 36430
rect 47406 36482 47458 36494
rect 47406 36418 47458 36430
rect 47966 36482 48018 36494
rect 47966 36418 48018 36430
rect 48190 36482 48242 36494
rect 48190 36418 48242 36430
rect 48526 36482 48578 36494
rect 48526 36418 48578 36430
rect 48750 36482 48802 36494
rect 50094 36482 50146 36494
rect 53006 36482 53058 36494
rect 53454 36482 53506 36494
rect 49634 36430 49646 36482
rect 49698 36430 49710 36482
rect 50866 36430 50878 36482
rect 50930 36430 50942 36482
rect 51426 36430 51438 36482
rect 51490 36430 51502 36482
rect 52210 36430 52222 36482
rect 52274 36430 52286 36482
rect 52658 36430 52670 36482
rect 52722 36430 52734 36482
rect 53218 36430 53230 36482
rect 53282 36430 53294 36482
rect 48750 36418 48802 36430
rect 50094 36418 50146 36430
rect 53006 36418 53058 36430
rect 53454 36418 53506 36430
rect 54350 36482 54402 36494
rect 54898 36430 54910 36482
rect 54962 36430 54974 36482
rect 56578 36430 56590 36482
rect 56642 36430 56654 36482
rect 57026 36430 57038 36482
rect 57090 36430 57102 36482
rect 57586 36430 57598 36482
rect 57650 36430 57662 36482
rect 54350 36418 54402 36430
rect 4958 36370 5010 36382
rect 4958 36306 5010 36318
rect 5966 36370 6018 36382
rect 5966 36306 6018 36318
rect 6414 36370 6466 36382
rect 6414 36306 6466 36318
rect 7534 36370 7586 36382
rect 12686 36370 12738 36382
rect 9874 36318 9886 36370
rect 9938 36318 9950 36370
rect 10546 36318 10558 36370
rect 10610 36318 10622 36370
rect 7534 36306 7586 36318
rect 12686 36306 12738 36318
rect 12798 36370 12850 36382
rect 12798 36306 12850 36318
rect 13918 36370 13970 36382
rect 13918 36306 13970 36318
rect 15038 36370 15090 36382
rect 20638 36370 20690 36382
rect 16706 36318 16718 36370
rect 16770 36318 16782 36370
rect 19954 36318 19966 36370
rect 20018 36318 20030 36370
rect 15038 36306 15090 36318
rect 20638 36306 20690 36318
rect 22654 36370 22706 36382
rect 22654 36306 22706 36318
rect 22766 36370 22818 36382
rect 22766 36306 22818 36318
rect 24558 36370 24610 36382
rect 24558 36306 24610 36318
rect 26798 36370 26850 36382
rect 26798 36306 26850 36318
rect 28142 36370 28194 36382
rect 35758 36370 35810 36382
rect 32386 36318 32398 36370
rect 32450 36318 32462 36370
rect 28142 36306 28194 36318
rect 35758 36306 35810 36318
rect 38894 36370 38946 36382
rect 38894 36306 38946 36318
rect 39118 36370 39170 36382
rect 39118 36306 39170 36318
rect 43150 36370 43202 36382
rect 43150 36306 43202 36318
rect 45166 36370 45218 36382
rect 46510 36370 46562 36382
rect 45490 36318 45502 36370
rect 45554 36318 45566 36370
rect 45166 36306 45218 36318
rect 46510 36306 46562 36318
rect 50430 36370 50482 36382
rect 53778 36318 53790 36370
rect 53842 36318 53854 36370
rect 55346 36318 55358 36370
rect 55410 36318 55422 36370
rect 50430 36306 50482 36318
rect 8206 36258 8258 36270
rect 6738 36206 6750 36258
rect 6802 36206 6814 36258
rect 8206 36194 8258 36206
rect 13022 36258 13074 36270
rect 14590 36258 14642 36270
rect 21310 36258 21362 36270
rect 13458 36206 13470 36258
rect 13522 36206 13534 36258
rect 16034 36206 16046 36258
rect 16098 36206 16110 36258
rect 13022 36194 13074 36206
rect 14590 36194 14642 36206
rect 21310 36194 21362 36206
rect 23550 36258 23602 36270
rect 23550 36194 23602 36206
rect 23662 36258 23714 36270
rect 23662 36194 23714 36206
rect 24446 36258 24498 36270
rect 24446 36194 24498 36206
rect 26686 36258 26738 36270
rect 26686 36194 26738 36206
rect 27806 36258 27858 36270
rect 27806 36194 27858 36206
rect 28030 36258 28082 36270
rect 28030 36194 28082 36206
rect 29150 36258 29202 36270
rect 29150 36194 29202 36206
rect 30270 36258 30322 36270
rect 30270 36194 30322 36206
rect 34862 36258 34914 36270
rect 34862 36194 34914 36206
rect 34974 36258 35026 36270
rect 34974 36194 35026 36206
rect 35086 36258 35138 36270
rect 35086 36194 35138 36206
rect 36206 36258 36258 36270
rect 36206 36194 36258 36206
rect 38110 36258 38162 36270
rect 38110 36194 38162 36206
rect 38222 36258 38274 36270
rect 38222 36194 38274 36206
rect 38334 36258 38386 36270
rect 38334 36194 38386 36206
rect 39230 36258 39282 36270
rect 39230 36194 39282 36206
rect 43598 36258 43650 36270
rect 43598 36194 43650 36206
rect 45838 36258 45890 36270
rect 45838 36194 45890 36206
rect 48302 36258 48354 36270
rect 48302 36194 48354 36206
rect 50318 36258 50370 36270
rect 50318 36194 50370 36206
rect 52670 36258 52722 36270
rect 54002 36206 54014 36258
rect 54066 36206 54078 36258
rect 52670 36194 52722 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 15374 35922 15426 35934
rect 19518 35922 19570 35934
rect 5282 35870 5294 35922
rect 5346 35870 5358 35922
rect 11218 35870 11230 35922
rect 11282 35870 11294 35922
rect 17938 35870 17950 35922
rect 18002 35870 18014 35922
rect 18722 35870 18734 35922
rect 18786 35870 18798 35922
rect 15374 35858 15426 35870
rect 19518 35858 19570 35870
rect 22542 35922 22594 35934
rect 22542 35858 22594 35870
rect 23998 35922 24050 35934
rect 32398 35922 32450 35934
rect 31378 35870 31390 35922
rect 31442 35870 31454 35922
rect 23998 35858 24050 35870
rect 32398 35858 32450 35870
rect 33630 35922 33682 35934
rect 33630 35858 33682 35870
rect 34078 35922 34130 35934
rect 37998 35922 38050 35934
rect 35746 35870 35758 35922
rect 35810 35870 35822 35922
rect 34078 35858 34130 35870
rect 37998 35858 38050 35870
rect 40910 35922 40962 35934
rect 40910 35858 40962 35870
rect 44270 35922 44322 35934
rect 44270 35858 44322 35870
rect 44382 35922 44434 35934
rect 44382 35858 44434 35870
rect 45390 35922 45442 35934
rect 45390 35858 45442 35870
rect 46286 35922 46338 35934
rect 46286 35858 46338 35870
rect 47182 35922 47234 35934
rect 47182 35858 47234 35870
rect 47742 35922 47794 35934
rect 47742 35858 47794 35870
rect 48078 35922 48130 35934
rect 48078 35858 48130 35870
rect 48190 35922 48242 35934
rect 48190 35858 48242 35870
rect 51550 35922 51602 35934
rect 51550 35858 51602 35870
rect 54910 35922 54962 35934
rect 54910 35858 54962 35870
rect 7870 35810 7922 35822
rect 14702 35810 14754 35822
rect 12114 35758 12126 35810
rect 12178 35758 12190 35810
rect 7870 35746 7922 35758
rect 14702 35746 14754 35758
rect 14814 35810 14866 35822
rect 14814 35746 14866 35758
rect 16718 35810 16770 35822
rect 16718 35746 16770 35758
rect 16830 35810 16882 35822
rect 16830 35746 16882 35758
rect 18286 35810 18338 35822
rect 33854 35810 33906 35822
rect 41134 35810 41186 35822
rect 26786 35758 26798 35810
rect 26850 35758 26862 35810
rect 27794 35758 27806 35810
rect 27858 35758 27870 35810
rect 35298 35758 35310 35810
rect 35362 35758 35374 35810
rect 36866 35758 36878 35810
rect 36930 35758 36942 35810
rect 40114 35758 40126 35810
rect 40178 35758 40190 35810
rect 18286 35746 18338 35758
rect 33854 35746 33906 35758
rect 41134 35746 41186 35758
rect 41246 35810 41298 35822
rect 41246 35746 41298 35758
rect 41582 35810 41634 35822
rect 41582 35746 41634 35758
rect 43934 35810 43986 35822
rect 43934 35746 43986 35758
rect 44494 35810 44546 35822
rect 44494 35746 44546 35758
rect 44718 35810 44770 35822
rect 44718 35746 44770 35758
rect 49870 35810 49922 35822
rect 49870 35746 49922 35758
rect 51438 35810 51490 35822
rect 51438 35746 51490 35758
rect 53230 35810 53282 35822
rect 53230 35746 53282 35758
rect 56590 35810 56642 35822
rect 56590 35746 56642 35758
rect 3054 35698 3106 35710
rect 2706 35646 2718 35698
rect 2770 35646 2782 35698
rect 3054 35634 3106 35646
rect 4398 35698 4450 35710
rect 4398 35634 4450 35646
rect 4734 35698 4786 35710
rect 4734 35634 4786 35646
rect 4958 35698 5010 35710
rect 7982 35698 8034 35710
rect 10670 35698 10722 35710
rect 6066 35646 6078 35698
rect 6130 35646 6142 35698
rect 8194 35646 8206 35698
rect 8258 35646 8270 35698
rect 4958 35634 5010 35646
rect 7982 35634 8034 35646
rect 10670 35634 10722 35646
rect 10894 35698 10946 35710
rect 15038 35698 15090 35710
rect 11778 35646 11790 35698
rect 11842 35646 11854 35698
rect 13458 35646 13470 35698
rect 13522 35646 13534 35698
rect 10894 35634 10946 35646
rect 15038 35634 15090 35646
rect 15598 35698 15650 35710
rect 15598 35634 15650 35646
rect 16494 35698 16546 35710
rect 28254 35698 28306 35710
rect 29822 35698 29874 35710
rect 37886 35698 37938 35710
rect 18946 35646 18958 35698
rect 19010 35646 19022 35698
rect 23538 35646 23550 35698
rect 23602 35646 23614 35698
rect 23762 35646 23774 35698
rect 23826 35646 23838 35698
rect 25666 35646 25678 35698
rect 25730 35646 25742 35698
rect 26674 35646 26686 35698
rect 26738 35646 26750 35698
rect 27682 35646 27694 35698
rect 27746 35646 27758 35698
rect 28578 35646 28590 35698
rect 28642 35646 28654 35698
rect 29474 35646 29486 35698
rect 29538 35646 29550 35698
rect 29922 35646 29934 35698
rect 29986 35646 29998 35698
rect 31154 35646 31166 35698
rect 31218 35646 31230 35698
rect 32162 35646 32174 35698
rect 32226 35646 32238 35698
rect 35186 35646 35198 35698
rect 35250 35646 35262 35698
rect 36194 35646 36206 35698
rect 36258 35646 36270 35698
rect 16494 35634 16546 35646
rect 28254 35634 28306 35646
rect 29822 35634 29874 35646
rect 37886 35634 37938 35646
rect 38334 35698 38386 35710
rect 38334 35634 38386 35646
rect 38894 35698 38946 35710
rect 42478 35698 42530 35710
rect 39218 35646 39230 35698
rect 39282 35646 39294 35698
rect 42018 35646 42030 35698
rect 42082 35646 42094 35698
rect 38894 35634 38946 35646
rect 42478 35634 42530 35646
rect 43038 35698 43090 35710
rect 45726 35698 45778 35710
rect 43250 35646 43262 35698
rect 43314 35646 43326 35698
rect 43038 35634 43090 35646
rect 45726 35634 45778 35646
rect 47966 35698 48018 35710
rect 52110 35698 52162 35710
rect 49186 35646 49198 35698
rect 49250 35646 49262 35698
rect 47966 35634 48018 35646
rect 52110 35634 52162 35646
rect 52222 35698 52274 35710
rect 52222 35634 52274 35646
rect 53342 35698 53394 35710
rect 53342 35634 53394 35646
rect 53566 35698 53618 35710
rect 54238 35698 54290 35710
rect 53778 35646 53790 35698
rect 53842 35646 53854 35698
rect 53566 35634 53618 35646
rect 54238 35634 54290 35646
rect 54686 35698 54738 35710
rect 54686 35634 54738 35646
rect 55582 35698 55634 35710
rect 55582 35634 55634 35646
rect 55806 35698 55858 35710
rect 57486 35698 57538 35710
rect 56018 35646 56030 35698
rect 56082 35646 56094 35698
rect 57026 35646 57038 35698
rect 57090 35646 57102 35698
rect 55806 35634 55858 35646
rect 57486 35634 57538 35646
rect 57934 35698 57986 35710
rect 57934 35634 57986 35646
rect 8654 35586 8706 35598
rect 15822 35586 15874 35598
rect 3938 35534 3950 35586
rect 4002 35534 4014 35586
rect 5730 35534 5742 35586
rect 5794 35534 5806 35586
rect 13906 35534 13918 35586
rect 13970 35534 13982 35586
rect 15474 35534 15486 35586
rect 15538 35534 15550 35586
rect 8654 35522 8706 35534
rect 15822 35522 15874 35534
rect 16270 35586 16322 35598
rect 16270 35522 16322 35534
rect 17390 35586 17442 35598
rect 17390 35522 17442 35534
rect 18398 35586 18450 35598
rect 18398 35522 18450 35534
rect 21198 35586 21250 35598
rect 21198 35522 21250 35534
rect 21646 35586 21698 35598
rect 33742 35586 33794 35598
rect 22642 35534 22654 35586
rect 22706 35534 22718 35586
rect 27458 35534 27470 35586
rect 27522 35534 27534 35586
rect 21646 35522 21698 35534
rect 33742 35522 33794 35534
rect 34638 35586 34690 35598
rect 50990 35586 51042 35598
rect 49522 35534 49534 35586
rect 49586 35534 49598 35586
rect 34638 35522 34690 35534
rect 50990 35522 51042 35534
rect 51662 35586 51714 35598
rect 51662 35522 51714 35534
rect 54798 35586 54850 35598
rect 54798 35522 54850 35534
rect 58046 35586 58098 35598
rect 58046 35522 58098 35534
rect 16046 35474 16098 35486
rect 3154 35422 3166 35474
rect 3218 35422 3230 35474
rect 7410 35422 7422 35474
rect 7474 35422 7486 35474
rect 16046 35410 16098 35422
rect 17614 35474 17666 35486
rect 17614 35410 17666 35422
rect 22318 35474 22370 35486
rect 22318 35410 22370 35422
rect 24110 35474 24162 35486
rect 32510 35474 32562 35486
rect 30370 35422 30382 35474
rect 30434 35422 30446 35474
rect 24110 35410 24162 35422
rect 32510 35410 32562 35422
rect 37998 35474 38050 35486
rect 37998 35410 38050 35422
rect 38558 35474 38610 35486
rect 38558 35410 38610 35422
rect 52446 35474 52498 35486
rect 52446 35410 52498 35422
rect 52558 35474 52610 35486
rect 55470 35474 55522 35486
rect 53778 35422 53790 35474
rect 53842 35422 53854 35474
rect 52558 35410 52610 35422
rect 55470 35410 55522 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 3166 35138 3218 35150
rect 3166 35074 3218 35086
rect 8206 35138 8258 35150
rect 8206 35074 8258 35086
rect 10110 35138 10162 35150
rect 10110 35074 10162 35086
rect 12798 35138 12850 35150
rect 12798 35074 12850 35086
rect 13582 35138 13634 35150
rect 13582 35074 13634 35086
rect 13806 35138 13858 35150
rect 13806 35074 13858 35086
rect 18958 35138 19010 35150
rect 18958 35074 19010 35086
rect 19294 35138 19346 35150
rect 19294 35074 19346 35086
rect 23662 35138 23714 35150
rect 23662 35074 23714 35086
rect 30270 35138 30322 35150
rect 53006 35138 53058 35150
rect 52658 35086 52670 35138
rect 52722 35086 52734 35138
rect 30270 35074 30322 35086
rect 53006 35074 53058 35086
rect 53902 35138 53954 35150
rect 53902 35074 53954 35086
rect 4846 35026 4898 35038
rect 32398 35026 32450 35038
rect 2818 34974 2830 35026
rect 2882 34974 2894 35026
rect 18050 34974 18062 35026
rect 18114 34974 18126 35026
rect 19842 34974 19854 35026
rect 19906 34974 19918 35026
rect 22194 34974 22206 35026
rect 22258 34974 22270 35026
rect 30594 34974 30606 35026
rect 30658 34974 30670 35026
rect 4846 34962 4898 34974
rect 32398 34962 32450 34974
rect 34414 35026 34466 35038
rect 38782 35026 38834 35038
rect 43934 35026 43986 35038
rect 51774 35026 51826 35038
rect 35186 34974 35198 35026
rect 35250 34974 35262 35026
rect 36418 34974 36430 35026
rect 36482 34974 36494 35026
rect 39666 34974 39678 35026
rect 39730 34974 39742 35026
rect 41346 34974 41358 35026
rect 41410 34974 41422 35026
rect 47842 34974 47854 35026
rect 47906 34974 47918 35026
rect 49970 34974 49982 35026
rect 50034 34974 50046 35026
rect 34414 34962 34466 34974
rect 38782 34962 38834 34974
rect 43934 34962 43986 34974
rect 51774 34962 51826 34974
rect 52110 35026 52162 35038
rect 55122 34974 55134 35026
rect 55186 34974 55198 35026
rect 57250 34974 57262 35026
rect 57314 34974 57326 35026
rect 52110 34962 52162 34974
rect 7198 34914 7250 34926
rect 6738 34862 6750 34914
rect 6802 34862 6814 34914
rect 7198 34850 7250 34862
rect 7646 34914 7698 34926
rect 7646 34850 7698 34862
rect 8430 34914 8482 34926
rect 8430 34850 8482 34862
rect 8654 34914 8706 34926
rect 8654 34850 8706 34862
rect 8878 34914 8930 34926
rect 14254 34914 14306 34926
rect 10658 34862 10670 34914
rect 10722 34862 10734 34914
rect 18622 34914 18674 34926
rect 8878 34850 8930 34862
rect 14254 34850 14306 34862
rect 15250 34850 15262 34902
rect 15314 34850 15326 34902
rect 18622 34850 18674 34862
rect 19518 34914 19570 34926
rect 19518 34850 19570 34862
rect 21310 34914 21362 34926
rect 22990 34914 23042 34926
rect 22418 34862 22430 34914
rect 22482 34862 22494 34914
rect 21310 34850 21362 34862
rect 22990 34850 23042 34862
rect 23438 34914 23490 34926
rect 23438 34850 23490 34862
rect 23886 34914 23938 34926
rect 23886 34850 23938 34862
rect 24334 34914 24386 34926
rect 24334 34850 24386 34862
rect 25678 34914 25730 34926
rect 27918 34914 27970 34926
rect 26450 34862 26462 34914
rect 26514 34862 26526 34914
rect 27122 34862 27134 34914
rect 27186 34862 27198 34914
rect 27346 34862 27358 34914
rect 27410 34862 27422 34914
rect 25678 34850 25730 34862
rect 27918 34850 27970 34862
rect 29150 34914 29202 34926
rect 29150 34850 29202 34862
rect 29374 34914 29426 34926
rect 29374 34850 29426 34862
rect 29710 34914 29762 34926
rect 29710 34850 29762 34862
rect 30830 34914 30882 34926
rect 30830 34850 30882 34862
rect 31502 34914 31554 34926
rect 31502 34850 31554 34862
rect 32174 34914 32226 34926
rect 32174 34850 32226 34862
rect 32846 34914 32898 34926
rect 35870 34914 35922 34926
rect 34850 34862 34862 34914
rect 34914 34862 34926 34914
rect 32846 34850 32898 34862
rect 35870 34850 35922 34862
rect 35982 34914 36034 34926
rect 40462 34914 40514 34926
rect 42254 34914 42306 34926
rect 38210 34862 38222 34914
rect 38274 34862 38286 34914
rect 38658 34862 38670 34914
rect 38722 34862 38734 34914
rect 39330 34862 39342 34914
rect 39394 34862 39406 34914
rect 40114 34862 40126 34914
rect 40178 34862 40190 34914
rect 41794 34862 41806 34914
rect 41858 34862 41870 34914
rect 35982 34850 36034 34862
rect 40462 34850 40514 34862
rect 42254 34850 42306 34862
rect 42702 34914 42754 34926
rect 42702 34850 42754 34862
rect 42814 34914 42866 34926
rect 42814 34850 42866 34862
rect 45054 34914 45106 34926
rect 50430 34914 50482 34926
rect 47058 34862 47070 34914
rect 47122 34862 47134 34914
rect 45054 34850 45106 34862
rect 50430 34850 50482 34862
rect 53230 34914 53282 34926
rect 53554 34862 53566 34914
rect 53618 34862 53630 34914
rect 54450 34862 54462 34914
rect 54514 34862 54526 34914
rect 53230 34850 53282 34862
rect 7870 34802 7922 34814
rect 6962 34750 6974 34802
rect 7026 34750 7038 34802
rect 7870 34738 7922 34750
rect 9886 34802 9938 34814
rect 9886 34738 9938 34750
rect 9998 34802 10050 34814
rect 9998 34738 10050 34750
rect 10446 34802 10498 34814
rect 10446 34738 10498 34750
rect 10894 34802 10946 34814
rect 12686 34802 12738 34814
rect 11442 34750 11454 34802
rect 11506 34750 11518 34802
rect 10894 34738 10946 34750
rect 12686 34738 12738 34750
rect 14366 34802 14418 34814
rect 19966 34802 20018 34814
rect 15922 34750 15934 34802
rect 15986 34750 15998 34802
rect 14366 34738 14418 34750
rect 19966 34738 20018 34750
rect 20190 34802 20242 34814
rect 20190 34738 20242 34750
rect 21422 34802 21474 34814
rect 31166 34802 31218 34814
rect 32622 34802 32674 34814
rect 26338 34750 26350 34802
rect 26402 34750 26414 34802
rect 28578 34750 28590 34802
rect 28642 34750 28654 34802
rect 31826 34750 31838 34802
rect 31890 34750 31902 34802
rect 21422 34738 21474 34750
rect 31166 34738 31218 34750
rect 32622 34738 32674 34750
rect 35758 34802 35810 34814
rect 40686 34802 40738 34814
rect 39778 34750 39790 34802
rect 39842 34750 39854 34802
rect 35758 34738 35810 34750
rect 40686 34738 40738 34750
rect 40798 34802 40850 34814
rect 40798 34738 40850 34750
rect 43038 34802 43090 34814
rect 43038 34738 43090 34750
rect 46398 34802 46450 34814
rect 46722 34750 46734 34802
rect 46786 34750 46798 34802
rect 46398 34738 46450 34750
rect 2942 34690 2994 34702
rect 2942 34626 2994 34638
rect 7422 34690 7474 34702
rect 7422 34626 7474 34638
rect 8766 34690 8818 34702
rect 8766 34626 8818 34638
rect 10334 34690 10386 34702
rect 10334 34626 10386 34638
rect 11790 34690 11842 34702
rect 11790 34626 11842 34638
rect 12798 34690 12850 34702
rect 12798 34626 12850 34638
rect 13470 34690 13522 34702
rect 13470 34626 13522 34638
rect 14814 34690 14866 34702
rect 14814 34626 14866 34638
rect 21646 34690 21698 34702
rect 21646 34626 21698 34638
rect 24110 34690 24162 34702
rect 24110 34626 24162 34638
rect 24222 34690 24274 34702
rect 24222 34626 24274 34638
rect 25342 34690 25394 34702
rect 25342 34626 25394 34638
rect 26798 34690 26850 34702
rect 26798 34626 26850 34638
rect 26910 34690 26962 34702
rect 26910 34626 26962 34638
rect 27582 34690 27634 34702
rect 27582 34626 27634 34638
rect 27806 34690 27858 34702
rect 27806 34626 27858 34638
rect 28254 34690 28306 34702
rect 28254 34626 28306 34638
rect 29598 34690 29650 34702
rect 29598 34626 29650 34638
rect 30494 34690 30546 34702
rect 30494 34626 30546 34638
rect 31054 34690 31106 34702
rect 31054 34626 31106 34638
rect 42590 34690 42642 34702
rect 42590 34626 42642 34638
rect 45390 34690 45442 34702
rect 45390 34626 45442 34638
rect 53790 34690 53842 34702
rect 53790 34626 53842 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 7422 34354 7474 34366
rect 8990 34354 9042 34366
rect 8082 34302 8094 34354
rect 8146 34302 8158 34354
rect 8642 34302 8654 34354
rect 8706 34351 8718 34354
rect 8866 34351 8878 34354
rect 8706 34305 8878 34351
rect 8706 34302 8718 34305
rect 8866 34302 8878 34305
rect 8930 34302 8942 34354
rect 7422 34290 7474 34302
rect 8990 34290 9042 34302
rect 9998 34354 10050 34366
rect 9998 34290 10050 34302
rect 10110 34354 10162 34366
rect 10110 34290 10162 34302
rect 13470 34354 13522 34366
rect 15150 34354 15202 34366
rect 14578 34302 14590 34354
rect 14642 34302 14654 34354
rect 13470 34290 13522 34302
rect 15150 34290 15202 34302
rect 16046 34354 16098 34366
rect 16046 34290 16098 34302
rect 17502 34354 17554 34366
rect 17502 34290 17554 34302
rect 19294 34354 19346 34366
rect 24558 34354 24610 34366
rect 21634 34302 21646 34354
rect 21698 34302 21710 34354
rect 19294 34290 19346 34302
rect 24558 34290 24610 34302
rect 25342 34354 25394 34366
rect 34190 34354 34242 34366
rect 28914 34302 28926 34354
rect 28978 34302 28990 34354
rect 25342 34290 25394 34302
rect 34190 34290 34242 34302
rect 35310 34354 35362 34366
rect 50206 34354 50258 34366
rect 43362 34302 43374 34354
rect 43426 34302 43438 34354
rect 35310 34290 35362 34302
rect 50206 34290 50258 34302
rect 7758 34242 7810 34254
rect 15038 34242 15090 34254
rect 2482 34190 2494 34242
rect 2546 34190 2558 34242
rect 7970 34190 7982 34242
rect 8034 34190 8046 34242
rect 10770 34190 10782 34242
rect 10834 34190 10846 34242
rect 7758 34178 7810 34190
rect 15038 34178 15090 34190
rect 15262 34242 15314 34254
rect 15262 34178 15314 34190
rect 16270 34242 16322 34254
rect 16270 34178 16322 34190
rect 21086 34242 21138 34254
rect 31278 34242 31330 34254
rect 26898 34190 26910 34242
rect 26962 34190 26974 34242
rect 27570 34190 27582 34242
rect 27634 34190 27646 34242
rect 28466 34190 28478 34242
rect 28530 34190 28542 34242
rect 29922 34190 29934 34242
rect 29986 34190 29998 34242
rect 30930 34190 30942 34242
rect 30994 34190 31006 34242
rect 21086 34178 21138 34190
rect 31278 34178 31330 34190
rect 31726 34242 31778 34254
rect 31726 34178 31778 34190
rect 37998 34242 38050 34254
rect 37998 34178 38050 34190
rect 40350 34242 40402 34254
rect 50766 34242 50818 34254
rect 42690 34190 42702 34242
rect 42754 34190 42766 34242
rect 53890 34190 53902 34242
rect 53954 34190 53966 34242
rect 40350 34178 40402 34190
rect 50766 34178 50818 34190
rect 5070 34130 5122 34142
rect 1810 34078 1822 34130
rect 1874 34078 1886 34130
rect 5070 34066 5122 34078
rect 5294 34130 5346 34142
rect 5294 34066 5346 34078
rect 5406 34130 5458 34142
rect 9886 34130 9938 34142
rect 13246 34130 13298 34142
rect 7186 34078 7198 34130
rect 7250 34078 7262 34130
rect 8530 34078 8542 34130
rect 8594 34078 8606 34130
rect 10434 34078 10446 34130
rect 10498 34078 10510 34130
rect 10994 34078 11006 34130
rect 11058 34078 11070 34130
rect 11554 34078 11566 34130
rect 11618 34078 11630 34130
rect 12002 34078 12014 34130
rect 12066 34078 12078 34130
rect 13010 34078 13022 34130
rect 13074 34078 13086 34130
rect 5406 34066 5458 34078
rect 9886 34066 9938 34078
rect 13246 34066 13298 34078
rect 13582 34130 13634 34142
rect 13582 34066 13634 34078
rect 14030 34130 14082 34142
rect 14030 34066 14082 34078
rect 15934 34130 15986 34142
rect 15934 34066 15986 34078
rect 16494 34130 16546 34142
rect 18958 34130 19010 34142
rect 18610 34078 18622 34130
rect 18674 34078 18686 34130
rect 16494 34066 16546 34078
rect 18958 34066 19010 34078
rect 19854 34130 19906 34142
rect 19854 34066 19906 34078
rect 21310 34130 21362 34142
rect 21310 34066 21362 34078
rect 22654 34130 22706 34142
rect 25230 34130 25282 34142
rect 23090 34078 23102 34130
rect 23154 34078 23166 34130
rect 24658 34078 24670 34130
rect 24722 34078 24734 34130
rect 22654 34066 22706 34078
rect 25230 34066 25282 34078
rect 25566 34130 25618 34142
rect 30606 34130 30658 34142
rect 26226 34078 26238 34130
rect 26290 34078 26302 34130
rect 26786 34078 26798 34130
rect 26850 34078 26862 34130
rect 27906 34078 27918 34130
rect 27970 34078 27982 34130
rect 28354 34078 28366 34130
rect 28418 34078 28430 34130
rect 29362 34078 29374 34130
rect 29426 34078 29438 34130
rect 25566 34066 25618 34078
rect 30606 34066 30658 34078
rect 31502 34130 31554 34142
rect 34414 34130 34466 34142
rect 31938 34078 31950 34130
rect 32002 34078 32014 34130
rect 31502 34066 31554 34078
rect 34414 34066 34466 34078
rect 34862 34130 34914 34142
rect 34862 34066 34914 34078
rect 37102 34130 37154 34142
rect 37102 34066 37154 34078
rect 37662 34130 37714 34142
rect 39454 34130 39506 34142
rect 43038 34130 43090 34142
rect 38434 34078 38446 34130
rect 38498 34078 38510 34130
rect 39778 34078 39790 34130
rect 39842 34078 39854 34130
rect 41122 34078 41134 34130
rect 41186 34078 41198 34130
rect 41682 34078 41694 34130
rect 41746 34078 41758 34130
rect 37662 34066 37714 34078
rect 39454 34066 39506 34078
rect 43038 34066 43090 34078
rect 49534 34130 49586 34142
rect 49534 34066 49586 34078
rect 49758 34130 49810 34142
rect 49758 34066 49810 34078
rect 50094 34130 50146 34142
rect 50094 34066 50146 34078
rect 50430 34130 50482 34142
rect 50430 34066 50482 34078
rect 51662 34130 51714 34142
rect 51662 34066 51714 34078
rect 52222 34130 52274 34142
rect 52222 34066 52274 34078
rect 52782 34130 52834 34142
rect 53218 34078 53230 34130
rect 53282 34078 53294 34130
rect 52782 34066 52834 34078
rect 13358 34018 13410 34030
rect 20750 34018 20802 34030
rect 31614 34018 31666 34030
rect 4610 33966 4622 34018
rect 4674 33966 4686 34018
rect 18498 33966 18510 34018
rect 18562 33966 18574 34018
rect 28018 33966 28030 34018
rect 28082 33966 28094 34018
rect 13358 33954 13410 33966
rect 20750 33954 20802 33966
rect 31614 33954 31666 33966
rect 34302 34018 34354 34030
rect 47406 34018 47458 34030
rect 38770 33966 38782 34018
rect 38834 33966 38846 34018
rect 56018 33966 56030 34018
rect 56082 33966 56094 34018
rect 34302 33954 34354 33966
rect 47406 33954 47458 33966
rect 4958 33906 5010 33918
rect 12014 33906 12066 33918
rect 8306 33854 8318 33906
rect 8370 33854 8382 33906
rect 4958 33842 5010 33854
rect 12014 33842 12066 33854
rect 14254 33906 14306 33918
rect 20078 33906 20130 33918
rect 19394 33854 19406 33906
rect 19458 33903 19470 33906
rect 19618 33903 19630 33906
rect 19458 33857 19630 33903
rect 19458 33854 19470 33857
rect 19618 33854 19630 33857
rect 19682 33854 19694 33906
rect 14254 33842 14306 33854
rect 20078 33842 20130 33854
rect 20302 33906 20354 33918
rect 20302 33842 20354 33854
rect 24222 33906 24274 33918
rect 24222 33842 24274 33854
rect 24446 33906 24498 33918
rect 51326 33906 51378 33918
rect 49186 33854 49198 33906
rect 49250 33854 49262 33906
rect 24446 33842 24498 33854
rect 51326 33842 51378 33854
rect 51438 33906 51490 33918
rect 51438 33842 51490 33854
rect 51774 33906 51826 33918
rect 51774 33842 51826 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 10782 33570 10834 33582
rect 4722 33518 4734 33570
rect 4786 33567 4798 33570
rect 4946 33567 4958 33570
rect 4786 33521 4958 33567
rect 4786 33518 4798 33521
rect 4946 33518 4958 33521
rect 5010 33518 5022 33570
rect 10782 33506 10834 33518
rect 12686 33570 12738 33582
rect 19966 33570 20018 33582
rect 16258 33518 16270 33570
rect 16322 33567 16334 33570
rect 16482 33567 16494 33570
rect 16322 33521 16494 33567
rect 16322 33518 16334 33521
rect 16482 33518 16494 33521
rect 16546 33518 16558 33570
rect 12686 33506 12738 33518
rect 19966 33506 20018 33518
rect 20190 33570 20242 33582
rect 20190 33506 20242 33518
rect 20638 33570 20690 33582
rect 20638 33506 20690 33518
rect 22654 33570 22706 33582
rect 22654 33506 22706 33518
rect 31950 33570 32002 33582
rect 31950 33506 32002 33518
rect 39342 33570 39394 33582
rect 39342 33506 39394 33518
rect 39902 33570 39954 33582
rect 54002 33518 54014 33570
rect 54066 33567 54078 33570
rect 55010 33567 55022 33570
rect 54066 33521 55022 33567
rect 54066 33518 54078 33521
rect 55010 33518 55022 33521
rect 55074 33518 55086 33570
rect 39902 33506 39954 33518
rect 4846 33458 4898 33470
rect 12126 33458 12178 33470
rect 5954 33406 5966 33458
rect 6018 33406 6030 33458
rect 8082 33406 8094 33458
rect 8146 33406 8158 33458
rect 4846 33394 4898 33406
rect 12126 33394 12178 33406
rect 14814 33458 14866 33470
rect 14814 33394 14866 33406
rect 16494 33458 16546 33470
rect 16494 33394 16546 33406
rect 17054 33458 17106 33470
rect 17054 33394 17106 33406
rect 20302 33458 20354 33470
rect 48414 33458 48466 33470
rect 52782 33458 52834 33470
rect 36418 33406 36430 33458
rect 36482 33406 36494 33458
rect 46162 33406 46174 33458
rect 46226 33406 46238 33458
rect 50978 33406 50990 33458
rect 51042 33406 51054 33458
rect 20302 33394 20354 33406
rect 48414 33394 48466 33406
rect 52782 33394 52834 33406
rect 54014 33458 54066 33470
rect 54014 33394 54066 33406
rect 54574 33458 54626 33470
rect 54574 33394 54626 33406
rect 54910 33458 54962 33470
rect 54910 33394 54962 33406
rect 10558 33346 10610 33358
rect 13694 33346 13746 33358
rect 8754 33294 8766 33346
rect 8818 33294 8830 33346
rect 11666 33294 11678 33346
rect 11730 33294 11742 33346
rect 10558 33282 10610 33294
rect 13694 33282 13746 33294
rect 14142 33346 14194 33358
rect 14142 33282 14194 33294
rect 19182 33346 19234 33358
rect 21982 33346 22034 33358
rect 25118 33346 25170 33358
rect 19730 33294 19742 33346
rect 19794 33294 19806 33346
rect 22306 33294 22318 33346
rect 22370 33294 22382 33346
rect 19182 33282 19234 33294
rect 21982 33282 22034 33294
rect 25118 33282 25170 33294
rect 25342 33346 25394 33358
rect 26686 33346 26738 33358
rect 26226 33294 26238 33346
rect 26290 33294 26302 33346
rect 25342 33282 25394 33294
rect 26686 33282 26738 33294
rect 26910 33346 26962 33358
rect 26910 33282 26962 33294
rect 27470 33346 27522 33358
rect 27470 33282 27522 33294
rect 30606 33346 30658 33358
rect 30606 33282 30658 33294
rect 30942 33346 30994 33358
rect 32510 33346 32562 33358
rect 32274 33294 32286 33346
rect 32338 33294 32350 33346
rect 30942 33282 30994 33294
rect 32510 33282 32562 33294
rect 33182 33346 33234 33358
rect 39454 33346 39506 33358
rect 33618 33294 33630 33346
rect 33682 33294 33694 33346
rect 33182 33282 33234 33294
rect 39454 33282 39506 33294
rect 39790 33346 39842 33358
rect 46622 33346 46674 33358
rect 45826 33294 45838 33346
rect 45890 33294 45902 33346
rect 39790 33282 39842 33294
rect 46622 33282 46674 33294
rect 47182 33346 47234 33358
rect 49310 33346 49362 33358
rect 51214 33346 51266 33358
rect 48850 33294 48862 33346
rect 48914 33294 48926 33346
rect 50642 33294 50654 33346
rect 50706 33294 50718 33346
rect 47182 33282 47234 33294
rect 49310 33282 49362 33294
rect 51214 33282 51266 33294
rect 12686 33234 12738 33246
rect 11442 33182 11454 33234
rect 11506 33182 11518 33234
rect 12686 33170 12738 33182
rect 12798 33234 12850 33246
rect 12798 33170 12850 33182
rect 14366 33234 14418 33246
rect 14366 33170 14418 33182
rect 18846 33234 18898 33246
rect 18846 33170 18898 33182
rect 20750 33234 20802 33246
rect 22542 33234 22594 33246
rect 21746 33182 21758 33234
rect 21810 33182 21822 33234
rect 20750 33170 20802 33182
rect 22542 33170 22594 33182
rect 25678 33234 25730 33246
rect 27358 33234 27410 33246
rect 26002 33182 26014 33234
rect 26066 33182 26078 33234
rect 25678 33170 25730 33182
rect 27358 33170 27410 33182
rect 29150 33234 29202 33246
rect 29150 33170 29202 33182
rect 32734 33234 32786 33246
rect 32734 33170 32786 33182
rect 32958 33234 33010 33246
rect 39342 33234 39394 33246
rect 34290 33182 34302 33234
rect 34354 33182 34366 33234
rect 32958 33170 33010 33182
rect 39342 33170 39394 33182
rect 47742 33234 47794 33246
rect 47742 33170 47794 33182
rect 47966 33234 48018 33246
rect 50082 33182 50094 33234
rect 50146 33182 50158 33234
rect 51650 33182 51662 33234
rect 51714 33182 51726 33234
rect 47966 33170 48018 33182
rect 9326 33122 9378 33134
rect 12238 33122 12290 33134
rect 11106 33070 11118 33122
rect 11170 33070 11182 33122
rect 9326 33058 9378 33070
rect 12238 33058 12290 33070
rect 13918 33122 13970 33134
rect 13918 33058 13970 33070
rect 15598 33122 15650 33134
rect 15598 33058 15650 33070
rect 17950 33122 18002 33134
rect 19070 33122 19122 33134
rect 18274 33070 18286 33122
rect 18338 33070 18350 33122
rect 17950 33058 18002 33070
rect 19070 33058 19122 33070
rect 19294 33122 19346 33134
rect 19294 33058 19346 33070
rect 21422 33122 21474 33134
rect 21422 33058 21474 33070
rect 25566 33122 25618 33134
rect 25566 33058 25618 33070
rect 27134 33122 27186 33134
rect 27134 33058 27186 33070
rect 27806 33122 27858 33134
rect 27806 33058 27858 33070
rect 29486 33122 29538 33134
rect 29486 33058 29538 33070
rect 30718 33122 30770 33134
rect 30718 33058 30770 33070
rect 32062 33122 32114 33134
rect 32062 33058 32114 33070
rect 37102 33122 37154 33134
rect 37102 33058 37154 33070
rect 37550 33122 37602 33134
rect 37550 33058 37602 33070
rect 41470 33122 41522 33134
rect 41470 33058 41522 33070
rect 47854 33122 47906 33134
rect 47854 33058 47906 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 6526 32786 6578 32798
rect 6526 32722 6578 32734
rect 14366 32786 14418 32798
rect 14366 32722 14418 32734
rect 17390 32786 17442 32798
rect 17390 32722 17442 32734
rect 19182 32786 19234 32798
rect 19182 32722 19234 32734
rect 25230 32786 25282 32798
rect 27358 32786 27410 32798
rect 26114 32734 26126 32786
rect 26178 32734 26190 32786
rect 29822 32786 29874 32798
rect 25230 32722 25282 32734
rect 27358 32722 27410 32734
rect 27582 32730 27634 32742
rect 14702 32674 14754 32686
rect 3938 32622 3950 32674
rect 4002 32622 4014 32674
rect 14702 32610 14754 32622
rect 15262 32674 15314 32686
rect 15262 32610 15314 32622
rect 15598 32674 15650 32686
rect 15598 32610 15650 32622
rect 15822 32674 15874 32686
rect 15822 32610 15874 32622
rect 18622 32674 18674 32686
rect 18622 32610 18674 32622
rect 18846 32674 18898 32686
rect 18846 32610 18898 32622
rect 19406 32674 19458 32686
rect 19406 32610 19458 32622
rect 20862 32674 20914 32686
rect 29822 32722 29874 32734
rect 30046 32786 30098 32798
rect 32286 32786 32338 32798
rect 30258 32734 30270 32786
rect 30322 32783 30334 32786
rect 30482 32783 30494 32786
rect 30322 32737 30494 32783
rect 30322 32734 30334 32737
rect 30482 32734 30494 32737
rect 30546 32734 30558 32786
rect 30046 32722 30098 32734
rect 32286 32722 32338 32734
rect 39790 32786 39842 32798
rect 39790 32722 39842 32734
rect 46286 32786 46338 32798
rect 46286 32722 46338 32734
rect 47518 32786 47570 32798
rect 47518 32722 47570 32734
rect 47966 32786 48018 32798
rect 50530 32734 50542 32786
rect 50594 32734 50606 32786
rect 47966 32722 48018 32734
rect 21858 32622 21870 32674
rect 21922 32622 21934 32674
rect 24546 32622 24558 32674
rect 24610 32622 24622 32674
rect 26338 32622 26350 32674
rect 26402 32671 26414 32674
rect 26674 32671 26686 32674
rect 26402 32625 26686 32671
rect 26402 32622 26414 32625
rect 26674 32622 26686 32625
rect 26738 32622 26750 32674
rect 27582 32666 27634 32678
rect 27694 32674 27746 32686
rect 20862 32610 20914 32622
rect 27694 32610 27746 32622
rect 28478 32674 28530 32686
rect 28478 32610 28530 32622
rect 30606 32674 30658 32686
rect 30606 32610 30658 32622
rect 33182 32674 33234 32686
rect 37662 32674 37714 32686
rect 41022 32674 41074 32686
rect 45726 32674 45778 32686
rect 35186 32622 35198 32674
rect 35250 32622 35262 32674
rect 39106 32622 39118 32674
rect 39170 32622 39182 32674
rect 44594 32622 44606 32674
rect 44658 32622 44670 32674
rect 33182 32610 33234 32622
rect 37662 32610 37714 32622
rect 41022 32610 41074 32622
rect 45726 32610 45778 32622
rect 48190 32674 48242 32686
rect 48190 32610 48242 32622
rect 48750 32674 48802 32686
rect 48750 32610 48802 32622
rect 49646 32674 49698 32686
rect 49646 32610 49698 32622
rect 51774 32674 51826 32686
rect 51774 32610 51826 32622
rect 16158 32562 16210 32574
rect 19518 32562 19570 32574
rect 25342 32562 25394 32574
rect 3266 32510 3278 32562
rect 3330 32510 3342 32562
rect 16594 32510 16606 32562
rect 16658 32510 16670 32562
rect 20402 32510 20414 32562
rect 20466 32510 20478 32562
rect 21298 32510 21310 32562
rect 21362 32510 21374 32562
rect 22418 32510 22430 32562
rect 22482 32510 22494 32562
rect 22978 32510 22990 32562
rect 23042 32510 23054 32562
rect 24322 32510 24334 32562
rect 24386 32510 24398 32562
rect 16158 32498 16210 32510
rect 19518 32498 19570 32510
rect 25342 32498 25394 32510
rect 25790 32562 25842 32574
rect 25790 32498 25842 32510
rect 26798 32562 26850 32574
rect 26798 32498 26850 32510
rect 28590 32562 28642 32574
rect 29262 32562 29314 32574
rect 28802 32510 28814 32562
rect 28866 32510 28878 32562
rect 28590 32498 28642 32510
rect 29262 32498 29314 32510
rect 29374 32562 29426 32574
rect 29374 32498 29426 32510
rect 30830 32562 30882 32574
rect 31838 32562 31890 32574
rect 31154 32510 31166 32562
rect 31218 32510 31230 32562
rect 30830 32498 30882 32510
rect 31838 32498 31890 32510
rect 32062 32562 32114 32574
rect 32062 32498 32114 32510
rect 32398 32562 32450 32574
rect 32398 32498 32450 32510
rect 33070 32562 33122 32574
rect 38782 32562 38834 32574
rect 34514 32510 34526 32562
rect 34578 32510 34590 32562
rect 33070 32498 33122 32510
rect 38782 32498 38834 32510
rect 39678 32562 39730 32574
rect 39678 32498 39730 32510
rect 41134 32562 41186 32574
rect 46734 32562 46786 32574
rect 42130 32510 42142 32562
rect 42194 32510 42206 32562
rect 45378 32510 45390 32562
rect 45442 32510 45454 32562
rect 41134 32498 41186 32510
rect 46734 32498 46786 32510
rect 48974 32562 49026 32574
rect 48974 32498 49026 32510
rect 49198 32562 49250 32574
rect 49198 32498 49250 32510
rect 49310 32562 49362 32574
rect 49310 32498 49362 32510
rect 50206 32562 50258 32574
rect 51662 32562 51714 32574
rect 51202 32510 51214 32562
rect 51266 32510 51278 32562
rect 51538 32510 51550 32562
rect 51602 32510 51614 32562
rect 54226 32510 54238 32562
rect 54290 32510 54302 32562
rect 55010 32510 55022 32562
rect 55074 32510 55086 32562
rect 50206 32498 50258 32510
rect 51662 32498 51714 32510
rect 10894 32450 10946 32462
rect 6066 32398 6078 32450
rect 6130 32398 6142 32450
rect 10894 32386 10946 32398
rect 13806 32450 13858 32462
rect 13806 32386 13858 32398
rect 15374 32450 15426 32462
rect 15374 32386 15426 32398
rect 17950 32450 18002 32462
rect 28254 32450 28306 32462
rect 18946 32398 18958 32450
rect 19010 32398 19022 32450
rect 20514 32398 20526 32450
rect 20578 32398 20590 32450
rect 21186 32398 21198 32450
rect 21250 32398 21262 32450
rect 21970 32398 21982 32450
rect 22034 32398 22046 32450
rect 27010 32398 27022 32450
rect 27074 32398 27086 32450
rect 17950 32386 18002 32398
rect 28254 32386 28306 32398
rect 29934 32450 29986 32462
rect 29934 32386 29986 32398
rect 31614 32450 31666 32462
rect 31614 32386 31666 32398
rect 31726 32450 31778 32462
rect 31726 32386 31778 32398
rect 33630 32450 33682 32462
rect 47406 32450 47458 32462
rect 48862 32450 48914 32462
rect 37314 32398 37326 32450
rect 37378 32398 37390 32450
rect 38098 32398 38110 32450
rect 38162 32398 38174 32450
rect 42466 32398 42478 32450
rect 42530 32398 42542 32450
rect 47842 32398 47854 32450
rect 47906 32398 47918 32450
rect 33630 32386 33682 32398
rect 47406 32386 47458 32398
rect 48862 32386 48914 32398
rect 49982 32450 50034 32462
rect 52098 32398 52110 32450
rect 52162 32398 52174 32450
rect 49982 32386 50034 32398
rect 14590 32338 14642 32350
rect 14130 32286 14142 32338
rect 14194 32335 14206 32338
rect 14354 32335 14366 32338
rect 14194 32289 14366 32335
rect 14194 32286 14206 32289
rect 14354 32286 14366 32289
rect 14418 32286 14430 32338
rect 14590 32274 14642 32286
rect 31390 32338 31442 32350
rect 31390 32274 31442 32286
rect 39790 32338 39842 32350
rect 39790 32274 39842 32286
rect 41022 32338 41074 32350
rect 41022 32274 41074 32286
rect 41806 32338 41858 32350
rect 41806 32274 41858 32286
rect 42142 32338 42194 32350
rect 42142 32274 42194 32286
rect 51326 32338 51378 32350
rect 51326 32274 51378 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 22082 31950 22094 32002
rect 22146 31950 22158 32002
rect 24994 31950 25006 32002
rect 25058 31950 25070 32002
rect 14702 31890 14754 31902
rect 8530 31838 8542 31890
rect 8594 31838 8606 31890
rect 10658 31838 10670 31890
rect 10722 31838 10734 31890
rect 14702 31826 14754 31838
rect 17838 31890 17890 31902
rect 17838 31826 17890 31838
rect 20302 31890 20354 31902
rect 25902 31890 25954 31902
rect 34638 31890 34690 31902
rect 52670 31890 52722 31902
rect 24658 31838 24670 31890
rect 24722 31838 24734 31890
rect 31602 31838 31614 31890
rect 31666 31838 31678 31890
rect 33730 31838 33742 31890
rect 33794 31838 33806 31890
rect 40338 31838 40350 31890
rect 40402 31838 40414 31890
rect 41346 31838 41358 31890
rect 41410 31838 41422 31890
rect 46498 31838 46510 31890
rect 46562 31838 46574 31890
rect 48626 31838 48638 31890
rect 48690 31838 48702 31890
rect 50418 31838 50430 31890
rect 50482 31838 50494 31890
rect 20302 31826 20354 31838
rect 25902 31826 25954 31838
rect 34638 31826 34690 31838
rect 52670 31826 52722 31838
rect 52782 31890 52834 31902
rect 52782 31826 52834 31838
rect 11006 31778 11058 31790
rect 7746 31726 7758 31778
rect 7810 31726 7822 31778
rect 11006 31714 11058 31726
rect 11566 31778 11618 31790
rect 12462 31778 12514 31790
rect 15262 31778 15314 31790
rect 19742 31778 19794 31790
rect 12002 31726 12014 31778
rect 12066 31726 12078 31778
rect 13458 31726 13470 31778
rect 13522 31726 13534 31778
rect 14130 31726 14142 31778
rect 14194 31726 14206 31778
rect 16034 31726 16046 31778
rect 16098 31726 16110 31778
rect 11566 31714 11618 31726
rect 12462 31714 12514 31726
rect 15262 31714 15314 31726
rect 19742 31714 19794 31726
rect 20414 31778 20466 31790
rect 21422 31778 21474 31790
rect 22542 31778 22594 31790
rect 20738 31726 20750 31778
rect 20802 31726 20814 31778
rect 21634 31726 21646 31778
rect 21698 31726 21710 31778
rect 20414 31714 20466 31726
rect 21422 31714 21474 31726
rect 22542 31714 22594 31726
rect 23214 31778 23266 31790
rect 25790 31778 25842 31790
rect 30046 31778 30098 31790
rect 23650 31726 23662 31778
rect 23714 31726 23726 31778
rect 24210 31726 24222 31778
rect 24274 31726 24286 31778
rect 24770 31726 24782 31778
rect 24834 31726 24846 31778
rect 26786 31726 26798 31778
rect 26850 31726 26862 31778
rect 27906 31726 27918 31778
rect 27970 31726 27982 31778
rect 23214 31714 23266 31726
rect 25790 31714 25842 31726
rect 30046 31714 30098 31726
rect 30270 31778 30322 31790
rect 30270 31714 30322 31726
rect 30606 31778 30658 31790
rect 34190 31778 34242 31790
rect 30930 31726 30942 31778
rect 30994 31726 31006 31778
rect 30606 31714 30658 31726
rect 34190 31714 34242 31726
rect 36990 31778 37042 31790
rect 36990 31714 37042 31726
rect 37886 31778 37938 31790
rect 38782 31778 38834 31790
rect 49422 31778 49474 31790
rect 38546 31726 38558 31778
rect 38610 31726 38622 31778
rect 39330 31726 39342 31778
rect 39394 31726 39406 31778
rect 39890 31726 39902 31778
rect 39954 31726 39966 31778
rect 40226 31726 40238 31778
rect 40290 31726 40302 31778
rect 43474 31726 43486 31778
rect 43538 31726 43550 31778
rect 44258 31726 44270 31778
rect 44322 31726 44334 31778
rect 45826 31726 45838 31778
rect 45890 31726 45902 31778
rect 37886 31714 37938 31726
rect 38782 31714 38834 31726
rect 49422 31714 49474 31726
rect 49646 31778 49698 31790
rect 49646 31714 49698 31726
rect 49982 31778 50034 31790
rect 51214 31778 51266 31790
rect 50754 31726 50766 31778
rect 50818 31726 50830 31778
rect 49982 31714 50034 31726
rect 51214 31714 51266 31726
rect 51774 31778 51826 31790
rect 51774 31714 51826 31726
rect 6302 31666 6354 31678
rect 6302 31602 6354 31614
rect 14814 31666 14866 31678
rect 14814 31602 14866 31614
rect 17166 31666 17218 31678
rect 17166 31602 17218 31614
rect 18622 31666 18674 31678
rect 18622 31602 18674 31614
rect 22654 31666 22706 31678
rect 22654 31602 22706 31614
rect 26238 31666 26290 31678
rect 27358 31666 27410 31678
rect 26450 31614 26462 31666
rect 26514 31614 26526 31666
rect 26238 31602 26290 31614
rect 27358 31602 27410 31614
rect 27470 31666 27522 31678
rect 27470 31602 27522 31614
rect 29150 31666 29202 31678
rect 29150 31602 29202 31614
rect 29262 31666 29314 31678
rect 29262 31602 29314 31614
rect 37214 31666 37266 31678
rect 37214 31602 37266 31614
rect 37326 31666 37378 31678
rect 37326 31602 37378 31614
rect 37662 31666 37714 31678
rect 37662 31602 37714 31614
rect 38894 31666 38946 31678
rect 51550 31666 51602 31678
rect 40786 31614 40798 31666
rect 40850 31614 40862 31666
rect 38894 31602 38946 31614
rect 51550 31602 51602 31614
rect 6190 31554 6242 31566
rect 6190 31490 6242 31502
rect 13694 31554 13746 31566
rect 13694 31490 13746 31502
rect 13806 31554 13858 31566
rect 13806 31490 13858 31502
rect 13918 31554 13970 31566
rect 13918 31490 13970 31502
rect 14590 31554 14642 31566
rect 14590 31490 14642 31502
rect 20190 31554 20242 31566
rect 20190 31490 20242 31502
rect 26574 31554 26626 31566
rect 26574 31490 26626 31502
rect 27134 31554 27186 31566
rect 27134 31490 27186 31502
rect 27246 31554 27298 31566
rect 27246 31490 27298 31502
rect 29486 31554 29538 31566
rect 29486 31490 29538 31502
rect 30270 31554 30322 31566
rect 44942 31554 44994 31566
rect 38210 31502 38222 31554
rect 38274 31502 38286 31554
rect 30270 31490 30322 31502
rect 44942 31490 44994 31502
rect 45390 31554 45442 31566
rect 45390 31490 45442 31502
rect 49758 31554 49810 31566
rect 52098 31502 52110 31554
rect 52162 31502 52174 31554
rect 49758 31490 49810 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 8542 31218 8594 31230
rect 8542 31154 8594 31166
rect 9102 31218 9154 31230
rect 9102 31154 9154 31166
rect 9662 31218 9714 31230
rect 9662 31154 9714 31166
rect 10334 31218 10386 31230
rect 10334 31154 10386 31166
rect 14926 31218 14978 31230
rect 14926 31154 14978 31166
rect 15822 31218 15874 31230
rect 15822 31154 15874 31166
rect 17390 31218 17442 31230
rect 17390 31154 17442 31166
rect 17502 31218 17554 31230
rect 19070 31218 19122 31230
rect 18386 31166 18398 31218
rect 18450 31166 18462 31218
rect 17502 31154 17554 31166
rect 19070 31154 19122 31166
rect 21086 31218 21138 31230
rect 21086 31154 21138 31166
rect 26014 31218 26066 31230
rect 26014 31154 26066 31166
rect 27694 31218 27746 31230
rect 27694 31154 27746 31166
rect 34638 31218 34690 31230
rect 34638 31154 34690 31166
rect 37550 31218 37602 31230
rect 37550 31154 37602 31166
rect 40014 31218 40066 31230
rect 40014 31154 40066 31166
rect 40238 31218 40290 31230
rect 40238 31154 40290 31166
rect 42142 31218 42194 31230
rect 42142 31154 42194 31166
rect 48190 31218 48242 31230
rect 48190 31154 48242 31166
rect 48862 31218 48914 31230
rect 48862 31154 48914 31166
rect 49422 31218 49474 31230
rect 51998 31218 52050 31230
rect 50530 31166 50542 31218
rect 50594 31166 50606 31218
rect 49422 31154 49474 31166
rect 51998 31154 52050 31166
rect 10558 31106 10610 31118
rect 5730 31054 5742 31106
rect 5794 31054 5806 31106
rect 8194 31054 8206 31106
rect 8258 31054 8270 31106
rect 10558 31042 10610 31054
rect 14478 31106 14530 31118
rect 14478 31042 14530 31054
rect 15262 31106 15314 31118
rect 15262 31042 15314 31054
rect 15710 31106 15762 31118
rect 17614 31106 17666 31118
rect 24558 31106 24610 31118
rect 33070 31106 33122 31118
rect 16594 31054 16606 31106
rect 16658 31054 16670 31106
rect 19842 31054 19854 31106
rect 19906 31054 19918 31106
rect 30146 31054 30158 31106
rect 30210 31054 30222 31106
rect 15710 31042 15762 31054
rect 17614 31042 17666 31054
rect 24558 31042 24610 31054
rect 33070 31042 33122 31054
rect 33294 31106 33346 31118
rect 33294 31042 33346 31054
rect 33966 31106 34018 31118
rect 33966 31042 34018 31054
rect 34078 31106 34130 31118
rect 34078 31042 34130 31054
rect 37326 31106 37378 31118
rect 37326 31042 37378 31054
rect 37774 31106 37826 31118
rect 37774 31042 37826 31054
rect 38110 31106 38162 31118
rect 38110 31042 38162 31054
rect 41918 31106 41970 31118
rect 41918 31042 41970 31054
rect 42366 31106 42418 31118
rect 50418 31054 50430 31106
rect 50482 31054 50494 31106
rect 42366 31042 42418 31054
rect 10894 30994 10946 31006
rect 5058 30942 5070 30994
rect 5122 30942 5134 30994
rect 10894 30930 10946 30942
rect 11118 30994 11170 31006
rect 11118 30930 11170 30942
rect 11342 30994 11394 31006
rect 11342 30930 11394 30942
rect 12014 30994 12066 31006
rect 12014 30930 12066 30942
rect 12574 30994 12626 31006
rect 12574 30930 12626 30942
rect 13806 30994 13858 31006
rect 13806 30930 13858 30942
rect 14254 30994 14306 31006
rect 16270 30994 16322 31006
rect 15474 30942 15486 30994
rect 15538 30942 15550 30994
rect 14254 30930 14306 30942
rect 16270 30930 16322 30942
rect 18062 30994 18114 31006
rect 18062 30930 18114 30942
rect 18734 30994 18786 31006
rect 19630 30994 19682 31006
rect 20974 30994 21026 31006
rect 19282 30942 19294 30994
rect 19346 30942 19358 30994
rect 20178 30942 20190 30994
rect 20242 30942 20254 30994
rect 18734 30930 18786 30942
rect 19630 30930 19682 30942
rect 20974 30930 21026 30942
rect 21198 30994 21250 31006
rect 21198 30930 21250 30942
rect 21422 30994 21474 31006
rect 21422 30930 21474 30942
rect 21646 30994 21698 31006
rect 25342 30994 25394 31006
rect 22306 30942 22318 30994
rect 22370 30942 22382 30994
rect 22754 30942 22766 30994
rect 22818 30942 22830 30994
rect 23314 30942 23326 30994
rect 23378 30942 23390 30994
rect 21646 30930 21698 30942
rect 25342 30930 25394 30942
rect 25790 30994 25842 31006
rect 25790 30930 25842 30942
rect 25902 30994 25954 31006
rect 33742 30994 33794 31006
rect 39118 30994 39170 31006
rect 40350 30994 40402 31006
rect 26674 30942 26686 30994
rect 26738 30942 26750 30994
rect 27010 30942 27022 30994
rect 27074 30942 27086 30994
rect 29474 30942 29486 30994
rect 29538 30942 29550 30994
rect 38322 30942 38334 30994
rect 38386 30942 38398 30994
rect 39442 30942 39454 30994
rect 39506 30942 39518 30994
rect 25902 30930 25954 30942
rect 33742 30930 33794 30942
rect 39118 30930 39170 30942
rect 40350 30930 40402 30942
rect 41022 30994 41074 31006
rect 42478 30994 42530 31006
rect 41234 30942 41246 30994
rect 41298 30942 41310 30994
rect 41022 30930 41074 30942
rect 42478 30930 42530 30942
rect 50094 30994 50146 31006
rect 50094 30930 50146 30942
rect 50654 30994 50706 31006
rect 50654 30930 50706 30942
rect 50878 30994 50930 31006
rect 50878 30930 50930 30942
rect 51102 30994 51154 31006
rect 51102 30930 51154 30942
rect 51438 30994 51490 31006
rect 51438 30930 51490 30942
rect 14030 30882 14082 30894
rect 7858 30830 7870 30882
rect 7922 30830 7934 30882
rect 14030 30818 14082 30830
rect 19406 30882 19458 30894
rect 23998 30882 24050 30894
rect 33518 30882 33570 30894
rect 49758 30882 49810 30894
rect 20514 30830 20526 30882
rect 20578 30830 20590 30882
rect 22194 30830 22206 30882
rect 22258 30830 22270 30882
rect 32274 30830 32286 30882
rect 32338 30830 32350 30882
rect 39554 30830 39566 30882
rect 39618 30830 39630 30882
rect 19406 30818 19458 30830
rect 23998 30818 24050 30830
rect 33518 30818 33570 30830
rect 49758 30818 49810 30830
rect 51550 30882 51602 30894
rect 51550 30818 51602 30830
rect 10222 30770 10274 30782
rect 10222 30706 10274 30718
rect 11790 30770 11842 30782
rect 11790 30706 11842 30718
rect 24334 30770 24386 30782
rect 34078 30770 34130 30782
rect 27010 30718 27022 30770
rect 27074 30718 27086 30770
rect 24334 30706 24386 30718
rect 34078 30706 34130 30718
rect 37886 30770 37938 30782
rect 37886 30706 37938 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 7310 30434 7362 30446
rect 7310 30370 7362 30382
rect 12238 30434 12290 30446
rect 12238 30370 12290 30382
rect 12350 30434 12402 30446
rect 12350 30370 12402 30382
rect 12574 30434 12626 30446
rect 12574 30370 12626 30382
rect 14926 30434 14978 30446
rect 14926 30370 14978 30382
rect 15598 30434 15650 30446
rect 21422 30434 21474 30446
rect 18386 30382 18398 30434
rect 18450 30382 18462 30434
rect 15598 30370 15650 30382
rect 21422 30370 21474 30382
rect 22990 30434 23042 30446
rect 22990 30370 23042 30382
rect 23326 30434 23378 30446
rect 23326 30370 23378 30382
rect 24782 30434 24834 30446
rect 24782 30370 24834 30382
rect 34750 30434 34802 30446
rect 34750 30370 34802 30382
rect 15710 30322 15762 30334
rect 41246 30322 41298 30334
rect 6962 30270 6974 30322
rect 7026 30270 7038 30322
rect 11106 30270 11118 30322
rect 11170 30270 11182 30322
rect 13794 30270 13806 30322
rect 13858 30270 13870 30322
rect 38210 30270 38222 30322
rect 38274 30270 38286 30322
rect 40114 30270 40126 30322
rect 40178 30270 40190 30322
rect 52098 30270 52110 30322
rect 52162 30270 52174 30322
rect 15710 30258 15762 30270
rect 41246 30258 41298 30270
rect 11790 30210 11842 30222
rect 8306 30158 8318 30210
rect 8370 30158 8382 30210
rect 8978 30158 8990 30210
rect 9042 30158 9054 30210
rect 11790 30146 11842 30158
rect 12798 30210 12850 30222
rect 12798 30146 12850 30158
rect 14478 30210 14530 30222
rect 14478 30146 14530 30158
rect 14702 30210 14754 30222
rect 17166 30210 17218 30222
rect 15026 30158 15038 30210
rect 15090 30158 15102 30210
rect 15922 30158 15934 30210
rect 15986 30158 15998 30210
rect 14702 30146 14754 30158
rect 17166 30146 17218 30158
rect 17502 30210 17554 30222
rect 17502 30146 17554 30158
rect 18174 30210 18226 30222
rect 18958 30210 19010 30222
rect 18610 30158 18622 30210
rect 18674 30158 18686 30210
rect 18174 30146 18226 30158
rect 18958 30146 19010 30158
rect 21534 30210 21586 30222
rect 21534 30146 21586 30158
rect 21982 30210 22034 30222
rect 21982 30146 22034 30158
rect 22318 30210 22370 30222
rect 23998 30210 24050 30222
rect 22978 30158 22990 30210
rect 23042 30158 23054 30210
rect 22318 30146 22370 30158
rect 23998 30146 24050 30158
rect 24334 30210 24386 30222
rect 24334 30146 24386 30158
rect 24894 30210 24946 30222
rect 24894 30146 24946 30158
rect 25230 30210 25282 30222
rect 25230 30146 25282 30158
rect 25342 30210 25394 30222
rect 28702 30210 28754 30222
rect 35870 30210 35922 30222
rect 38782 30210 38834 30222
rect 39790 30210 39842 30222
rect 48862 30210 48914 30222
rect 25778 30158 25790 30210
rect 25842 30158 25854 30210
rect 29138 30158 29150 30210
rect 29202 30158 29214 30210
rect 37762 30158 37774 30210
rect 37826 30158 37838 30210
rect 39106 30158 39118 30210
rect 39170 30158 39182 30210
rect 40226 30158 40238 30210
rect 40290 30158 40302 30210
rect 49298 30158 49310 30210
rect 49362 30158 49374 30210
rect 49970 30158 49982 30210
rect 50034 30158 50046 30210
rect 25342 30146 25394 30158
rect 28702 30146 28754 30158
rect 35870 30146 35922 30158
rect 38782 30146 38834 30158
rect 39790 30146 39842 30158
rect 48862 30146 48914 30158
rect 13470 30098 13522 30110
rect 13470 30034 13522 30046
rect 15262 30098 15314 30110
rect 15262 30034 15314 30046
rect 17390 30098 17442 30110
rect 17390 30034 17442 30046
rect 17838 30098 17890 30110
rect 17838 30034 17890 30046
rect 22654 30098 22706 30110
rect 36430 30098 36482 30110
rect 26674 30046 26686 30098
rect 26738 30046 26750 30098
rect 32834 30046 32846 30098
rect 32898 30046 32910 30098
rect 22654 30034 22706 30046
rect 36430 30034 36482 30046
rect 37326 30098 37378 30110
rect 37326 30034 37378 30046
rect 41470 30098 41522 30110
rect 41470 30034 41522 30046
rect 7086 29986 7138 29998
rect 7086 29922 7138 29934
rect 12686 29986 12738 29998
rect 12686 29922 12738 29934
rect 13694 29986 13746 29998
rect 13694 29922 13746 29934
rect 13918 29986 13970 29998
rect 13918 29922 13970 29934
rect 14142 29986 14194 29998
rect 14142 29922 14194 29934
rect 14366 29986 14418 29998
rect 14366 29922 14418 29934
rect 17950 29986 18002 29998
rect 17950 29922 18002 29934
rect 19518 29986 19570 29998
rect 19518 29922 19570 29934
rect 21422 29986 21474 29998
rect 21422 29922 21474 29934
rect 22542 29986 22594 29998
rect 22542 29922 22594 29934
rect 24110 29986 24162 29998
rect 24110 29922 24162 29934
rect 24782 29986 24834 29998
rect 24782 29922 24834 29934
rect 27022 29986 27074 29998
rect 27022 29922 27074 29934
rect 34862 29986 34914 29998
rect 34862 29922 34914 29934
rect 34974 29986 35026 29998
rect 34974 29922 35026 29934
rect 40910 29986 40962 29998
rect 40910 29922 40962 29934
rect 41358 29986 41410 29998
rect 41358 29922 41410 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 11230 29650 11282 29662
rect 11230 29586 11282 29598
rect 12014 29650 12066 29662
rect 12014 29586 12066 29598
rect 18622 29650 18674 29662
rect 18622 29586 18674 29598
rect 20526 29650 20578 29662
rect 20526 29586 20578 29598
rect 22094 29650 22146 29662
rect 23550 29650 23602 29662
rect 28366 29650 28418 29662
rect 22866 29598 22878 29650
rect 22930 29598 22942 29650
rect 27458 29598 27470 29650
rect 27522 29598 27534 29650
rect 22094 29586 22146 29598
rect 23550 29586 23602 29598
rect 28366 29586 28418 29598
rect 28702 29650 28754 29662
rect 28702 29586 28754 29598
rect 35758 29650 35810 29662
rect 35758 29586 35810 29598
rect 13134 29538 13186 29550
rect 15038 29538 15090 29550
rect 6850 29486 6862 29538
rect 6914 29486 6926 29538
rect 13346 29486 13358 29538
rect 13410 29486 13422 29538
rect 13134 29474 13186 29486
rect 15038 29474 15090 29486
rect 15150 29538 15202 29550
rect 15150 29474 15202 29486
rect 19070 29538 19122 29550
rect 19070 29474 19122 29486
rect 20862 29538 20914 29550
rect 20862 29474 20914 29486
rect 23662 29538 23714 29550
rect 23662 29474 23714 29486
rect 29598 29538 29650 29550
rect 32286 29538 32338 29550
rect 37438 29538 37490 29550
rect 29922 29486 29934 29538
rect 29986 29486 29998 29538
rect 34290 29486 34302 29538
rect 34354 29486 34366 29538
rect 29598 29474 29650 29486
rect 32286 29474 32338 29486
rect 37438 29474 37490 29486
rect 40350 29538 40402 29550
rect 43362 29486 43374 29538
rect 43426 29486 43438 29538
rect 40350 29474 40402 29486
rect 12686 29426 12738 29438
rect 6178 29374 6190 29426
rect 6242 29374 6254 29426
rect 12686 29362 12738 29374
rect 13806 29426 13858 29438
rect 13806 29362 13858 29374
rect 14254 29426 14306 29438
rect 17502 29426 17554 29438
rect 15810 29374 15822 29426
rect 15874 29374 15886 29426
rect 16482 29374 16494 29426
rect 16546 29374 16558 29426
rect 14254 29362 14306 29374
rect 17502 29362 17554 29374
rect 17950 29426 18002 29438
rect 17950 29362 18002 29374
rect 22542 29426 22594 29438
rect 27806 29426 27858 29438
rect 26450 29374 26462 29426
rect 26514 29374 26526 29426
rect 26898 29374 26910 29426
rect 26962 29374 26974 29426
rect 22542 29362 22594 29374
rect 27806 29362 27858 29374
rect 29262 29426 29314 29438
rect 32510 29426 32562 29438
rect 33406 29426 33458 29438
rect 31938 29374 31950 29426
rect 32002 29374 32014 29426
rect 33058 29374 33070 29426
rect 33122 29374 33134 29426
rect 29262 29362 29314 29374
rect 32510 29362 32562 29374
rect 33406 29362 33458 29374
rect 33518 29426 33570 29438
rect 33518 29362 33570 29374
rect 33630 29426 33682 29438
rect 33630 29362 33682 29374
rect 35870 29426 35922 29438
rect 35870 29362 35922 29374
rect 36318 29426 36370 29438
rect 40238 29426 40290 29438
rect 44606 29426 44658 29438
rect 39666 29374 39678 29426
rect 39730 29374 39742 29426
rect 44034 29374 44046 29426
rect 44098 29374 44110 29426
rect 36318 29362 36370 29374
rect 40238 29362 40290 29374
rect 44606 29362 44658 29374
rect 9774 29314 9826 29326
rect 13470 29314 13522 29326
rect 8978 29262 8990 29314
rect 9042 29262 9054 29314
rect 11554 29262 11566 29314
rect 11618 29262 11630 29314
rect 9774 29250 9826 29262
rect 13470 29250 13522 29262
rect 16606 29314 16658 29326
rect 16606 29250 16658 29262
rect 20974 29314 21026 29326
rect 20974 29250 21026 29262
rect 25454 29314 25506 29326
rect 25454 29250 25506 29262
rect 25902 29314 25954 29326
rect 25902 29250 25954 29262
rect 27134 29314 27186 29326
rect 27134 29250 27186 29262
rect 32398 29314 32450 29326
rect 32398 29250 32450 29262
rect 38894 29314 38946 29326
rect 41234 29262 41246 29314
rect 41298 29262 41310 29314
rect 38894 29250 38946 29262
rect 12462 29202 12514 29214
rect 15038 29202 15090 29214
rect 14466 29150 14478 29202
rect 14530 29150 14542 29202
rect 12462 29138 12514 29150
rect 15038 29138 15090 29150
rect 15598 29202 15650 29214
rect 19182 29202 19234 29214
rect 38670 29202 38722 29214
rect 17266 29150 17278 29202
rect 17330 29199 17342 29202
rect 17938 29199 17950 29202
rect 17330 29153 17950 29199
rect 17330 29150 17342 29153
rect 17938 29150 17950 29153
rect 18002 29150 18014 29202
rect 38322 29150 38334 29202
rect 38386 29150 38398 29202
rect 15598 29138 15650 29150
rect 19182 29138 19234 29150
rect 38670 29138 38722 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 13694 28866 13746 28878
rect 13694 28802 13746 28814
rect 14814 28866 14866 28878
rect 14814 28802 14866 28814
rect 16158 28866 16210 28878
rect 16158 28802 16210 28814
rect 23438 28866 23490 28878
rect 23438 28802 23490 28814
rect 32398 28866 32450 28878
rect 32398 28802 32450 28814
rect 42142 28866 42194 28878
rect 42142 28802 42194 28814
rect 6974 28754 7026 28766
rect 6974 28690 7026 28702
rect 14702 28754 14754 28766
rect 19966 28754 20018 28766
rect 18386 28702 18398 28754
rect 18450 28702 18462 28754
rect 14702 28690 14754 28702
rect 19966 28690 20018 28702
rect 24446 28754 24498 28766
rect 24446 28690 24498 28702
rect 27470 28754 27522 28766
rect 27470 28690 27522 28702
rect 28366 28754 28418 28766
rect 36990 28754 37042 28766
rect 32050 28702 32062 28754
rect 32114 28702 32126 28754
rect 33842 28702 33854 28754
rect 33906 28702 33918 28754
rect 35970 28702 35982 28754
rect 36034 28702 36046 28754
rect 38434 28702 38446 28754
rect 38498 28702 38510 28754
rect 28366 28690 28418 28702
rect 36990 28690 37042 28702
rect 6526 28642 6578 28654
rect 6526 28578 6578 28590
rect 13470 28642 13522 28654
rect 13470 28578 13522 28590
rect 17054 28642 17106 28654
rect 17054 28578 17106 28590
rect 17278 28642 17330 28654
rect 18958 28642 19010 28654
rect 18274 28590 18286 28642
rect 18338 28590 18350 28642
rect 17278 28578 17330 28590
rect 18958 28578 19010 28590
rect 19070 28642 19122 28654
rect 19070 28578 19122 28590
rect 19182 28642 19234 28654
rect 19182 28578 19234 28590
rect 19406 28642 19458 28654
rect 19406 28578 19458 28590
rect 20302 28642 20354 28654
rect 20302 28578 20354 28590
rect 21422 28642 21474 28654
rect 21422 28578 21474 28590
rect 22094 28642 22146 28654
rect 22094 28578 22146 28590
rect 22654 28642 22706 28654
rect 22654 28578 22706 28590
rect 23102 28642 23154 28654
rect 23102 28578 23154 28590
rect 25678 28642 25730 28654
rect 26910 28642 26962 28654
rect 26338 28590 26350 28642
rect 26402 28590 26414 28642
rect 25678 28578 25730 28590
rect 26910 28578 26962 28590
rect 27022 28642 27074 28654
rect 27022 28578 27074 28590
rect 27358 28642 27410 28654
rect 39790 28642 39842 28654
rect 27682 28590 27694 28642
rect 27746 28590 27758 28642
rect 29250 28590 29262 28642
rect 29314 28590 29326 28642
rect 33170 28590 33182 28642
rect 33234 28590 33246 28642
rect 37426 28590 37438 28642
rect 37490 28590 37502 28642
rect 37986 28590 37998 28642
rect 38050 28590 38062 28642
rect 38882 28590 38894 28642
rect 38946 28590 38958 28642
rect 27358 28578 27410 28590
rect 39790 28578 39842 28590
rect 40126 28642 40178 28654
rect 40126 28578 40178 28590
rect 41806 28642 41858 28654
rect 41806 28578 41858 28590
rect 41918 28642 41970 28654
rect 41918 28578 41970 28590
rect 16046 28530 16098 28542
rect 18622 28530 18674 28542
rect 22430 28530 22482 28542
rect 16706 28478 16718 28530
rect 16770 28478 16782 28530
rect 20626 28478 20638 28530
rect 20690 28478 20702 28530
rect 16046 28466 16098 28478
rect 18622 28466 18674 28478
rect 22430 28466 22482 28478
rect 23326 28530 23378 28542
rect 23326 28466 23378 28478
rect 23438 28530 23490 28542
rect 32622 28530 32674 28542
rect 25330 28478 25342 28530
rect 25394 28478 25406 28530
rect 29922 28478 29934 28530
rect 29986 28478 29998 28530
rect 23438 28466 23490 28478
rect 32622 28466 32674 28478
rect 36430 28530 36482 28542
rect 39454 28530 39506 28542
rect 38098 28478 38110 28530
rect 38162 28478 38174 28530
rect 36430 28466 36482 28478
rect 39454 28466 39506 28478
rect 39566 28530 39618 28542
rect 39566 28466 39618 28478
rect 42254 28530 42306 28542
rect 42254 28466 42306 28478
rect 16158 28418 16210 28430
rect 6178 28366 6190 28418
rect 6242 28366 6254 28418
rect 14018 28366 14030 28418
rect 14082 28366 14094 28418
rect 16158 28354 16210 28366
rect 17726 28418 17778 28430
rect 17726 28354 17778 28366
rect 17838 28418 17890 28430
rect 17838 28354 17890 28366
rect 17950 28418 18002 28430
rect 17950 28354 18002 28366
rect 21870 28418 21922 28430
rect 21870 28354 21922 28366
rect 21982 28418 22034 28430
rect 21982 28354 22034 28366
rect 22542 28418 22594 28430
rect 22542 28354 22594 28366
rect 24110 28418 24162 28430
rect 24110 28354 24162 28366
rect 32510 28418 32562 28430
rect 32510 28354 32562 28366
rect 40238 28418 40290 28430
rect 40238 28354 40290 28366
rect 40462 28418 40514 28430
rect 40462 28354 40514 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 8206 28082 8258 28094
rect 8206 28018 8258 28030
rect 16046 28082 16098 28094
rect 16046 28018 16098 28030
rect 16606 28082 16658 28094
rect 16606 28018 16658 28030
rect 24782 28082 24834 28094
rect 24782 28018 24834 28030
rect 25454 28082 25506 28094
rect 25454 28018 25506 28030
rect 29598 28082 29650 28094
rect 29598 28018 29650 28030
rect 30046 28082 30098 28094
rect 30046 28018 30098 28030
rect 30606 28082 30658 28094
rect 30606 28018 30658 28030
rect 36430 28082 36482 28094
rect 37650 28030 37662 28082
rect 37714 28030 37726 28082
rect 37986 28030 37998 28082
rect 38050 28030 38062 28082
rect 36430 28018 36482 28030
rect 16718 27970 16770 27982
rect 30158 27970 30210 27982
rect 37102 27970 37154 27982
rect 10210 27918 10222 27970
rect 10274 27918 10286 27970
rect 18162 27918 18174 27970
rect 18226 27918 18238 27970
rect 22754 27918 22766 27970
rect 22818 27918 22830 27970
rect 33842 27918 33854 27970
rect 33906 27918 33918 27970
rect 16718 27906 16770 27918
rect 30158 27906 30210 27918
rect 37102 27906 37154 27918
rect 40126 27970 40178 27982
rect 41682 27918 41694 27970
rect 41746 27918 41758 27970
rect 40126 27906 40178 27918
rect 10558 27858 10610 27870
rect 4946 27806 4958 27858
rect 5010 27806 5022 27858
rect 9874 27806 9886 27858
rect 9938 27806 9950 27858
rect 10558 27794 10610 27806
rect 13134 27858 13186 27870
rect 13134 27794 13186 27806
rect 13358 27858 13410 27870
rect 32286 27858 32338 27870
rect 37326 27858 37378 27870
rect 13570 27806 13582 27858
rect 13634 27806 13646 27858
rect 17490 27806 17502 27858
rect 17554 27806 17566 27858
rect 23426 27806 23438 27858
rect 23490 27806 23502 27858
rect 29810 27806 29822 27858
rect 29874 27806 29886 27858
rect 33170 27806 33182 27858
rect 33234 27806 33246 27858
rect 13358 27794 13410 27806
rect 32286 27794 32338 27806
rect 37326 27794 37378 27806
rect 38334 27858 38386 27870
rect 38334 27794 38386 27806
rect 38558 27858 38610 27870
rect 38558 27794 38610 27806
rect 38894 27858 38946 27870
rect 39330 27806 39342 27858
rect 39394 27806 39406 27858
rect 39778 27806 39790 27858
rect 39842 27806 39854 27858
rect 40786 27806 40798 27858
rect 40850 27806 40862 27858
rect 41906 27806 41918 27858
rect 41970 27806 41982 27858
rect 38894 27794 38946 27806
rect 15150 27746 15202 27758
rect 5618 27694 5630 27746
rect 5682 27694 5694 27746
rect 7746 27694 7758 27746
rect 7810 27694 7822 27746
rect 15150 27682 15202 27694
rect 15598 27746 15650 27758
rect 24334 27746 24386 27758
rect 20290 27694 20302 27746
rect 20354 27694 20366 27746
rect 20626 27694 20638 27746
rect 20690 27694 20702 27746
rect 35970 27694 35982 27746
rect 36034 27694 36046 27746
rect 41458 27694 41470 27746
rect 41522 27694 41534 27746
rect 15598 27682 15650 27694
rect 24334 27682 24386 27694
rect 9550 27634 9602 27646
rect 9550 27570 9602 27582
rect 9886 27634 9938 27646
rect 9886 27570 9938 27582
rect 13022 27634 13074 27646
rect 25230 27634 25282 27646
rect 15138 27582 15150 27634
rect 15202 27631 15214 27634
rect 16258 27631 16270 27634
rect 15202 27585 16270 27631
rect 15202 27582 15214 27585
rect 16258 27582 16270 27585
rect 16322 27582 16334 27634
rect 13022 27570 13074 27582
rect 25230 27570 25282 27582
rect 25566 27634 25618 27646
rect 25566 27570 25618 27582
rect 30494 27634 30546 27646
rect 30494 27570 30546 27582
rect 30830 27634 30882 27646
rect 30830 27570 30882 27582
rect 39790 27634 39842 27646
rect 39790 27570 39842 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 5742 27298 5794 27310
rect 5742 27234 5794 27246
rect 12462 27298 12514 27310
rect 41458 27246 41470 27298
rect 41522 27246 41534 27298
rect 12462 27234 12514 27246
rect 6078 27186 6130 27198
rect 6078 27122 6130 27134
rect 6526 27186 6578 27198
rect 14702 27186 14754 27198
rect 18734 27186 18786 27198
rect 9538 27134 9550 27186
rect 9602 27134 9614 27186
rect 10210 27134 10222 27186
rect 10274 27134 10286 27186
rect 15810 27134 15822 27186
rect 15874 27134 15886 27186
rect 17938 27134 17950 27186
rect 18002 27134 18014 27186
rect 6526 27122 6578 27134
rect 14702 27122 14754 27134
rect 18734 27122 18786 27134
rect 19294 27186 19346 27198
rect 19294 27122 19346 27134
rect 22430 27186 22482 27198
rect 36430 27186 36482 27198
rect 25666 27134 25678 27186
rect 25730 27134 25742 27186
rect 29922 27134 29934 27186
rect 29986 27134 29998 27186
rect 32050 27134 32062 27186
rect 32114 27134 32126 27186
rect 33394 27134 33406 27186
rect 33458 27134 33470 27186
rect 35522 27134 35534 27186
rect 35586 27134 35598 27186
rect 39890 27134 39902 27186
rect 39954 27134 39966 27186
rect 40786 27134 40798 27186
rect 40850 27134 40862 27186
rect 22430 27122 22482 27134
rect 36430 27122 36482 27134
rect 7982 27074 8034 27086
rect 11454 27074 11506 27086
rect 8866 27022 8878 27074
rect 8930 27022 8942 27074
rect 9650 27022 9662 27074
rect 9714 27022 9726 27074
rect 10434 27022 10446 27074
rect 10498 27022 10510 27074
rect 7982 27010 8034 27022
rect 11454 27010 11506 27022
rect 12238 27074 12290 27086
rect 35870 27074 35922 27086
rect 41806 27074 41858 27086
rect 15026 27022 15038 27074
rect 15090 27022 15102 27074
rect 22866 27022 22878 27074
rect 22930 27022 22942 27074
rect 23538 27022 23550 27074
rect 23602 27022 23614 27074
rect 29250 27022 29262 27074
rect 29314 27022 29326 27074
rect 32722 27022 32734 27074
rect 32786 27022 32798 27074
rect 36978 27022 36990 27074
rect 37042 27022 37054 27074
rect 40674 27022 40686 27074
rect 40738 27022 40750 27074
rect 12238 27010 12290 27022
rect 35870 27010 35922 27022
rect 41806 27010 41858 27022
rect 42142 27074 42194 27086
rect 42142 27010 42194 27022
rect 5854 26962 5906 26974
rect 8542 26962 8594 26974
rect 11118 26962 11170 26974
rect 14254 26962 14306 26974
rect 42030 26962 42082 26974
rect 7634 26910 7646 26962
rect 7698 26910 7710 26962
rect 9314 26910 9326 26962
rect 9378 26910 9390 26962
rect 11554 26910 11566 26962
rect 11618 26910 11630 26962
rect 11890 26910 11902 26962
rect 11954 26910 11966 26962
rect 37762 26910 37774 26962
rect 37826 26910 37838 26962
rect 5854 26898 5906 26910
rect 8542 26898 8594 26910
rect 11118 26898 11170 26910
rect 14254 26898 14306 26910
rect 42030 26898 42082 26910
rect 42478 26962 42530 26974
rect 42478 26898 42530 26910
rect 14590 26850 14642 26862
rect 14590 26786 14642 26798
rect 18622 26850 18674 26862
rect 18622 26786 18674 26798
rect 20526 26850 20578 26862
rect 20526 26786 20578 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 7198 26514 7250 26526
rect 7198 26450 7250 26462
rect 9998 26514 10050 26526
rect 9998 26450 10050 26462
rect 14590 26514 14642 26526
rect 14590 26450 14642 26462
rect 15822 26514 15874 26526
rect 15822 26450 15874 26462
rect 16494 26514 16546 26526
rect 16494 26450 16546 26462
rect 20974 26514 21026 26526
rect 20974 26450 21026 26462
rect 35534 26514 35586 26526
rect 35534 26450 35586 26462
rect 35982 26514 36034 26526
rect 35982 26450 36034 26462
rect 36430 26514 36482 26526
rect 36430 26450 36482 26462
rect 39678 26514 39730 26526
rect 39678 26450 39730 26462
rect 39902 26514 39954 26526
rect 39902 26450 39954 26462
rect 40462 26514 40514 26526
rect 40462 26450 40514 26462
rect 41358 26514 41410 26526
rect 41358 26450 41410 26462
rect 41470 26514 41522 26526
rect 41470 26450 41522 26462
rect 42142 26514 42194 26526
rect 42142 26450 42194 26462
rect 8878 26402 8930 26414
rect 14366 26402 14418 26414
rect 12226 26350 12238 26402
rect 12290 26350 12302 26402
rect 13122 26350 13134 26402
rect 13186 26350 13198 26402
rect 8878 26338 8930 26350
rect 14366 26338 14418 26350
rect 17502 26402 17554 26414
rect 17502 26338 17554 26350
rect 18622 26402 18674 26414
rect 18622 26338 18674 26350
rect 19854 26402 19906 26414
rect 31054 26402 31106 26414
rect 26002 26350 26014 26402
rect 26066 26350 26078 26402
rect 19854 26338 19906 26350
rect 31054 26338 31106 26350
rect 36766 26402 36818 26414
rect 36766 26338 36818 26350
rect 7310 26290 7362 26302
rect 8766 26290 8818 26302
rect 9774 26290 9826 26302
rect 10894 26290 10946 26302
rect 15038 26290 15090 26302
rect 16046 26290 16098 26302
rect 3490 26238 3502 26290
rect 3554 26238 3566 26290
rect 8418 26238 8430 26290
rect 8482 26238 8494 26290
rect 9538 26238 9550 26290
rect 9602 26238 9614 26290
rect 10210 26238 10222 26290
rect 10274 26238 10286 26290
rect 13346 26238 13358 26290
rect 13410 26238 13422 26290
rect 15250 26238 15262 26290
rect 15314 26238 15326 26290
rect 15810 26238 15822 26290
rect 15874 26238 15886 26290
rect 7310 26226 7362 26238
rect 8766 26226 8818 26238
rect 9774 26226 9826 26238
rect 10894 26226 10946 26238
rect 15038 26226 15090 26238
rect 16046 26226 16098 26238
rect 16718 26290 16770 26302
rect 36878 26290 36930 26302
rect 18274 26238 18286 26290
rect 18338 26238 18350 26290
rect 18834 26238 18846 26290
rect 18898 26238 18910 26290
rect 19170 26238 19182 26290
rect 19234 26238 19246 26290
rect 25330 26238 25342 26290
rect 25394 26238 25406 26290
rect 30594 26238 30606 26290
rect 30658 26238 30670 26290
rect 16718 26226 16770 26238
rect 36878 26226 36930 26238
rect 37102 26290 37154 26302
rect 39566 26290 39618 26302
rect 41246 26290 41298 26302
rect 37314 26238 37326 26290
rect 37378 26238 37390 26290
rect 40898 26238 40910 26290
rect 40962 26238 40974 26290
rect 37102 26226 37154 26238
rect 39566 26226 39618 26238
rect 41246 26226 41298 26238
rect 41806 26290 41858 26302
rect 41806 26226 41858 26238
rect 6750 26178 6802 26190
rect 16606 26178 16658 26190
rect 4162 26126 4174 26178
rect 4226 26126 4238 26178
rect 6290 26126 6302 26178
rect 6354 26126 6366 26178
rect 9650 26126 9662 26178
rect 9714 26126 9726 26178
rect 13234 26126 13246 26178
rect 13298 26126 13310 26178
rect 6750 26114 6802 26126
rect 16606 26114 16658 26126
rect 18734 26178 18786 26190
rect 18734 26114 18786 26126
rect 20302 26178 20354 26190
rect 20302 26114 20354 26126
rect 24670 26178 24722 26190
rect 24670 26114 24722 26126
rect 28142 26178 28194 26190
rect 31390 26178 31442 26190
rect 30818 26126 30830 26178
rect 30882 26126 30894 26178
rect 28142 26114 28194 26126
rect 31390 26114 31442 26126
rect 31614 26178 31666 26190
rect 31614 26114 31666 26126
rect 32398 26178 32450 26190
rect 32398 26114 32450 26126
rect 7198 26066 7250 26078
rect 7198 26002 7250 26014
rect 14702 26066 14754 26078
rect 14702 26002 14754 26014
rect 15486 26066 15538 26078
rect 15486 26002 15538 26014
rect 17390 26066 17442 26078
rect 17390 26002 17442 26014
rect 17950 26066 18002 26078
rect 17950 26002 18002 26014
rect 18286 26066 18338 26078
rect 18286 26002 18338 26014
rect 19070 26066 19122 26078
rect 31938 26014 31950 26066
rect 32002 26014 32014 26066
rect 19070 26002 19122 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 5630 25730 5682 25742
rect 5630 25666 5682 25678
rect 5966 25730 6018 25742
rect 5966 25666 6018 25678
rect 14926 25730 14978 25742
rect 14926 25666 14978 25678
rect 30718 25730 30770 25742
rect 30718 25666 30770 25678
rect 7646 25618 7698 25630
rect 11230 25618 11282 25630
rect 30494 25618 30546 25630
rect 7186 25566 7198 25618
rect 7250 25566 7262 25618
rect 10322 25566 10334 25618
rect 10386 25566 10398 25618
rect 12338 25566 12350 25618
rect 12402 25566 12414 25618
rect 12786 25566 12798 25618
rect 12850 25566 12862 25618
rect 17266 25566 17278 25618
rect 17330 25566 17342 25618
rect 18610 25566 18622 25618
rect 18674 25566 18686 25618
rect 20738 25566 20750 25618
rect 20802 25566 20814 25618
rect 22082 25566 22094 25618
rect 22146 25566 22158 25618
rect 24210 25566 24222 25618
rect 24274 25566 24286 25618
rect 28578 25566 28590 25618
rect 28642 25566 28654 25618
rect 7646 25554 7698 25566
rect 11230 25554 11282 25566
rect 30494 25554 30546 25566
rect 36542 25618 36594 25630
rect 42814 25618 42866 25630
rect 39442 25566 39454 25618
rect 39506 25566 39518 25618
rect 41570 25566 41582 25618
rect 41634 25566 41646 25618
rect 36542 25554 36594 25566
rect 42814 25554 42866 25566
rect 9550 25506 9602 25518
rect 14478 25506 14530 25518
rect 15934 25506 15986 25518
rect 5618 25454 5630 25506
rect 5682 25454 5694 25506
rect 7298 25454 7310 25506
rect 7362 25454 7374 25506
rect 10770 25454 10782 25506
rect 10834 25454 10846 25506
rect 12226 25454 12238 25506
rect 12290 25454 12302 25506
rect 13010 25454 13022 25506
rect 13074 25454 13086 25506
rect 14690 25454 14702 25506
rect 14754 25454 14766 25506
rect 15138 25454 15150 25506
rect 15202 25454 15214 25506
rect 16594 25454 16606 25506
rect 16658 25454 16670 25506
rect 17378 25454 17390 25506
rect 17442 25454 17454 25506
rect 17826 25454 17838 25506
rect 17890 25454 17902 25506
rect 21298 25454 21310 25506
rect 21362 25454 21374 25506
rect 25778 25454 25790 25506
rect 25842 25454 25854 25506
rect 42354 25454 42366 25506
rect 42418 25454 42430 25506
rect 9550 25442 9602 25454
rect 14478 25442 14530 25454
rect 15934 25442 15986 25454
rect 9662 25394 9714 25406
rect 8754 25342 8766 25394
rect 8818 25342 8830 25394
rect 9314 25342 9326 25394
rect 9378 25342 9390 25394
rect 14130 25342 14142 25394
rect 14194 25342 14206 25394
rect 17490 25342 17502 25394
rect 17554 25342 17566 25394
rect 26450 25342 26462 25394
rect 26514 25342 26526 25394
rect 9662 25330 9714 25342
rect 13806 25282 13858 25294
rect 13806 25218 13858 25230
rect 14590 25282 14642 25294
rect 14590 25218 14642 25230
rect 16046 25282 16098 25294
rect 16046 25218 16098 25230
rect 24670 25282 24722 25294
rect 24670 25218 24722 25230
rect 25342 25282 25394 25294
rect 33630 25282 33682 25294
rect 31042 25230 31054 25282
rect 31106 25230 31118 25282
rect 25342 25218 25394 25230
rect 33630 25218 33682 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 10782 24946 10834 24958
rect 10782 24882 10834 24894
rect 11006 24946 11058 24958
rect 11006 24882 11058 24894
rect 36430 24946 36482 24958
rect 36430 24882 36482 24894
rect 36878 24946 36930 24958
rect 36878 24882 36930 24894
rect 10334 24834 10386 24846
rect 7858 24782 7870 24834
rect 7922 24782 7934 24834
rect 10334 24770 10386 24782
rect 10670 24834 10722 24846
rect 14590 24834 14642 24846
rect 13458 24782 13470 24834
rect 13522 24782 13534 24834
rect 10670 24770 10722 24782
rect 14590 24770 14642 24782
rect 16830 24834 16882 24846
rect 20862 24834 20914 24846
rect 17826 24782 17838 24834
rect 17890 24782 17902 24834
rect 20066 24782 20078 24834
rect 20130 24782 20142 24834
rect 16830 24770 16882 24782
rect 20862 24770 20914 24782
rect 28926 24834 28978 24846
rect 28926 24770 28978 24782
rect 32510 24834 32562 24846
rect 33842 24782 33854 24834
rect 33906 24782 33918 24834
rect 32510 24770 32562 24782
rect 18062 24722 18114 24734
rect 9762 24670 9774 24722
rect 9826 24670 9838 24722
rect 14242 24670 14254 24722
rect 14306 24670 14318 24722
rect 15026 24670 15038 24722
rect 15090 24670 15102 24722
rect 17602 24670 17614 24722
rect 17666 24670 17678 24722
rect 18062 24658 18114 24670
rect 18510 24722 18562 24734
rect 18510 24658 18562 24670
rect 18734 24722 18786 24734
rect 18734 24658 18786 24670
rect 19070 24722 19122 24734
rect 19070 24658 19122 24670
rect 19294 24722 19346 24734
rect 19294 24658 19346 24670
rect 20414 24722 20466 24734
rect 20414 24658 20466 24670
rect 20750 24722 20802 24734
rect 20750 24658 20802 24670
rect 21086 24722 21138 24734
rect 21086 24658 21138 24670
rect 32174 24722 32226 24734
rect 33170 24670 33182 24722
rect 33234 24670 33246 24722
rect 32174 24658 32226 24670
rect 18286 24610 18338 24622
rect 7634 24558 7646 24610
rect 7698 24558 7710 24610
rect 9650 24558 9662 24610
rect 9714 24558 9726 24610
rect 11330 24558 11342 24610
rect 11394 24558 11406 24610
rect 15474 24558 15486 24610
rect 15538 24558 15550 24610
rect 16370 24558 16382 24610
rect 16434 24558 16446 24610
rect 18286 24546 18338 24558
rect 26910 24610 26962 24622
rect 38222 24610 38274 24622
rect 35970 24558 35982 24610
rect 36034 24558 36046 24610
rect 26910 24546 26962 24558
rect 38222 24546 38274 24558
rect 38670 24610 38722 24622
rect 38670 24546 38722 24558
rect 8654 24498 8706 24510
rect 26798 24498 26850 24510
rect 19618 24446 19630 24498
rect 19682 24446 19694 24498
rect 8654 24434 8706 24446
rect 26798 24434 26850 24446
rect 28814 24498 28866 24510
rect 28814 24434 28866 24446
rect 38110 24498 38162 24510
rect 38110 24434 38162 24446
rect 38558 24498 38610 24510
rect 38558 24434 38610 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 9326 24162 9378 24174
rect 9326 24098 9378 24110
rect 14590 24162 14642 24174
rect 14590 24098 14642 24110
rect 32062 24162 32114 24174
rect 32062 24098 32114 24110
rect 14030 24050 14082 24062
rect 8754 23998 8766 24050
rect 8818 23998 8830 24050
rect 12898 23998 12910 24050
rect 12962 23998 12974 24050
rect 18386 23998 18398 24050
rect 18450 23998 18462 24050
rect 26898 23998 26910 24050
rect 26962 23998 26974 24050
rect 29474 23998 29486 24050
rect 29538 23998 29550 24050
rect 35970 23998 35982 24050
rect 36034 23998 36046 24050
rect 39890 23998 39902 24050
rect 39954 23998 39966 24050
rect 14030 23986 14082 23998
rect 7310 23938 7362 23950
rect 13470 23938 13522 23950
rect 5618 23886 5630 23938
rect 5682 23886 5694 23938
rect 8530 23886 8542 23938
rect 8594 23886 8606 23938
rect 10098 23886 10110 23938
rect 10162 23886 10174 23938
rect 7310 23874 7362 23886
rect 13470 23874 13522 23886
rect 14814 23938 14866 23950
rect 15822 23938 15874 23950
rect 15026 23886 15038 23938
rect 15090 23886 15102 23938
rect 14814 23874 14866 23886
rect 15822 23874 15874 23886
rect 15934 23938 15986 23950
rect 15934 23874 15986 23886
rect 16046 23938 16098 23950
rect 16046 23874 16098 23886
rect 16494 23938 16546 23950
rect 32398 23938 32450 23950
rect 18162 23886 18174 23938
rect 18226 23886 18238 23938
rect 19730 23886 19742 23938
rect 19794 23886 19806 23938
rect 20402 23886 20414 23938
rect 20466 23886 20478 23938
rect 20626 23886 20638 23938
rect 20690 23886 20702 23938
rect 23986 23886 23998 23938
rect 24050 23886 24062 23938
rect 33618 23886 33630 23938
rect 33682 23886 33694 23938
rect 36978 23886 36990 23938
rect 37042 23886 37054 23938
rect 16494 23874 16546 23886
rect 32398 23874 32450 23886
rect 5966 23826 6018 23838
rect 5966 23762 6018 23774
rect 6974 23826 7026 23838
rect 6974 23762 7026 23774
rect 7086 23826 7138 23838
rect 7086 23762 7138 23774
rect 7534 23826 7586 23838
rect 7534 23762 7586 23774
rect 7870 23826 7922 23838
rect 7870 23762 7922 23774
rect 9214 23826 9266 23838
rect 14478 23826 14530 23838
rect 18958 23826 19010 23838
rect 21310 23826 21362 23838
rect 10770 23774 10782 23826
rect 10834 23774 10846 23826
rect 16818 23774 16830 23826
rect 16882 23774 16894 23826
rect 17378 23774 17390 23826
rect 17442 23774 17454 23826
rect 20290 23774 20302 23826
rect 20354 23774 20366 23826
rect 9214 23762 9266 23774
rect 14478 23762 14530 23774
rect 18958 23762 19010 23774
rect 21310 23762 21362 23774
rect 23550 23826 23602 23838
rect 27470 23826 27522 23838
rect 24770 23774 24782 23826
rect 24834 23774 24846 23826
rect 23550 23762 23602 23774
rect 27470 23762 27522 23774
rect 27694 23826 27746 23838
rect 27694 23762 27746 23774
rect 28030 23826 28082 23838
rect 28030 23762 28082 23774
rect 29150 23826 29202 23838
rect 32610 23774 32622 23826
rect 32674 23774 32686 23826
rect 33170 23774 33182 23826
rect 33234 23774 33246 23826
rect 37762 23774 37774 23826
rect 37826 23774 37838 23826
rect 29150 23762 29202 23774
rect 5854 23714 5906 23726
rect 5854 23650 5906 23662
rect 7198 23714 7250 23726
rect 19070 23714 19122 23726
rect 22206 23714 22258 23726
rect 15362 23662 15374 23714
rect 15426 23662 15438 23714
rect 21634 23662 21646 23714
rect 21698 23662 21710 23714
rect 7198 23650 7250 23662
rect 19070 23650 19122 23662
rect 22206 23650 22258 23662
rect 23214 23714 23266 23726
rect 23214 23650 23266 23662
rect 23662 23714 23714 23726
rect 23662 23650 23714 23662
rect 27806 23714 27858 23726
rect 27806 23650 27858 23662
rect 29374 23714 29426 23726
rect 29374 23650 29426 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 7310 23378 7362 23390
rect 7310 23314 7362 23326
rect 7534 23378 7586 23390
rect 7534 23314 7586 23326
rect 7646 23378 7698 23390
rect 25566 23378 25618 23390
rect 13570 23326 13582 23378
rect 13634 23326 13646 23378
rect 21410 23326 21422 23378
rect 21474 23326 21486 23378
rect 7646 23314 7698 23326
rect 25566 23314 25618 23326
rect 8318 23266 8370 23278
rect 15150 23266 15202 23278
rect 3938 23214 3950 23266
rect 4002 23214 4014 23266
rect 14242 23214 14254 23266
rect 14306 23214 14318 23266
rect 8318 23202 8370 23214
rect 15150 23202 15202 23214
rect 15374 23266 15426 23278
rect 18398 23266 18450 23278
rect 16482 23214 16494 23266
rect 16546 23214 16558 23266
rect 15374 23202 15426 23214
rect 18398 23202 18450 23214
rect 20750 23266 20802 23278
rect 20750 23202 20802 23214
rect 20862 23266 20914 23278
rect 20862 23202 20914 23214
rect 27246 23266 27298 23278
rect 27246 23202 27298 23214
rect 31726 23266 31778 23278
rect 31726 23202 31778 23214
rect 32062 23266 32114 23278
rect 32062 23202 32114 23214
rect 33182 23266 33234 23278
rect 34862 23266 34914 23278
rect 33730 23214 33742 23266
rect 33794 23214 33806 23266
rect 34066 23214 34078 23266
rect 34130 23214 34142 23266
rect 33182 23202 33234 23214
rect 34862 23202 34914 23214
rect 7422 23154 7474 23166
rect 8206 23154 8258 23166
rect 20974 23154 21026 23166
rect 25230 23154 25282 23166
rect 3266 23102 3278 23154
rect 3330 23102 3342 23154
rect 7858 23102 7870 23154
rect 7922 23102 7934 23154
rect 10098 23102 10110 23154
rect 10162 23102 10174 23154
rect 11442 23102 11454 23154
rect 11506 23102 11518 23154
rect 12898 23102 12910 23154
rect 12962 23102 12974 23154
rect 13458 23102 13470 23154
rect 13522 23102 13534 23154
rect 16706 23102 16718 23154
rect 16770 23102 16782 23154
rect 17378 23102 17390 23154
rect 17442 23102 17454 23154
rect 24658 23102 24670 23154
rect 24722 23102 24734 23154
rect 7422 23090 7474 23102
rect 8206 23090 8258 23102
rect 20974 23090 21026 23102
rect 25230 23090 25282 23102
rect 25566 23154 25618 23166
rect 25566 23090 25618 23102
rect 25902 23154 25954 23166
rect 25902 23090 25954 23102
rect 26126 23154 26178 23166
rect 31054 23154 31106 23166
rect 26450 23102 26462 23154
rect 26514 23102 26526 23154
rect 27682 23102 27694 23154
rect 27746 23102 27758 23154
rect 35858 23102 35870 23154
rect 35922 23102 35934 23154
rect 26126 23090 26178 23102
rect 31054 23090 31106 23102
rect 6526 23042 6578 23054
rect 10782 23042 10834 23054
rect 6066 22990 6078 23042
rect 6130 22990 6142 23042
rect 10322 22990 10334 23042
rect 10386 22990 10398 23042
rect 6526 22978 6578 22990
rect 10782 22978 10834 22990
rect 19182 23042 19234 23054
rect 19182 22978 19234 22990
rect 19742 23042 19794 23054
rect 26238 23042 26290 23054
rect 32510 23042 32562 23054
rect 21746 22990 21758 23042
rect 21810 22990 21822 23042
rect 23874 22990 23886 23042
rect 23938 22990 23950 23042
rect 27346 22990 27358 23042
rect 27410 22990 27422 23042
rect 28466 22990 28478 23042
rect 28530 22990 28542 23042
rect 30594 22990 30606 23042
rect 30658 22990 30670 23042
rect 19742 22978 19794 22990
rect 26238 22978 26290 22990
rect 32510 22978 32562 22990
rect 35310 23042 35362 23054
rect 36530 22990 36542 23042
rect 36594 22990 36606 23042
rect 38658 22990 38670 23042
rect 38722 22990 38734 23042
rect 35310 22978 35362 22990
rect 15486 22930 15538 22942
rect 15486 22866 15538 22878
rect 16718 22930 16770 22942
rect 16718 22866 16770 22878
rect 27022 22930 27074 22942
rect 27022 22866 27074 22878
rect 30942 22930 30994 22942
rect 30942 22866 30994 22878
rect 33518 22930 33570 22942
rect 33518 22866 33570 22878
rect 34750 22930 34802 22942
rect 34750 22866 34802 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 14142 22594 14194 22606
rect 14142 22530 14194 22542
rect 14926 22594 14978 22606
rect 14926 22530 14978 22542
rect 20414 22594 20466 22606
rect 20414 22530 20466 22542
rect 21310 22594 21362 22606
rect 21310 22530 21362 22542
rect 21982 22594 22034 22606
rect 21982 22530 22034 22542
rect 24782 22594 24834 22606
rect 24782 22530 24834 22542
rect 25118 22594 25170 22606
rect 25118 22530 25170 22542
rect 8990 22482 9042 22494
rect 8530 22430 8542 22482
rect 8594 22430 8606 22482
rect 8990 22418 9042 22430
rect 12910 22482 12962 22494
rect 12910 22418 12962 22430
rect 13806 22482 13858 22494
rect 13806 22418 13858 22430
rect 14254 22482 14306 22494
rect 14254 22418 14306 22430
rect 15150 22482 15202 22494
rect 15150 22418 15202 22430
rect 20190 22482 20242 22494
rect 20190 22418 20242 22430
rect 27358 22482 27410 22494
rect 27358 22418 27410 22430
rect 29262 22482 29314 22494
rect 35086 22482 35138 22494
rect 31714 22430 31726 22482
rect 31778 22430 31790 22482
rect 33842 22430 33854 22482
rect 33906 22430 33918 22482
rect 29262 22418 29314 22430
rect 35086 22418 35138 22430
rect 35982 22482 36034 22494
rect 35982 22418 36034 22430
rect 37438 22482 37490 22494
rect 42926 22482 42978 22494
rect 42466 22430 42478 22482
rect 42530 22430 42542 22482
rect 37438 22418 37490 22430
rect 42926 22418 42978 22430
rect 43374 22482 43426 22494
rect 43374 22418 43426 22430
rect 11118 22370 11170 22382
rect 17390 22370 17442 22382
rect 5730 22318 5742 22370
rect 5794 22318 5806 22370
rect 15698 22318 15710 22370
rect 15762 22318 15774 22370
rect 11118 22306 11170 22318
rect 17390 22306 17442 22318
rect 19070 22370 19122 22382
rect 19070 22306 19122 22318
rect 23438 22370 23490 22382
rect 23438 22306 23490 22318
rect 23662 22370 23714 22382
rect 23662 22306 23714 22318
rect 24222 22370 24274 22382
rect 29038 22370 29090 22382
rect 25106 22318 25118 22370
rect 25170 22318 25182 22370
rect 24222 22306 24274 22318
rect 29038 22306 29090 22318
rect 29374 22370 29426 22382
rect 29374 22306 29426 22318
rect 29598 22370 29650 22382
rect 35646 22370 35698 22382
rect 31042 22318 31054 22370
rect 31106 22318 31118 22370
rect 36978 22318 36990 22370
rect 37042 22318 37054 22370
rect 39666 22318 39678 22370
rect 39730 22318 39742 22370
rect 29598 22306 29650 22318
rect 35646 22306 35698 22318
rect 11678 22258 11730 22270
rect 18286 22258 18338 22270
rect 6402 22206 6414 22258
rect 6466 22206 6478 22258
rect 16818 22206 16830 22258
rect 16882 22206 16894 22258
rect 11678 22194 11730 22206
rect 18286 22194 18338 22206
rect 21534 22258 21586 22270
rect 21534 22194 21586 22206
rect 22206 22258 22258 22270
rect 22206 22194 22258 22206
rect 23102 22258 23154 22270
rect 23102 22194 23154 22206
rect 23998 22258 24050 22270
rect 23998 22194 24050 22206
rect 35310 22258 35362 22270
rect 35310 22194 35362 22206
rect 35870 22258 35922 22270
rect 35870 22194 35922 22206
rect 37550 22258 37602 22270
rect 37550 22194 37602 22206
rect 37886 22258 37938 22270
rect 40338 22206 40350 22258
rect 40402 22206 40414 22258
rect 37886 22194 37938 22206
rect 19630 22146 19682 22158
rect 21422 22146 21474 22158
rect 14578 22094 14590 22146
rect 14642 22094 14654 22146
rect 20738 22094 20750 22146
rect 20802 22094 20814 22146
rect 19630 22082 19682 22094
rect 21422 22082 21474 22094
rect 22094 22146 22146 22158
rect 22094 22082 22146 22094
rect 22878 22146 22930 22158
rect 22878 22082 22930 22094
rect 23214 22146 23266 22158
rect 23214 22082 23266 22094
rect 23886 22146 23938 22158
rect 23886 22082 23938 22094
rect 25566 22146 25618 22158
rect 25566 22082 25618 22094
rect 34302 22146 34354 22158
rect 34302 22082 34354 22094
rect 35422 22146 35474 22158
rect 35422 22082 35474 22094
rect 36094 22146 36146 22158
rect 36094 22082 36146 22094
rect 36318 22146 36370 22158
rect 36318 22082 36370 22094
rect 37326 22146 37378 22158
rect 37326 22082 37378 22094
rect 37998 22146 38050 22158
rect 37998 22082 38050 22094
rect 38222 22146 38274 22158
rect 38222 22082 38274 22094
rect 42814 22146 42866 22158
rect 42814 22082 42866 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 5854 21810 5906 21822
rect 5854 21746 5906 21758
rect 6750 21810 6802 21822
rect 6750 21746 6802 21758
rect 7310 21810 7362 21822
rect 28030 21810 28082 21822
rect 21074 21758 21086 21810
rect 21138 21758 21150 21810
rect 21970 21758 21982 21810
rect 22034 21758 22046 21810
rect 7310 21746 7362 21758
rect 28030 21746 28082 21758
rect 28590 21810 28642 21822
rect 40238 21810 40290 21822
rect 35186 21758 35198 21810
rect 35250 21758 35262 21810
rect 28590 21746 28642 21758
rect 40238 21746 40290 21758
rect 6526 21698 6578 21710
rect 6066 21646 6078 21698
rect 6130 21695 6142 21698
rect 6402 21695 6414 21698
rect 6130 21649 6414 21695
rect 6130 21646 6142 21649
rect 6402 21646 6414 21649
rect 6466 21646 6478 21698
rect 6526 21634 6578 21646
rect 7534 21698 7586 21710
rect 20526 21698 20578 21710
rect 29486 21698 29538 21710
rect 11330 21646 11342 21698
rect 11394 21646 11406 21698
rect 17490 21646 17502 21698
rect 17554 21646 17566 21698
rect 21858 21646 21870 21698
rect 21922 21646 21934 21698
rect 7534 21634 7586 21646
rect 20526 21634 20578 21646
rect 29486 21634 29538 21646
rect 33182 21698 33234 21710
rect 33182 21634 33234 21646
rect 33854 21698 33906 21710
rect 33854 21634 33906 21646
rect 39342 21698 39394 21710
rect 39342 21634 39394 21646
rect 5966 21586 6018 21598
rect 16606 21586 16658 21598
rect 27918 21586 27970 21598
rect 5618 21534 5630 21586
rect 5682 21534 5694 21586
rect 10210 21534 10222 21586
rect 10274 21534 10286 21586
rect 12114 21534 12126 21586
rect 12178 21534 12190 21586
rect 15922 21534 15934 21586
rect 15986 21534 15998 21586
rect 17378 21534 17390 21586
rect 17442 21534 17454 21586
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 21970 21534 21982 21586
rect 22034 21534 22046 21586
rect 22642 21534 22654 21586
rect 22706 21534 22718 21586
rect 23986 21534 23998 21586
rect 24050 21534 24062 21586
rect 24658 21534 24670 21586
rect 24722 21534 24734 21586
rect 5966 21522 6018 21534
rect 16606 21522 16658 21534
rect 27918 21522 27970 21534
rect 29374 21586 29426 21598
rect 29374 21522 29426 21534
rect 29710 21586 29762 21598
rect 29710 21522 29762 21534
rect 32286 21586 32338 21598
rect 32286 21522 32338 21534
rect 33518 21586 33570 21598
rect 33518 21522 33570 21534
rect 34638 21586 34690 21598
rect 39790 21586 39842 21598
rect 35746 21534 35758 21586
rect 35810 21534 35822 21586
rect 34638 21522 34690 21534
rect 39790 21522 39842 21534
rect 40126 21586 40178 21598
rect 40126 21522 40178 21534
rect 40350 21586 40402 21598
rect 40898 21534 40910 21586
rect 40962 21534 40974 21586
rect 40350 21522 40402 21534
rect 12574 21474 12626 21486
rect 16382 21474 16434 21486
rect 23774 21474 23826 21486
rect 7186 21422 7198 21474
rect 7250 21422 7262 21474
rect 13010 21422 13022 21474
rect 13074 21422 13086 21474
rect 15138 21422 15150 21474
rect 15202 21422 15214 21474
rect 22978 21422 22990 21474
rect 23042 21422 23054 21474
rect 12574 21410 12626 21422
rect 16382 21410 16434 21422
rect 23774 21410 23826 21422
rect 25342 21474 25394 21486
rect 25342 21410 25394 21422
rect 30046 21474 30098 21486
rect 30046 21410 30098 21422
rect 34414 21474 34466 21486
rect 44270 21474 44322 21486
rect 36530 21422 36542 21474
rect 36594 21422 36606 21474
rect 38658 21422 38670 21474
rect 38722 21422 38734 21474
rect 39442 21422 39454 21474
rect 39506 21422 39518 21474
rect 41682 21422 41694 21474
rect 41746 21422 41758 21474
rect 43810 21422 43822 21474
rect 43874 21422 43886 21474
rect 34414 21410 34466 21422
rect 44270 21410 44322 21422
rect 6862 21362 6914 21374
rect 6862 21298 6914 21310
rect 16270 21362 16322 21374
rect 16270 21298 16322 21310
rect 16718 21362 16770 21374
rect 16718 21298 16770 21310
rect 23662 21362 23714 21374
rect 23662 21298 23714 21310
rect 24334 21362 24386 21374
rect 24334 21298 24386 21310
rect 24670 21362 24722 21374
rect 24670 21298 24722 21310
rect 28030 21362 28082 21374
rect 28030 21298 28082 21310
rect 33070 21362 33122 21374
rect 33070 21298 33122 21310
rect 34862 21362 34914 21374
rect 34862 21298 34914 21310
rect 39118 21362 39170 21374
rect 39118 21298 39170 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 6302 21026 6354 21038
rect 6302 20962 6354 20974
rect 14926 20914 14978 20926
rect 19182 20914 19234 20926
rect 37102 20914 37154 20926
rect 10770 20862 10782 20914
rect 10834 20862 10846 20914
rect 12450 20862 12462 20914
rect 12514 20862 12526 20914
rect 13570 20862 13582 20914
rect 13634 20862 13646 20914
rect 15586 20862 15598 20914
rect 15650 20862 15662 20914
rect 20514 20862 20526 20914
rect 20578 20862 20590 20914
rect 25330 20862 25342 20914
rect 25394 20862 25406 20914
rect 28578 20862 28590 20914
rect 28642 20862 28654 20914
rect 32050 20862 32062 20914
rect 32114 20862 32126 20914
rect 35634 20862 35646 20914
rect 35698 20862 35710 20914
rect 14926 20850 14978 20862
rect 19182 20850 19234 20862
rect 37102 20850 37154 20862
rect 37998 20914 38050 20926
rect 37998 20850 38050 20862
rect 39678 20914 39730 20926
rect 39678 20850 39730 20862
rect 40574 20914 40626 20926
rect 40574 20850 40626 20862
rect 42366 20914 42418 20926
rect 42366 20850 42418 20862
rect 14030 20802 14082 20814
rect 6626 20750 6638 20802
rect 6690 20750 6702 20802
rect 7970 20750 7982 20802
rect 8034 20750 8046 20802
rect 12562 20750 12574 20802
rect 12626 20750 12638 20802
rect 14030 20738 14082 20750
rect 14366 20802 14418 20814
rect 14366 20738 14418 20750
rect 16606 20802 16658 20814
rect 17502 20802 17554 20814
rect 36430 20802 36482 20814
rect 16930 20750 16942 20802
rect 16994 20750 17006 20802
rect 20402 20750 20414 20802
rect 20466 20750 20478 20802
rect 22418 20750 22430 20802
rect 22482 20750 22494 20802
rect 25666 20750 25678 20802
rect 25730 20750 25742 20802
rect 29250 20750 29262 20802
rect 29314 20750 29326 20802
rect 32610 20750 32622 20802
rect 32674 20750 32686 20802
rect 33282 20750 33294 20802
rect 33346 20750 33358 20802
rect 16606 20738 16658 20750
rect 17502 20738 17554 20750
rect 36430 20738 36482 20750
rect 36878 20802 36930 20814
rect 36878 20738 36930 20750
rect 39006 20802 39058 20814
rect 39006 20738 39058 20750
rect 40126 20802 40178 20814
rect 40126 20738 40178 20750
rect 40462 20802 40514 20814
rect 40462 20738 40514 20750
rect 11454 20690 11506 20702
rect 8642 20638 8654 20690
rect 8706 20638 8718 20690
rect 11454 20626 11506 20638
rect 11790 20690 11842 20702
rect 16718 20690 16770 20702
rect 15362 20638 15374 20690
rect 15426 20638 15438 20690
rect 11790 20626 11842 20638
rect 16718 20626 16770 20638
rect 18398 20690 18450 20702
rect 18398 20626 18450 20638
rect 21870 20690 21922 20702
rect 21870 20626 21922 20638
rect 21982 20690 22034 20702
rect 37326 20690 37378 20702
rect 23202 20638 23214 20690
rect 23266 20638 23278 20690
rect 26450 20638 26462 20690
rect 26514 20638 26526 20690
rect 29922 20638 29934 20690
rect 29986 20638 29998 20690
rect 21982 20626 22034 20638
rect 37326 20626 37378 20638
rect 37550 20690 37602 20702
rect 37550 20626 37602 20638
rect 38334 20690 38386 20702
rect 38334 20626 38386 20638
rect 38446 20690 38498 20702
rect 38446 20626 38498 20638
rect 38670 20690 38722 20702
rect 38670 20626 38722 20638
rect 39790 20690 39842 20702
rect 39790 20626 39842 20638
rect 40686 20690 40738 20702
rect 40686 20626 40738 20638
rect 42254 20690 42306 20702
rect 42254 20626 42306 20638
rect 6414 20578 6466 20590
rect 6414 20514 6466 20526
rect 11230 20578 11282 20590
rect 11230 20514 11282 20526
rect 11342 20578 11394 20590
rect 11342 20514 11394 20526
rect 18958 20578 19010 20590
rect 18958 20514 19010 20526
rect 21534 20578 21586 20590
rect 21534 20514 21586 20526
rect 22206 20578 22258 20590
rect 36094 20578 36146 20590
rect 32386 20526 32398 20578
rect 32450 20526 32462 20578
rect 22206 20514 22258 20526
rect 36094 20514 36146 20526
rect 36318 20578 36370 20590
rect 36318 20514 36370 20526
rect 37886 20578 37938 20590
rect 37886 20514 37938 20526
rect 39566 20578 39618 20590
rect 39566 20514 39618 20526
rect 41246 20578 41298 20590
rect 41246 20514 41298 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 13358 20242 13410 20254
rect 13358 20178 13410 20190
rect 16718 20242 16770 20254
rect 16718 20178 16770 20190
rect 19742 20242 19794 20254
rect 27582 20242 27634 20254
rect 27234 20190 27246 20242
rect 27298 20190 27310 20242
rect 19742 20178 19794 20190
rect 27582 20178 27634 20190
rect 28030 20242 28082 20254
rect 28030 20178 28082 20190
rect 29374 20242 29426 20254
rect 29374 20178 29426 20190
rect 29486 20242 29538 20254
rect 29486 20178 29538 20190
rect 40238 20242 40290 20254
rect 40238 20178 40290 20190
rect 11006 20130 11058 20142
rect 11006 20066 11058 20078
rect 13134 20130 13186 20142
rect 13134 20066 13186 20078
rect 13470 20130 13522 20142
rect 13470 20066 13522 20078
rect 15822 20130 15874 20142
rect 15822 20066 15874 20078
rect 18398 20130 18450 20142
rect 18398 20066 18450 20078
rect 24222 20130 24274 20142
rect 24222 20066 24274 20078
rect 24670 20130 24722 20142
rect 24670 20066 24722 20078
rect 25566 20130 25618 20142
rect 25566 20066 25618 20078
rect 27694 20130 27746 20142
rect 27694 20066 27746 20078
rect 28590 20130 28642 20142
rect 28590 20066 28642 20078
rect 30942 20130 30994 20142
rect 30942 20066 30994 20078
rect 31278 20130 31330 20142
rect 31278 20066 31330 20078
rect 31614 20130 31666 20142
rect 31614 20066 31666 20078
rect 31950 20130 32002 20142
rect 31950 20066 32002 20078
rect 32286 20130 32338 20142
rect 36766 20130 36818 20142
rect 35074 20078 35086 20130
rect 35138 20078 35150 20130
rect 32286 20066 32338 20078
rect 36766 20066 36818 20078
rect 37662 20130 37714 20142
rect 37662 20066 37714 20078
rect 38670 20130 38722 20142
rect 38670 20066 38722 20078
rect 38782 20130 38834 20142
rect 38782 20066 38834 20078
rect 39678 20130 39730 20142
rect 39678 20066 39730 20078
rect 40014 20130 40066 20142
rect 40014 20066 40066 20078
rect 15038 20018 15090 20030
rect 12338 19966 12350 20018
rect 12402 19966 12414 20018
rect 15038 19954 15090 19966
rect 16718 20018 16770 20030
rect 23662 20018 23714 20030
rect 17378 19966 17390 20018
rect 17442 19966 17454 20018
rect 20402 19966 20414 20018
rect 20466 19966 20478 20018
rect 16718 19954 16770 19966
rect 23662 19954 23714 19966
rect 23998 20018 24050 20030
rect 23998 19954 24050 19966
rect 24446 20018 24498 20030
rect 24446 19954 24498 19966
rect 25454 20018 25506 20030
rect 25454 19954 25506 19966
rect 27806 20018 27858 20030
rect 27806 19954 27858 19966
rect 29598 20018 29650 20030
rect 29598 19954 29650 19966
rect 30046 20018 30098 20030
rect 30046 19954 30098 19966
rect 30830 20018 30882 20030
rect 30830 19954 30882 19966
rect 33070 20018 33122 20030
rect 33070 19954 33122 19966
rect 34190 20018 34242 20030
rect 35870 20018 35922 20030
rect 35298 19966 35310 20018
rect 35362 19966 35374 20018
rect 34190 19954 34242 19966
rect 35870 19954 35922 19966
rect 36206 20018 36258 20030
rect 36206 19954 36258 19966
rect 36542 20018 36594 20030
rect 36542 19954 36594 19966
rect 39006 20018 39058 20030
rect 41122 19966 41134 20018
rect 41186 19966 41198 20018
rect 39006 19954 39058 19966
rect 12910 19906 12962 19918
rect 12114 19854 12126 19906
rect 12178 19854 12190 19906
rect 12910 19842 12962 19854
rect 19182 19906 19234 19918
rect 26350 19906 26402 19918
rect 21074 19854 21086 19906
rect 21138 19854 21150 19906
rect 23202 19854 23214 19906
rect 23266 19854 23278 19906
rect 19182 19842 19234 19854
rect 26350 19842 26402 19854
rect 26686 19906 26738 19918
rect 26686 19842 26738 19854
rect 26910 19906 26962 19918
rect 26910 19842 26962 19854
rect 28478 19906 28530 19918
rect 36654 19906 36706 19918
rect 33506 19854 33518 19906
rect 33570 19854 33582 19906
rect 34626 19854 34638 19906
rect 34690 19854 34702 19906
rect 28478 19842 28530 19854
rect 36654 19842 36706 19854
rect 37214 19906 37266 19918
rect 37214 19842 37266 19854
rect 38334 19906 38386 19918
rect 40226 19854 40238 19906
rect 40290 19854 40302 19906
rect 42242 19854 42254 19906
rect 42306 19854 42318 19906
rect 38334 19842 38386 19854
rect 23550 19794 23602 19806
rect 23550 19730 23602 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 12126 19458 12178 19470
rect 12126 19394 12178 19406
rect 12462 19458 12514 19470
rect 32834 19406 32846 19458
rect 32898 19455 32910 19458
rect 33506 19455 33518 19458
rect 32898 19409 33518 19455
rect 32898 19406 32910 19409
rect 33506 19406 33518 19409
rect 33570 19406 33582 19458
rect 12462 19394 12514 19406
rect 10670 19346 10722 19358
rect 8082 19294 8094 19346
rect 8146 19294 8158 19346
rect 10210 19294 10222 19346
rect 10274 19294 10286 19346
rect 10670 19282 10722 19294
rect 16158 19346 16210 19358
rect 16158 19282 16210 19294
rect 19518 19346 19570 19358
rect 19518 19282 19570 19294
rect 20750 19346 20802 19358
rect 20750 19282 20802 19294
rect 22094 19346 22146 19358
rect 22094 19282 22146 19294
rect 23998 19346 24050 19358
rect 23998 19282 24050 19294
rect 33406 19346 33458 19358
rect 33406 19282 33458 19294
rect 35982 19346 36034 19358
rect 37762 19294 37774 19346
rect 37826 19294 37838 19346
rect 39890 19294 39902 19346
rect 39954 19294 39966 19346
rect 42802 19294 42814 19346
rect 42866 19294 42878 19346
rect 35982 19282 36034 19294
rect 14478 19234 14530 19246
rect 21646 19234 21698 19246
rect 7410 19182 7422 19234
rect 7474 19182 7486 19234
rect 12114 19182 12126 19234
rect 12178 19182 12190 19234
rect 15026 19182 15038 19234
rect 15090 19182 15102 19234
rect 17714 19182 17726 19234
rect 17778 19182 17790 19234
rect 14478 19170 14530 19182
rect 21646 19170 21698 19182
rect 21982 19234 22034 19246
rect 21982 19170 22034 19182
rect 22318 19234 22370 19246
rect 22318 19170 22370 19182
rect 22542 19234 22594 19246
rect 29934 19234 29986 19246
rect 22866 19182 22878 19234
rect 22930 19182 22942 19234
rect 27570 19182 27582 19234
rect 27634 19182 27646 19234
rect 22542 19170 22594 19182
rect 29934 19170 29986 19182
rect 33742 19234 33794 19246
rect 33742 19170 33794 19182
rect 35086 19234 35138 19246
rect 35746 19182 35758 19234
rect 35810 19182 35822 19234
rect 37090 19182 37102 19234
rect 37154 19182 37166 19234
rect 41010 19182 41022 19234
rect 41074 19182 41086 19234
rect 35086 19170 35138 19182
rect 18286 19122 18338 19134
rect 24446 19122 24498 19134
rect 15250 19070 15262 19122
rect 15314 19070 15326 19122
rect 22978 19070 22990 19122
rect 23042 19070 23054 19122
rect 18286 19058 18338 19070
rect 24446 19058 24498 19070
rect 32958 19122 33010 19134
rect 32958 19058 33010 19070
rect 34526 19122 34578 19134
rect 34526 19058 34578 19070
rect 34750 19122 34802 19134
rect 36094 19122 36146 19134
rect 35410 19070 35422 19122
rect 35474 19070 35486 19122
rect 34750 19058 34802 19070
rect 36094 19058 36146 19070
rect 43486 19122 43538 19134
rect 43486 19058 43538 19070
rect 14142 19010 14194 19022
rect 26126 19010 26178 19022
rect 19618 18958 19630 19010
rect 19682 18958 19694 19010
rect 21298 18958 21310 19010
rect 21362 18958 21374 19010
rect 23426 18958 23438 19010
rect 23490 18958 23502 19010
rect 14142 18946 14194 18958
rect 26126 18946 26178 18958
rect 27358 19010 27410 19022
rect 27358 18946 27410 18958
rect 29598 19010 29650 19022
rect 29598 18946 29650 18958
rect 29822 19010 29874 19022
rect 34638 19010 34690 19022
rect 34066 18958 34078 19010
rect 34130 18958 34142 19010
rect 29822 18946 29874 18958
rect 34638 18946 34690 18958
rect 43374 19010 43426 19022
rect 43374 18946 43426 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 22542 18674 22594 18686
rect 22542 18610 22594 18622
rect 26350 18674 26402 18686
rect 26350 18610 26402 18622
rect 32398 18674 32450 18686
rect 32398 18610 32450 18622
rect 35422 18674 35474 18686
rect 35422 18610 35474 18622
rect 35870 18674 35922 18686
rect 35870 18610 35922 18622
rect 38782 18674 38834 18686
rect 38782 18610 38834 18622
rect 44270 18674 44322 18686
rect 44270 18610 44322 18622
rect 18510 18562 18562 18574
rect 23662 18562 23714 18574
rect 11778 18510 11790 18562
rect 11842 18510 11854 18562
rect 17490 18510 17502 18562
rect 17554 18510 17566 18562
rect 23314 18510 23326 18562
rect 23378 18510 23390 18562
rect 18510 18498 18562 18510
rect 23662 18498 23714 18510
rect 24670 18562 24722 18574
rect 24670 18498 24722 18510
rect 25230 18562 25282 18574
rect 25230 18498 25282 18510
rect 27358 18562 27410 18574
rect 27358 18498 27410 18510
rect 27470 18562 27522 18574
rect 27470 18498 27522 18510
rect 27806 18562 27858 18574
rect 27806 18498 27858 18510
rect 29262 18562 29314 18574
rect 29262 18498 29314 18510
rect 32510 18562 32562 18574
rect 32510 18498 32562 18510
rect 33294 18562 33346 18574
rect 33294 18498 33346 18510
rect 39118 18562 39170 18574
rect 39118 18498 39170 18510
rect 39790 18562 39842 18574
rect 39790 18498 39842 18510
rect 9662 18450 9714 18462
rect 17838 18450 17890 18462
rect 23998 18450 24050 18462
rect 6066 18398 6078 18450
rect 6130 18398 6142 18450
rect 6738 18398 6750 18450
rect 6802 18398 6814 18450
rect 11890 18398 11902 18450
rect 11954 18398 11966 18450
rect 12338 18398 12350 18450
rect 12402 18398 12414 18450
rect 18274 18398 18286 18450
rect 18338 18398 18350 18450
rect 18834 18398 18846 18450
rect 18898 18398 18910 18450
rect 23090 18398 23102 18450
rect 23154 18398 23166 18450
rect 9662 18386 9714 18398
rect 17838 18386 17890 18398
rect 23998 18386 24050 18398
rect 24334 18450 24386 18462
rect 24334 18386 24386 18398
rect 25566 18450 25618 18462
rect 26574 18450 26626 18462
rect 26002 18398 26014 18450
rect 26066 18398 26078 18450
rect 25566 18386 25618 18398
rect 26574 18386 26626 18398
rect 27022 18450 27074 18462
rect 27022 18386 27074 18398
rect 28030 18450 28082 18462
rect 28030 18386 28082 18398
rect 28366 18450 28418 18462
rect 28366 18386 28418 18398
rect 28814 18450 28866 18462
rect 28814 18386 28866 18398
rect 29038 18450 29090 18462
rect 29038 18386 29090 18398
rect 29710 18450 29762 18462
rect 29710 18386 29762 18398
rect 29822 18450 29874 18462
rect 29822 18386 29874 18398
rect 30270 18450 30322 18462
rect 30270 18386 30322 18398
rect 30494 18450 30546 18462
rect 30494 18386 30546 18398
rect 30718 18450 30770 18462
rect 30718 18386 30770 18398
rect 31166 18450 31218 18462
rect 31166 18386 31218 18398
rect 33070 18450 33122 18462
rect 33070 18386 33122 18398
rect 33630 18450 33682 18462
rect 33630 18386 33682 18398
rect 34414 18450 34466 18462
rect 34414 18386 34466 18398
rect 34638 18450 34690 18462
rect 34638 18386 34690 18398
rect 35086 18450 35138 18462
rect 35086 18386 35138 18398
rect 36094 18450 36146 18462
rect 36094 18386 36146 18398
rect 38110 18450 38162 18462
rect 40014 18450 40066 18462
rect 39442 18398 39454 18450
rect 39506 18398 39518 18450
rect 38110 18386 38162 18398
rect 40014 18386 40066 18398
rect 40350 18450 40402 18462
rect 40898 18398 40910 18450
rect 40962 18398 40974 18450
rect 40350 18386 40402 18398
rect 15710 18338 15762 18350
rect 25342 18338 25394 18350
rect 8866 18286 8878 18338
rect 8930 18286 8942 18338
rect 13122 18286 13134 18338
rect 13186 18286 13198 18338
rect 15250 18286 15262 18338
rect 15314 18286 15326 18338
rect 19618 18286 19630 18338
rect 19682 18286 19694 18338
rect 21746 18286 21758 18338
rect 21810 18286 21822 18338
rect 15710 18274 15762 18286
rect 25342 18274 25394 18286
rect 26462 18338 26514 18350
rect 26462 18274 26514 18286
rect 27918 18338 27970 18350
rect 27918 18274 27970 18286
rect 29150 18338 29202 18350
rect 29150 18274 29202 18286
rect 30046 18338 30098 18350
rect 30046 18274 30098 18286
rect 30942 18338 30994 18350
rect 30942 18274 30994 18286
rect 33518 18338 33570 18350
rect 33518 18274 33570 18286
rect 34862 18338 34914 18350
rect 34862 18274 34914 18286
rect 35982 18338 36034 18350
rect 35982 18274 36034 18286
rect 37998 18338 38050 18350
rect 37998 18274 38050 18286
rect 39902 18338 39954 18350
rect 41682 18286 41694 18338
rect 41746 18286 41758 18338
rect 43810 18286 43822 18338
rect 43874 18286 43886 18338
rect 39902 18274 39954 18286
rect 10782 18226 10834 18238
rect 10782 18162 10834 18174
rect 11118 18226 11170 18238
rect 11118 18162 11170 18174
rect 25678 18226 25730 18238
rect 25678 18162 25730 18174
rect 27358 18226 27410 18238
rect 27358 18162 27410 18174
rect 32398 18226 32450 18238
rect 32398 18162 32450 18174
rect 39454 18226 39506 18238
rect 39454 18162 39506 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 14478 17890 14530 17902
rect 14478 17826 14530 17838
rect 19294 17890 19346 17902
rect 19294 17826 19346 17838
rect 24782 17890 24834 17902
rect 24782 17826 24834 17838
rect 36094 17890 36146 17902
rect 36094 17826 36146 17838
rect 12014 17778 12066 17790
rect 11330 17726 11342 17778
rect 11394 17726 11406 17778
rect 12014 17714 12066 17726
rect 12462 17778 12514 17790
rect 18846 17778 18898 17790
rect 36206 17778 36258 17790
rect 18274 17726 18286 17778
rect 18338 17726 18350 17778
rect 21522 17726 21534 17778
rect 21586 17726 21598 17778
rect 27794 17726 27806 17778
rect 27858 17726 27870 17778
rect 12462 17714 12514 17726
rect 18846 17714 18898 17726
rect 36206 17714 36258 17726
rect 39006 17778 39058 17790
rect 40562 17726 40574 17778
rect 40626 17726 40638 17778
rect 42690 17726 42702 17778
rect 42754 17726 42766 17778
rect 39006 17714 39058 17726
rect 13806 17666 13858 17678
rect 19630 17666 19682 17678
rect 25902 17666 25954 17678
rect 7858 17614 7870 17666
rect 7922 17614 7934 17666
rect 8418 17614 8430 17666
rect 8482 17614 8494 17666
rect 15474 17614 15486 17666
rect 15538 17614 15550 17666
rect 23874 17614 23886 17666
rect 23938 17614 23950 17666
rect 24770 17614 24782 17666
rect 24834 17614 24846 17666
rect 13806 17602 13858 17614
rect 19630 17602 19682 17614
rect 25902 17602 25954 17614
rect 27022 17666 27074 17678
rect 27022 17602 27074 17614
rect 29486 17666 29538 17678
rect 29486 17602 29538 17614
rect 32846 17666 32898 17678
rect 32846 17602 32898 17614
rect 33518 17666 33570 17678
rect 33518 17602 33570 17614
rect 34078 17666 34130 17678
rect 34078 17602 34130 17614
rect 35086 17666 35138 17678
rect 35086 17602 35138 17614
rect 35534 17666 35586 17678
rect 35534 17602 35586 17614
rect 36878 17666 36930 17678
rect 36878 17602 36930 17614
rect 37438 17666 37490 17678
rect 37438 17602 37490 17614
rect 38894 17666 38946 17678
rect 38894 17602 38946 17614
rect 39118 17666 39170 17678
rect 39118 17602 39170 17614
rect 39454 17666 39506 17678
rect 39890 17614 39902 17666
rect 39954 17614 39966 17666
rect 39454 17602 39506 17614
rect 13470 17554 13522 17566
rect 24446 17554 24498 17566
rect 9202 17502 9214 17554
rect 9266 17502 9278 17554
rect 16146 17502 16158 17554
rect 16210 17502 16222 17554
rect 19842 17502 19854 17554
rect 19906 17502 19918 17554
rect 20178 17502 20190 17554
rect 20242 17502 20254 17554
rect 13470 17490 13522 17502
rect 24446 17490 24498 17502
rect 26238 17554 26290 17566
rect 27358 17554 27410 17566
rect 29822 17554 29874 17566
rect 33294 17554 33346 17566
rect 26338 17502 26350 17554
rect 26402 17502 26414 17554
rect 27458 17502 27470 17554
rect 27522 17502 27534 17554
rect 31042 17502 31054 17554
rect 31106 17502 31118 17554
rect 32050 17502 32062 17554
rect 32114 17502 32126 17554
rect 26238 17490 26290 17502
rect 27358 17490 27410 17502
rect 29822 17490 29874 17502
rect 33294 17490 33346 17502
rect 34526 17554 34578 17566
rect 34526 17490 34578 17502
rect 35198 17554 35250 17566
rect 35198 17490 35250 17502
rect 36318 17554 36370 17566
rect 36318 17490 36370 17502
rect 37326 17554 37378 17566
rect 37326 17490 37378 17502
rect 8094 17442 8146 17454
rect 8094 17378 8146 17390
rect 14590 17442 14642 17454
rect 14590 17378 14642 17390
rect 14702 17442 14754 17454
rect 14702 17378 14754 17390
rect 25230 17442 25282 17454
rect 26014 17442 26066 17454
rect 25554 17390 25566 17442
rect 25618 17390 25630 17442
rect 25230 17378 25282 17390
rect 26014 17378 26066 17390
rect 26126 17442 26178 17454
rect 26126 17378 26178 17390
rect 27246 17442 27298 17454
rect 27246 17378 27298 17390
rect 31390 17442 31442 17454
rect 31390 17378 31442 17390
rect 31726 17442 31778 17454
rect 31726 17378 31778 17390
rect 33182 17442 33234 17454
rect 33182 17378 33234 17390
rect 33742 17442 33794 17454
rect 33742 17378 33794 17390
rect 33966 17442 34018 17454
rect 33966 17378 34018 17390
rect 34414 17442 34466 17454
rect 34414 17378 34466 17390
rect 35310 17442 35362 17454
rect 35310 17378 35362 17390
rect 37102 17442 37154 17454
rect 37102 17378 37154 17390
rect 43150 17442 43202 17454
rect 43150 17378 43202 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 9550 17106 9602 17118
rect 9550 17042 9602 17054
rect 16494 17106 16546 17118
rect 16494 17042 16546 17054
rect 20974 17106 21026 17118
rect 20974 17042 21026 17054
rect 22094 17106 22146 17118
rect 26350 17106 26402 17118
rect 22754 17054 22766 17106
rect 22818 17054 22830 17106
rect 22094 17042 22146 17054
rect 26350 17042 26402 17054
rect 28030 17106 28082 17118
rect 28030 17042 28082 17054
rect 29710 17106 29762 17118
rect 39678 17106 39730 17118
rect 30370 17054 30382 17106
rect 30434 17054 30446 17106
rect 29710 17042 29762 17054
rect 39678 17042 39730 17054
rect 16830 16994 16882 17006
rect 16830 16930 16882 16942
rect 17502 16994 17554 17006
rect 21310 16994 21362 17006
rect 18386 16942 18398 16994
rect 18450 16942 18462 16994
rect 19170 16942 19182 16994
rect 19234 16942 19246 16994
rect 19618 16942 19630 16994
rect 19682 16942 19694 16994
rect 17502 16930 17554 16942
rect 21310 16930 21362 16942
rect 22542 16994 22594 17006
rect 22542 16930 22594 16942
rect 26574 16994 26626 17006
rect 26574 16930 26626 16942
rect 27022 16994 27074 17006
rect 27022 16930 27074 16942
rect 27806 16994 27858 17006
rect 27806 16930 27858 16942
rect 28254 16994 28306 17006
rect 31054 16994 31106 17006
rect 30034 16942 30046 16994
rect 30098 16942 30110 16994
rect 28254 16930 28306 16942
rect 31054 16930 31106 16942
rect 31390 16994 31442 17006
rect 42030 16994 42082 17006
rect 32162 16942 32174 16994
rect 32226 16942 32238 16994
rect 33842 16942 33854 16994
rect 33906 16942 33918 16994
rect 37090 16942 37102 16994
rect 37154 16942 37166 16994
rect 31390 16930 31442 16942
rect 42030 16930 42082 16942
rect 9886 16882 9938 16894
rect 17838 16882 17890 16894
rect 22206 16882 22258 16894
rect 13122 16830 13134 16882
rect 13186 16830 13198 16882
rect 16034 16830 16046 16882
rect 16098 16830 16110 16882
rect 18610 16830 18622 16882
rect 18674 16830 18686 16882
rect 19282 16830 19294 16882
rect 19346 16830 19358 16882
rect 21522 16830 21534 16882
rect 21586 16830 21598 16882
rect 9886 16818 9938 16830
rect 17838 16818 17890 16830
rect 22206 16818 22258 16830
rect 22878 16882 22930 16894
rect 24110 16882 24162 16894
rect 23314 16830 23326 16882
rect 23378 16830 23390 16882
rect 23650 16830 23662 16882
rect 23714 16830 23726 16882
rect 22878 16818 22930 16830
rect 24110 16818 24162 16830
rect 24334 16882 24386 16894
rect 24334 16818 24386 16830
rect 24446 16882 24498 16894
rect 24446 16818 24498 16830
rect 25230 16882 25282 16894
rect 25230 16818 25282 16830
rect 25454 16882 25506 16894
rect 26014 16882 26066 16894
rect 25778 16830 25790 16882
rect 25842 16830 25854 16882
rect 25454 16818 25506 16830
rect 26014 16818 26066 16830
rect 26910 16882 26962 16894
rect 26910 16818 26962 16830
rect 27134 16882 27186 16894
rect 27134 16818 27186 16830
rect 27582 16882 27634 16894
rect 27582 16818 27634 16830
rect 30718 16882 30770 16894
rect 30718 16818 30770 16830
rect 31838 16882 31890 16894
rect 41918 16882 41970 16894
rect 33058 16830 33070 16882
rect 33122 16830 33134 16882
rect 36418 16830 36430 16882
rect 36482 16830 36494 16882
rect 31838 16818 31890 16830
rect 41918 16818 41970 16830
rect 22990 16770 23042 16782
rect 12002 16718 12014 16770
rect 12066 16718 12078 16770
rect 14914 16718 14926 16770
rect 14978 16718 14990 16770
rect 22990 16706 23042 16718
rect 25342 16770 25394 16782
rect 35970 16718 35982 16770
rect 36034 16718 36046 16770
rect 39218 16718 39230 16770
rect 39282 16718 39294 16770
rect 25342 16706 25394 16718
rect 22094 16658 22146 16670
rect 22094 16594 22146 16606
rect 23998 16658 24050 16670
rect 23998 16594 24050 16606
rect 26238 16658 26290 16670
rect 26238 16594 26290 16606
rect 27918 16658 27970 16670
rect 27918 16594 27970 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 11230 16322 11282 16334
rect 11230 16258 11282 16270
rect 11566 16322 11618 16334
rect 11566 16258 11618 16270
rect 14702 16322 14754 16334
rect 14702 16258 14754 16270
rect 16270 16322 16322 16334
rect 16270 16258 16322 16270
rect 12910 16210 12962 16222
rect 8642 16158 8654 16210
rect 8706 16158 8718 16210
rect 10770 16158 10782 16210
rect 10834 16158 10846 16210
rect 12910 16146 12962 16158
rect 16718 16210 16770 16222
rect 30718 16210 30770 16222
rect 22754 16158 22766 16210
rect 22818 16158 22830 16210
rect 16718 16146 16770 16158
rect 30718 16146 30770 16158
rect 38222 16210 38274 16222
rect 38222 16146 38274 16158
rect 18958 16098 19010 16110
rect 7970 16046 7982 16098
rect 8034 16046 8046 16098
rect 15138 16046 15150 16098
rect 15202 16046 15214 16098
rect 18958 16034 19010 16046
rect 19294 16098 19346 16110
rect 24558 16098 24610 16110
rect 25006 16098 25058 16110
rect 23874 16046 23886 16098
rect 23938 16046 23950 16098
rect 24434 16046 24446 16098
rect 24498 16046 24510 16098
rect 24770 16046 24782 16098
rect 24834 16046 24846 16098
rect 19294 16034 19346 16046
rect 24558 16034 24610 16046
rect 25006 16034 25058 16046
rect 29598 16098 29650 16110
rect 34302 16098 34354 16110
rect 31826 16046 31838 16098
rect 31890 16046 31902 16098
rect 29598 16034 29650 16046
rect 34302 16034 34354 16046
rect 34526 16098 34578 16110
rect 34526 16034 34578 16046
rect 34862 16098 34914 16110
rect 34862 16034 34914 16046
rect 13918 15986 13970 15998
rect 11890 15934 11902 15986
rect 11954 15934 11966 15986
rect 12114 15934 12126 15986
rect 12178 15934 12190 15986
rect 13918 15922 13970 15934
rect 14366 15986 14418 15998
rect 15934 15986 15986 15998
rect 15474 15934 15486 15986
rect 15538 15934 15550 15986
rect 14366 15922 14418 15934
rect 15934 15922 15986 15934
rect 16158 15986 16210 15998
rect 16158 15922 16210 15934
rect 13582 15874 13634 15886
rect 13582 15810 13634 15822
rect 18734 15874 18786 15886
rect 18734 15810 18786 15822
rect 19182 15874 19234 15886
rect 25902 15874 25954 15886
rect 24546 15822 24558 15874
rect 24610 15822 24622 15874
rect 19182 15810 19234 15822
rect 25902 15810 25954 15822
rect 29934 15874 29986 15886
rect 34638 15874 34690 15886
rect 32050 15822 32062 15874
rect 32114 15822 32126 15874
rect 29934 15810 29986 15822
rect 34638 15810 34690 15822
rect 36206 15874 36258 15886
rect 36206 15810 36258 15822
rect 38110 15874 38162 15886
rect 38110 15810 38162 15822
rect 43822 15874 43874 15886
rect 43822 15810 43874 15822
rect 44270 15874 44322 15886
rect 44270 15810 44322 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 16046 15538 16098 15550
rect 16046 15474 16098 15486
rect 23326 15538 23378 15550
rect 23326 15474 23378 15486
rect 24222 15538 24274 15550
rect 36542 15538 36594 15550
rect 28466 15486 28478 15538
rect 28530 15486 28542 15538
rect 24222 15474 24274 15486
rect 36542 15474 36594 15486
rect 38782 15538 38834 15550
rect 38782 15474 38834 15486
rect 17614 15426 17666 15438
rect 6738 15374 6750 15426
rect 6802 15374 6814 15426
rect 11890 15374 11902 15426
rect 11954 15374 11966 15426
rect 13458 15374 13470 15426
rect 13522 15374 13534 15426
rect 17614 15362 17666 15374
rect 18398 15426 18450 15438
rect 26126 15426 26178 15438
rect 28030 15426 28082 15438
rect 30158 15426 30210 15438
rect 19282 15374 19294 15426
rect 19346 15374 19358 15426
rect 20738 15374 20750 15426
rect 20802 15374 20814 15426
rect 26450 15374 26462 15426
rect 26514 15374 26526 15426
rect 29922 15374 29934 15426
rect 29986 15374 29998 15426
rect 18398 15362 18450 15374
rect 26126 15362 26178 15374
rect 28030 15362 28082 15374
rect 30158 15362 30210 15374
rect 37326 15426 37378 15438
rect 37326 15362 37378 15374
rect 39678 15426 39730 15438
rect 39678 15362 39730 15374
rect 10558 15314 10610 15326
rect 18734 15314 18786 15326
rect 6066 15262 6078 15314
rect 6130 15262 6142 15314
rect 12002 15262 12014 15314
rect 12066 15262 12078 15314
rect 12786 15262 12798 15314
rect 12850 15262 12862 15314
rect 10558 15250 10610 15262
rect 18734 15250 18786 15262
rect 19630 15314 19682 15326
rect 25230 15314 25282 15326
rect 20066 15262 20078 15314
rect 20130 15262 20142 15314
rect 19630 15250 19682 15262
rect 25230 15250 25282 15262
rect 25454 15314 25506 15326
rect 25454 15250 25506 15262
rect 25790 15314 25842 15326
rect 25790 15250 25842 15262
rect 28366 15314 28418 15326
rect 36990 15314 37042 15326
rect 28802 15262 28814 15314
rect 28866 15262 28878 15314
rect 29586 15262 29598 15314
rect 29650 15262 29662 15314
rect 36530 15262 36542 15314
rect 36594 15262 36606 15314
rect 39442 15262 39454 15314
rect 39506 15262 39518 15314
rect 40898 15262 40910 15314
rect 40962 15262 40974 15314
rect 44258 15262 44270 15314
rect 44322 15262 44334 15314
rect 28366 15250 28418 15262
rect 36990 15250 37042 15262
rect 9662 15202 9714 15214
rect 8866 15150 8878 15202
rect 8930 15150 8942 15202
rect 9662 15138 9714 15150
rect 11342 15202 11394 15214
rect 17390 15202 17442 15214
rect 25342 15202 25394 15214
rect 15586 15150 15598 15202
rect 15650 15150 15662 15202
rect 22866 15150 22878 15202
rect 22930 15150 22942 15202
rect 11342 15138 11394 15150
rect 17390 15138 17442 15150
rect 25342 15138 25394 15150
rect 30046 15202 30098 15214
rect 38658 15150 38670 15202
rect 38722 15150 38734 15202
rect 41682 15150 41694 15202
rect 41746 15150 41758 15202
rect 43810 15150 43822 15202
rect 43874 15150 43886 15202
rect 44930 15150 44942 15202
rect 44994 15150 45006 15202
rect 47058 15150 47070 15202
rect 47122 15150 47134 15202
rect 30046 15138 30098 15150
rect 11006 15090 11058 15102
rect 11006 15026 11058 15038
rect 17726 15090 17778 15102
rect 36878 15090 36930 15102
rect 28578 15038 28590 15090
rect 28642 15038 28654 15090
rect 29586 15038 29598 15090
rect 29650 15038 29662 15090
rect 36082 15038 36094 15090
rect 36146 15087 36158 15090
rect 36418 15087 36430 15090
rect 36146 15041 36430 15087
rect 36146 15038 36158 15041
rect 36418 15038 36430 15041
rect 36482 15038 36494 15090
rect 17726 15026 17778 15038
rect 36878 15026 36930 15038
rect 39006 15090 39058 15102
rect 39006 15026 39058 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 21422 14754 21474 14766
rect 21422 14690 21474 14702
rect 21758 14754 21810 14766
rect 21758 14690 21810 14702
rect 24334 14754 24386 14766
rect 24334 14690 24386 14702
rect 35982 14754 36034 14766
rect 35982 14690 36034 14702
rect 42478 14754 42530 14766
rect 42478 14690 42530 14702
rect 11790 14642 11842 14654
rect 20750 14642 20802 14654
rect 11330 14590 11342 14642
rect 11394 14590 11406 14642
rect 18162 14590 18174 14642
rect 18226 14590 18238 14642
rect 20290 14590 20302 14642
rect 20354 14590 20366 14642
rect 27010 14590 27022 14642
rect 27074 14590 27086 14642
rect 28130 14590 28142 14642
rect 28194 14590 28206 14642
rect 31938 14590 31950 14642
rect 32002 14590 32014 14642
rect 37874 14590 37886 14642
rect 37938 14590 37950 14642
rect 40002 14590 40014 14642
rect 40066 14590 40078 14642
rect 11790 14578 11842 14590
rect 20750 14578 20802 14590
rect 25902 14530 25954 14542
rect 8530 14478 8542 14530
rect 8594 14478 8606 14530
rect 16594 14478 16606 14530
rect 16658 14478 16670 14530
rect 17378 14478 17390 14530
rect 17442 14478 17454 14530
rect 24098 14478 24110 14530
rect 24162 14478 24174 14530
rect 24434 14478 24446 14530
rect 24498 14478 24510 14530
rect 25442 14478 25454 14530
rect 25506 14478 25518 14530
rect 25902 14466 25954 14478
rect 26686 14530 26738 14542
rect 35310 14530 35362 14542
rect 36094 14530 36146 14542
rect 27458 14478 27470 14530
rect 27522 14478 27534 14530
rect 28354 14478 28366 14530
rect 28418 14478 28430 14530
rect 29138 14478 29150 14530
rect 29202 14478 29214 14530
rect 30146 14478 30158 14530
rect 30210 14478 30222 14530
rect 31042 14478 31054 14530
rect 31106 14478 31118 14530
rect 35634 14478 35646 14530
rect 35698 14478 35710 14530
rect 40786 14478 40798 14530
rect 40850 14478 40862 14530
rect 41458 14478 41470 14530
rect 41522 14478 41534 14530
rect 43922 14478 43934 14530
rect 43986 14478 43998 14530
rect 26686 14466 26738 14478
rect 35310 14466 35362 14478
rect 36094 14466 36146 14478
rect 23886 14418 23938 14430
rect 9202 14366 9214 14418
rect 9266 14366 9278 14418
rect 16370 14366 16382 14418
rect 16434 14366 16446 14418
rect 16930 14366 16942 14418
rect 16994 14366 17006 14418
rect 21970 14366 21982 14418
rect 22034 14366 22046 14418
rect 22306 14366 22318 14418
rect 22370 14366 22382 14418
rect 23886 14354 23938 14366
rect 26126 14418 26178 14430
rect 26126 14354 26178 14366
rect 26462 14418 26514 14430
rect 26462 14354 26514 14366
rect 26910 14418 26962 14430
rect 32398 14418 32450 14430
rect 27906 14366 27918 14418
rect 27970 14366 27982 14418
rect 30258 14366 30270 14418
rect 30322 14366 30334 14418
rect 31154 14366 31166 14418
rect 31218 14366 31230 14418
rect 26910 14354 26962 14366
rect 32398 14354 32450 14366
rect 33182 14418 33234 14430
rect 33182 14354 33234 14366
rect 34862 14418 34914 14430
rect 34862 14354 34914 14366
rect 35086 14418 35138 14430
rect 35086 14354 35138 14366
rect 36430 14418 36482 14430
rect 36430 14354 36482 14366
rect 41694 14418 41746 14430
rect 41694 14354 41746 14366
rect 42142 14418 42194 14430
rect 44158 14418 44210 14430
rect 42690 14366 42702 14418
rect 42754 14366 42766 14418
rect 43250 14366 43262 14418
rect 43314 14366 43326 14418
rect 42142 14354 42194 14366
rect 44158 14354 44210 14366
rect 23998 14306 24050 14318
rect 23998 14242 24050 14254
rect 25678 14306 25730 14318
rect 25678 14242 25730 14254
rect 25790 14306 25842 14318
rect 25790 14242 25842 14254
rect 27022 14306 27074 14318
rect 27022 14242 27074 14254
rect 29038 14306 29090 14318
rect 29038 14242 29090 14254
rect 31950 14306 32002 14318
rect 31950 14242 32002 14254
rect 32174 14306 32226 14318
rect 32174 14242 32226 14254
rect 32622 14306 32674 14318
rect 32622 14242 32674 14254
rect 32734 14306 32786 14318
rect 32734 14242 32786 14254
rect 32958 14306 33010 14318
rect 32958 14242 33010 14254
rect 35198 14306 35250 14318
rect 35970 14254 35982 14306
rect 36034 14254 36046 14306
rect 35198 14242 35250 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 9550 13970 9602 13982
rect 9550 13906 9602 13918
rect 19742 13970 19794 13982
rect 19742 13906 19794 13918
rect 21310 13970 21362 13982
rect 21310 13906 21362 13918
rect 23326 13970 23378 13982
rect 26014 13970 26066 13982
rect 24098 13918 24110 13970
rect 24162 13918 24174 13970
rect 23326 13906 23378 13918
rect 26014 13906 26066 13918
rect 28814 13970 28866 13982
rect 28814 13906 28866 13918
rect 32062 13970 32114 13982
rect 32062 13906 32114 13918
rect 32174 13970 32226 13982
rect 32174 13906 32226 13918
rect 34302 13970 34354 13982
rect 34302 13906 34354 13918
rect 35310 13970 35362 13982
rect 35310 13906 35362 13918
rect 36430 13970 36482 13982
rect 36430 13906 36482 13918
rect 37662 13970 37714 13982
rect 37662 13906 37714 13918
rect 38222 13970 38274 13982
rect 38222 13906 38274 13918
rect 39902 13970 39954 13982
rect 39902 13906 39954 13918
rect 41022 13970 41074 13982
rect 41022 13906 41074 13918
rect 41918 13970 41970 13982
rect 41918 13906 41970 13918
rect 44718 13970 44770 13982
rect 44718 13906 44770 13918
rect 8990 13858 9042 13870
rect 6402 13806 6414 13858
rect 6466 13806 6478 13858
rect 8990 13794 9042 13806
rect 10222 13858 10274 13870
rect 10222 13794 10274 13806
rect 10558 13858 10610 13870
rect 15486 13858 15538 13870
rect 25342 13858 25394 13870
rect 12002 13806 12014 13858
rect 12066 13806 12078 13858
rect 13682 13806 13694 13858
rect 13746 13806 13758 13858
rect 16482 13806 16494 13858
rect 16546 13806 16558 13858
rect 17602 13806 17614 13858
rect 17666 13806 17678 13858
rect 20626 13806 20638 13858
rect 20690 13806 20702 13858
rect 23874 13806 23886 13858
rect 23938 13806 23950 13858
rect 10558 13794 10610 13806
rect 15486 13794 15538 13806
rect 25342 13794 25394 13806
rect 25566 13858 25618 13870
rect 33294 13858 33346 13870
rect 27906 13806 27918 13858
rect 27970 13806 27982 13858
rect 30258 13806 30270 13858
rect 30322 13806 30334 13858
rect 30818 13806 30830 13858
rect 30882 13806 30894 13858
rect 25566 13794 25618 13806
rect 33294 13794 33346 13806
rect 33406 13858 33458 13870
rect 37214 13858 37266 13870
rect 35858 13806 35870 13858
rect 35922 13806 35934 13858
rect 36978 13806 36990 13858
rect 37042 13806 37054 13858
rect 33406 13794 33458 13806
rect 37214 13794 37266 13806
rect 38110 13858 38162 13870
rect 38110 13794 38162 13806
rect 38446 13858 38498 13870
rect 38882 13806 38894 13858
rect 38946 13806 38958 13858
rect 42578 13806 42590 13858
rect 42642 13806 42654 13858
rect 42802 13806 42814 13858
rect 42866 13806 42878 13858
rect 43586 13806 43598 13858
rect 43650 13806 43662 13858
rect 38446 13794 38498 13806
rect 9886 13746 9938 13758
rect 5730 13694 5742 13746
rect 5794 13694 5806 13746
rect 9886 13682 9938 13694
rect 11118 13746 11170 13758
rect 11118 13682 11170 13694
rect 11454 13746 11506 13758
rect 15822 13746 15874 13758
rect 18622 13746 18674 13758
rect 12226 13694 12238 13746
rect 12290 13694 12302 13746
rect 13570 13694 13582 13746
rect 13634 13694 13646 13746
rect 16594 13694 16606 13746
rect 16658 13694 16670 13746
rect 17714 13694 17726 13746
rect 17778 13694 17790 13746
rect 11454 13682 11506 13694
rect 15822 13682 15874 13694
rect 18622 13682 18674 13694
rect 20078 13746 20130 13758
rect 22542 13746 22594 13758
rect 22990 13746 23042 13758
rect 23662 13746 23714 13758
rect 26574 13746 26626 13758
rect 31950 13746 32002 13758
rect 33070 13746 33122 13758
rect 34190 13746 34242 13758
rect 20850 13694 20862 13746
rect 20914 13694 20926 13746
rect 22754 13694 22766 13746
rect 22818 13694 22830 13746
rect 23314 13694 23326 13746
rect 23378 13694 23390 13746
rect 24434 13694 24446 13746
rect 24498 13694 24510 13746
rect 27458 13694 27470 13746
rect 27522 13694 27534 13746
rect 28354 13694 28366 13746
rect 28418 13694 28430 13746
rect 29250 13694 29262 13746
rect 29314 13694 29326 13746
rect 29922 13694 29934 13746
rect 29986 13694 29998 13746
rect 31042 13694 31054 13746
rect 31106 13694 31118 13746
rect 32498 13694 32510 13746
rect 32562 13694 32574 13746
rect 33842 13694 33854 13746
rect 33906 13694 33918 13746
rect 20078 13682 20130 13694
rect 22542 13682 22594 13694
rect 22990 13682 23042 13694
rect 23662 13682 23714 13694
rect 26574 13682 26626 13694
rect 31950 13682 32002 13694
rect 33070 13682 33122 13694
rect 34190 13682 34242 13694
rect 34414 13746 34466 13758
rect 36094 13746 36146 13758
rect 39566 13746 39618 13758
rect 34738 13694 34750 13746
rect 34802 13694 34814 13746
rect 35410 13694 35422 13746
rect 35474 13694 35486 13746
rect 36530 13694 36542 13746
rect 36594 13694 36606 13746
rect 38770 13694 38782 13746
rect 38834 13694 38846 13746
rect 34414 13682 34466 13694
rect 36094 13682 36146 13694
rect 39566 13682 39618 13694
rect 42254 13746 42306 13758
rect 44382 13746 44434 13758
rect 43810 13694 43822 13746
rect 43874 13694 43886 13746
rect 42254 13682 42306 13694
rect 44382 13682 44434 13694
rect 19182 13634 19234 13646
rect 27246 13634 27298 13646
rect 45278 13634 45330 13646
rect 8530 13582 8542 13634
rect 8594 13582 8606 13634
rect 21746 13582 21758 13634
rect 21810 13582 21822 13634
rect 27794 13582 27806 13634
rect 27858 13582 27870 13634
rect 33282 13582 33294 13634
rect 33346 13582 33358 13634
rect 19182 13570 19234 13582
rect 27246 13570 27298 13582
rect 45278 13570 45330 13582
rect 14366 13522 14418 13534
rect 14366 13458 14418 13470
rect 14702 13522 14754 13534
rect 14702 13458 14754 13470
rect 16718 13522 16770 13534
rect 16718 13458 16770 13470
rect 18286 13522 18338 13534
rect 25678 13522 25730 13534
rect 24210 13470 24222 13522
rect 24274 13470 24286 13522
rect 18286 13458 18338 13470
rect 25678 13458 25730 13470
rect 35646 13522 35698 13534
rect 35646 13458 35698 13470
rect 36766 13522 36818 13534
rect 36766 13458 36818 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 18062 13186 18114 13198
rect 26350 13186 26402 13198
rect 24546 13134 24558 13186
rect 24610 13134 24622 13186
rect 18062 13122 18114 13134
rect 26350 13122 26402 13134
rect 26686 13186 26738 13198
rect 26686 13122 26738 13134
rect 42142 13186 42194 13198
rect 42142 13122 42194 13134
rect 11566 13074 11618 13086
rect 25342 13074 25394 13086
rect 29262 13074 29314 13086
rect 35534 13074 35586 13086
rect 8978 13022 8990 13074
rect 9042 13022 9054 13074
rect 11106 13022 11118 13074
rect 11170 13022 11182 13074
rect 15138 13022 15150 13074
rect 15202 13022 15214 13074
rect 17266 13022 17278 13074
rect 17330 13022 17342 13074
rect 25778 13022 25790 13074
rect 25842 13022 25854 13074
rect 31378 13022 31390 13074
rect 31442 13022 31454 13074
rect 33394 13022 33406 13074
rect 33458 13022 33470 13074
rect 11566 13010 11618 13022
rect 25342 13010 25394 13022
rect 29262 13010 29314 13022
rect 35534 13010 35586 13022
rect 37774 13074 37826 13086
rect 37774 13010 37826 13022
rect 38222 13074 38274 13086
rect 47730 13022 47742 13074
rect 47794 13022 47806 13074
rect 38222 13010 38274 13022
rect 17726 12962 17778 12974
rect 23998 12962 24050 12974
rect 34862 12962 34914 12974
rect 8306 12910 8318 12962
rect 8370 12910 8382 12962
rect 14354 12910 14366 12962
rect 14418 12910 14430 12962
rect 18498 12910 18510 12962
rect 18562 12910 18574 12962
rect 21522 12910 21534 12962
rect 21586 12910 21598 12962
rect 23538 12910 23550 12962
rect 23602 12910 23614 12962
rect 24546 12910 24558 12962
rect 24610 12910 24622 12962
rect 25890 12910 25902 12962
rect 25954 12910 25966 12962
rect 29474 12910 29486 12962
rect 29538 12910 29550 12962
rect 17726 12898 17778 12910
rect 23998 12898 24050 12910
rect 34862 12898 34914 12910
rect 34974 12962 35026 12974
rect 34974 12898 35026 12910
rect 35758 12962 35810 12974
rect 35758 12898 35810 12910
rect 35982 12962 36034 12974
rect 35982 12898 36034 12910
rect 39342 12962 39394 12974
rect 39342 12898 39394 12910
rect 42478 12962 42530 12974
rect 44034 12910 44046 12962
rect 44098 12910 44110 12962
rect 44818 12910 44830 12962
rect 44882 12910 44894 12962
rect 42478 12898 42530 12910
rect 23326 12850 23378 12862
rect 25566 12850 25618 12862
rect 18722 12798 18734 12850
rect 18786 12798 18798 12850
rect 24210 12798 24222 12850
rect 24274 12798 24286 12850
rect 23326 12786 23378 12798
rect 25566 12786 25618 12798
rect 26574 12850 26626 12862
rect 26574 12786 26626 12798
rect 27582 12850 27634 12862
rect 27582 12786 27634 12798
rect 28254 12850 28306 12862
rect 29150 12850 29202 12862
rect 28578 12798 28590 12850
rect 28642 12798 28654 12850
rect 28254 12786 28306 12798
rect 29150 12786 29202 12798
rect 30942 12850 30994 12862
rect 32958 12850 33010 12862
rect 34638 12850 34690 12862
rect 32162 12798 32174 12850
rect 32226 12798 32238 12850
rect 33170 12798 33182 12850
rect 33234 12798 33246 12850
rect 30942 12786 30994 12798
rect 32958 12786 33010 12798
rect 34638 12786 34690 12798
rect 35422 12850 35474 12862
rect 35422 12786 35474 12798
rect 39006 12850 39058 12862
rect 39006 12786 39058 12798
rect 39118 12850 39170 12862
rect 39118 12786 39170 12798
rect 39678 12850 39730 12862
rect 44270 12850 44322 12862
rect 42690 12798 42702 12850
rect 42754 12798 42766 12850
rect 43250 12798 43262 12850
rect 43314 12798 43326 12850
rect 45602 12798 45614 12850
rect 45666 12798 45678 12850
rect 39678 12786 39730 12798
rect 44270 12786 44322 12798
rect 21310 12738 21362 12750
rect 21310 12674 21362 12686
rect 22542 12738 22594 12750
rect 22542 12674 22594 12686
rect 22990 12738 23042 12750
rect 22990 12674 23042 12686
rect 24782 12738 24834 12750
rect 24782 12674 24834 12686
rect 27246 12738 27298 12750
rect 27246 12674 27298 12686
rect 27918 12738 27970 12750
rect 27918 12674 27970 12686
rect 30606 12738 30658 12750
rect 30606 12674 30658 12686
rect 31838 12738 31890 12750
rect 31838 12674 31890 12686
rect 32622 12738 32674 12750
rect 32622 12674 32674 12686
rect 32846 12738 32898 12750
rect 32846 12674 32898 12686
rect 35086 12738 35138 12750
rect 35086 12674 35138 12686
rect 38670 12738 38722 12750
rect 38670 12674 38722 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 17502 12402 17554 12414
rect 23998 12402 24050 12414
rect 23202 12350 23214 12402
rect 23266 12350 23278 12402
rect 17502 12338 17554 12350
rect 23998 12338 24050 12350
rect 25902 12402 25954 12414
rect 25902 12338 25954 12350
rect 27470 12402 27522 12414
rect 27470 12338 27522 12350
rect 27694 12402 27746 12414
rect 27694 12338 27746 12350
rect 28814 12402 28866 12414
rect 34750 12402 34802 12414
rect 31042 12350 31054 12402
rect 31106 12350 31118 12402
rect 32050 12350 32062 12402
rect 32114 12350 32126 12402
rect 28814 12338 28866 12350
rect 34750 12338 34802 12350
rect 35534 12402 35586 12414
rect 35534 12338 35586 12350
rect 36206 12402 36258 12414
rect 36206 12338 36258 12350
rect 37998 12402 38050 12414
rect 37998 12338 38050 12350
rect 38222 12402 38274 12414
rect 38222 12338 38274 12350
rect 44942 12402 44994 12414
rect 44942 12338 44994 12350
rect 24222 12290 24274 12302
rect 15250 12238 15262 12290
rect 15314 12238 15326 12290
rect 20626 12238 20638 12290
rect 20690 12238 20702 12290
rect 24222 12226 24274 12238
rect 25230 12290 25282 12302
rect 33854 12290 33906 12302
rect 30370 12238 30382 12290
rect 30434 12238 30446 12290
rect 25230 12226 25282 12238
rect 33854 12226 33906 12238
rect 34302 12290 34354 12302
rect 34302 12226 34354 12238
rect 35198 12290 35250 12302
rect 35198 12226 35250 12238
rect 35422 12290 35474 12302
rect 35422 12226 35474 12238
rect 37326 12290 37378 12302
rect 39218 12238 39230 12290
rect 39282 12238 39294 12290
rect 39666 12238 39678 12290
rect 39730 12238 39742 12290
rect 42690 12238 42702 12290
rect 42754 12238 42766 12290
rect 43138 12238 43150 12290
rect 43202 12238 43214 12290
rect 43922 12238 43934 12290
rect 43986 12238 43998 12290
rect 37326 12226 37378 12238
rect 14590 12178 14642 12190
rect 23886 12178 23938 12190
rect 10994 12126 11006 12178
rect 11058 12126 11070 12178
rect 15362 12126 15374 12178
rect 15426 12126 15438 12178
rect 19842 12126 19854 12178
rect 19906 12126 19918 12178
rect 23426 12126 23438 12178
rect 23490 12126 23502 12178
rect 14590 12114 14642 12126
rect 23886 12114 23938 12126
rect 24446 12178 24498 12190
rect 24446 12114 24498 12126
rect 25342 12178 25394 12190
rect 25342 12114 25394 12126
rect 27246 12178 27298 12190
rect 28478 12178 28530 12190
rect 28926 12178 28978 12190
rect 28354 12126 28366 12178
rect 28418 12126 28430 12178
rect 28690 12126 28702 12178
rect 28754 12126 28766 12178
rect 27246 12114 27298 12126
rect 28478 12114 28530 12126
rect 28926 12114 28978 12126
rect 29262 12178 29314 12190
rect 31390 12178 31442 12190
rect 29474 12126 29486 12178
rect 29538 12126 29550 12178
rect 30034 12126 30046 12178
rect 30098 12126 30110 12178
rect 30594 12126 30606 12178
rect 30658 12126 30670 12178
rect 29262 12114 29314 12126
rect 31390 12114 31442 12126
rect 31726 12178 31778 12190
rect 34638 12178 34690 12190
rect 33618 12126 33630 12178
rect 33682 12126 33694 12178
rect 31726 12114 31778 12126
rect 34638 12114 34690 12126
rect 34974 12178 35026 12190
rect 34974 12114 35026 12126
rect 35870 12178 35922 12190
rect 35870 12114 35922 12126
rect 35982 12178 36034 12190
rect 35982 12114 36034 12126
rect 36430 12178 36482 12190
rect 36430 12114 36482 12126
rect 36542 12178 36594 12190
rect 36542 12114 36594 12126
rect 37886 12178 37938 12190
rect 44606 12178 44658 12190
rect 43810 12126 43822 12178
rect 43874 12126 43886 12178
rect 37886 12114 37938 12126
rect 44606 12114 44658 12126
rect 27358 12066 27410 12078
rect 11666 12014 11678 12066
rect 11730 12014 11742 12066
rect 13794 12014 13806 12066
rect 13858 12014 13870 12066
rect 22754 12014 22766 12066
rect 22818 12014 22830 12066
rect 27358 12002 27410 12014
rect 29374 12066 29426 12078
rect 37202 12014 37214 12066
rect 37266 12014 37278 12066
rect 29374 12002 29426 12014
rect 14254 11954 14306 11966
rect 37550 11954 37602 11966
rect 29810 11902 29822 11954
rect 29874 11902 29886 11954
rect 14254 11890 14306 11902
rect 37550 11890 37602 11902
rect 38558 11954 38610 11966
rect 38558 11890 38610 11902
rect 38894 11954 38946 11966
rect 38894 11890 38946 11902
rect 42142 11954 42194 11966
rect 42142 11890 42194 11902
rect 42478 11954 42530 11966
rect 42478 11890 42530 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 21422 11618 21474 11630
rect 21422 11554 21474 11566
rect 21758 11618 21810 11630
rect 21758 11554 21810 11566
rect 23102 11618 23154 11630
rect 23102 11554 23154 11566
rect 14030 11506 14082 11518
rect 20638 11506 20690 11518
rect 20178 11454 20190 11506
rect 20242 11454 20254 11506
rect 14030 11442 14082 11454
rect 20638 11442 20690 11454
rect 30270 11506 30322 11518
rect 36430 11506 36482 11518
rect 41022 11506 41074 11518
rect 31042 11454 31054 11506
rect 31106 11454 31118 11506
rect 33842 11454 33854 11506
rect 33906 11454 33918 11506
rect 35970 11454 35982 11506
rect 36034 11454 36046 11506
rect 37650 11454 37662 11506
rect 37714 11454 37726 11506
rect 44258 11454 44270 11506
rect 44322 11454 44334 11506
rect 30270 11442 30322 11454
rect 36430 11442 36482 11454
rect 41022 11442 41074 11454
rect 12462 11394 12514 11406
rect 12462 11330 12514 11342
rect 15710 11394 15762 11406
rect 22990 11394 23042 11406
rect 17266 11342 17278 11394
rect 17330 11342 17342 11394
rect 15710 11330 15762 11342
rect 22990 11330 23042 11342
rect 23886 11394 23938 11406
rect 23886 11330 23938 11342
rect 24334 11394 24386 11406
rect 24334 11330 24386 11342
rect 24446 11394 24498 11406
rect 24446 11330 24498 11342
rect 24782 11394 24834 11406
rect 24782 11330 24834 11342
rect 27470 11394 27522 11406
rect 27470 11330 27522 11342
rect 27806 11394 27858 11406
rect 27806 11330 27858 11342
rect 28142 11394 28194 11406
rect 31838 11394 31890 11406
rect 30706 11342 30718 11394
rect 30770 11342 30782 11394
rect 33170 11342 33182 11394
rect 33234 11342 33246 11394
rect 40562 11342 40574 11394
rect 40626 11342 40638 11394
rect 41346 11342 41358 11394
rect 41410 11342 41422 11394
rect 28142 11330 28194 11342
rect 31838 11330 31890 11342
rect 12126 11282 12178 11294
rect 24222 11282 24274 11294
rect 18050 11230 18062 11282
rect 18114 11230 18126 11282
rect 21970 11230 21982 11282
rect 22034 11230 22046 11282
rect 22306 11230 22318 11282
rect 22370 11230 22382 11282
rect 12126 11218 12178 11230
rect 24222 11218 24274 11230
rect 25118 11282 25170 11294
rect 25118 11218 25170 11230
rect 25454 11282 25506 11294
rect 39778 11230 39790 11282
rect 39842 11230 39854 11282
rect 42130 11230 42142 11282
rect 42194 11230 42206 11282
rect 25454 11218 25506 11230
rect 16270 11170 16322 11182
rect 16270 11106 16322 11118
rect 23102 11170 23154 11182
rect 23102 11106 23154 11118
rect 23550 11170 23602 11182
rect 23550 11106 23602 11118
rect 25902 11170 25954 11182
rect 25902 11106 25954 11118
rect 27022 11170 27074 11182
rect 27022 11106 27074 11118
rect 27694 11170 27746 11182
rect 27694 11106 27746 11118
rect 31502 11170 31554 11182
rect 31502 11106 31554 11118
rect 37326 11170 37378 11182
rect 37326 11106 37378 11118
rect 44942 11170 44994 11182
rect 44942 11106 44994 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 15038 10834 15090 10846
rect 15038 10770 15090 10782
rect 18622 10834 18674 10846
rect 18622 10770 18674 10782
rect 24222 10834 24274 10846
rect 24222 10770 24274 10782
rect 26126 10834 26178 10846
rect 26126 10770 26178 10782
rect 33406 10834 33458 10846
rect 33406 10770 33458 10782
rect 33854 10834 33906 10846
rect 33854 10770 33906 10782
rect 35870 10834 35922 10846
rect 35870 10770 35922 10782
rect 38670 10834 38722 10846
rect 38670 10770 38722 10782
rect 42030 10834 42082 10846
rect 42030 10770 42082 10782
rect 25342 10722 25394 10734
rect 27582 10722 27634 10734
rect 14130 10670 14142 10722
rect 14194 10670 14206 10722
rect 14466 10670 14478 10722
rect 14530 10670 14542 10722
rect 20514 10670 20526 10722
rect 20578 10670 20590 10722
rect 22306 10670 22318 10722
rect 22370 10670 22382 10722
rect 26562 10670 26574 10722
rect 26626 10670 26638 10722
rect 25342 10658 25394 10670
rect 27582 10658 27634 10670
rect 28814 10722 28866 10734
rect 28814 10658 28866 10670
rect 31390 10722 31442 10734
rect 40014 10722 40066 10734
rect 34962 10670 34974 10722
rect 35026 10670 35038 10722
rect 36418 10670 36430 10722
rect 36482 10670 36494 10722
rect 36866 10670 36878 10722
rect 36930 10670 36942 10722
rect 31390 10658 31442 10670
rect 40014 10658 40066 10670
rect 18958 10610 19010 10622
rect 10434 10558 10446 10610
rect 10498 10558 10510 10610
rect 17826 10558 17838 10610
rect 17890 10558 17902 10610
rect 18958 10546 19010 10558
rect 19630 10610 19682 10622
rect 19630 10546 19682 10558
rect 19966 10610 20018 10622
rect 34190 10610 34242 10622
rect 36206 10610 36258 10622
rect 20738 10558 20750 10610
rect 20802 10558 20814 10610
rect 22082 10558 22094 10610
rect 22146 10558 22158 10610
rect 23202 10558 23214 10610
rect 23266 10558 23278 10610
rect 26450 10558 26462 10610
rect 26514 10558 26526 10610
rect 27794 10558 27806 10610
rect 27858 10558 27870 10610
rect 31154 10558 31166 10610
rect 31218 10558 31230 10610
rect 34738 10558 34750 10610
rect 34802 10558 34814 10610
rect 38434 10558 38446 10610
rect 38498 10558 38510 10610
rect 39778 10558 39790 10610
rect 39842 10558 39854 10610
rect 42242 10558 42254 10610
rect 42306 10558 42318 10610
rect 19966 10546 20018 10558
rect 34190 10546 34242 10558
rect 36206 10546 36258 10558
rect 14702 10498 14754 10510
rect 11106 10446 11118 10498
rect 11170 10446 11182 10498
rect 13234 10446 13246 10498
rect 13298 10446 13310 10498
rect 14702 10434 14754 10446
rect 18286 10498 18338 10510
rect 18286 10434 18338 10446
rect 22766 10498 22818 10510
rect 23538 10446 23550 10498
rect 23602 10446 23614 10498
rect 25218 10446 25230 10498
rect 25282 10446 25294 10498
rect 27010 10446 27022 10498
rect 27074 10446 27086 10498
rect 22766 10434 22818 10446
rect 25566 10386 25618 10398
rect 25566 10322 25618 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 14366 10050 14418 10062
rect 14366 9986 14418 9998
rect 25902 10050 25954 10062
rect 25902 9986 25954 9998
rect 27358 10050 27410 10062
rect 27358 9986 27410 9998
rect 29486 10050 29538 10062
rect 31938 9998 31950 10050
rect 32002 10047 32014 10050
rect 33170 10047 33182 10050
rect 32002 10001 33182 10047
rect 32002 9998 32014 10001
rect 33170 9998 33182 10001
rect 33234 9998 33246 10050
rect 29486 9986 29538 9998
rect 13582 9938 13634 9950
rect 13582 9874 13634 9886
rect 17054 9938 17106 9950
rect 17054 9874 17106 9886
rect 22430 9938 22482 9950
rect 27694 9938 27746 9950
rect 23986 9886 23998 9938
rect 24050 9886 24062 9938
rect 22430 9874 22482 9886
rect 27694 9874 27746 9886
rect 31950 9938 32002 9950
rect 42814 9938 42866 9950
rect 39442 9886 39454 9938
rect 39506 9886 39518 9938
rect 41570 9886 41582 9938
rect 41634 9886 41646 9938
rect 31950 9874 32002 9886
rect 42814 9874 42866 9886
rect 17502 9826 17554 9838
rect 14802 9774 14814 9826
rect 14866 9774 14878 9826
rect 17502 9762 17554 9774
rect 18062 9826 18114 9838
rect 18062 9762 18114 9774
rect 18734 9826 18786 9838
rect 18734 9762 18786 9774
rect 19294 9826 19346 9838
rect 19294 9762 19346 9774
rect 22094 9826 22146 9838
rect 22094 9762 22146 9774
rect 22654 9826 22706 9838
rect 32398 9826 32450 9838
rect 24322 9774 24334 9826
rect 24386 9774 24398 9826
rect 22654 9762 22706 9774
rect 32398 9762 32450 9774
rect 33406 9826 33458 9838
rect 33406 9762 33458 9774
rect 33630 9826 33682 9838
rect 42242 9774 42254 9826
rect 42306 9774 42318 9826
rect 33630 9762 33682 9774
rect 11342 9714 11394 9726
rect 11342 9650 11394 9662
rect 11678 9714 11730 9726
rect 11678 9650 11730 9662
rect 14030 9714 14082 9726
rect 17390 9714 17442 9726
rect 14914 9662 14926 9714
rect 14978 9662 14990 9714
rect 14030 9650 14082 9662
rect 17390 9650 17442 9662
rect 17950 9714 18002 9726
rect 17950 9650 18002 9662
rect 19182 9714 19234 9726
rect 19182 9650 19234 9662
rect 19742 9714 19794 9726
rect 25118 9714 25170 9726
rect 22978 9662 22990 9714
rect 23042 9662 23054 9714
rect 19742 9650 19794 9662
rect 25118 9650 25170 9662
rect 25566 9714 25618 9726
rect 29150 9714 29202 9726
rect 26114 9662 26126 9714
rect 26178 9662 26190 9714
rect 26450 9662 26462 9714
rect 26514 9662 26526 9714
rect 27906 9662 27918 9714
rect 27970 9662 27982 9714
rect 28466 9662 28478 9714
rect 28530 9662 28542 9714
rect 38658 9662 38670 9714
rect 38722 9662 38734 9714
rect 25566 9650 25618 9662
rect 29150 9650 29202 9662
rect 17166 9602 17218 9614
rect 17166 9538 17218 9550
rect 17726 9602 17778 9614
rect 17726 9538 17778 9550
rect 18398 9602 18450 9614
rect 18398 9538 18450 9550
rect 18622 9602 18674 9614
rect 18622 9538 18674 9550
rect 18958 9602 19010 9614
rect 18958 9538 19010 9550
rect 20190 9602 20242 9614
rect 20190 9538 20242 9550
rect 21646 9602 21698 9614
rect 21646 9538 21698 9550
rect 24782 9602 24834 9614
rect 24782 9538 24834 9550
rect 29374 9602 29426 9614
rect 29374 9538 29426 9550
rect 32846 9602 32898 9614
rect 35758 9602 35810 9614
rect 33954 9550 33966 9602
rect 34018 9550 34030 9602
rect 32846 9538 32898 9550
rect 35758 9538 35810 9550
rect 36206 9602 36258 9614
rect 36206 9538 36258 9550
rect 37998 9602 38050 9614
rect 37998 9538 38050 9550
rect 38334 9602 38386 9614
rect 38334 9538 38386 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 16718 9266 16770 9278
rect 16718 9202 16770 9214
rect 18622 9266 18674 9278
rect 23662 9266 23714 9278
rect 21186 9214 21198 9266
rect 21250 9214 21262 9266
rect 18622 9202 18674 9214
rect 23662 9202 23714 9214
rect 34302 9266 34354 9278
rect 34302 9202 34354 9214
rect 36430 9266 36482 9278
rect 36430 9202 36482 9214
rect 36990 9266 37042 9278
rect 36990 9202 37042 9214
rect 37998 9266 38050 9278
rect 37998 9202 38050 9214
rect 40238 9266 40290 9278
rect 40238 9202 40290 9214
rect 17614 9154 17666 9166
rect 22654 9154 22706 9166
rect 14914 9102 14926 9154
rect 14978 9102 14990 9154
rect 15586 9102 15598 9154
rect 15650 9102 15662 9154
rect 16034 9102 16046 9154
rect 16098 9102 16110 9154
rect 19618 9102 19630 9154
rect 19682 9102 19694 9154
rect 21858 9102 21870 9154
rect 21922 9102 21934 9154
rect 17614 9090 17666 9102
rect 22654 9090 22706 9102
rect 22766 9154 22818 9166
rect 33182 9154 33234 9166
rect 27122 9102 27134 9154
rect 27186 9102 27198 9154
rect 22766 9090 22818 9102
rect 33182 9090 33234 9102
rect 33294 9154 33346 9166
rect 33294 9090 33346 9102
rect 33742 9154 33794 9166
rect 33742 9090 33794 9102
rect 33854 9154 33906 9166
rect 36542 9154 36594 9166
rect 35298 9102 35310 9154
rect 35362 9102 35374 9154
rect 35858 9102 35870 9154
rect 35922 9102 35934 9154
rect 33854 9090 33906 9102
rect 36542 9090 36594 9102
rect 38446 9154 38498 9166
rect 38446 9090 38498 9102
rect 38558 9154 38610 9166
rect 39330 9102 39342 9154
rect 39394 9102 39406 9154
rect 38558 9090 38610 9102
rect 14254 9042 14306 9054
rect 17950 9042 18002 9054
rect 21534 9042 21586 9054
rect 10546 8990 10558 9042
rect 10610 8990 10622 9042
rect 15026 8990 15038 9042
rect 15090 8990 15102 9042
rect 19394 8990 19406 9042
rect 19458 8990 19470 9042
rect 14254 8978 14306 8990
rect 17950 8978 18002 8990
rect 21534 8978 21586 8990
rect 22206 9042 22258 9054
rect 22206 8978 22258 8990
rect 22430 9042 22482 9054
rect 33518 9042 33570 9054
rect 26338 8990 26350 9042
rect 26402 8990 26414 9042
rect 29698 8990 29710 9042
rect 29762 8990 29774 9042
rect 22430 8978 22482 8990
rect 33518 8978 33570 8990
rect 36206 9042 36258 9054
rect 36206 8978 36258 8990
rect 37438 9042 37490 9054
rect 37438 8978 37490 8990
rect 38782 9042 38834 9054
rect 39902 9042 39954 9054
rect 39106 8990 39118 9042
rect 39170 8990 39182 9042
rect 38782 8978 38834 8990
rect 39902 8978 39954 8990
rect 19070 8930 19122 8942
rect 11330 8878 11342 8930
rect 11394 8878 11406 8930
rect 13458 8878 13470 8930
rect 13522 8878 13534 8930
rect 19070 8866 19122 8878
rect 23214 8930 23266 8942
rect 23214 8866 23266 8878
rect 26014 8930 26066 8942
rect 29250 8878 29262 8930
rect 29314 8878 29326 8930
rect 30370 8878 30382 8930
rect 30434 8878 30446 8930
rect 32498 8878 32510 8930
rect 32562 8878 32574 8930
rect 26014 8866 26066 8878
rect 13918 8818 13970 8830
rect 13918 8754 13970 8766
rect 16382 8818 16434 8830
rect 20190 8818 20242 8830
rect 18722 8766 18734 8818
rect 18786 8815 18798 8818
rect 19058 8815 19070 8818
rect 18786 8769 19070 8815
rect 18786 8766 18798 8769
rect 19058 8766 19070 8769
rect 19122 8766 19134 8818
rect 16382 8754 16434 8766
rect 20190 8754 20242 8766
rect 20526 8818 20578 8830
rect 20526 8754 20578 8766
rect 33182 8818 33234 8830
rect 33182 8754 33234 8766
rect 34750 8818 34802 8830
rect 34750 8754 34802 8766
rect 35086 8818 35138 8830
rect 35086 8754 35138 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 32286 8482 32338 8494
rect 32286 8418 32338 8430
rect 15150 8370 15202 8382
rect 20638 8370 20690 8382
rect 17378 8318 17390 8370
rect 17442 8318 17454 8370
rect 19506 8318 19518 8370
rect 19570 8318 19582 8370
rect 15150 8306 15202 8318
rect 20638 8306 20690 8318
rect 23550 8370 23602 8382
rect 33742 8370 33794 8382
rect 24658 8318 24670 8370
rect 24722 8318 24734 8370
rect 26786 8318 26798 8370
rect 26850 8318 26862 8370
rect 23550 8306 23602 8318
rect 33742 8306 33794 8318
rect 34190 8370 34242 8382
rect 34190 8306 34242 8318
rect 34526 8370 34578 8382
rect 34526 8306 34578 8318
rect 37102 8370 37154 8382
rect 37102 8306 37154 8318
rect 37438 8370 37490 8382
rect 37438 8306 37490 8318
rect 11902 8258 11954 8270
rect 34862 8258 34914 8270
rect 15922 8206 15934 8258
rect 15986 8206 15998 8258
rect 16706 8206 16718 8258
rect 16770 8206 16782 8258
rect 19954 8206 19966 8258
rect 20018 8206 20030 8258
rect 23874 8206 23886 8258
rect 23938 8206 23950 8258
rect 33058 8206 33070 8258
rect 33122 8206 33134 8258
rect 11902 8194 11954 8206
rect 34862 8194 34914 8206
rect 36094 8258 36146 8270
rect 36094 8194 36146 8206
rect 39342 8258 39394 8270
rect 39342 8194 39394 8206
rect 11566 8146 11618 8158
rect 21982 8146 22034 8158
rect 15810 8094 15822 8146
rect 15874 8094 15886 8146
rect 11566 8082 11618 8094
rect 21982 8082 22034 8094
rect 30942 8146 30994 8158
rect 30942 8082 30994 8094
rect 31278 8146 31330 8158
rect 31278 8082 31330 8094
rect 31950 8146 32002 8158
rect 32834 8094 32846 8146
rect 32898 8094 32910 8146
rect 37650 8094 37662 8146
rect 37714 8094 37726 8146
rect 38210 8094 38222 8146
rect 38274 8094 38286 8146
rect 39554 8094 39566 8146
rect 39618 8094 39630 8146
rect 39890 8094 39902 8146
rect 39954 8094 39966 8146
rect 31950 8082 32002 8094
rect 13694 8034 13746 8046
rect 13694 7970 13746 7982
rect 14814 8034 14866 8046
rect 14814 7970 14866 7982
rect 20190 8034 20242 8046
rect 22654 8034 22706 8046
rect 22306 7982 22318 8034
rect 22370 7982 22382 8034
rect 20190 7970 20242 7982
rect 22654 7970 22706 7982
rect 23102 8034 23154 8046
rect 23102 7970 23154 7982
rect 35198 8034 35250 8046
rect 39006 8034 39058 8046
rect 35746 7982 35758 8034
rect 35810 7982 35822 8034
rect 35198 7970 35250 7982
rect 39006 7970 39058 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 17838 7698 17890 7710
rect 17838 7634 17890 7646
rect 24558 7698 24610 7710
rect 24558 7634 24610 7646
rect 28814 7698 28866 7710
rect 28814 7634 28866 7646
rect 33406 7698 33458 7710
rect 33406 7634 33458 7646
rect 33742 7698 33794 7710
rect 33742 7634 33794 7646
rect 37886 7698 37938 7710
rect 37886 7634 37938 7646
rect 38446 7586 38498 7598
rect 39454 7586 39506 7598
rect 18834 7534 18846 7586
rect 18898 7534 18910 7586
rect 20178 7534 20190 7586
rect 20242 7534 20254 7586
rect 22642 7534 22654 7586
rect 22706 7534 22718 7586
rect 23538 7534 23550 7586
rect 23602 7534 23614 7586
rect 27794 7534 27806 7586
rect 27858 7534 27870 7586
rect 28242 7534 28254 7586
rect 28306 7534 28318 7586
rect 35298 7534 35310 7586
rect 35362 7534 35374 7586
rect 39106 7534 39118 7586
rect 39170 7534 39182 7586
rect 38446 7522 38498 7534
rect 39454 7522 39506 7534
rect 39790 7586 39842 7598
rect 39790 7522 39842 7534
rect 18174 7474 18226 7486
rect 22990 7474 23042 7486
rect 38782 7474 38834 7486
rect 12226 7422 12238 7474
rect 12290 7422 12302 7474
rect 18946 7422 18958 7474
rect 19010 7422 19022 7474
rect 19394 7422 19406 7474
rect 19458 7422 19470 7474
rect 23426 7422 23438 7474
rect 23490 7422 23502 7474
rect 29698 7422 29710 7474
rect 29762 7422 29774 7474
rect 34626 7422 34638 7474
rect 34690 7422 34702 7474
rect 18174 7410 18226 7422
rect 22990 7410 23042 7422
rect 38782 7410 38834 7422
rect 15486 7362 15538 7374
rect 12898 7310 12910 7362
rect 12962 7310 12974 7362
rect 15026 7310 15038 7362
rect 15090 7310 15102 7362
rect 22306 7310 22318 7362
rect 22370 7310 22382 7362
rect 30370 7310 30382 7362
rect 30434 7310 30446 7362
rect 32498 7310 32510 7362
rect 32562 7310 32574 7362
rect 37426 7310 37438 7362
rect 37490 7310 37502 7362
rect 15486 7298 15538 7310
rect 24222 7250 24274 7262
rect 24222 7186 24274 7198
rect 28478 7250 28530 7262
rect 28478 7186 28530 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 15486 6914 15538 6926
rect 15486 6850 15538 6862
rect 32398 6914 32450 6926
rect 32398 6850 32450 6862
rect 23998 6802 24050 6814
rect 27234 6750 27246 6802
rect 27298 6750 27310 6802
rect 38210 6750 38222 6802
rect 38274 6750 38286 6802
rect 23998 6738 24050 6750
rect 13806 6690 13858 6702
rect 22542 6690 22594 6702
rect 41582 6690 41634 6702
rect 16258 6638 16270 6690
rect 16322 6638 16334 6690
rect 24322 6638 24334 6690
rect 24386 6638 24398 6690
rect 29362 6638 29374 6690
rect 29426 6638 29438 6690
rect 33058 6638 33070 6690
rect 33122 6638 33134 6690
rect 41122 6638 41134 6690
rect 41186 6638 41198 6690
rect 13806 6626 13858 6638
rect 22542 6626 22594 6638
rect 41582 6626 41634 6638
rect 13470 6578 13522 6590
rect 23214 6578 23266 6590
rect 29934 6578 29986 6590
rect 16034 6526 16046 6578
rect 16098 6526 16110 6578
rect 25106 6526 25118 6578
rect 25170 6526 25182 6578
rect 13470 6514 13522 6526
rect 23214 6514 23266 6526
rect 29934 6514 29986 6526
rect 30942 6578 30994 6590
rect 30942 6514 30994 6526
rect 31278 6578 31330 6590
rect 31278 6514 31330 6526
rect 32062 6578 32114 6590
rect 32946 6526 32958 6578
rect 33010 6526 33022 6578
rect 40338 6526 40350 6578
rect 40402 6526 40414 6578
rect 32062 6514 32114 6526
rect 15150 6466 15202 6478
rect 29138 6414 29150 6466
rect 29202 6414 29214 6466
rect 15150 6402 15202 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 23886 6130 23938 6142
rect 23886 6066 23938 6078
rect 25566 6130 25618 6142
rect 25566 6066 25618 6078
rect 29262 6130 29314 6142
rect 29262 6066 29314 6078
rect 19070 6018 19122 6030
rect 18386 5966 18398 6018
rect 18450 5966 18462 6018
rect 19070 5954 19122 5966
rect 20638 6018 20690 6030
rect 30270 6018 30322 6030
rect 21970 5966 21982 6018
rect 22034 5966 22046 6018
rect 22978 5966 22990 6018
rect 23042 5966 23054 6018
rect 23314 5966 23326 6018
rect 23378 5966 23390 6018
rect 27010 5966 27022 6018
rect 27074 5966 27086 6018
rect 27570 5966 27582 6018
rect 27634 5966 27646 6018
rect 28242 5966 28254 6018
rect 28306 5966 28318 6018
rect 28690 5966 28702 6018
rect 28754 5966 28766 6018
rect 32162 5966 32174 6018
rect 32226 5966 32238 6018
rect 33842 5966 33854 6018
rect 33906 5966 33918 6018
rect 34290 5966 34302 6018
rect 34354 5966 34366 6018
rect 35410 5966 35422 6018
rect 35474 5966 35486 6018
rect 35970 5966 35982 6018
rect 36034 5966 36046 6018
rect 20638 5954 20690 5966
rect 30270 5954 30322 5966
rect 19406 5906 19458 5918
rect 25902 5906 25954 5918
rect 13346 5854 13358 5906
rect 13410 5854 13422 5906
rect 18274 5854 18286 5906
rect 18338 5854 18350 5906
rect 20402 5854 20414 5906
rect 20466 5854 20478 5906
rect 22194 5854 22206 5906
rect 22258 5854 22270 5906
rect 19406 5842 19458 5854
rect 25902 5842 25954 5854
rect 26462 5906 26514 5918
rect 26462 5842 26514 5854
rect 26798 5906 26850 5918
rect 26798 5842 26850 5854
rect 30606 5906 30658 5918
rect 30606 5842 30658 5854
rect 31278 5906 31330 5918
rect 31278 5842 31330 5854
rect 31614 5906 31666 5918
rect 33518 5906 33570 5918
rect 32386 5854 32398 5906
rect 32450 5854 32462 5906
rect 31614 5842 31666 5854
rect 33518 5842 33570 5854
rect 36206 5906 36258 5918
rect 36206 5842 36258 5854
rect 16606 5794 16658 5806
rect 14018 5742 14030 5794
rect 14082 5742 14094 5794
rect 16146 5742 16158 5794
rect 16210 5742 16222 5794
rect 16606 5730 16658 5742
rect 17838 5794 17890 5806
rect 17838 5730 17890 5742
rect 21086 5794 21138 5806
rect 21086 5730 21138 5742
rect 28926 5794 28978 5806
rect 28926 5730 28978 5742
rect 17502 5682 17554 5694
rect 17502 5618 17554 5630
rect 21422 5682 21474 5694
rect 21422 5618 21474 5630
rect 23550 5682 23602 5694
rect 23550 5618 23602 5630
rect 33182 5682 33234 5694
rect 33182 5618 33234 5630
rect 36542 5682 36594 5694
rect 36542 5618 36594 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 34974 5346 35026 5358
rect 34974 5282 35026 5294
rect 22318 5234 22370 5246
rect 34078 5234 34130 5246
rect 40350 5234 40402 5246
rect 18498 5182 18510 5234
rect 18562 5182 18574 5234
rect 20626 5182 20638 5234
rect 20690 5182 20702 5234
rect 26002 5182 26014 5234
rect 26066 5182 26078 5234
rect 31490 5182 31502 5234
rect 31554 5182 31566 5234
rect 33618 5182 33630 5234
rect 33682 5182 33694 5234
rect 36978 5182 36990 5234
rect 37042 5182 37054 5234
rect 22318 5170 22370 5182
rect 34078 5170 34130 5182
rect 40350 5170 40402 5182
rect 27694 5122 27746 5134
rect 14466 5070 14478 5122
rect 14530 5070 14542 5122
rect 17714 5070 17726 5122
rect 17778 5070 17790 5122
rect 23202 5070 23214 5122
rect 23266 5070 23278 5122
rect 30146 5070 30158 5122
rect 30210 5070 30222 5122
rect 30818 5070 30830 5122
rect 30882 5070 30894 5122
rect 35746 5070 35758 5122
rect 35810 5070 35822 5122
rect 39106 5070 39118 5122
rect 39170 5070 39182 5122
rect 39890 5070 39902 5122
rect 39954 5070 39966 5122
rect 27694 5058 27746 5070
rect 14254 5010 14306 5022
rect 30382 5010 30434 5022
rect 21746 4958 21758 5010
rect 21810 4958 21822 5010
rect 22082 4958 22094 5010
rect 22146 4958 22158 5010
rect 23874 4958 23886 5010
rect 23938 4958 23950 5010
rect 27906 4958 27918 5010
rect 27970 4958 27982 5010
rect 28354 4958 28366 5010
rect 28418 4958 28430 5010
rect 35522 4958 35534 5010
rect 35586 4958 35598 5010
rect 14254 4946 14306 4958
rect 30382 4946 30434 4958
rect 22654 4898 22706 4910
rect 22654 4834 22706 4846
rect 27358 4898 27410 4910
rect 27358 4834 27410 4846
rect 34638 4898 34690 4910
rect 34638 4834 34690 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 19630 4562 19682 4574
rect 19630 4498 19682 4510
rect 23886 4562 23938 4574
rect 23886 4498 23938 4510
rect 24334 4562 24386 4574
rect 24334 4498 24386 4510
rect 25566 4562 25618 4574
rect 25566 4498 25618 4510
rect 32510 4562 32562 4574
rect 32510 4498 32562 4510
rect 37326 4562 37378 4574
rect 37326 4498 37378 4510
rect 37774 4562 37826 4574
rect 37774 4498 37826 4510
rect 17390 4450 17442 4462
rect 23550 4450 23602 4462
rect 36990 4450 37042 4462
rect 14690 4398 14702 4450
rect 14754 4398 14766 4450
rect 18722 4398 18734 4450
rect 18786 4398 18798 4450
rect 21074 4398 21086 4450
rect 21138 4398 21150 4450
rect 29922 4398 29934 4450
rect 29986 4398 29998 4450
rect 17390 4386 17442 4398
rect 23550 4386 23602 4398
rect 36990 4386 37042 4398
rect 19294 4338 19346 4350
rect 14018 4286 14030 4338
rect 14082 4286 14094 4338
rect 17602 4286 17614 4338
rect 17666 4286 17678 4338
rect 18498 4286 18510 4338
rect 18562 4286 18574 4338
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 26002 4286 26014 4338
rect 26066 4286 26078 4338
rect 29250 4286 29262 4338
rect 29314 4286 29326 4338
rect 36642 4286 36654 4338
rect 36706 4286 36718 4338
rect 19294 4274 19346 4286
rect 16818 4174 16830 4226
rect 16882 4174 16894 4226
rect 23202 4174 23214 4226
rect 23266 4174 23278 4226
rect 26674 4174 26686 4226
rect 26738 4174 26750 4226
rect 28802 4174 28814 4226
rect 28866 4174 28878 4226
rect 32050 4174 32062 4226
rect 32114 4174 32126 4226
rect 33730 4174 33742 4226
rect 33794 4174 33806 4226
rect 35858 4174 35870 4226
rect 35922 4174 35934 4226
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 17166 3666 17218 3678
rect 17166 3602 17218 3614
rect 20974 3666 21026 3678
rect 20974 3602 21026 3614
rect 22878 3666 22930 3678
rect 22878 3602 22930 3614
rect 27358 3554 27410 3566
rect 34514 3502 34526 3554
rect 34578 3502 34590 3554
rect 27358 3490 27410 3502
rect 27022 3442 27074 3454
rect 27022 3378 27074 3390
rect 34750 3442 34802 3454
rect 34750 3378 34802 3390
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 12574 56814 12626 56866
rect 13358 56814 13410 56866
rect 54238 56814 54290 56866
rect 55022 56814 55074 56866
rect 13470 56590 13522 56642
rect 14814 56590 14866 56642
rect 20190 56590 20242 56642
rect 20750 56590 20802 56642
rect 23662 56590 23714 56642
rect 24670 56590 24722 56642
rect 28702 56590 28754 56642
rect 29374 56590 29426 56642
rect 35422 56590 35474 56642
rect 36766 56590 36818 56642
rect 43038 56590 43090 56642
rect 43598 56590 43650 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4622 56254 4674 56306
rect 5518 56254 5570 56306
rect 6190 56254 6242 56306
rect 7422 56254 7474 56306
rect 8654 56254 8706 56306
rect 10110 56254 10162 56306
rect 11230 56254 11282 56306
rect 12126 56254 12178 56306
rect 14366 56254 14418 56306
rect 18734 56254 18786 56306
rect 31054 56254 31106 56306
rect 35310 56254 35362 56306
rect 36766 56254 36818 56306
rect 39118 56254 39170 56306
rect 40574 56254 40626 56306
rect 41134 56254 41186 56306
rect 44046 56254 44098 56306
rect 45054 56254 45106 56306
rect 46398 56254 46450 56306
rect 47854 56254 47906 56306
rect 49086 56254 49138 56306
rect 50430 56254 50482 56306
rect 51774 56254 51826 56306
rect 53118 56254 53170 56306
rect 55022 56254 55074 56306
rect 55918 56254 55970 56306
rect 5854 56142 5906 56194
rect 15038 56142 15090 56194
rect 17838 56142 17890 56194
rect 23662 56142 23714 56194
rect 41358 56142 41410 56194
rect 41694 56142 41746 56194
rect 42366 56142 42418 56194
rect 14814 56030 14866 56082
rect 15486 56030 15538 56082
rect 15934 56030 15986 56082
rect 18734 56030 18786 56082
rect 21198 56030 21250 56082
rect 22766 56030 22818 56082
rect 24670 56030 24722 56082
rect 28702 56030 28754 56082
rect 30270 56030 30322 56082
rect 32286 56030 32338 56082
rect 34302 56030 34354 56082
rect 36094 56030 36146 56082
rect 37550 56030 37602 56082
rect 39790 56030 39842 56082
rect 42030 56030 42082 56082
rect 4958 55918 5010 55970
rect 6974 55918 7026 55970
rect 8206 55918 8258 55970
rect 9662 55918 9714 55970
rect 10782 55918 10834 55970
rect 11678 55918 11730 55970
rect 12574 55918 12626 55970
rect 13470 55918 13522 55970
rect 13918 55918 13970 55970
rect 16494 55918 16546 55970
rect 19070 55918 19122 55970
rect 20750 55918 20802 55970
rect 21982 55918 22034 55970
rect 25342 55918 25394 55970
rect 27470 55918 27522 55970
rect 29374 55918 29426 55970
rect 32622 55918 32674 55970
rect 34638 55918 34690 55970
rect 37998 55918 38050 55970
rect 42702 55918 42754 55970
rect 43598 55918 43650 55970
rect 44606 55918 44658 55970
rect 45950 55918 46002 55970
rect 47406 55918 47458 55970
rect 48638 55918 48690 55970
rect 49982 55918 50034 55970
rect 51326 55918 51378 55970
rect 52670 55918 52722 55970
rect 54014 55918 54066 55970
rect 55470 55918 55522 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 17054 55470 17106 55522
rect 17614 55470 17666 55522
rect 19630 55470 19682 55522
rect 42254 55470 42306 55522
rect 5070 55358 5122 55410
rect 11678 55358 11730 55410
rect 14702 55358 14754 55410
rect 16494 55358 16546 55410
rect 16718 55358 16770 55410
rect 24222 55358 24274 55410
rect 28590 55358 28642 55410
rect 29598 55358 29650 55410
rect 34302 55358 34354 55410
rect 35086 55358 35138 55410
rect 39902 55358 39954 55410
rect 40686 55358 40738 55410
rect 41582 55358 41634 55410
rect 2158 55246 2210 55298
rect 8766 55246 8818 55298
rect 15374 55246 15426 55298
rect 15598 55246 15650 55298
rect 15934 55246 15986 55298
rect 18398 55246 18450 55298
rect 18958 55246 19010 55298
rect 19854 55246 19906 55298
rect 20302 55246 20354 55298
rect 21422 55246 21474 55298
rect 25678 55246 25730 55298
rect 31502 55246 31554 55298
rect 34750 55246 34802 55298
rect 37102 55246 37154 55298
rect 40238 55246 40290 55298
rect 2942 55134 2994 55186
rect 9550 55134 9602 55186
rect 13694 55134 13746 55186
rect 15038 55134 15090 55186
rect 17502 55134 17554 55186
rect 18846 55134 18898 55186
rect 20638 55134 20690 55186
rect 22094 55134 22146 55186
rect 24558 55134 24610 55186
rect 25342 55134 25394 55186
rect 26462 55134 26514 55186
rect 30942 55134 30994 55186
rect 32174 55134 32226 55186
rect 36206 55134 36258 55186
rect 37774 55134 37826 55186
rect 41806 55134 41858 55186
rect 42702 55134 42754 55186
rect 5966 55022 6018 55074
rect 6302 55022 6354 55074
rect 30382 55022 30434 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 7310 54686 7362 54738
rect 15486 54686 15538 54738
rect 16718 54686 16770 54738
rect 17614 54686 17666 54738
rect 21534 54686 21586 54738
rect 21982 54686 22034 54738
rect 22654 54686 22706 54738
rect 22990 54686 23042 54738
rect 23438 54686 23490 54738
rect 24670 54686 24722 54738
rect 25230 54686 25282 54738
rect 27806 54686 27858 54738
rect 28590 54686 28642 54738
rect 32174 54686 32226 54738
rect 33070 54686 33122 54738
rect 38894 54686 38946 54738
rect 39342 54686 39394 54738
rect 9886 54574 9938 54626
rect 10670 54574 10722 54626
rect 16606 54574 16658 54626
rect 16942 54574 16994 54626
rect 17838 54574 17890 54626
rect 18398 54574 18450 54626
rect 20750 54574 20802 54626
rect 21086 54574 21138 54626
rect 1822 54462 1874 54514
rect 6302 54462 6354 54514
rect 10446 54462 10498 54514
rect 10782 54462 10834 54514
rect 16382 54462 16434 54514
rect 17390 54462 17442 54514
rect 18958 54462 19010 54514
rect 19294 54462 19346 54514
rect 19518 54462 19570 54514
rect 19854 54462 19906 54514
rect 24222 54462 24274 54514
rect 25566 54462 25618 54514
rect 26350 54462 26402 54514
rect 28142 54462 28194 54514
rect 31838 54462 31890 54514
rect 32398 54462 32450 54514
rect 35758 54462 35810 54514
rect 40910 54462 40962 54514
rect 47070 54462 47122 54514
rect 2494 54350 2546 54402
rect 4622 54350 4674 54402
rect 6190 54350 6242 54402
rect 9774 54350 9826 54402
rect 15822 54350 15874 54402
rect 19406 54350 19458 54402
rect 20302 54350 20354 54402
rect 26686 54350 26738 54402
rect 28926 54350 28978 54402
rect 31054 54350 31106 54402
rect 36430 54350 36482 54402
rect 38558 54350 38610 54402
rect 41694 54350 41746 54402
rect 43822 54350 43874 54402
rect 44158 54350 44210 54402
rect 46286 54350 46338 54402
rect 5518 54238 5570 54290
rect 6974 54238 7026 54290
rect 7198 54238 7250 54290
rect 7310 54238 7362 54290
rect 10110 54238 10162 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 17726 53902 17778 53954
rect 19070 53902 19122 53954
rect 21870 53902 21922 53954
rect 2494 53790 2546 53842
rect 3726 53790 3778 53842
rect 5966 53790 6018 53842
rect 8094 53790 8146 53842
rect 9998 53790 10050 53842
rect 16382 53790 16434 53842
rect 18846 53790 18898 53842
rect 20526 53790 20578 53842
rect 23662 53790 23714 53842
rect 34750 53790 34802 53842
rect 37102 53790 37154 53842
rect 41694 53790 41746 53842
rect 42478 53790 42530 53842
rect 44830 53790 44882 53842
rect 50990 53790 51042 53842
rect 3838 53678 3890 53730
rect 8766 53678 8818 53730
rect 12798 53678 12850 53730
rect 13582 53678 13634 53730
rect 21870 53678 21922 53730
rect 22878 53678 22930 53730
rect 23438 53678 23490 53730
rect 24334 53678 24386 53730
rect 24894 53678 24946 53730
rect 29710 53678 29762 53730
rect 30382 53678 30434 53730
rect 31950 53678 32002 53730
rect 36990 53678 37042 53730
rect 38782 53678 38834 53730
rect 42366 53678 42418 53730
rect 43038 53678 43090 53730
rect 43486 53678 43538 53730
rect 47742 53678 47794 53730
rect 48190 53678 48242 53730
rect 2606 53566 2658 53618
rect 2942 53566 2994 53618
rect 12126 53566 12178 53618
rect 14254 53566 14306 53618
rect 18174 53566 18226 53618
rect 19854 53566 19906 53618
rect 21534 53566 21586 53618
rect 27134 53566 27186 53618
rect 28478 53566 28530 53618
rect 29934 53566 29986 53618
rect 30606 53566 30658 53618
rect 32622 53566 32674 53618
rect 35646 53566 35698 53618
rect 35982 53566 36034 53618
rect 39566 53566 39618 53618
rect 46958 53566 47010 53618
rect 48862 53566 48914 53618
rect 2382 53454 2434 53506
rect 16718 53454 16770 53506
rect 17054 53454 17106 53506
rect 23102 53454 23154 53506
rect 23998 53454 24050 53506
rect 29374 53454 29426 53506
rect 42590 53454 42642 53506
rect 43934 53454 43986 53506
rect 51550 53454 51602 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 3278 53118 3330 53170
rect 6638 53118 6690 53170
rect 7198 53118 7250 53170
rect 11678 53118 11730 53170
rect 16046 53118 16098 53170
rect 22430 53118 22482 53170
rect 28366 53118 28418 53170
rect 30494 53118 30546 53170
rect 31278 53118 31330 53170
rect 41470 53118 41522 53170
rect 44158 53118 44210 53170
rect 47070 53118 47122 53170
rect 47518 53118 47570 53170
rect 48078 53118 48130 53170
rect 3502 53006 3554 53058
rect 6078 53006 6130 53058
rect 6190 53006 6242 53058
rect 10110 53006 10162 53058
rect 23662 53006 23714 53058
rect 23886 53006 23938 53058
rect 30718 53006 30770 53058
rect 41358 53006 41410 53058
rect 41582 53006 41634 53058
rect 42030 53006 42082 53058
rect 44382 53006 44434 53058
rect 44494 53006 44546 53058
rect 44830 53006 44882 53058
rect 47966 53006 48018 53058
rect 48750 53006 48802 53058
rect 49870 53006 49922 53058
rect 5854 52894 5906 52946
rect 6862 52894 6914 52946
rect 7310 52894 7362 52946
rect 7422 52894 7474 52946
rect 10558 52894 10610 52946
rect 11454 52894 11506 52946
rect 11678 52894 11730 52946
rect 11902 52894 11954 52946
rect 15822 52894 15874 52946
rect 16158 52894 16210 52946
rect 16606 52894 16658 52946
rect 18286 52894 18338 52946
rect 19182 52894 19234 52946
rect 22878 52894 22930 52946
rect 28030 52894 28082 52946
rect 28590 52894 28642 52946
rect 28926 52894 28978 52946
rect 29150 52894 29202 52946
rect 29598 52894 29650 52946
rect 33182 52894 33234 52946
rect 39006 52894 39058 52946
rect 42142 52894 42194 52946
rect 48974 52894 49026 52946
rect 49422 52894 49474 52946
rect 50206 52894 50258 52946
rect 53790 52894 53842 52946
rect 3166 52782 3218 52834
rect 5182 52782 5234 52834
rect 10446 52782 10498 52834
rect 13134 52782 13186 52834
rect 17950 52782 18002 52834
rect 18734 52782 18786 52834
rect 19854 52782 19906 52834
rect 21982 52782 22034 52834
rect 27806 52782 27858 52834
rect 28814 52782 28866 52834
rect 33854 52782 33906 52834
rect 35982 52782 36034 52834
rect 39454 52782 39506 52834
rect 40462 52782 40514 52834
rect 48190 52782 48242 52834
rect 48862 52782 48914 52834
rect 50878 52782 50930 52834
rect 53006 52782 53058 52834
rect 5070 52670 5122 52722
rect 5406 52670 5458 52722
rect 5518 52670 5570 52722
rect 16270 52670 16322 52722
rect 22990 52670 23042 52722
rect 24222 52670 24274 52722
rect 24558 52670 24610 52722
rect 29822 52670 29874 52722
rect 30046 52670 30098 52722
rect 30942 52670 30994 52722
rect 42030 52670 42082 52722
rect 44942 52670 44994 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 6414 52334 6466 52386
rect 6974 52334 7026 52386
rect 7086 52334 7138 52386
rect 7422 52334 7474 52386
rect 17950 52334 18002 52386
rect 19406 52334 19458 52386
rect 19742 52334 19794 52386
rect 27918 52334 27970 52386
rect 30046 52334 30098 52386
rect 30382 52334 30434 52386
rect 2494 52222 2546 52274
rect 4622 52222 4674 52274
rect 11342 52222 11394 52274
rect 11790 52222 11842 52274
rect 16158 52222 16210 52274
rect 18510 52222 18562 52274
rect 24894 52222 24946 52274
rect 26910 52222 26962 52274
rect 30270 52222 30322 52274
rect 31054 52222 31106 52274
rect 34078 52222 34130 52274
rect 34974 52222 35026 52274
rect 39006 52222 39058 52274
rect 40798 52222 40850 52274
rect 46734 52222 46786 52274
rect 50766 52222 50818 52274
rect 52782 52222 52834 52274
rect 1822 52110 1874 52162
rect 5630 52110 5682 52162
rect 5854 52110 5906 52162
rect 7310 52110 7362 52162
rect 7758 52110 7810 52162
rect 7870 52110 7922 52162
rect 8430 52110 8482 52162
rect 15710 52110 15762 52162
rect 16270 52110 16322 52162
rect 16606 52110 16658 52162
rect 17054 52110 17106 52162
rect 17838 52110 17890 52162
rect 19742 52110 19794 52162
rect 21870 52110 21922 52162
rect 22766 52110 22818 52162
rect 23998 52110 24050 52162
rect 24446 52110 24498 52162
rect 26462 52110 26514 52162
rect 27134 52110 27186 52162
rect 27358 52110 27410 52162
rect 29150 52110 29202 52162
rect 29374 52110 29426 52162
rect 29598 52110 29650 52162
rect 31278 52110 31330 52162
rect 31502 52110 31554 52162
rect 34302 52110 34354 52162
rect 38894 52110 38946 52162
rect 40126 52110 40178 52162
rect 40910 52110 40962 52162
rect 41358 52110 41410 52162
rect 41582 52110 41634 52162
rect 41806 52110 41858 52162
rect 42142 52110 42194 52162
rect 44046 52110 44098 52162
rect 44942 52110 44994 52162
rect 45166 52110 45218 52162
rect 46622 52110 46674 52162
rect 47742 52110 47794 52162
rect 48078 52110 48130 52162
rect 48526 52110 48578 52162
rect 49310 52110 49362 52162
rect 49646 52110 49698 52162
rect 50542 52110 50594 52162
rect 50878 52110 50930 52162
rect 51326 52110 51378 52162
rect 51886 52110 51938 52162
rect 5966 51998 6018 52050
rect 9214 51998 9266 52050
rect 11902 51998 11954 52050
rect 15486 51998 15538 52050
rect 16046 51998 16098 52050
rect 17950 51998 18002 52050
rect 21982 51998 22034 52050
rect 24670 51998 24722 52050
rect 33294 51998 33346 52050
rect 39454 51998 39506 52050
rect 40350 51998 40402 52050
rect 42702 51998 42754 52050
rect 45838 51998 45890 52050
rect 46398 51998 46450 52050
rect 48974 51998 49026 52050
rect 49870 51998 49922 52050
rect 51438 51998 51490 52050
rect 11678 51886 11730 51938
rect 12126 51886 12178 51938
rect 15598 51886 15650 51938
rect 17278 51886 17330 51938
rect 17502 51886 17554 51938
rect 17614 51886 17666 51938
rect 18398 51886 18450 51938
rect 22654 51886 22706 51938
rect 25902 51886 25954 51938
rect 32286 51886 32338 51938
rect 33630 51886 33682 51938
rect 39790 51886 39842 51938
rect 41694 51886 41746 51938
rect 43262 51886 43314 51938
rect 44270 51886 44322 51938
rect 49534 51886 49586 51938
rect 51214 51886 51266 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 5070 51550 5122 51602
rect 6974 51550 7026 51602
rect 7198 51550 7250 51602
rect 9998 51550 10050 51602
rect 11006 51550 11058 51602
rect 16494 51550 16546 51602
rect 22542 51550 22594 51602
rect 27246 51550 27298 51602
rect 28926 51550 28978 51602
rect 32174 51550 32226 51602
rect 33182 51550 33234 51602
rect 33406 51550 33458 51602
rect 33854 51550 33906 51602
rect 34190 51550 34242 51602
rect 39902 51550 39954 51602
rect 41694 51550 41746 51602
rect 43150 51550 43202 51602
rect 46846 51550 46898 51602
rect 48750 51550 48802 51602
rect 4622 51438 4674 51490
rect 5182 51438 5234 51490
rect 6750 51438 6802 51490
rect 10782 51438 10834 51490
rect 12350 51438 12402 51490
rect 16718 51438 16770 51490
rect 16830 51438 16882 51490
rect 23214 51438 23266 51490
rect 23326 51438 23378 51490
rect 23886 51438 23938 51490
rect 25454 51438 25506 51490
rect 25566 51438 25618 51490
rect 26462 51438 26514 51490
rect 27134 51438 27186 51490
rect 27694 51438 27746 51490
rect 28702 51438 28754 51490
rect 31838 51438 31890 51490
rect 32398 51438 32450 51490
rect 36206 51438 36258 51490
rect 37102 51438 37154 51490
rect 39678 51438 39730 51490
rect 40350 51438 40402 51490
rect 40910 51438 40962 51490
rect 41022 51438 41074 51490
rect 43710 51438 43762 51490
rect 47294 51438 47346 51490
rect 51662 51438 51714 51490
rect 51998 51438 52050 51490
rect 4846 51326 4898 51378
rect 5630 51326 5682 51378
rect 5854 51326 5906 51378
rect 6078 51326 6130 51378
rect 9886 51326 9938 51378
rect 10222 51326 10274 51378
rect 10446 51326 10498 51378
rect 11454 51326 11506 51378
rect 12462 51326 12514 51378
rect 13134 51326 13186 51378
rect 17614 51326 17666 51378
rect 18062 51326 18114 51378
rect 19294 51326 19346 51378
rect 23550 51326 23602 51378
rect 23774 51326 23826 51378
rect 28254 51326 28306 51378
rect 31726 51326 31778 51378
rect 32510 51326 32562 51378
rect 33070 51326 33122 51378
rect 35870 51326 35922 51378
rect 36542 51326 36594 51378
rect 37438 51326 37490 51378
rect 37886 51326 37938 51378
rect 38110 51326 38162 51378
rect 39454 51326 39506 51378
rect 40126 51326 40178 51378
rect 41246 51326 41298 51378
rect 41918 51326 41970 51378
rect 42142 51326 42194 51378
rect 42366 51326 42418 51378
rect 42926 51326 42978 51378
rect 43262 51326 43314 51378
rect 45278 51326 45330 51378
rect 45726 51326 45778 51378
rect 48862 51326 48914 51378
rect 49198 51326 49250 51378
rect 49534 51326 49586 51378
rect 50766 51326 50818 51378
rect 51886 51326 51938 51378
rect 53902 51326 53954 51378
rect 13918 51214 13970 51266
rect 16046 51214 16098 51266
rect 17390 51214 17442 51266
rect 19966 51214 20018 51266
rect 22094 51214 22146 51266
rect 26350 51214 26402 51266
rect 27806 51214 27858 51266
rect 29038 51214 29090 51266
rect 39230 51214 39282 51266
rect 41806 51214 41858 51266
rect 47966 51214 48018 51266
rect 50094 51214 50146 51266
rect 50878 51214 50930 51266
rect 52558 51214 52610 51266
rect 53342 51214 53394 51266
rect 6190 51102 6242 51154
rect 7310 51102 7362 51154
rect 23886 51102 23938 51154
rect 25566 51102 25618 51154
rect 26686 51102 26738 51154
rect 27358 51102 27410 51154
rect 28030 51102 28082 51154
rect 31838 51102 31890 51154
rect 37662 51102 37714 51154
rect 38558 51102 38610 51154
rect 39902 51102 39954 51154
rect 49086 51102 49138 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 15598 50766 15650 50818
rect 16046 50766 16098 50818
rect 16830 50766 16882 50818
rect 25566 50766 25618 50818
rect 25902 50766 25954 50818
rect 27134 50766 27186 50818
rect 27470 50766 27522 50818
rect 28142 50766 28194 50818
rect 28590 50766 28642 50818
rect 30382 50766 30434 50818
rect 38670 50766 38722 50818
rect 39006 50766 39058 50818
rect 50766 50766 50818 50818
rect 4622 50654 4674 50706
rect 6414 50654 6466 50706
rect 11342 50654 11394 50706
rect 15934 50654 15986 50706
rect 18174 50654 18226 50706
rect 20078 50654 20130 50706
rect 22766 50654 22818 50706
rect 28478 50654 28530 50706
rect 31838 50654 31890 50706
rect 32510 50654 32562 50706
rect 36430 50654 36482 50706
rect 37998 50654 38050 50706
rect 40238 50654 40290 50706
rect 46734 50654 46786 50706
rect 49422 50654 49474 50706
rect 54462 50654 54514 50706
rect 1822 50542 1874 50594
rect 5742 50542 5794 50594
rect 10894 50542 10946 50594
rect 11230 50542 11282 50594
rect 11454 50542 11506 50594
rect 11902 50542 11954 50594
rect 12238 50542 12290 50594
rect 16270 50542 16322 50594
rect 16606 50542 16658 50594
rect 17054 50542 17106 50594
rect 17726 50542 17778 50594
rect 18958 50542 19010 50594
rect 19966 50542 20018 50594
rect 21534 50542 21586 50594
rect 22654 50542 22706 50594
rect 23774 50542 23826 50594
rect 23998 50542 24050 50594
rect 24110 50542 24162 50594
rect 26798 50542 26850 50594
rect 27134 50542 27186 50594
rect 28254 50542 28306 50594
rect 29710 50542 29762 50594
rect 30270 50542 30322 50594
rect 31278 50542 31330 50594
rect 32174 50542 32226 50594
rect 33630 50542 33682 50594
rect 40014 50542 40066 50594
rect 40686 50542 40738 50594
rect 41694 50542 41746 50594
rect 42478 50542 42530 50594
rect 44158 50542 44210 50594
rect 46510 50542 46562 50594
rect 46846 50542 46898 50594
rect 50878 50542 50930 50594
rect 51102 50542 51154 50594
rect 51326 50542 51378 50594
rect 52782 50542 52834 50594
rect 53006 50542 53058 50594
rect 54574 50542 54626 50594
rect 54910 50542 54962 50594
rect 2494 50430 2546 50482
rect 9774 50430 9826 50482
rect 10110 50430 10162 50482
rect 10782 50430 10834 50482
rect 12462 50430 12514 50482
rect 17390 50430 17442 50482
rect 18846 50430 18898 50482
rect 19294 50430 19346 50482
rect 22430 50430 22482 50482
rect 24558 50430 24610 50482
rect 25342 50430 25394 50482
rect 26238 50430 26290 50482
rect 29150 50430 29202 50482
rect 29934 50430 29986 50482
rect 30494 50430 30546 50482
rect 30942 50430 30994 50482
rect 31502 50430 31554 50482
rect 33182 50430 33234 50482
rect 34302 50430 34354 50482
rect 37550 50430 37602 50482
rect 38446 50430 38498 50482
rect 39566 50430 39618 50482
rect 39790 50430 39842 50482
rect 40350 50430 40402 50482
rect 41918 50430 41970 50482
rect 42702 50430 42754 50482
rect 43262 50430 43314 50482
rect 43822 50430 43874 50482
rect 44046 50430 44098 50482
rect 45390 50430 45442 50482
rect 47406 50430 47458 50482
rect 49534 50430 49586 50482
rect 49870 50430 49922 50482
rect 50318 50430 50370 50482
rect 51774 50430 51826 50482
rect 8654 50318 8706 50370
rect 16382 50318 16434 50370
rect 21310 50318 21362 50370
rect 22878 50318 22930 50370
rect 29262 50318 29314 50370
rect 30718 50318 30770 50370
rect 31726 50318 31778 50370
rect 31838 50318 31890 50370
rect 32510 50318 32562 50370
rect 32734 50318 32786 50370
rect 33070 50318 33122 50370
rect 41806 50318 41858 50370
rect 43598 50318 43650 50370
rect 49086 50318 49138 50370
rect 49310 50318 49362 50370
rect 49982 50318 50034 50370
rect 50094 50318 50146 50370
rect 53342 50318 53394 50370
rect 55022 50318 55074 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 2046 49982 2098 50034
rect 2158 49982 2210 50034
rect 6302 49982 6354 50034
rect 7646 49982 7698 50034
rect 9662 49982 9714 50034
rect 17390 49982 17442 50034
rect 19070 49982 19122 50034
rect 22430 49982 22482 50034
rect 26574 49982 26626 50034
rect 28814 49982 28866 50034
rect 29486 49982 29538 50034
rect 32622 49982 32674 50034
rect 33070 49982 33122 50034
rect 33182 49982 33234 50034
rect 40238 49982 40290 50034
rect 40798 49982 40850 50034
rect 42702 49982 42754 50034
rect 46286 49982 46338 50034
rect 4958 49870 5010 49922
rect 6414 49870 6466 49922
rect 9550 49870 9602 49922
rect 10670 49870 10722 49922
rect 16606 49870 16658 49922
rect 19518 49870 19570 49922
rect 22542 49870 22594 49922
rect 23886 49870 23938 49922
rect 24446 49870 24498 49922
rect 24782 49870 24834 49922
rect 27358 49870 27410 49922
rect 27582 49870 27634 49922
rect 28030 49870 28082 49922
rect 30382 49870 30434 49922
rect 31278 49870 31330 49922
rect 33294 49870 33346 49922
rect 33406 49870 33458 49922
rect 33630 49870 33682 49922
rect 36542 49870 36594 49922
rect 37326 49870 37378 49922
rect 40126 49870 40178 49922
rect 42590 49870 42642 49922
rect 43150 49870 43202 49922
rect 44606 49870 44658 49922
rect 45278 49870 45330 49922
rect 45614 49870 45666 49922
rect 47966 49870 48018 49922
rect 50206 49870 50258 49922
rect 56702 49870 56754 49922
rect 2270 49758 2322 49810
rect 2606 49758 2658 49810
rect 3502 49758 3554 49810
rect 4846 49758 4898 49810
rect 5854 49758 5906 49810
rect 6974 49758 7026 49810
rect 7086 49758 7138 49810
rect 7198 49758 7250 49810
rect 11006 49758 11058 49810
rect 11566 49758 11618 49810
rect 11902 49758 11954 49810
rect 12350 49758 12402 49810
rect 12462 49758 12514 49810
rect 12574 49758 12626 49810
rect 12798 49758 12850 49810
rect 16830 49758 16882 49810
rect 17726 49758 17778 49810
rect 18734 49758 18786 49810
rect 18958 49758 19010 49810
rect 19182 49758 19234 49810
rect 19742 49758 19794 49810
rect 20078 49758 20130 49810
rect 20638 49758 20690 49810
rect 21310 49758 21362 49810
rect 21646 49758 21698 49810
rect 21870 49758 21922 49810
rect 22206 49758 22258 49810
rect 23662 49758 23714 49810
rect 26126 49758 26178 49810
rect 26238 49758 26290 49810
rect 27470 49758 27522 49810
rect 28254 49758 28306 49810
rect 28702 49758 28754 49810
rect 28926 49758 28978 49810
rect 29374 49758 29426 49810
rect 29598 49758 29650 49810
rect 30046 49758 30098 49810
rect 30606 49758 30658 49810
rect 31166 49758 31218 49810
rect 32062 49758 32114 49810
rect 34414 49758 34466 49810
rect 37886 49758 37938 49810
rect 38670 49758 38722 49810
rect 41470 49758 41522 49810
rect 41806 49758 41858 49810
rect 43598 49758 43650 49810
rect 44046 49758 44098 49810
rect 45950 49758 46002 49810
rect 46286 49758 46338 49810
rect 46622 49758 46674 49810
rect 46846 49758 46898 49810
rect 46958 49758 47010 49810
rect 47070 49758 47122 49810
rect 47518 49758 47570 49810
rect 48750 49758 48802 49810
rect 49310 49758 49362 49810
rect 49646 49758 49698 49810
rect 51550 49758 51602 49810
rect 51774 49758 51826 49810
rect 52670 49758 52722 49810
rect 53118 49758 53170 49810
rect 53790 49758 53842 49810
rect 54574 49758 54626 49810
rect 54686 49758 54738 49810
rect 55246 49758 55298 49810
rect 56478 49758 56530 49810
rect 56814 49758 56866 49810
rect 3390 49646 3442 49698
rect 17950 49646 18002 49698
rect 19966 49646 20018 49698
rect 26686 49646 26738 49698
rect 34190 49646 34242 49698
rect 36654 49646 36706 49698
rect 39230 49646 39282 49698
rect 41918 49646 41970 49698
rect 44158 49646 44210 49698
rect 48078 49646 48130 49698
rect 50094 49646 50146 49698
rect 50878 49646 50930 49698
rect 52782 49646 52834 49698
rect 54126 49646 54178 49698
rect 54462 49646 54514 49698
rect 9662 49534 9714 49586
rect 11454 49534 11506 49586
rect 11790 49534 11842 49586
rect 16494 49534 16546 49586
rect 36318 49534 36370 49586
rect 40350 49534 40402 49586
rect 48190 49534 48242 49586
rect 48862 49534 48914 49586
rect 49086 49534 49138 49586
rect 49870 49534 49922 49586
rect 53006 49534 53058 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 2718 49198 2770 49250
rect 18846 49198 18898 49250
rect 20190 49198 20242 49250
rect 23662 49198 23714 49250
rect 26574 49198 26626 49250
rect 27806 49198 27858 49250
rect 29262 49198 29314 49250
rect 45502 49198 45554 49250
rect 47294 49198 47346 49250
rect 52894 49198 52946 49250
rect 5742 49086 5794 49138
rect 10334 49086 10386 49138
rect 17166 49086 17218 49138
rect 26798 49086 26850 49138
rect 28590 49086 28642 49138
rect 29822 49086 29874 49138
rect 30830 49086 30882 49138
rect 32174 49086 32226 49138
rect 37214 49086 37266 49138
rect 40238 49086 40290 49138
rect 42590 49086 42642 49138
rect 47182 49086 47234 49138
rect 48750 49086 48802 49138
rect 51102 49086 51154 49138
rect 51662 49086 51714 49138
rect 51998 49086 52050 49138
rect 56702 49086 56754 49138
rect 57486 49086 57538 49138
rect 4734 48974 4786 49026
rect 5966 48974 6018 49026
rect 6190 48974 6242 49026
rect 9774 48974 9826 49026
rect 9998 48974 10050 49026
rect 12014 48974 12066 49026
rect 12238 48974 12290 49026
rect 12798 48974 12850 49026
rect 14366 48974 14418 49026
rect 18622 48974 18674 49026
rect 19070 48974 19122 49026
rect 19518 48974 19570 49026
rect 19630 48974 19682 49026
rect 19742 48974 19794 49026
rect 21310 48974 21362 49026
rect 21534 48974 21586 49026
rect 21870 48974 21922 49026
rect 22094 48974 22146 49026
rect 22990 48974 23042 49026
rect 25678 48974 25730 49026
rect 26238 48974 26290 49026
rect 26910 48974 26962 49026
rect 27134 48974 27186 49026
rect 28254 48974 28306 49026
rect 29934 48974 29986 49026
rect 31390 48974 31442 49026
rect 31726 48974 31778 49026
rect 31950 48974 32002 49026
rect 32286 48974 32338 49026
rect 32734 48974 32786 49026
rect 36542 48974 36594 49026
rect 39006 48974 39058 49026
rect 40014 48974 40066 49026
rect 40350 48974 40402 49026
rect 42142 48974 42194 49026
rect 42478 48974 42530 49026
rect 43822 48974 43874 49026
rect 43934 48974 43986 49026
rect 44382 48974 44434 49026
rect 44942 48974 44994 49026
rect 45614 48974 45666 49026
rect 46286 48974 46338 49026
rect 46622 48974 46674 49026
rect 47966 48974 48018 49026
rect 48414 48974 48466 49026
rect 50542 48974 50594 49026
rect 52110 48974 52162 49026
rect 52670 48974 52722 49026
rect 53118 48974 53170 49026
rect 53454 48974 53506 49026
rect 53902 48974 53954 49026
rect 57038 48974 57090 49026
rect 2942 48862 2994 48914
rect 3502 48862 3554 48914
rect 4398 48862 4450 48914
rect 5630 48862 5682 48914
rect 10670 48862 10722 48914
rect 10894 48862 10946 48914
rect 11902 48862 11954 48914
rect 15038 48862 15090 48914
rect 18510 48862 18562 48914
rect 22430 48862 22482 48914
rect 22878 48862 22930 48914
rect 23998 48862 24050 48914
rect 28030 48862 28082 48914
rect 29374 48862 29426 48914
rect 30158 48862 30210 48914
rect 30942 48862 30994 48914
rect 36206 48862 36258 48914
rect 36318 48862 36370 48914
rect 41246 48862 41298 48914
rect 45166 48862 45218 48914
rect 46174 48862 46226 48914
rect 53342 48862 53394 48914
rect 54574 48862 54626 48914
rect 2830 48750 2882 48802
rect 3838 48750 3890 48802
rect 10782 48750 10834 48802
rect 11454 48750 11506 48802
rect 12574 48750 12626 48802
rect 17502 48750 17554 48802
rect 17838 48750 17890 48802
rect 20750 48750 20802 48802
rect 21422 48750 21474 48802
rect 22318 48750 22370 48802
rect 27470 48750 27522 48802
rect 27694 48750 27746 48802
rect 28478 48750 28530 48802
rect 29262 48750 29314 48802
rect 29710 48750 29762 48802
rect 30606 48750 30658 48802
rect 30830 48750 30882 48802
rect 32958 48750 33010 48802
rect 35870 48750 35922 48802
rect 44158 48750 44210 48802
rect 45726 48750 45778 48802
rect 46062 48750 46114 48802
rect 47070 48750 47122 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 6974 48414 7026 48466
rect 11118 48414 11170 48466
rect 20974 48414 21026 48466
rect 26238 48414 26290 48466
rect 26574 48414 26626 48466
rect 32062 48414 32114 48466
rect 39678 48414 39730 48466
rect 44382 48414 44434 48466
rect 45166 48414 45218 48466
rect 45726 48414 45778 48466
rect 46062 48414 46114 48466
rect 46174 48414 46226 48466
rect 48862 48414 48914 48466
rect 49310 48414 49362 48466
rect 49870 48414 49922 48466
rect 50542 48414 50594 48466
rect 2494 48302 2546 48354
rect 6638 48302 6690 48354
rect 7982 48302 8034 48354
rect 8094 48302 8146 48354
rect 8766 48302 8818 48354
rect 13582 48302 13634 48354
rect 16046 48302 16098 48354
rect 20526 48302 20578 48354
rect 22542 48302 22594 48354
rect 27022 48302 27074 48354
rect 28254 48302 28306 48354
rect 31950 48302 32002 48354
rect 39230 48302 39282 48354
rect 40350 48302 40402 48354
rect 42478 48302 42530 48354
rect 45054 48302 45106 48354
rect 49646 48302 49698 48354
rect 54014 48302 54066 48354
rect 1822 48190 1874 48242
rect 5630 48190 5682 48242
rect 5854 48190 5906 48242
rect 8318 48190 8370 48242
rect 9998 48190 10050 48242
rect 14366 48190 14418 48242
rect 14814 48190 14866 48242
rect 16158 48190 16210 48242
rect 16382 48190 16434 48242
rect 16606 48190 16658 48242
rect 17950 48190 18002 48242
rect 20862 48190 20914 48242
rect 21086 48190 21138 48242
rect 21870 48190 21922 48242
rect 27358 48190 27410 48242
rect 28142 48190 28194 48242
rect 31054 48190 31106 48242
rect 31614 48190 31666 48242
rect 37998 48190 38050 48242
rect 39006 48190 39058 48242
rect 39118 48190 39170 48242
rect 40126 48190 40178 48242
rect 40910 48190 40962 48242
rect 42142 48190 42194 48242
rect 42702 48190 42754 48242
rect 43822 48190 43874 48242
rect 44158 48190 44210 48242
rect 44382 48190 44434 48242
rect 44606 48190 44658 48242
rect 45950 48190 46002 48242
rect 46622 48190 46674 48242
rect 47182 48190 47234 48242
rect 50990 48190 51042 48242
rect 51326 48190 51378 48242
rect 52334 48190 52386 48242
rect 52782 48190 52834 48242
rect 53566 48190 53618 48242
rect 53790 48190 53842 48242
rect 57038 48190 57090 48242
rect 4622 48078 4674 48130
rect 8878 48078 8930 48130
rect 9886 48078 9938 48130
rect 10558 48078 10610 48130
rect 11454 48078 11506 48130
rect 19742 48078 19794 48130
rect 24670 48078 24722 48130
rect 27246 48078 27298 48130
rect 29038 48078 29090 48130
rect 35646 48078 35698 48130
rect 36206 48078 36258 48130
rect 45278 48078 45330 48130
rect 48078 48078 48130 48130
rect 51886 48078 51938 48130
rect 53230 48078 53282 48130
rect 53678 48078 53730 48130
rect 54574 48078 54626 48130
rect 56590 48078 56642 48130
rect 6190 47966 6242 48018
rect 8990 47966 9042 48018
rect 9550 47966 9602 48018
rect 9662 47966 9714 48018
rect 10782 47966 10834 48018
rect 21086 47966 21138 48018
rect 32062 47966 32114 48018
rect 49982 47966 50034 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 5070 47630 5122 47682
rect 10894 47630 10946 47682
rect 20190 47630 20242 47682
rect 20526 47630 20578 47682
rect 21646 47630 21698 47682
rect 22206 47630 22258 47682
rect 22542 47630 22594 47682
rect 28254 47630 28306 47682
rect 28590 47630 28642 47682
rect 31278 47630 31330 47682
rect 49534 47630 49586 47682
rect 50206 47630 50258 47682
rect 50318 47630 50370 47682
rect 50542 47630 50594 47682
rect 50654 47630 50706 47682
rect 51102 47630 51154 47682
rect 51438 47630 51490 47682
rect 51774 47630 51826 47682
rect 5742 47518 5794 47570
rect 7758 47518 7810 47570
rect 9886 47518 9938 47570
rect 11230 47518 11282 47570
rect 11790 47518 11842 47570
rect 17278 47518 17330 47570
rect 19406 47518 19458 47570
rect 19854 47518 19906 47570
rect 30830 47518 30882 47570
rect 31166 47518 31218 47570
rect 36318 47518 36370 47570
rect 38558 47518 38610 47570
rect 39566 47518 39618 47570
rect 42142 47518 42194 47570
rect 43038 47518 43090 47570
rect 43374 47518 43426 47570
rect 43822 47518 43874 47570
rect 44158 47518 44210 47570
rect 45502 47518 45554 47570
rect 47966 47518 48018 47570
rect 51998 47518 52050 47570
rect 57598 47518 57650 47570
rect 4958 47406 5010 47458
rect 5966 47406 6018 47458
rect 6078 47406 6130 47458
rect 6974 47406 7026 47458
rect 11006 47406 11058 47458
rect 12014 47406 12066 47458
rect 12238 47406 12290 47458
rect 12574 47406 12626 47458
rect 15934 47406 15986 47458
rect 16606 47406 16658 47458
rect 20750 47406 20802 47458
rect 21422 47406 21474 47458
rect 21758 47406 21810 47458
rect 28030 47406 28082 47458
rect 29262 47406 29314 47458
rect 29822 47406 29874 47458
rect 33518 47406 33570 47458
rect 37102 47406 37154 47458
rect 37438 47406 37490 47458
rect 38894 47406 38946 47458
rect 40014 47406 40066 47458
rect 41022 47406 41074 47458
rect 42926 47406 42978 47458
rect 44270 47406 44322 47458
rect 45838 47406 45890 47458
rect 46174 47406 46226 47458
rect 46286 47406 46338 47458
rect 47070 47406 47122 47458
rect 48078 47406 48130 47458
rect 48750 47406 48802 47458
rect 48974 47406 49026 47458
rect 49310 47406 49362 47458
rect 49758 47406 49810 47458
rect 52110 47406 52162 47458
rect 52670 47406 52722 47458
rect 53006 47406 53058 47458
rect 53230 47406 53282 47458
rect 54798 47406 54850 47458
rect 4846 47294 4898 47346
rect 5630 47294 5682 47346
rect 11342 47294 11394 47346
rect 11678 47294 11730 47346
rect 16158 47294 16210 47346
rect 22318 47294 22370 47346
rect 34190 47294 34242 47346
rect 40350 47294 40402 47346
rect 41246 47294 41298 47346
rect 41806 47294 41858 47346
rect 47742 47294 47794 47346
rect 53790 47294 53842 47346
rect 55470 47294 55522 47346
rect 12686 47182 12738 47234
rect 12798 47182 12850 47234
rect 21758 47182 21810 47234
rect 22990 47182 23042 47234
rect 44942 47182 44994 47234
rect 46398 47182 46450 47234
rect 48526 47182 48578 47234
rect 48862 47182 48914 47234
rect 49422 47182 49474 47234
rect 51326 47182 51378 47234
rect 52894 47182 52946 47234
rect 53454 47182 53506 47234
rect 53678 47182 53730 47234
rect 54238 47182 54290 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 8990 46846 9042 46898
rect 15262 46846 15314 46898
rect 20302 46846 20354 46898
rect 20638 46846 20690 46898
rect 37102 46846 37154 46898
rect 37550 46846 37602 46898
rect 39678 46846 39730 46898
rect 39790 46846 39842 46898
rect 41918 46846 41970 46898
rect 42478 46846 42530 46898
rect 44382 46846 44434 46898
rect 45054 46846 45106 46898
rect 45278 46846 45330 46898
rect 52110 46846 52162 46898
rect 2942 46734 2994 46786
rect 6862 46734 6914 46786
rect 7310 46734 7362 46786
rect 14030 46734 14082 46786
rect 23662 46734 23714 46786
rect 31726 46734 31778 46786
rect 36766 46734 36818 46786
rect 38334 46734 38386 46786
rect 38670 46734 38722 46786
rect 39006 46734 39058 46786
rect 39230 46734 39282 46786
rect 41246 46734 41298 46786
rect 51662 46734 51714 46786
rect 2270 46622 2322 46674
rect 5518 46622 5570 46674
rect 5966 46622 6018 46674
rect 6302 46622 6354 46674
rect 7646 46622 7698 46674
rect 8430 46622 8482 46674
rect 8654 46622 8706 46674
rect 10222 46622 10274 46674
rect 10558 46622 10610 46674
rect 14814 46622 14866 46674
rect 17950 46622 18002 46674
rect 24334 46622 24386 46674
rect 28142 46622 28194 46674
rect 31390 46622 31442 46674
rect 32062 46622 32114 46674
rect 35870 46622 35922 46674
rect 36318 46622 36370 46674
rect 37550 46622 37602 46674
rect 37998 46622 38050 46674
rect 39566 46622 39618 46674
rect 40238 46622 40290 46674
rect 40910 46622 40962 46674
rect 41806 46622 41858 46674
rect 42702 46622 42754 46674
rect 42926 46622 42978 46674
rect 43262 46622 43314 46674
rect 44606 46622 44658 46674
rect 45614 46622 45666 46674
rect 49646 46622 49698 46674
rect 50206 46622 50258 46674
rect 51102 46622 51154 46674
rect 51886 46622 51938 46674
rect 52222 46622 52274 46674
rect 52558 46622 52610 46674
rect 52894 46622 52946 46674
rect 53230 46622 53282 46674
rect 53454 46622 53506 46674
rect 53678 46622 53730 46674
rect 54126 46622 54178 46674
rect 55358 46622 55410 46674
rect 57710 46622 57762 46674
rect 5070 46510 5122 46562
rect 8094 46510 8146 46562
rect 9774 46510 9826 46562
rect 11902 46510 11954 46562
rect 19630 46510 19682 46562
rect 21310 46510 21362 46562
rect 21534 46510 21586 46562
rect 25230 46510 25282 46562
rect 27358 46510 27410 46562
rect 28590 46510 28642 46562
rect 31054 46510 31106 46562
rect 32286 46510 32338 46562
rect 35534 46510 35586 46562
rect 37886 46510 37938 46562
rect 38782 46510 38834 46562
rect 42814 46510 42866 46562
rect 43710 46510 43762 46562
rect 45166 46510 45218 46562
rect 47966 46510 48018 46562
rect 49870 46510 49922 46562
rect 50766 46510 50818 46562
rect 53006 46510 53058 46562
rect 53902 46510 53954 46562
rect 54462 46510 54514 46562
rect 54910 46510 54962 46562
rect 57150 46510 57202 46562
rect 5406 46398 5458 46450
rect 5742 46398 5794 46450
rect 6526 46398 6578 46450
rect 7646 46398 7698 46450
rect 10334 46398 10386 46450
rect 32398 46398 32450 46450
rect 35982 46398 36034 46450
rect 36430 46398 36482 46450
rect 50654 46398 50706 46450
rect 54350 46398 54402 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 5070 46062 5122 46114
rect 17278 46062 17330 46114
rect 25790 46062 25842 46114
rect 38446 46062 38498 46114
rect 39566 46062 39618 46114
rect 4958 45950 5010 46002
rect 6974 45950 7026 46002
rect 10110 45950 10162 46002
rect 16942 45950 16994 46002
rect 17614 45950 17666 46002
rect 17838 45950 17890 46002
rect 18622 45950 18674 46002
rect 20414 45950 20466 46002
rect 32622 45950 32674 46002
rect 34750 45950 34802 46002
rect 35198 45950 35250 46002
rect 36542 45950 36594 46002
rect 37214 45950 37266 46002
rect 40014 45950 40066 46002
rect 43934 45950 43986 46002
rect 48638 45950 48690 46002
rect 50206 45950 50258 46002
rect 52670 45950 52722 46002
rect 57822 45950 57874 46002
rect 8766 45838 8818 45890
rect 9774 45838 9826 45890
rect 12238 45838 12290 45890
rect 14142 45838 14194 45890
rect 18958 45838 19010 45890
rect 19518 45838 19570 45890
rect 25790 45838 25842 45890
rect 29822 45838 29874 45890
rect 31950 45838 32002 45890
rect 37326 45838 37378 45890
rect 37550 45838 37602 45890
rect 37774 45838 37826 45890
rect 38670 45838 38722 45890
rect 39230 45838 39282 45890
rect 41806 45838 41858 45890
rect 42142 45838 42194 45890
rect 42478 45838 42530 45890
rect 43038 45838 43090 45890
rect 45614 45838 45666 45890
rect 45726 45838 45778 45890
rect 46286 45838 46338 45890
rect 49534 45838 49586 45890
rect 50094 45838 50146 45890
rect 50766 45838 50818 45890
rect 50878 45838 50930 45890
rect 51102 45838 51154 45890
rect 51326 45838 51378 45890
rect 53454 45838 53506 45890
rect 53902 45838 53954 45890
rect 54126 45838 54178 45890
rect 54350 45838 54402 45890
rect 54910 45838 54962 45890
rect 4846 45726 4898 45778
rect 9662 45726 9714 45778
rect 10670 45726 10722 45778
rect 14814 45726 14866 45778
rect 25454 45726 25506 45778
rect 30158 45726 30210 45778
rect 38110 45726 38162 45778
rect 39006 45726 39058 45778
rect 41582 45726 41634 45778
rect 45838 45726 45890 45778
rect 53006 45726 53058 45778
rect 53678 45726 53730 45778
rect 55694 45726 55746 45778
rect 19070 45614 19122 45666
rect 19182 45614 19234 45666
rect 20078 45614 20130 45666
rect 21422 45614 21474 45666
rect 21870 45614 21922 45666
rect 25118 45614 25170 45666
rect 26238 45614 26290 45666
rect 26686 45614 26738 45666
rect 37102 45614 37154 45666
rect 40462 45614 40514 45666
rect 41246 45614 41298 45666
rect 42142 45614 42194 45666
rect 42814 45614 42866 45666
rect 44270 45614 44322 45666
rect 45166 45614 45218 45666
rect 50542 45614 50594 45666
rect 51774 45614 51826 45666
rect 52782 45614 52834 45666
rect 54462 45614 54514 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 8878 45278 8930 45330
rect 9662 45278 9714 45330
rect 11118 45278 11170 45330
rect 25902 45278 25954 45330
rect 33182 45278 33234 45330
rect 34638 45278 34690 45330
rect 37886 45278 37938 45330
rect 37998 45278 38050 45330
rect 38782 45278 38834 45330
rect 41246 45278 41298 45330
rect 42142 45278 42194 45330
rect 42366 45278 42418 45330
rect 43150 45278 43202 45330
rect 43486 45278 43538 45330
rect 44270 45278 44322 45330
rect 45950 45278 46002 45330
rect 48862 45278 48914 45330
rect 49758 45278 49810 45330
rect 5070 45166 5122 45218
rect 10222 45166 10274 45218
rect 13358 45166 13410 45218
rect 18734 45166 18786 45218
rect 34862 45166 34914 45218
rect 38670 45166 38722 45218
rect 49982 45166 50034 45218
rect 50766 45166 50818 45218
rect 55582 45166 55634 45218
rect 56590 45166 56642 45218
rect 4398 45054 4450 45106
rect 8094 45054 8146 45106
rect 8430 45054 8482 45106
rect 14142 45054 14194 45106
rect 14590 45054 14642 45106
rect 18062 45054 18114 45106
rect 21198 45054 21250 45106
rect 26350 45054 26402 45106
rect 29598 45054 29650 45106
rect 34414 45054 34466 45106
rect 34526 45054 34578 45106
rect 35310 45054 35362 45106
rect 37774 45054 37826 45106
rect 38446 45054 38498 45106
rect 39006 45054 39058 45106
rect 41022 45054 41074 45106
rect 42254 45054 42306 45106
rect 42814 45054 42866 45106
rect 43038 45054 43090 45106
rect 43262 45054 43314 45106
rect 44158 45054 44210 45106
rect 44494 45054 44546 45106
rect 44718 45054 44770 45106
rect 44942 45054 44994 45106
rect 45166 45054 45218 45106
rect 45390 45054 45442 45106
rect 51102 45054 51154 45106
rect 52670 45054 52722 45106
rect 53566 45054 53618 45106
rect 53790 45054 53842 45106
rect 54126 45054 54178 45106
rect 55358 45054 55410 45106
rect 57150 45054 57202 45106
rect 7198 44942 7250 44994
rect 8542 44942 8594 44994
rect 17502 44942 17554 44994
rect 20862 44942 20914 44994
rect 21982 44942 22034 44994
rect 24110 44942 24162 44994
rect 25342 44942 25394 44994
rect 27134 44942 27186 44994
rect 29262 44942 29314 44994
rect 30382 44942 30434 44994
rect 32510 44942 32562 44994
rect 36878 44942 36930 44994
rect 39454 44942 39506 44994
rect 45278 44942 45330 44994
rect 46398 44942 46450 44994
rect 48750 44942 48802 44994
rect 49646 44942 49698 44994
rect 51214 44942 51266 44994
rect 54686 44942 54738 44994
rect 55022 44942 55074 44994
rect 57374 44942 57426 44994
rect 25678 44830 25730 44882
rect 26014 44830 26066 44882
rect 35422 44830 35474 44882
rect 49086 44830 49138 44882
rect 52894 44830 52946 44882
rect 53342 44830 53394 44882
rect 54350 44830 54402 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 11790 44494 11842 44546
rect 53342 44494 53394 44546
rect 55582 44494 55634 44546
rect 7422 44382 7474 44434
rect 9550 44382 9602 44434
rect 12126 44382 12178 44434
rect 12798 44382 12850 44434
rect 14814 44382 14866 44434
rect 19518 44382 19570 44434
rect 21422 44382 21474 44434
rect 22206 44382 22258 44434
rect 25454 44382 25506 44434
rect 27582 44382 27634 44434
rect 31054 44382 31106 44434
rect 32510 44382 32562 44434
rect 38222 44382 38274 44434
rect 43038 44382 43090 44434
rect 43374 44382 43426 44434
rect 57262 44382 57314 44434
rect 7310 44270 7362 44322
rect 7870 44270 7922 44322
rect 8318 44270 8370 44322
rect 10334 44270 10386 44322
rect 15150 44270 15202 44322
rect 16046 44270 16098 44322
rect 16718 44270 16770 44322
rect 20414 44270 20466 44322
rect 22430 44270 22482 44322
rect 23326 44270 23378 44322
rect 28366 44270 28418 44322
rect 31390 44270 31442 44322
rect 32174 44270 32226 44322
rect 33294 44270 33346 44322
rect 34302 44270 34354 44322
rect 34862 44270 34914 44322
rect 35198 44270 35250 44322
rect 35982 44270 36034 44322
rect 37102 44270 37154 44322
rect 37662 44270 37714 44322
rect 37774 44270 37826 44322
rect 38670 44270 38722 44322
rect 40798 44270 40850 44322
rect 42478 44270 42530 44322
rect 43934 44270 43986 44322
rect 46062 44270 46114 44322
rect 48078 44270 48130 44322
rect 49310 44270 49362 44322
rect 50430 44270 50482 44322
rect 53118 44270 53170 44322
rect 53678 44270 53730 44322
rect 53902 44270 53954 44322
rect 54798 44270 54850 44322
rect 55358 44270 55410 44322
rect 56366 44270 56418 44322
rect 56814 44270 56866 44322
rect 57486 44270 57538 44322
rect 57598 44270 57650 44322
rect 7198 44158 7250 44210
rect 9886 44158 9938 44210
rect 10558 44158 10610 44210
rect 12350 44158 12402 44210
rect 16270 44158 16322 44210
rect 17390 44158 17442 44210
rect 19854 44158 19906 44210
rect 20190 44158 20242 44210
rect 22094 44158 22146 44210
rect 22990 44158 23042 44210
rect 32846 44158 32898 44210
rect 34638 44158 34690 44210
rect 35310 44158 35362 44210
rect 38110 44158 38162 44210
rect 38446 44158 38498 44210
rect 43486 44158 43538 44210
rect 43822 44158 43874 44210
rect 45726 44158 45778 44210
rect 48974 44158 49026 44210
rect 50318 44158 50370 44210
rect 50766 44158 50818 44210
rect 50878 44158 50930 44210
rect 51102 44158 51154 44210
rect 55022 44158 55074 44210
rect 56254 44158 56306 44210
rect 56590 44158 56642 44210
rect 57150 44158 57202 44210
rect 15486 44046 15538 44098
rect 20078 44046 20130 44098
rect 23102 44046 23154 44098
rect 29262 44046 29314 44098
rect 33518 44046 33570 44098
rect 37550 44046 37602 44098
rect 39118 44046 39170 44098
rect 41022 44046 41074 44098
rect 44382 44046 44434 44098
rect 46174 44046 46226 44098
rect 50094 44046 50146 44098
rect 51438 44046 51490 44098
rect 52222 44046 52274 44098
rect 52894 44046 52946 44098
rect 53566 44046 53618 44098
rect 54350 44046 54402 44098
rect 55918 44046 55970 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 10110 43710 10162 43762
rect 37998 43710 38050 43762
rect 40014 43710 40066 43762
rect 45502 43710 45554 43762
rect 48638 43710 48690 43762
rect 9774 43598 9826 43650
rect 11454 43598 11506 43650
rect 18062 43598 18114 43650
rect 18510 43598 18562 43650
rect 18958 43598 19010 43650
rect 21310 43598 21362 43650
rect 27246 43598 27298 43650
rect 27918 43598 27970 43650
rect 28254 43598 28306 43650
rect 28702 43598 28754 43650
rect 30158 43598 30210 43650
rect 30494 43598 30546 43650
rect 33966 43598 34018 43650
rect 35646 43598 35698 43650
rect 36654 43598 36706 43650
rect 39790 43598 39842 43650
rect 43038 43598 43090 43650
rect 52446 43598 52498 43650
rect 52782 43598 52834 43650
rect 53006 43598 53058 43650
rect 53790 43598 53842 43650
rect 56030 43598 56082 43650
rect 57038 43598 57090 43650
rect 6974 43486 7026 43538
rect 9550 43486 9602 43538
rect 10558 43486 10610 43538
rect 11006 43486 11058 43538
rect 11678 43486 11730 43538
rect 12238 43486 12290 43538
rect 17838 43486 17890 43538
rect 20862 43486 20914 43538
rect 21198 43486 21250 43538
rect 21422 43486 21474 43538
rect 24558 43486 24610 43538
rect 27582 43486 27634 43538
rect 33630 43486 33682 43538
rect 34414 43486 34466 43538
rect 34862 43486 34914 43538
rect 35870 43486 35922 43538
rect 36094 43486 36146 43538
rect 36206 43486 36258 43538
rect 36542 43486 36594 43538
rect 36878 43486 36930 43538
rect 38782 43486 38834 43538
rect 39230 43486 39282 43538
rect 42478 43486 42530 43538
rect 42814 43486 42866 43538
rect 46174 43486 46226 43538
rect 46510 43486 46562 43538
rect 47294 43486 47346 43538
rect 47630 43486 47682 43538
rect 48190 43486 48242 43538
rect 49422 43486 49474 43538
rect 49646 43486 49698 43538
rect 50318 43486 50370 43538
rect 51774 43486 51826 43538
rect 52110 43486 52162 43538
rect 55470 43486 55522 43538
rect 55806 43486 55858 43538
rect 56590 43486 56642 43538
rect 56814 43486 56866 43538
rect 7534 43374 7586 43426
rect 12910 43374 12962 43426
rect 15038 43374 15090 43426
rect 19742 43374 19794 43426
rect 21758 43374 21810 43426
rect 23886 43374 23938 43426
rect 28590 43374 28642 43426
rect 33406 43374 33458 43426
rect 35310 43374 35362 43426
rect 39006 43374 39058 43426
rect 39342 43374 39394 43426
rect 42926 43374 42978 43426
rect 45838 43374 45890 43426
rect 49534 43374 49586 43426
rect 51326 43374 51378 43426
rect 53118 43374 53170 43426
rect 55918 43374 55970 43426
rect 18846 43262 18898 43314
rect 28926 43262 28978 43314
rect 38558 43262 38610 43314
rect 40126 43262 40178 43314
rect 47406 43262 47458 43314
rect 50542 43262 50594 43314
rect 50878 43262 50930 43314
rect 53566 43262 53618 43314
rect 53902 43262 53954 43314
rect 57374 43262 57426 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 22654 42926 22706 42978
rect 37550 42926 37602 42978
rect 40462 42926 40514 42978
rect 43822 42926 43874 42978
rect 9550 42814 9602 42866
rect 17054 42814 17106 42866
rect 17838 42814 17890 42866
rect 21758 42814 21810 42866
rect 22318 42814 22370 42866
rect 24334 42814 24386 42866
rect 26462 42814 26514 42866
rect 33742 42814 33794 42866
rect 34638 42814 34690 42866
rect 36318 42814 36370 42866
rect 38670 42814 38722 42866
rect 38782 42814 38834 42866
rect 40574 42814 40626 42866
rect 42478 42814 42530 42866
rect 45838 42814 45890 42866
rect 48974 42814 49026 42866
rect 53118 42814 53170 42866
rect 55694 42814 55746 42866
rect 57822 42814 57874 42866
rect 6750 42702 6802 42754
rect 14926 42702 14978 42754
rect 16270 42702 16322 42754
rect 18062 42702 18114 42754
rect 18286 42702 18338 42754
rect 18846 42702 18898 42754
rect 23550 42702 23602 42754
rect 31278 42702 31330 42754
rect 31950 42702 32002 42754
rect 32510 42702 32562 42754
rect 34302 42702 34354 42754
rect 35870 42702 35922 42754
rect 36206 42702 36258 42754
rect 37662 42702 37714 42754
rect 38110 42702 38162 42754
rect 39230 42702 39282 42754
rect 40126 42702 40178 42754
rect 42814 42702 42866 42754
rect 43150 42702 43202 42754
rect 43598 42702 43650 42754
rect 43934 42702 43986 42754
rect 44270 42702 44322 42754
rect 44942 42702 44994 42754
rect 46286 42702 46338 42754
rect 47182 42702 47234 42754
rect 50990 42702 51042 42754
rect 51662 42702 51714 42754
rect 52558 42702 52610 42754
rect 53006 42702 53058 42754
rect 54910 42702 54962 42754
rect 7422 42590 7474 42642
rect 17390 42590 17442 42642
rect 17614 42590 17666 42642
rect 21310 42590 21362 42642
rect 22542 42590 22594 42642
rect 30606 42590 30658 42642
rect 30830 42590 30882 42642
rect 38446 42590 38498 42642
rect 42366 42590 42418 42642
rect 42926 42590 42978 42642
rect 45166 42590 45218 42642
rect 46734 42590 46786 42642
rect 47294 42590 47346 42642
rect 50878 42590 50930 42642
rect 53230 42590 53282 42642
rect 9998 42478 10050 42530
rect 10782 42478 10834 42530
rect 11790 42478 11842 42530
rect 14590 42478 14642 42530
rect 16382 42478 16434 42530
rect 17726 42478 17778 42530
rect 18622 42478 18674 42530
rect 21534 42478 21586 42530
rect 21758 42478 21810 42530
rect 21870 42478 21922 42530
rect 23214 42478 23266 42530
rect 27806 42478 27858 42530
rect 31054 42478 31106 42530
rect 37550 42478 37602 42530
rect 41470 42478 41522 42530
rect 44158 42478 44210 42530
rect 51438 42478 51490 42530
rect 51774 42478 51826 42530
rect 51886 42478 51938 42530
rect 53678 42478 53730 42530
rect 54126 42478 54178 42530
rect 54574 42478 54626 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 9886 42142 9938 42194
rect 10670 42142 10722 42194
rect 10894 42142 10946 42194
rect 21422 42142 21474 42194
rect 22094 42142 22146 42194
rect 37998 42142 38050 42194
rect 40126 42142 40178 42194
rect 43710 42142 43762 42194
rect 47294 42142 47346 42194
rect 47854 42142 47906 42194
rect 48750 42142 48802 42194
rect 55806 42142 55858 42194
rect 10222 42030 10274 42082
rect 14478 42030 14530 42082
rect 14814 42030 14866 42082
rect 15822 42030 15874 42082
rect 19630 42030 19682 42082
rect 19966 42030 20018 42082
rect 31278 42030 31330 42082
rect 37886 42030 37938 42082
rect 39454 42030 39506 42082
rect 39566 42030 39618 42082
rect 40238 42030 40290 42082
rect 45838 42030 45890 42082
rect 49534 42030 49586 42082
rect 56702 42030 56754 42082
rect 6078 41918 6130 41970
rect 10558 41918 10610 41970
rect 11118 41918 11170 41970
rect 14366 41918 14418 41970
rect 15262 41918 15314 41970
rect 16046 41918 16098 41970
rect 17726 41918 17778 41970
rect 17950 41918 18002 41970
rect 18174 41918 18226 41970
rect 18398 41918 18450 41970
rect 18734 41918 18786 41970
rect 18846 41918 18898 41970
rect 19070 41918 19122 41970
rect 19294 41918 19346 41970
rect 20974 41918 21026 41970
rect 21198 41918 21250 41970
rect 21310 41918 21362 41970
rect 21534 41918 21586 41970
rect 25566 41918 25618 41970
rect 25902 41918 25954 41970
rect 31950 41918 32002 41970
rect 32510 41918 32562 41970
rect 34526 41918 34578 41970
rect 34862 41918 34914 41970
rect 38222 41918 38274 41970
rect 39006 41918 39058 41970
rect 39790 41918 39842 41970
rect 41022 41918 41074 41970
rect 41582 41918 41634 41970
rect 41806 41918 41858 41970
rect 42030 41918 42082 41970
rect 42142 41918 42194 41970
rect 42366 41918 42418 41970
rect 43038 41918 43090 41970
rect 43598 41918 43650 41970
rect 45278 41918 45330 41970
rect 45502 41918 45554 41970
rect 46958 41918 47010 41970
rect 47630 41918 47682 41970
rect 48302 41918 48354 41970
rect 48974 41918 49026 41970
rect 49198 41918 49250 41970
rect 51326 41918 51378 41970
rect 52222 41918 52274 41970
rect 52446 41918 52498 41970
rect 53118 41918 53170 41970
rect 53454 41918 53506 41970
rect 56030 41918 56082 41970
rect 57038 41918 57090 41970
rect 6862 41806 6914 41858
rect 8990 41806 9042 41858
rect 11902 41806 11954 41858
rect 14030 41806 14082 41858
rect 15486 41806 15538 41858
rect 26686 41806 26738 41858
rect 28814 41806 28866 41858
rect 29150 41806 29202 41858
rect 34302 41806 34354 41858
rect 38446 41806 38498 41858
rect 43262 41806 43314 41858
rect 46622 41806 46674 41858
rect 47742 41806 47794 41858
rect 50206 41806 50258 41858
rect 51102 41806 51154 41858
rect 52894 41806 52946 41858
rect 53006 41806 53058 41858
rect 53566 41806 53618 41858
rect 54014 41806 54066 41858
rect 54462 41806 54514 41858
rect 54910 41806 54962 41858
rect 55694 41806 55746 41858
rect 57262 41806 57314 41858
rect 38670 41694 38722 41746
rect 40126 41694 40178 41746
rect 40910 41694 40962 41746
rect 42814 41694 42866 41746
rect 49086 41694 49138 41746
rect 52670 41694 52722 41746
rect 54014 41694 54066 41746
rect 54238 41694 54290 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 17278 41358 17330 41410
rect 18062 41358 18114 41410
rect 19518 41358 19570 41410
rect 51662 41358 51714 41410
rect 9886 41246 9938 41298
rect 14254 41246 14306 41298
rect 16718 41246 16770 41298
rect 19854 41246 19906 41298
rect 21422 41246 21474 41298
rect 22430 41246 22482 41298
rect 25678 41246 25730 41298
rect 30606 41246 30658 41298
rect 34638 41246 34690 41298
rect 40126 41246 40178 41298
rect 41918 41246 41970 41298
rect 46174 41246 46226 41298
rect 50654 41246 50706 41298
rect 51550 41246 51602 41298
rect 53454 41246 53506 41298
rect 55582 41246 55634 41298
rect 57262 41246 57314 41298
rect 10110 41134 10162 41186
rect 13582 41134 13634 41186
rect 14366 41134 14418 41186
rect 14814 41134 14866 41186
rect 15038 41134 15090 41186
rect 15262 41134 15314 41186
rect 16270 41134 16322 41186
rect 16942 41134 16994 41186
rect 18286 41134 18338 41186
rect 19294 41134 19346 41186
rect 19742 41134 19794 41186
rect 25342 41134 25394 41186
rect 28590 41134 28642 41186
rect 29262 41134 29314 41186
rect 31390 41134 31442 41186
rect 31726 41134 31778 41186
rect 39230 41134 39282 41186
rect 39790 41134 39842 41186
rect 39902 41134 39954 41186
rect 40350 41134 40402 41186
rect 44942 41134 44994 41186
rect 48974 41134 49026 41186
rect 49982 41134 50034 41186
rect 50094 41134 50146 41186
rect 50542 41134 50594 41186
rect 50990 41134 51042 41186
rect 51886 41134 51938 41186
rect 52670 41134 52722 41186
rect 57598 41134 57650 41186
rect 15934 41022 15986 41074
rect 17614 41022 17666 41074
rect 17838 41022 17890 41074
rect 18510 41022 18562 41074
rect 19070 41022 19122 41074
rect 19966 41022 20018 41074
rect 20638 41022 20690 41074
rect 24558 41022 24610 41074
rect 27806 41022 27858 41074
rect 30830 41022 30882 41074
rect 31054 41022 31106 41074
rect 31166 41022 31218 41074
rect 32510 41022 32562 41074
rect 35086 41022 35138 41074
rect 35198 41022 35250 41074
rect 39454 41022 39506 41074
rect 40910 41022 40962 41074
rect 41358 41022 41410 41074
rect 41470 41022 41522 41074
rect 43038 41022 43090 41074
rect 45166 41022 45218 41074
rect 48302 41022 48354 41074
rect 50206 41022 50258 41074
rect 50878 41022 50930 41074
rect 51998 41022 52050 41074
rect 56702 41022 56754 41074
rect 5070 40910 5122 40962
rect 9214 40910 9266 40962
rect 10446 40910 10498 40962
rect 13806 40910 13858 40962
rect 14142 40910 14194 40962
rect 15150 40910 15202 40962
rect 15486 40910 15538 40962
rect 16046 40910 16098 40962
rect 17950 40910 18002 40962
rect 20302 40910 20354 40962
rect 21310 40910 21362 40962
rect 21534 40910 21586 40962
rect 21758 40910 21810 40962
rect 34862 40910 34914 40962
rect 35646 40910 35698 40962
rect 36094 40910 36146 40962
rect 37550 40910 37602 40962
rect 39790 40910 39842 40962
rect 40574 40910 40626 40962
rect 40798 40910 40850 40962
rect 41134 40910 41186 40962
rect 42702 40910 42754 40962
rect 43374 40910 43426 40962
rect 43822 40910 43874 40962
rect 49758 40910 49810 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 8094 40574 8146 40626
rect 8878 40574 8930 40626
rect 7646 40462 7698 40514
rect 9886 40462 9938 40514
rect 10110 40462 10162 40514
rect 11230 40518 11282 40570
rect 12014 40574 12066 40626
rect 13470 40574 13522 40626
rect 14814 40574 14866 40626
rect 16382 40574 16434 40626
rect 19294 40574 19346 40626
rect 20638 40574 20690 40626
rect 22318 40574 22370 40626
rect 23214 40574 23266 40626
rect 26462 40574 26514 40626
rect 27918 40574 27970 40626
rect 33518 40574 33570 40626
rect 39678 40574 39730 40626
rect 41022 40574 41074 40626
rect 41806 40574 41858 40626
rect 42030 40574 42082 40626
rect 43038 40574 43090 40626
rect 43598 40574 43650 40626
rect 47294 40574 47346 40626
rect 47854 40574 47906 40626
rect 48750 40574 48802 40626
rect 49534 40574 49586 40626
rect 56926 40574 56978 40626
rect 10558 40462 10610 40514
rect 10894 40462 10946 40514
rect 11342 40462 11394 40514
rect 15934 40462 15986 40514
rect 16270 40462 16322 40514
rect 18510 40462 18562 40514
rect 24222 40462 24274 40514
rect 24558 40462 24610 40514
rect 27582 40462 27634 40514
rect 31166 40462 31218 40514
rect 36542 40462 36594 40514
rect 39902 40462 39954 40514
rect 40126 40462 40178 40514
rect 44046 40462 44098 40514
rect 47630 40462 47682 40514
rect 49086 40462 49138 40514
rect 50878 40462 50930 40514
rect 54686 40462 54738 40514
rect 55022 40462 55074 40514
rect 57038 40462 57090 40514
rect 57374 40462 57426 40514
rect 4062 40350 4114 40402
rect 4846 40350 4898 40402
rect 7310 40350 7362 40402
rect 8542 40350 8594 40402
rect 10222 40350 10274 40402
rect 12014 40350 12066 40402
rect 12462 40350 12514 40402
rect 12798 40350 12850 40402
rect 13582 40350 13634 40402
rect 13806 40350 13858 40402
rect 14254 40350 14306 40402
rect 14478 40350 14530 40402
rect 15710 40350 15762 40402
rect 18846 40350 18898 40402
rect 19518 40350 19570 40402
rect 20862 40350 20914 40402
rect 21086 40350 21138 40402
rect 22542 40350 22594 40402
rect 26350 40350 26402 40402
rect 26574 40350 26626 40402
rect 26910 40350 26962 40402
rect 30942 40350 30994 40402
rect 32062 40350 32114 40402
rect 32510 40350 32562 40402
rect 33070 40350 33122 40402
rect 33406 40350 33458 40402
rect 33742 40350 33794 40402
rect 37214 40350 37266 40402
rect 37886 40350 37938 40402
rect 38782 40350 38834 40402
rect 39454 40350 39506 40402
rect 42254 40350 42306 40402
rect 42926 40350 42978 40402
rect 43262 40350 43314 40402
rect 43374 40350 43426 40402
rect 43822 40350 43874 40402
rect 44382 40350 44434 40402
rect 44718 40350 44770 40402
rect 44942 40350 44994 40402
rect 45502 40350 45554 40402
rect 46062 40350 46114 40402
rect 50206 40350 50258 40402
rect 51662 40350 51714 40402
rect 51886 40350 51938 40402
rect 54014 40350 54066 40402
rect 54350 40350 54402 40402
rect 55694 40350 55746 40402
rect 55918 40350 55970 40402
rect 56590 40350 56642 40402
rect 3278 40238 3330 40290
rect 6974 40238 7026 40290
rect 9774 40238 9826 40290
rect 20974 40238 21026 40290
rect 23214 40238 23266 40290
rect 31614 40238 31666 40290
rect 34414 40238 34466 40290
rect 38110 40238 38162 40290
rect 42142 40238 42194 40290
rect 44494 40238 44546 40290
rect 47966 40238 48018 40290
rect 53678 40238 53730 40290
rect 53902 40238 53954 40290
rect 2942 40126 2994 40178
rect 3054 40126 3106 40178
rect 3390 40126 3442 40178
rect 8766 40126 8818 40178
rect 8878 40126 8930 40178
rect 11342 40126 11394 40178
rect 12350 40126 12402 40178
rect 13470 40126 13522 40178
rect 22990 40126 23042 40178
rect 44830 40126 44882 40178
rect 45838 40126 45890 40178
rect 50990 40126 51042 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 10110 39790 10162 39842
rect 41022 39790 41074 39842
rect 50878 39790 50930 39842
rect 2494 39678 2546 39730
rect 5742 39678 5794 39730
rect 7982 39678 8034 39730
rect 9326 39678 9378 39730
rect 11118 39678 11170 39730
rect 13582 39678 13634 39730
rect 16158 39678 16210 39730
rect 17166 39678 17218 39730
rect 17502 39678 17554 39730
rect 18846 39678 18898 39730
rect 19294 39678 19346 39730
rect 26350 39678 26402 39730
rect 26910 39678 26962 39730
rect 27582 39678 27634 39730
rect 30494 39678 30546 39730
rect 38222 39678 38274 39730
rect 41246 39678 41298 39730
rect 43486 39678 43538 39730
rect 44942 39678 44994 39730
rect 51326 39678 51378 39730
rect 54126 39678 54178 39730
rect 55806 39678 55858 39730
rect 57934 39678 57986 39730
rect 1822 39566 1874 39618
rect 6078 39566 6130 39618
rect 6414 39566 6466 39618
rect 7422 39566 7474 39618
rect 8318 39566 8370 39618
rect 9662 39566 9714 39618
rect 9886 39566 9938 39618
rect 11006 39566 11058 39618
rect 13470 39566 13522 39618
rect 13694 39566 13746 39618
rect 14030 39566 14082 39618
rect 15486 39566 15538 39618
rect 15822 39566 15874 39618
rect 16606 39566 16658 39618
rect 17838 39566 17890 39618
rect 18286 39566 18338 39618
rect 18510 39566 18562 39618
rect 22094 39566 22146 39618
rect 23438 39566 23490 39618
rect 26574 39566 26626 39618
rect 27806 39566 27858 39618
rect 28030 39566 28082 39618
rect 30718 39566 30770 39618
rect 36094 39566 36146 39618
rect 37774 39566 37826 39618
rect 38110 39566 38162 39618
rect 40014 39566 40066 39618
rect 41134 39566 41186 39618
rect 42926 39566 42978 39618
rect 45166 39566 45218 39618
rect 45390 39566 45442 39618
rect 51102 39566 51154 39618
rect 51438 39566 51490 39618
rect 55022 39566 55074 39618
rect 5630 39454 5682 39506
rect 5854 39454 5906 39506
rect 7086 39454 7138 39506
rect 8766 39454 8818 39506
rect 10446 39454 10498 39506
rect 12910 39454 12962 39506
rect 17726 39454 17778 39506
rect 20078 39454 20130 39506
rect 21534 39454 21586 39506
rect 23774 39454 23826 39506
rect 40126 39454 40178 39506
rect 44830 39454 44882 39506
rect 52894 39454 52946 39506
rect 53006 39454 53058 39506
rect 53118 39454 53170 39506
rect 54350 39454 54402 39506
rect 4734 39342 4786 39394
rect 9214 39342 9266 39394
rect 9438 39342 9490 39394
rect 10558 39342 10610 39394
rect 10782 39342 10834 39394
rect 11566 39342 11618 39394
rect 12798 39342 12850 39394
rect 20190 39342 20242 39394
rect 23662 39342 23714 39394
rect 26238 39342 26290 39394
rect 26462 39342 26514 39394
rect 31054 39342 31106 39394
rect 36430 39342 36482 39394
rect 44046 39342 44098 39394
rect 48414 39342 48466 39394
rect 50430 39342 50482 39394
rect 52670 39342 52722 39394
rect 52782 39342 52834 39394
rect 53790 39342 53842 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 3502 39006 3554 39058
rect 3950 39006 4002 39058
rect 7198 39006 7250 39058
rect 8542 39006 8594 39058
rect 10334 39006 10386 39058
rect 11566 39006 11618 39058
rect 11902 39006 11954 39058
rect 13470 39006 13522 39058
rect 15934 39006 15986 39058
rect 19742 39006 19794 39058
rect 24446 39006 24498 39058
rect 2942 38894 2994 38946
rect 10222 38894 10274 38946
rect 10670 38894 10722 38946
rect 12798 38894 12850 38946
rect 13582 38894 13634 38946
rect 14926 38894 14978 38946
rect 15374 38894 15426 38946
rect 17614 38894 17666 38946
rect 17726 38950 17778 39002
rect 24558 39006 24610 39058
rect 27022 39006 27074 39058
rect 27806 39006 27858 39058
rect 28030 39006 28082 39058
rect 30046 39006 30098 39058
rect 30942 39006 30994 39058
rect 34302 39006 34354 39058
rect 34638 39006 34690 39058
rect 36990 39006 37042 39058
rect 37214 39006 37266 39058
rect 37774 39006 37826 39058
rect 40238 39006 40290 39058
rect 40462 39006 40514 39058
rect 41022 39006 41074 39058
rect 44382 39006 44434 39058
rect 48078 39006 48130 39058
rect 50990 39006 51042 39058
rect 51438 39006 51490 39058
rect 53678 39006 53730 39058
rect 55022 39006 55074 39058
rect 55470 39006 55522 39058
rect 57150 39006 57202 39058
rect 57486 39006 57538 39058
rect 18286 38894 18338 38946
rect 19182 38894 19234 38946
rect 21534 38894 21586 38946
rect 21758 38894 21810 38946
rect 23550 38894 23602 38946
rect 25230 38894 25282 38946
rect 27582 38894 27634 38946
rect 28366 38894 28418 38946
rect 28926 38894 28978 38946
rect 29710 38894 29762 38946
rect 36654 38894 36706 38946
rect 39566 38894 39618 38946
rect 40126 38894 40178 38946
rect 41358 38894 41410 38946
rect 43598 38894 43650 38946
rect 43822 38894 43874 38946
rect 46846 38894 46898 38946
rect 50654 38894 50706 38946
rect 51326 38894 51378 38946
rect 53118 38894 53170 38946
rect 53230 38894 53282 38946
rect 55918 38894 55970 38946
rect 2718 38782 2770 38834
rect 3054 38782 3106 38834
rect 3726 38782 3778 38834
rect 4174 38782 4226 38834
rect 4286 38782 4338 38834
rect 4734 38782 4786 38834
rect 5182 38782 5234 38834
rect 6078 38782 6130 38834
rect 6302 38782 6354 38834
rect 6414 38782 6466 38834
rect 7534 38782 7586 38834
rect 8318 38782 8370 38834
rect 8542 38782 8594 38834
rect 8766 38782 8818 38834
rect 8990 38782 9042 38834
rect 9662 38782 9714 38834
rect 9998 38782 10050 38834
rect 10894 38782 10946 38834
rect 11342 38782 11394 38834
rect 12350 38782 12402 38834
rect 13022 38782 13074 38834
rect 13694 38782 13746 38834
rect 14142 38782 14194 38834
rect 14254 38782 14306 38834
rect 14590 38782 14642 38834
rect 15486 38782 15538 38834
rect 16382 38782 16434 38834
rect 16830 38782 16882 38834
rect 18510 38782 18562 38834
rect 18734 38782 18786 38834
rect 19406 38782 19458 38834
rect 20302 38782 20354 38834
rect 20862 38782 20914 38834
rect 21086 38782 21138 38834
rect 21870 38782 21922 38834
rect 22094 38782 22146 38834
rect 22878 38782 22930 38834
rect 24110 38782 24162 38834
rect 24334 38782 24386 38834
rect 25342 38782 25394 38834
rect 26686 38782 26738 38834
rect 27470 38782 27522 38834
rect 29262 38782 29314 38834
rect 31390 38782 31442 38834
rect 31838 38782 31890 38834
rect 35198 38782 35250 38834
rect 35758 38782 35810 38834
rect 37326 38782 37378 38834
rect 37662 38782 37714 38834
rect 37998 38782 38050 38834
rect 38558 38782 38610 38834
rect 39230 38782 39282 38834
rect 39454 38782 39506 38834
rect 41694 38782 41746 38834
rect 41918 38782 41970 38834
rect 42366 38782 42418 38834
rect 42702 38782 42754 38834
rect 42926 38782 42978 38834
rect 44158 38782 44210 38834
rect 47630 38782 47682 38834
rect 48862 38782 48914 38834
rect 50430 38782 50482 38834
rect 52222 38782 52274 38834
rect 52894 38782 52946 38834
rect 56702 38782 56754 38834
rect 4846 38670 4898 38722
rect 6862 38670 6914 38722
rect 10558 38670 10610 38722
rect 13134 38670 13186 38722
rect 14478 38670 14530 38722
rect 18174 38670 18226 38722
rect 20078 38670 20130 38722
rect 22766 38670 22818 38722
rect 26462 38670 26514 38722
rect 30382 38670 30434 38722
rect 36094 38670 36146 38722
rect 41470 38670 41522 38722
rect 42590 38670 42642 38722
rect 44718 38670 44770 38722
rect 49198 38670 49250 38722
rect 52334 38670 52386 38722
rect 54126 38670 54178 38722
rect 54574 38670 54626 38722
rect 56590 38670 56642 38722
rect 5406 38558 5458 38610
rect 5742 38558 5794 38610
rect 12574 38558 12626 38610
rect 15374 38558 15426 38610
rect 17614 38558 17666 38610
rect 20638 38558 20690 38610
rect 23886 38558 23938 38610
rect 41806 38558 41858 38610
rect 44158 38558 44210 38610
rect 52446 38558 52498 38610
rect 54014 38558 54066 38610
rect 54462 38558 54514 38610
rect 55022 38558 55074 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 4062 38222 4114 38274
rect 20526 38222 20578 38274
rect 20638 38222 20690 38274
rect 36318 38222 36370 38274
rect 37326 38222 37378 38274
rect 37662 38222 37714 38274
rect 38110 38222 38162 38274
rect 39566 38222 39618 38274
rect 14142 38110 14194 38162
rect 15710 38110 15762 38162
rect 19630 38110 19682 38162
rect 28478 38110 28530 38162
rect 34750 38110 34802 38162
rect 40574 38110 40626 38162
rect 42702 38110 42754 38162
rect 43934 38110 43986 38162
rect 45950 38110 46002 38162
rect 48414 38110 48466 38162
rect 51326 38110 51378 38162
rect 53342 38110 53394 38162
rect 56814 38110 56866 38162
rect 4846 37998 4898 38050
rect 5854 37998 5906 38050
rect 7646 37998 7698 38050
rect 10222 37998 10274 38050
rect 10558 37998 10610 38050
rect 11118 37998 11170 38050
rect 11566 37998 11618 38050
rect 12686 37998 12738 38050
rect 13806 37998 13858 38050
rect 14030 37998 14082 38050
rect 14366 37998 14418 38050
rect 15822 37998 15874 38050
rect 17502 37998 17554 38050
rect 18846 37998 18898 38050
rect 19742 37998 19794 38050
rect 24558 37998 24610 38050
rect 24894 37998 24946 38050
rect 25230 37998 25282 38050
rect 25678 37998 25730 38050
rect 26238 37998 26290 38050
rect 29150 37998 29202 38050
rect 30046 37998 30098 38050
rect 31278 37998 31330 38050
rect 31950 37998 32002 38050
rect 35422 37998 35474 38050
rect 36206 37998 36258 38050
rect 37662 37998 37714 38050
rect 37886 37998 37938 38050
rect 38782 37998 38834 38050
rect 43486 37998 43538 38050
rect 45054 37998 45106 38050
rect 45502 37998 45554 38050
rect 49870 37998 49922 38050
rect 51438 37998 51490 38050
rect 51662 37998 51714 38050
rect 53118 37998 53170 38050
rect 53566 37998 53618 38050
rect 54014 37998 54066 38050
rect 57374 37998 57426 38050
rect 3502 37886 3554 37938
rect 3950 37886 4002 37938
rect 6862 37886 6914 37938
rect 10446 37886 10498 37938
rect 11678 37886 11730 37938
rect 12798 37886 12850 37938
rect 16046 37886 16098 37938
rect 19966 37886 20018 37938
rect 22206 37886 22258 37938
rect 22542 37886 22594 37938
rect 23662 37886 23714 37938
rect 23998 37886 24050 37938
rect 24222 37886 24274 37938
rect 27694 37886 27746 37938
rect 27806 37886 27858 37938
rect 28366 37886 28418 37938
rect 29262 37886 29314 37938
rect 31502 37886 31554 37938
rect 32622 37886 32674 37938
rect 39790 37886 39842 37938
rect 44830 37886 44882 37938
rect 46734 37886 46786 37938
rect 50206 37886 50258 37938
rect 50318 37886 50370 37938
rect 50542 37886 50594 37938
rect 52670 37886 52722 37938
rect 52894 37886 52946 37938
rect 54686 37886 54738 37938
rect 3726 37774 3778 37826
rect 4510 37774 4562 37826
rect 5070 37774 5122 37826
rect 8206 37774 8258 37826
rect 9214 37774 9266 37826
rect 13022 37774 13074 37826
rect 14254 37774 14306 37826
rect 14926 37774 14978 37826
rect 15262 37774 15314 37826
rect 20190 37774 20242 37826
rect 21310 37774 21362 37826
rect 21646 37774 21698 37826
rect 23886 37774 23938 37826
rect 24894 37774 24946 37826
rect 25902 37774 25954 37826
rect 26350 37774 26402 37826
rect 26574 37774 26626 37826
rect 27470 37774 27522 37826
rect 30046 37774 30098 37826
rect 35086 37774 35138 37826
rect 35870 37774 35922 37826
rect 36318 37774 36370 37826
rect 43822 37774 43874 37826
rect 46398 37774 46450 37826
rect 51998 37774 52050 37826
rect 53678 37774 53730 37826
rect 57038 37774 57090 37826
rect 57262 37774 57314 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 2382 37438 2434 37490
rect 9550 37438 9602 37490
rect 17390 37438 17442 37490
rect 17726 37438 17778 37490
rect 23102 37438 23154 37490
rect 28254 37438 28306 37490
rect 35982 37438 36034 37490
rect 40126 37438 40178 37490
rect 44606 37438 44658 37490
rect 45502 37438 45554 37490
rect 48862 37438 48914 37490
rect 51102 37438 51154 37490
rect 55694 37438 55746 37490
rect 55806 37438 55858 37490
rect 2718 37326 2770 37378
rect 4510 37326 4562 37378
rect 5294 37326 5346 37378
rect 7758 37326 7810 37378
rect 12350 37326 12402 37378
rect 13582 37326 13634 37378
rect 18286 37326 18338 37378
rect 20526 37326 20578 37378
rect 22542 37326 22594 37378
rect 23326 37326 23378 37378
rect 27582 37326 27634 37378
rect 34750 37326 34802 37378
rect 34974 37326 35026 37378
rect 36430 37326 36482 37378
rect 42702 37326 42754 37378
rect 46398 37326 46450 37378
rect 49758 37326 49810 37378
rect 52222 37326 52274 37378
rect 54126 37326 54178 37378
rect 54910 37326 54962 37378
rect 55582 37326 55634 37378
rect 2158 37214 2210 37266
rect 3054 37214 3106 37266
rect 3502 37214 3554 37266
rect 4622 37214 4674 37266
rect 5182 37214 5234 37266
rect 8878 37214 8930 37266
rect 10894 37214 10946 37266
rect 11230 37214 11282 37266
rect 11790 37214 11842 37266
rect 14926 37214 14978 37266
rect 15934 37214 15986 37266
rect 16718 37214 16770 37266
rect 18510 37214 18562 37266
rect 19854 37214 19906 37266
rect 20302 37214 20354 37266
rect 21310 37214 21362 37266
rect 21534 37214 21586 37266
rect 21982 37214 22034 37266
rect 22206 37214 22258 37266
rect 22766 37214 22818 37266
rect 25790 37214 25842 37266
rect 26462 37214 26514 37266
rect 27358 37214 27410 37266
rect 27694 37214 27746 37266
rect 28478 37214 28530 37266
rect 28926 37214 28978 37266
rect 31838 37214 31890 37266
rect 35534 37214 35586 37266
rect 36654 37214 36706 37266
rect 37438 37214 37490 37266
rect 37774 37214 37826 37266
rect 38782 37214 38834 37266
rect 39454 37214 39506 37266
rect 42366 37214 42418 37266
rect 42590 37214 42642 37266
rect 45166 37214 45218 37266
rect 46062 37214 46114 37266
rect 46734 37214 46786 37266
rect 51326 37214 51378 37266
rect 53454 37214 53506 37266
rect 53790 37214 53842 37266
rect 54238 37214 54290 37266
rect 54350 37214 54402 37266
rect 54686 37214 54738 37266
rect 55246 37214 55298 37266
rect 57262 37214 57314 37266
rect 3614 37102 3666 37154
rect 8318 37102 8370 37154
rect 9662 37102 9714 37154
rect 10334 37102 10386 37154
rect 15038 37102 15090 37154
rect 15710 37102 15762 37154
rect 16270 37102 16322 37154
rect 20190 37102 20242 37154
rect 22430 37102 22482 37154
rect 26350 37102 26402 37154
rect 28366 37102 28418 37154
rect 31502 37102 31554 37154
rect 39230 37102 39282 37154
rect 43710 37102 43762 37154
rect 47406 37102 47458 37154
rect 55134 37102 55186 37154
rect 57150 37102 57202 37154
rect 57598 37102 57650 37154
rect 3838 36990 3890 37042
rect 3950 36990 4002 37042
rect 4734 36990 4786 37042
rect 11342 36990 11394 37042
rect 15598 36990 15650 37042
rect 22990 36990 23042 37042
rect 26798 36990 26850 37042
rect 35086 36990 35138 37042
rect 36990 36990 37042 37042
rect 39678 36990 39730 37042
rect 42030 36990 42082 37042
rect 42142 36990 42194 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 5070 36654 5122 36706
rect 7646 36654 7698 36706
rect 7982 36654 8034 36706
rect 8318 36654 8370 36706
rect 10222 36654 10274 36706
rect 14478 36654 14530 36706
rect 15486 36654 15538 36706
rect 36318 36654 36370 36706
rect 51326 36654 51378 36706
rect 2494 36542 2546 36594
rect 4622 36542 4674 36594
rect 11566 36542 11618 36594
rect 21422 36542 21474 36594
rect 28590 36542 28642 36594
rect 29262 36542 29314 36594
rect 30158 36542 30210 36594
rect 34526 36542 34578 36594
rect 44158 36542 44210 36594
rect 49534 36542 49586 36594
rect 56142 36542 56194 36594
rect 1822 36430 1874 36482
rect 6190 36430 6242 36482
rect 8654 36430 8706 36482
rect 9438 36430 9490 36482
rect 10110 36430 10162 36482
rect 10670 36430 10722 36482
rect 14030 36430 14082 36482
rect 14142 36430 14194 36482
rect 14814 36430 14866 36482
rect 15374 36430 15426 36482
rect 16046 36430 16098 36482
rect 17614 36430 17666 36482
rect 19630 36430 19682 36482
rect 20414 36430 20466 36482
rect 20750 36430 20802 36482
rect 21534 36430 21586 36482
rect 21982 36430 22034 36482
rect 22990 36430 23042 36482
rect 23438 36430 23490 36482
rect 24110 36430 24162 36482
rect 24334 36430 24386 36482
rect 26238 36430 26290 36482
rect 26462 36430 26514 36482
rect 26910 36430 26962 36482
rect 28478 36430 28530 36482
rect 29598 36430 29650 36482
rect 29822 36430 29874 36482
rect 30046 36430 30098 36482
rect 31726 36430 31778 36482
rect 35534 36430 35586 36482
rect 35982 36430 36034 36482
rect 37998 36430 38050 36482
rect 38446 36430 38498 36482
rect 39566 36430 39618 36482
rect 43374 36430 43426 36482
rect 43822 36430 43874 36482
rect 44942 36430 44994 36482
rect 46286 36430 46338 36482
rect 46846 36430 46898 36482
rect 47406 36430 47458 36482
rect 47966 36430 48018 36482
rect 48190 36430 48242 36482
rect 48526 36430 48578 36482
rect 48750 36430 48802 36482
rect 49646 36430 49698 36482
rect 50094 36430 50146 36482
rect 50878 36430 50930 36482
rect 51438 36430 51490 36482
rect 52222 36430 52274 36482
rect 52670 36430 52722 36482
rect 53006 36430 53058 36482
rect 53230 36430 53282 36482
rect 53454 36430 53506 36482
rect 54350 36430 54402 36482
rect 54910 36430 54962 36482
rect 56590 36430 56642 36482
rect 57038 36430 57090 36482
rect 57598 36430 57650 36482
rect 4958 36318 5010 36370
rect 5966 36318 6018 36370
rect 6414 36318 6466 36370
rect 7534 36318 7586 36370
rect 9886 36318 9938 36370
rect 10558 36318 10610 36370
rect 12686 36318 12738 36370
rect 12798 36318 12850 36370
rect 13918 36318 13970 36370
rect 15038 36318 15090 36370
rect 16718 36318 16770 36370
rect 19966 36318 20018 36370
rect 20638 36318 20690 36370
rect 22654 36318 22706 36370
rect 22766 36318 22818 36370
rect 24558 36318 24610 36370
rect 26798 36318 26850 36370
rect 28142 36318 28194 36370
rect 32398 36318 32450 36370
rect 35758 36318 35810 36370
rect 38894 36318 38946 36370
rect 39118 36318 39170 36370
rect 43150 36318 43202 36370
rect 45166 36318 45218 36370
rect 45502 36318 45554 36370
rect 46510 36318 46562 36370
rect 50430 36318 50482 36370
rect 53790 36318 53842 36370
rect 55358 36318 55410 36370
rect 6750 36206 6802 36258
rect 8206 36206 8258 36258
rect 13022 36206 13074 36258
rect 13470 36206 13522 36258
rect 14590 36206 14642 36258
rect 16046 36206 16098 36258
rect 21310 36206 21362 36258
rect 23550 36206 23602 36258
rect 23662 36206 23714 36258
rect 24446 36206 24498 36258
rect 26686 36206 26738 36258
rect 27806 36206 27858 36258
rect 28030 36206 28082 36258
rect 29150 36206 29202 36258
rect 30270 36206 30322 36258
rect 34862 36206 34914 36258
rect 34974 36206 35026 36258
rect 35086 36206 35138 36258
rect 36206 36206 36258 36258
rect 38110 36206 38162 36258
rect 38222 36206 38274 36258
rect 38334 36206 38386 36258
rect 39230 36206 39282 36258
rect 43598 36206 43650 36258
rect 45838 36206 45890 36258
rect 48302 36206 48354 36258
rect 50318 36206 50370 36258
rect 52670 36206 52722 36258
rect 54014 36206 54066 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 5294 35870 5346 35922
rect 11230 35870 11282 35922
rect 15374 35870 15426 35922
rect 17950 35870 18002 35922
rect 18734 35870 18786 35922
rect 19518 35870 19570 35922
rect 22542 35870 22594 35922
rect 23998 35870 24050 35922
rect 31390 35870 31442 35922
rect 32398 35870 32450 35922
rect 33630 35870 33682 35922
rect 34078 35870 34130 35922
rect 35758 35870 35810 35922
rect 37998 35870 38050 35922
rect 40910 35870 40962 35922
rect 44270 35870 44322 35922
rect 44382 35870 44434 35922
rect 45390 35870 45442 35922
rect 46286 35870 46338 35922
rect 47182 35870 47234 35922
rect 47742 35870 47794 35922
rect 48078 35870 48130 35922
rect 48190 35870 48242 35922
rect 51550 35870 51602 35922
rect 54910 35870 54962 35922
rect 7870 35758 7922 35810
rect 12126 35758 12178 35810
rect 14702 35758 14754 35810
rect 14814 35758 14866 35810
rect 16718 35758 16770 35810
rect 16830 35758 16882 35810
rect 18286 35758 18338 35810
rect 26798 35758 26850 35810
rect 27806 35758 27858 35810
rect 33854 35758 33906 35810
rect 35310 35758 35362 35810
rect 36878 35758 36930 35810
rect 40126 35758 40178 35810
rect 41134 35758 41186 35810
rect 41246 35758 41298 35810
rect 41582 35758 41634 35810
rect 43934 35758 43986 35810
rect 44494 35758 44546 35810
rect 44718 35758 44770 35810
rect 49870 35758 49922 35810
rect 51438 35758 51490 35810
rect 53230 35758 53282 35810
rect 56590 35758 56642 35810
rect 2718 35646 2770 35698
rect 3054 35646 3106 35698
rect 4398 35646 4450 35698
rect 4734 35646 4786 35698
rect 4958 35646 5010 35698
rect 6078 35646 6130 35698
rect 7982 35646 8034 35698
rect 8206 35646 8258 35698
rect 10670 35646 10722 35698
rect 10894 35646 10946 35698
rect 11790 35646 11842 35698
rect 13470 35646 13522 35698
rect 15038 35646 15090 35698
rect 15598 35646 15650 35698
rect 16494 35646 16546 35698
rect 18958 35646 19010 35698
rect 23550 35646 23602 35698
rect 23774 35646 23826 35698
rect 25678 35646 25730 35698
rect 26686 35646 26738 35698
rect 27694 35646 27746 35698
rect 28254 35646 28306 35698
rect 28590 35646 28642 35698
rect 29486 35646 29538 35698
rect 29822 35646 29874 35698
rect 29934 35646 29986 35698
rect 31166 35646 31218 35698
rect 32174 35646 32226 35698
rect 35198 35646 35250 35698
rect 36206 35646 36258 35698
rect 37886 35646 37938 35698
rect 38334 35646 38386 35698
rect 38894 35646 38946 35698
rect 39230 35646 39282 35698
rect 42030 35646 42082 35698
rect 42478 35646 42530 35698
rect 43038 35646 43090 35698
rect 43262 35646 43314 35698
rect 45726 35646 45778 35698
rect 47966 35646 48018 35698
rect 49198 35646 49250 35698
rect 52110 35646 52162 35698
rect 52222 35646 52274 35698
rect 53342 35646 53394 35698
rect 53566 35646 53618 35698
rect 53790 35646 53842 35698
rect 54238 35646 54290 35698
rect 54686 35646 54738 35698
rect 55582 35646 55634 35698
rect 55806 35646 55858 35698
rect 56030 35646 56082 35698
rect 57038 35646 57090 35698
rect 57486 35646 57538 35698
rect 57934 35646 57986 35698
rect 3950 35534 4002 35586
rect 5742 35534 5794 35586
rect 8654 35534 8706 35586
rect 13918 35534 13970 35586
rect 15486 35534 15538 35586
rect 15822 35534 15874 35586
rect 16270 35534 16322 35586
rect 17390 35534 17442 35586
rect 18398 35534 18450 35586
rect 21198 35534 21250 35586
rect 21646 35534 21698 35586
rect 22654 35534 22706 35586
rect 27470 35534 27522 35586
rect 33742 35534 33794 35586
rect 34638 35534 34690 35586
rect 49534 35534 49586 35586
rect 50990 35534 51042 35586
rect 51662 35534 51714 35586
rect 54798 35534 54850 35586
rect 58046 35534 58098 35586
rect 3166 35422 3218 35474
rect 7422 35422 7474 35474
rect 16046 35422 16098 35474
rect 17614 35422 17666 35474
rect 22318 35422 22370 35474
rect 24110 35422 24162 35474
rect 30382 35422 30434 35474
rect 32510 35422 32562 35474
rect 37998 35422 38050 35474
rect 38558 35422 38610 35474
rect 52446 35422 52498 35474
rect 52558 35422 52610 35474
rect 53790 35422 53842 35474
rect 55470 35422 55522 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 3166 35086 3218 35138
rect 8206 35086 8258 35138
rect 10110 35086 10162 35138
rect 12798 35086 12850 35138
rect 13582 35086 13634 35138
rect 13806 35086 13858 35138
rect 18958 35086 19010 35138
rect 19294 35086 19346 35138
rect 23662 35086 23714 35138
rect 30270 35086 30322 35138
rect 52670 35086 52722 35138
rect 53006 35086 53058 35138
rect 53902 35086 53954 35138
rect 2830 34974 2882 35026
rect 4846 34974 4898 35026
rect 18062 34974 18114 35026
rect 19854 34974 19906 35026
rect 22206 34974 22258 35026
rect 30606 34974 30658 35026
rect 32398 34974 32450 35026
rect 34414 34974 34466 35026
rect 35198 34974 35250 35026
rect 36430 34974 36482 35026
rect 38782 34974 38834 35026
rect 39678 34974 39730 35026
rect 41358 34974 41410 35026
rect 43934 34974 43986 35026
rect 47854 34974 47906 35026
rect 49982 34974 50034 35026
rect 51774 34974 51826 35026
rect 52110 34974 52162 35026
rect 55134 34974 55186 35026
rect 57262 34974 57314 35026
rect 6750 34862 6802 34914
rect 7198 34862 7250 34914
rect 7646 34862 7698 34914
rect 8430 34862 8482 34914
rect 8654 34862 8706 34914
rect 8878 34862 8930 34914
rect 10670 34862 10722 34914
rect 14254 34862 14306 34914
rect 15262 34850 15314 34902
rect 18622 34862 18674 34914
rect 19518 34862 19570 34914
rect 21310 34862 21362 34914
rect 22430 34862 22482 34914
rect 22990 34862 23042 34914
rect 23438 34862 23490 34914
rect 23886 34862 23938 34914
rect 24334 34862 24386 34914
rect 25678 34862 25730 34914
rect 26462 34862 26514 34914
rect 27134 34862 27186 34914
rect 27358 34862 27410 34914
rect 27918 34862 27970 34914
rect 29150 34862 29202 34914
rect 29374 34862 29426 34914
rect 29710 34862 29762 34914
rect 30830 34862 30882 34914
rect 31502 34862 31554 34914
rect 32174 34862 32226 34914
rect 32846 34862 32898 34914
rect 34862 34862 34914 34914
rect 35870 34862 35922 34914
rect 35982 34862 36034 34914
rect 38222 34862 38274 34914
rect 38670 34862 38722 34914
rect 39342 34862 39394 34914
rect 40126 34862 40178 34914
rect 40462 34862 40514 34914
rect 41806 34862 41858 34914
rect 42254 34862 42306 34914
rect 42702 34862 42754 34914
rect 42814 34862 42866 34914
rect 45054 34862 45106 34914
rect 47070 34862 47122 34914
rect 50430 34862 50482 34914
rect 53230 34862 53282 34914
rect 53566 34862 53618 34914
rect 54462 34862 54514 34914
rect 6974 34750 7026 34802
rect 7870 34750 7922 34802
rect 9886 34750 9938 34802
rect 9998 34750 10050 34802
rect 10446 34750 10498 34802
rect 10894 34750 10946 34802
rect 11454 34750 11506 34802
rect 12686 34750 12738 34802
rect 14366 34750 14418 34802
rect 15934 34750 15986 34802
rect 19966 34750 20018 34802
rect 20190 34750 20242 34802
rect 21422 34750 21474 34802
rect 26350 34750 26402 34802
rect 28590 34750 28642 34802
rect 31166 34750 31218 34802
rect 31838 34750 31890 34802
rect 32622 34750 32674 34802
rect 35758 34750 35810 34802
rect 39790 34750 39842 34802
rect 40686 34750 40738 34802
rect 40798 34750 40850 34802
rect 43038 34750 43090 34802
rect 46398 34750 46450 34802
rect 46734 34750 46786 34802
rect 2942 34638 2994 34690
rect 7422 34638 7474 34690
rect 8766 34638 8818 34690
rect 10334 34638 10386 34690
rect 11790 34638 11842 34690
rect 12798 34638 12850 34690
rect 13470 34638 13522 34690
rect 14814 34638 14866 34690
rect 21646 34638 21698 34690
rect 24110 34638 24162 34690
rect 24222 34638 24274 34690
rect 25342 34638 25394 34690
rect 26798 34638 26850 34690
rect 26910 34638 26962 34690
rect 27582 34638 27634 34690
rect 27806 34638 27858 34690
rect 28254 34638 28306 34690
rect 29598 34638 29650 34690
rect 30494 34638 30546 34690
rect 31054 34638 31106 34690
rect 42590 34638 42642 34690
rect 45390 34638 45442 34690
rect 53790 34638 53842 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 7422 34302 7474 34354
rect 8094 34302 8146 34354
rect 8654 34302 8706 34354
rect 8878 34302 8930 34354
rect 8990 34302 9042 34354
rect 9998 34302 10050 34354
rect 10110 34302 10162 34354
rect 13470 34302 13522 34354
rect 14590 34302 14642 34354
rect 15150 34302 15202 34354
rect 16046 34302 16098 34354
rect 17502 34302 17554 34354
rect 19294 34302 19346 34354
rect 21646 34302 21698 34354
rect 24558 34302 24610 34354
rect 25342 34302 25394 34354
rect 28926 34302 28978 34354
rect 34190 34302 34242 34354
rect 35310 34302 35362 34354
rect 43374 34302 43426 34354
rect 50206 34302 50258 34354
rect 2494 34190 2546 34242
rect 7758 34190 7810 34242
rect 7982 34190 8034 34242
rect 10782 34190 10834 34242
rect 15038 34190 15090 34242
rect 15262 34190 15314 34242
rect 16270 34190 16322 34242
rect 21086 34190 21138 34242
rect 26910 34190 26962 34242
rect 27582 34190 27634 34242
rect 28478 34190 28530 34242
rect 29934 34190 29986 34242
rect 30942 34190 30994 34242
rect 31278 34190 31330 34242
rect 31726 34190 31778 34242
rect 37998 34190 38050 34242
rect 40350 34190 40402 34242
rect 42702 34190 42754 34242
rect 50766 34190 50818 34242
rect 53902 34190 53954 34242
rect 1822 34078 1874 34130
rect 5070 34078 5122 34130
rect 5294 34078 5346 34130
rect 5406 34078 5458 34130
rect 7198 34078 7250 34130
rect 8542 34078 8594 34130
rect 9886 34078 9938 34130
rect 10446 34078 10498 34130
rect 11006 34078 11058 34130
rect 11566 34078 11618 34130
rect 12014 34078 12066 34130
rect 13022 34078 13074 34130
rect 13246 34078 13298 34130
rect 13582 34078 13634 34130
rect 14030 34078 14082 34130
rect 15934 34078 15986 34130
rect 16494 34078 16546 34130
rect 18622 34078 18674 34130
rect 18958 34078 19010 34130
rect 19854 34078 19906 34130
rect 21310 34078 21362 34130
rect 22654 34078 22706 34130
rect 23102 34078 23154 34130
rect 24670 34078 24722 34130
rect 25230 34078 25282 34130
rect 25566 34078 25618 34130
rect 26238 34078 26290 34130
rect 26798 34078 26850 34130
rect 27918 34078 27970 34130
rect 28366 34078 28418 34130
rect 29374 34078 29426 34130
rect 30606 34078 30658 34130
rect 31502 34078 31554 34130
rect 31950 34078 32002 34130
rect 34414 34078 34466 34130
rect 34862 34078 34914 34130
rect 37102 34078 37154 34130
rect 37662 34078 37714 34130
rect 38446 34078 38498 34130
rect 39454 34078 39506 34130
rect 39790 34078 39842 34130
rect 41134 34078 41186 34130
rect 41694 34078 41746 34130
rect 43038 34078 43090 34130
rect 49534 34078 49586 34130
rect 49758 34078 49810 34130
rect 50094 34078 50146 34130
rect 50430 34078 50482 34130
rect 51662 34078 51714 34130
rect 52222 34078 52274 34130
rect 52782 34078 52834 34130
rect 53230 34078 53282 34130
rect 4622 33966 4674 34018
rect 13358 33966 13410 34018
rect 18510 33966 18562 34018
rect 20750 33966 20802 34018
rect 28030 33966 28082 34018
rect 31614 33966 31666 34018
rect 34302 33966 34354 34018
rect 38782 33966 38834 34018
rect 47406 33966 47458 34018
rect 56030 33966 56082 34018
rect 4958 33854 5010 33906
rect 8318 33854 8370 33906
rect 12014 33854 12066 33906
rect 14254 33854 14306 33906
rect 19406 33854 19458 33906
rect 19630 33854 19682 33906
rect 20078 33854 20130 33906
rect 20302 33854 20354 33906
rect 24222 33854 24274 33906
rect 24446 33854 24498 33906
rect 49198 33854 49250 33906
rect 51326 33854 51378 33906
rect 51438 33854 51490 33906
rect 51774 33854 51826 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 4734 33518 4786 33570
rect 4958 33518 5010 33570
rect 10782 33518 10834 33570
rect 12686 33518 12738 33570
rect 16270 33518 16322 33570
rect 16494 33518 16546 33570
rect 19966 33518 20018 33570
rect 20190 33518 20242 33570
rect 20638 33518 20690 33570
rect 22654 33518 22706 33570
rect 31950 33518 32002 33570
rect 39342 33518 39394 33570
rect 39902 33518 39954 33570
rect 54014 33518 54066 33570
rect 55022 33518 55074 33570
rect 4846 33406 4898 33458
rect 5966 33406 6018 33458
rect 8094 33406 8146 33458
rect 12126 33406 12178 33458
rect 14814 33406 14866 33458
rect 16494 33406 16546 33458
rect 17054 33406 17106 33458
rect 20302 33406 20354 33458
rect 36430 33406 36482 33458
rect 46174 33406 46226 33458
rect 48414 33406 48466 33458
rect 50990 33406 51042 33458
rect 52782 33406 52834 33458
rect 54014 33406 54066 33458
rect 54574 33406 54626 33458
rect 54910 33406 54962 33458
rect 8766 33294 8818 33346
rect 10558 33294 10610 33346
rect 11678 33294 11730 33346
rect 13694 33294 13746 33346
rect 14142 33294 14194 33346
rect 19182 33294 19234 33346
rect 19742 33294 19794 33346
rect 21982 33294 22034 33346
rect 22318 33294 22370 33346
rect 25118 33294 25170 33346
rect 25342 33294 25394 33346
rect 26238 33294 26290 33346
rect 26686 33294 26738 33346
rect 26910 33294 26962 33346
rect 27470 33294 27522 33346
rect 30606 33294 30658 33346
rect 30942 33294 30994 33346
rect 32286 33294 32338 33346
rect 32510 33294 32562 33346
rect 33182 33294 33234 33346
rect 33630 33294 33682 33346
rect 39454 33294 39506 33346
rect 39790 33294 39842 33346
rect 45838 33294 45890 33346
rect 46622 33294 46674 33346
rect 47182 33294 47234 33346
rect 48862 33294 48914 33346
rect 49310 33294 49362 33346
rect 50654 33294 50706 33346
rect 51214 33294 51266 33346
rect 11454 33182 11506 33234
rect 12686 33182 12738 33234
rect 12798 33182 12850 33234
rect 14366 33182 14418 33234
rect 18846 33182 18898 33234
rect 20750 33182 20802 33234
rect 21758 33182 21810 33234
rect 22542 33182 22594 33234
rect 25678 33182 25730 33234
rect 26014 33182 26066 33234
rect 27358 33182 27410 33234
rect 29150 33182 29202 33234
rect 32734 33182 32786 33234
rect 32958 33182 33010 33234
rect 34302 33182 34354 33234
rect 39342 33182 39394 33234
rect 47742 33182 47794 33234
rect 47966 33182 48018 33234
rect 50094 33182 50146 33234
rect 51662 33182 51714 33234
rect 9326 33070 9378 33122
rect 11118 33070 11170 33122
rect 12238 33070 12290 33122
rect 13918 33070 13970 33122
rect 15598 33070 15650 33122
rect 17950 33070 18002 33122
rect 18286 33070 18338 33122
rect 19070 33070 19122 33122
rect 19294 33070 19346 33122
rect 21422 33070 21474 33122
rect 25566 33070 25618 33122
rect 27134 33070 27186 33122
rect 27806 33070 27858 33122
rect 29486 33070 29538 33122
rect 30718 33070 30770 33122
rect 32062 33070 32114 33122
rect 37102 33070 37154 33122
rect 37550 33070 37602 33122
rect 41470 33070 41522 33122
rect 47854 33070 47906 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 6526 32734 6578 32786
rect 14366 32734 14418 32786
rect 17390 32734 17442 32786
rect 19182 32734 19234 32786
rect 25230 32734 25282 32786
rect 26126 32734 26178 32786
rect 27358 32734 27410 32786
rect 3950 32622 4002 32674
rect 14702 32622 14754 32674
rect 15262 32622 15314 32674
rect 15598 32622 15650 32674
rect 15822 32622 15874 32674
rect 18622 32622 18674 32674
rect 18846 32622 18898 32674
rect 19406 32622 19458 32674
rect 27582 32678 27634 32730
rect 29822 32734 29874 32786
rect 30046 32734 30098 32786
rect 30270 32734 30322 32786
rect 30494 32734 30546 32786
rect 32286 32734 32338 32786
rect 39790 32734 39842 32786
rect 46286 32734 46338 32786
rect 47518 32734 47570 32786
rect 47966 32734 48018 32786
rect 50542 32734 50594 32786
rect 20862 32622 20914 32674
rect 21870 32622 21922 32674
rect 24558 32622 24610 32674
rect 26350 32622 26402 32674
rect 26686 32622 26738 32674
rect 27694 32622 27746 32674
rect 28478 32622 28530 32674
rect 30606 32622 30658 32674
rect 33182 32622 33234 32674
rect 35198 32622 35250 32674
rect 37662 32622 37714 32674
rect 39118 32622 39170 32674
rect 41022 32622 41074 32674
rect 44606 32622 44658 32674
rect 45726 32622 45778 32674
rect 48190 32622 48242 32674
rect 48750 32622 48802 32674
rect 49646 32622 49698 32674
rect 51774 32622 51826 32674
rect 3278 32510 3330 32562
rect 16158 32510 16210 32562
rect 16606 32510 16658 32562
rect 19518 32510 19570 32562
rect 20414 32510 20466 32562
rect 21310 32510 21362 32562
rect 22430 32510 22482 32562
rect 22990 32510 23042 32562
rect 24334 32510 24386 32562
rect 25342 32510 25394 32562
rect 25790 32510 25842 32562
rect 26798 32510 26850 32562
rect 28590 32510 28642 32562
rect 28814 32510 28866 32562
rect 29262 32510 29314 32562
rect 29374 32510 29426 32562
rect 30830 32510 30882 32562
rect 31166 32510 31218 32562
rect 31838 32510 31890 32562
rect 32062 32510 32114 32562
rect 32398 32510 32450 32562
rect 33070 32510 33122 32562
rect 34526 32510 34578 32562
rect 38782 32510 38834 32562
rect 39678 32510 39730 32562
rect 41134 32510 41186 32562
rect 42142 32510 42194 32562
rect 45390 32510 45442 32562
rect 46734 32510 46786 32562
rect 48974 32510 49026 32562
rect 49198 32510 49250 32562
rect 49310 32510 49362 32562
rect 50206 32510 50258 32562
rect 51214 32510 51266 32562
rect 51550 32510 51602 32562
rect 51662 32510 51714 32562
rect 54238 32510 54290 32562
rect 55022 32510 55074 32562
rect 6078 32398 6130 32450
rect 10894 32398 10946 32450
rect 13806 32398 13858 32450
rect 15374 32398 15426 32450
rect 17950 32398 18002 32450
rect 18958 32398 19010 32450
rect 20526 32398 20578 32450
rect 21198 32398 21250 32450
rect 21982 32398 22034 32450
rect 27022 32398 27074 32450
rect 28254 32398 28306 32450
rect 29934 32398 29986 32450
rect 31614 32398 31666 32450
rect 31726 32398 31778 32450
rect 33630 32398 33682 32450
rect 37326 32398 37378 32450
rect 38110 32398 38162 32450
rect 42478 32398 42530 32450
rect 47406 32398 47458 32450
rect 47854 32398 47906 32450
rect 48862 32398 48914 32450
rect 49982 32398 50034 32450
rect 52110 32398 52162 32450
rect 14142 32286 14194 32338
rect 14366 32286 14418 32338
rect 14590 32286 14642 32338
rect 31390 32286 31442 32338
rect 39790 32286 39842 32338
rect 41022 32286 41074 32338
rect 41806 32286 41858 32338
rect 42142 32286 42194 32338
rect 51326 32286 51378 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 22094 31950 22146 32002
rect 25006 31950 25058 32002
rect 8542 31838 8594 31890
rect 10670 31838 10722 31890
rect 14702 31838 14754 31890
rect 17838 31838 17890 31890
rect 20302 31838 20354 31890
rect 24670 31838 24722 31890
rect 25902 31838 25954 31890
rect 31614 31838 31666 31890
rect 33742 31838 33794 31890
rect 34638 31838 34690 31890
rect 40350 31838 40402 31890
rect 41358 31838 41410 31890
rect 46510 31838 46562 31890
rect 48638 31838 48690 31890
rect 50430 31838 50482 31890
rect 52670 31838 52722 31890
rect 52782 31838 52834 31890
rect 7758 31726 7810 31778
rect 11006 31726 11058 31778
rect 11566 31726 11618 31778
rect 12014 31726 12066 31778
rect 12462 31726 12514 31778
rect 13470 31726 13522 31778
rect 14142 31726 14194 31778
rect 15262 31726 15314 31778
rect 16046 31726 16098 31778
rect 19742 31726 19794 31778
rect 20414 31726 20466 31778
rect 20750 31726 20802 31778
rect 21422 31726 21474 31778
rect 21646 31726 21698 31778
rect 22542 31726 22594 31778
rect 23214 31726 23266 31778
rect 23662 31726 23714 31778
rect 24222 31726 24274 31778
rect 24782 31726 24834 31778
rect 25790 31726 25842 31778
rect 26798 31726 26850 31778
rect 27918 31726 27970 31778
rect 30046 31726 30098 31778
rect 30270 31726 30322 31778
rect 30606 31726 30658 31778
rect 30942 31726 30994 31778
rect 34190 31726 34242 31778
rect 36990 31726 37042 31778
rect 37886 31726 37938 31778
rect 38558 31726 38610 31778
rect 38782 31726 38834 31778
rect 39342 31726 39394 31778
rect 39902 31726 39954 31778
rect 40238 31726 40290 31778
rect 43486 31726 43538 31778
rect 44270 31726 44322 31778
rect 45838 31726 45890 31778
rect 49422 31726 49474 31778
rect 49646 31726 49698 31778
rect 49982 31726 50034 31778
rect 50766 31726 50818 31778
rect 51214 31726 51266 31778
rect 51774 31726 51826 31778
rect 6302 31614 6354 31666
rect 14814 31614 14866 31666
rect 17166 31614 17218 31666
rect 18622 31614 18674 31666
rect 22654 31614 22706 31666
rect 26238 31614 26290 31666
rect 26462 31614 26514 31666
rect 27358 31614 27410 31666
rect 27470 31614 27522 31666
rect 29150 31614 29202 31666
rect 29262 31614 29314 31666
rect 37214 31614 37266 31666
rect 37326 31614 37378 31666
rect 37662 31614 37714 31666
rect 38894 31614 38946 31666
rect 40798 31614 40850 31666
rect 51550 31614 51602 31666
rect 6190 31502 6242 31554
rect 13694 31502 13746 31554
rect 13806 31502 13858 31554
rect 13918 31502 13970 31554
rect 14590 31502 14642 31554
rect 20190 31502 20242 31554
rect 26574 31502 26626 31554
rect 27134 31502 27186 31554
rect 27246 31502 27298 31554
rect 29486 31502 29538 31554
rect 30270 31502 30322 31554
rect 38222 31502 38274 31554
rect 44942 31502 44994 31554
rect 45390 31502 45442 31554
rect 49758 31502 49810 31554
rect 52110 31502 52162 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 8542 31166 8594 31218
rect 9102 31166 9154 31218
rect 9662 31166 9714 31218
rect 10334 31166 10386 31218
rect 14926 31166 14978 31218
rect 15822 31166 15874 31218
rect 17390 31166 17442 31218
rect 17502 31166 17554 31218
rect 18398 31166 18450 31218
rect 19070 31166 19122 31218
rect 21086 31166 21138 31218
rect 26014 31166 26066 31218
rect 27694 31166 27746 31218
rect 34638 31166 34690 31218
rect 37550 31166 37602 31218
rect 40014 31166 40066 31218
rect 40238 31166 40290 31218
rect 42142 31166 42194 31218
rect 48190 31166 48242 31218
rect 48862 31166 48914 31218
rect 49422 31166 49474 31218
rect 50542 31166 50594 31218
rect 51998 31166 52050 31218
rect 5742 31054 5794 31106
rect 8206 31054 8258 31106
rect 10558 31054 10610 31106
rect 14478 31054 14530 31106
rect 15262 31054 15314 31106
rect 15710 31054 15762 31106
rect 16606 31054 16658 31106
rect 17614 31054 17666 31106
rect 19854 31054 19906 31106
rect 24558 31054 24610 31106
rect 30158 31054 30210 31106
rect 33070 31054 33122 31106
rect 33294 31054 33346 31106
rect 33966 31054 34018 31106
rect 34078 31054 34130 31106
rect 37326 31054 37378 31106
rect 37774 31054 37826 31106
rect 38110 31054 38162 31106
rect 41918 31054 41970 31106
rect 42366 31054 42418 31106
rect 50430 31054 50482 31106
rect 5070 30942 5122 30994
rect 10894 30942 10946 30994
rect 11118 30942 11170 30994
rect 11342 30942 11394 30994
rect 12014 30942 12066 30994
rect 12574 30942 12626 30994
rect 13806 30942 13858 30994
rect 14254 30942 14306 30994
rect 15486 30942 15538 30994
rect 16270 30942 16322 30994
rect 18062 30942 18114 30994
rect 18734 30942 18786 30994
rect 19294 30942 19346 30994
rect 19630 30942 19682 30994
rect 20190 30942 20242 30994
rect 20974 30942 21026 30994
rect 21198 30942 21250 30994
rect 21422 30942 21474 30994
rect 21646 30942 21698 30994
rect 22318 30942 22370 30994
rect 22766 30942 22818 30994
rect 23326 30942 23378 30994
rect 25342 30942 25394 30994
rect 25790 30942 25842 30994
rect 25902 30942 25954 30994
rect 26686 30942 26738 30994
rect 27022 30942 27074 30994
rect 29486 30942 29538 30994
rect 33742 30942 33794 30994
rect 38334 30942 38386 30994
rect 39118 30942 39170 30994
rect 39454 30942 39506 30994
rect 40350 30942 40402 30994
rect 41022 30942 41074 30994
rect 41246 30942 41298 30994
rect 42478 30942 42530 30994
rect 50094 30942 50146 30994
rect 50654 30942 50706 30994
rect 50878 30942 50930 30994
rect 51102 30942 51154 30994
rect 51438 30942 51490 30994
rect 7870 30830 7922 30882
rect 14030 30830 14082 30882
rect 19406 30830 19458 30882
rect 20526 30830 20578 30882
rect 22206 30830 22258 30882
rect 23998 30830 24050 30882
rect 32286 30830 32338 30882
rect 33518 30830 33570 30882
rect 39566 30830 39618 30882
rect 49758 30830 49810 30882
rect 51550 30830 51602 30882
rect 10222 30718 10274 30770
rect 11790 30718 11842 30770
rect 24334 30718 24386 30770
rect 27022 30718 27074 30770
rect 34078 30718 34130 30770
rect 37886 30718 37938 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 7310 30382 7362 30434
rect 12238 30382 12290 30434
rect 12350 30382 12402 30434
rect 12574 30382 12626 30434
rect 14926 30382 14978 30434
rect 15598 30382 15650 30434
rect 18398 30382 18450 30434
rect 21422 30382 21474 30434
rect 22990 30382 23042 30434
rect 23326 30382 23378 30434
rect 24782 30382 24834 30434
rect 34750 30382 34802 30434
rect 6974 30270 7026 30322
rect 11118 30270 11170 30322
rect 13806 30270 13858 30322
rect 15710 30270 15762 30322
rect 38222 30270 38274 30322
rect 40126 30270 40178 30322
rect 41246 30270 41298 30322
rect 52110 30270 52162 30322
rect 8318 30158 8370 30210
rect 8990 30158 9042 30210
rect 11790 30158 11842 30210
rect 12798 30158 12850 30210
rect 14478 30158 14530 30210
rect 14702 30158 14754 30210
rect 15038 30158 15090 30210
rect 15934 30158 15986 30210
rect 17166 30158 17218 30210
rect 17502 30158 17554 30210
rect 18174 30158 18226 30210
rect 18622 30158 18674 30210
rect 18958 30158 19010 30210
rect 21534 30158 21586 30210
rect 21982 30158 22034 30210
rect 22318 30158 22370 30210
rect 22990 30158 23042 30210
rect 23998 30158 24050 30210
rect 24334 30158 24386 30210
rect 24894 30158 24946 30210
rect 25230 30158 25282 30210
rect 25342 30158 25394 30210
rect 25790 30158 25842 30210
rect 28702 30158 28754 30210
rect 29150 30158 29202 30210
rect 35870 30158 35922 30210
rect 37774 30158 37826 30210
rect 38782 30158 38834 30210
rect 39118 30158 39170 30210
rect 39790 30158 39842 30210
rect 40238 30158 40290 30210
rect 48862 30158 48914 30210
rect 49310 30158 49362 30210
rect 49982 30158 50034 30210
rect 13470 30046 13522 30098
rect 15262 30046 15314 30098
rect 17390 30046 17442 30098
rect 17838 30046 17890 30098
rect 22654 30046 22706 30098
rect 26686 30046 26738 30098
rect 32846 30046 32898 30098
rect 36430 30046 36482 30098
rect 37326 30046 37378 30098
rect 41470 30046 41522 30098
rect 7086 29934 7138 29986
rect 12686 29934 12738 29986
rect 13694 29934 13746 29986
rect 13918 29934 13970 29986
rect 14142 29934 14194 29986
rect 14366 29934 14418 29986
rect 17950 29934 18002 29986
rect 19518 29934 19570 29986
rect 21422 29934 21474 29986
rect 22542 29934 22594 29986
rect 24110 29934 24162 29986
rect 24782 29934 24834 29986
rect 27022 29934 27074 29986
rect 34862 29934 34914 29986
rect 34974 29934 35026 29986
rect 40910 29934 40962 29986
rect 41358 29934 41410 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 11230 29598 11282 29650
rect 12014 29598 12066 29650
rect 18622 29598 18674 29650
rect 20526 29598 20578 29650
rect 22094 29598 22146 29650
rect 22878 29598 22930 29650
rect 23550 29598 23602 29650
rect 27470 29598 27522 29650
rect 28366 29598 28418 29650
rect 28702 29598 28754 29650
rect 35758 29598 35810 29650
rect 6862 29486 6914 29538
rect 13134 29486 13186 29538
rect 13358 29486 13410 29538
rect 15038 29486 15090 29538
rect 15150 29486 15202 29538
rect 19070 29486 19122 29538
rect 20862 29486 20914 29538
rect 23662 29486 23714 29538
rect 29598 29486 29650 29538
rect 29934 29486 29986 29538
rect 32286 29486 32338 29538
rect 34302 29486 34354 29538
rect 37438 29486 37490 29538
rect 40350 29486 40402 29538
rect 43374 29486 43426 29538
rect 6190 29374 6242 29426
rect 12686 29374 12738 29426
rect 13806 29374 13858 29426
rect 14254 29374 14306 29426
rect 15822 29374 15874 29426
rect 16494 29374 16546 29426
rect 17502 29374 17554 29426
rect 17950 29374 18002 29426
rect 22542 29374 22594 29426
rect 26462 29374 26514 29426
rect 26910 29374 26962 29426
rect 27806 29374 27858 29426
rect 29262 29374 29314 29426
rect 31950 29374 32002 29426
rect 32510 29374 32562 29426
rect 33070 29374 33122 29426
rect 33406 29374 33458 29426
rect 33518 29374 33570 29426
rect 33630 29374 33682 29426
rect 35870 29374 35922 29426
rect 36318 29374 36370 29426
rect 39678 29374 39730 29426
rect 40238 29374 40290 29426
rect 44046 29374 44098 29426
rect 44606 29374 44658 29426
rect 8990 29262 9042 29314
rect 9774 29262 9826 29314
rect 11566 29262 11618 29314
rect 13470 29262 13522 29314
rect 16606 29262 16658 29314
rect 20974 29262 21026 29314
rect 25454 29262 25506 29314
rect 25902 29262 25954 29314
rect 27134 29262 27186 29314
rect 32398 29262 32450 29314
rect 38894 29262 38946 29314
rect 41246 29262 41298 29314
rect 12462 29150 12514 29202
rect 14478 29150 14530 29202
rect 15038 29150 15090 29202
rect 15598 29150 15650 29202
rect 17278 29150 17330 29202
rect 17950 29150 18002 29202
rect 19182 29150 19234 29202
rect 38334 29150 38386 29202
rect 38670 29150 38722 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 13694 28814 13746 28866
rect 14814 28814 14866 28866
rect 16158 28814 16210 28866
rect 23438 28814 23490 28866
rect 32398 28814 32450 28866
rect 42142 28814 42194 28866
rect 6974 28702 7026 28754
rect 14702 28702 14754 28754
rect 18398 28702 18450 28754
rect 19966 28702 20018 28754
rect 24446 28702 24498 28754
rect 27470 28702 27522 28754
rect 28366 28702 28418 28754
rect 32062 28702 32114 28754
rect 33854 28702 33906 28754
rect 35982 28702 36034 28754
rect 36990 28702 37042 28754
rect 38446 28702 38498 28754
rect 6526 28590 6578 28642
rect 13470 28590 13522 28642
rect 17054 28590 17106 28642
rect 17278 28590 17330 28642
rect 18286 28590 18338 28642
rect 18958 28590 19010 28642
rect 19070 28590 19122 28642
rect 19182 28590 19234 28642
rect 19406 28590 19458 28642
rect 20302 28590 20354 28642
rect 21422 28590 21474 28642
rect 22094 28590 22146 28642
rect 22654 28590 22706 28642
rect 23102 28590 23154 28642
rect 25678 28590 25730 28642
rect 26350 28590 26402 28642
rect 26910 28590 26962 28642
rect 27022 28590 27074 28642
rect 27358 28590 27410 28642
rect 27694 28590 27746 28642
rect 29262 28590 29314 28642
rect 33182 28590 33234 28642
rect 37438 28590 37490 28642
rect 37998 28590 38050 28642
rect 38894 28590 38946 28642
rect 39790 28590 39842 28642
rect 40126 28590 40178 28642
rect 41806 28590 41858 28642
rect 41918 28590 41970 28642
rect 16046 28478 16098 28530
rect 16718 28478 16770 28530
rect 18622 28478 18674 28530
rect 20638 28478 20690 28530
rect 22430 28478 22482 28530
rect 23326 28478 23378 28530
rect 23438 28478 23490 28530
rect 25342 28478 25394 28530
rect 29934 28478 29986 28530
rect 32622 28478 32674 28530
rect 36430 28478 36482 28530
rect 38110 28478 38162 28530
rect 39454 28478 39506 28530
rect 39566 28478 39618 28530
rect 42254 28478 42306 28530
rect 6190 28366 6242 28418
rect 14030 28366 14082 28418
rect 16158 28366 16210 28418
rect 17726 28366 17778 28418
rect 17838 28366 17890 28418
rect 17950 28366 18002 28418
rect 21870 28366 21922 28418
rect 21982 28366 22034 28418
rect 22542 28366 22594 28418
rect 24110 28366 24162 28418
rect 32510 28366 32562 28418
rect 40238 28366 40290 28418
rect 40462 28366 40514 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 8206 28030 8258 28082
rect 16046 28030 16098 28082
rect 16606 28030 16658 28082
rect 24782 28030 24834 28082
rect 25454 28030 25506 28082
rect 29598 28030 29650 28082
rect 30046 28030 30098 28082
rect 30606 28030 30658 28082
rect 36430 28030 36482 28082
rect 37662 28030 37714 28082
rect 37998 28030 38050 28082
rect 10222 27918 10274 27970
rect 16718 27918 16770 27970
rect 18174 27918 18226 27970
rect 22766 27918 22818 27970
rect 30158 27918 30210 27970
rect 33854 27918 33906 27970
rect 37102 27918 37154 27970
rect 40126 27918 40178 27970
rect 41694 27918 41746 27970
rect 4958 27806 5010 27858
rect 9886 27806 9938 27858
rect 10558 27806 10610 27858
rect 13134 27806 13186 27858
rect 13358 27806 13410 27858
rect 13582 27806 13634 27858
rect 17502 27806 17554 27858
rect 23438 27806 23490 27858
rect 29822 27806 29874 27858
rect 32286 27806 32338 27858
rect 33182 27806 33234 27858
rect 37326 27806 37378 27858
rect 38334 27806 38386 27858
rect 38558 27806 38610 27858
rect 38894 27806 38946 27858
rect 39342 27806 39394 27858
rect 39790 27806 39842 27858
rect 40798 27806 40850 27858
rect 41918 27806 41970 27858
rect 5630 27694 5682 27746
rect 7758 27694 7810 27746
rect 15150 27694 15202 27746
rect 15598 27694 15650 27746
rect 20302 27694 20354 27746
rect 20638 27694 20690 27746
rect 24334 27694 24386 27746
rect 35982 27694 36034 27746
rect 41470 27694 41522 27746
rect 9550 27582 9602 27634
rect 9886 27582 9938 27634
rect 13022 27582 13074 27634
rect 15150 27582 15202 27634
rect 16270 27582 16322 27634
rect 25230 27582 25282 27634
rect 25566 27582 25618 27634
rect 30494 27582 30546 27634
rect 30830 27582 30882 27634
rect 39790 27582 39842 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 5742 27246 5794 27298
rect 12462 27246 12514 27298
rect 41470 27246 41522 27298
rect 6078 27134 6130 27186
rect 6526 27134 6578 27186
rect 9550 27134 9602 27186
rect 10222 27134 10274 27186
rect 14702 27134 14754 27186
rect 15822 27134 15874 27186
rect 17950 27134 18002 27186
rect 18734 27134 18786 27186
rect 19294 27134 19346 27186
rect 22430 27134 22482 27186
rect 25678 27134 25730 27186
rect 29934 27134 29986 27186
rect 32062 27134 32114 27186
rect 33406 27134 33458 27186
rect 35534 27134 35586 27186
rect 36430 27134 36482 27186
rect 39902 27134 39954 27186
rect 40798 27134 40850 27186
rect 7982 27022 8034 27074
rect 8878 27022 8930 27074
rect 9662 27022 9714 27074
rect 10446 27022 10498 27074
rect 11454 27022 11506 27074
rect 12238 27022 12290 27074
rect 15038 27022 15090 27074
rect 22878 27022 22930 27074
rect 23550 27022 23602 27074
rect 29262 27022 29314 27074
rect 32734 27022 32786 27074
rect 35870 27022 35922 27074
rect 36990 27022 37042 27074
rect 40686 27022 40738 27074
rect 41806 27022 41858 27074
rect 42142 27022 42194 27074
rect 5854 26910 5906 26962
rect 7646 26910 7698 26962
rect 8542 26910 8594 26962
rect 9326 26910 9378 26962
rect 11118 26910 11170 26962
rect 11566 26910 11618 26962
rect 11902 26910 11954 26962
rect 14254 26910 14306 26962
rect 37774 26910 37826 26962
rect 42030 26910 42082 26962
rect 42478 26910 42530 26962
rect 14590 26798 14642 26850
rect 18622 26798 18674 26850
rect 20526 26798 20578 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 7198 26462 7250 26514
rect 9998 26462 10050 26514
rect 14590 26462 14642 26514
rect 15822 26462 15874 26514
rect 16494 26462 16546 26514
rect 20974 26462 21026 26514
rect 35534 26462 35586 26514
rect 35982 26462 36034 26514
rect 36430 26462 36482 26514
rect 39678 26462 39730 26514
rect 39902 26462 39954 26514
rect 40462 26462 40514 26514
rect 41358 26462 41410 26514
rect 41470 26462 41522 26514
rect 42142 26462 42194 26514
rect 8878 26350 8930 26402
rect 12238 26350 12290 26402
rect 13134 26350 13186 26402
rect 14366 26350 14418 26402
rect 17502 26350 17554 26402
rect 18622 26350 18674 26402
rect 19854 26350 19906 26402
rect 26014 26350 26066 26402
rect 31054 26350 31106 26402
rect 36766 26350 36818 26402
rect 3502 26238 3554 26290
rect 7310 26238 7362 26290
rect 8430 26238 8482 26290
rect 8766 26238 8818 26290
rect 9550 26238 9602 26290
rect 9774 26238 9826 26290
rect 10222 26238 10274 26290
rect 10894 26238 10946 26290
rect 13358 26238 13410 26290
rect 15038 26238 15090 26290
rect 15262 26238 15314 26290
rect 15822 26238 15874 26290
rect 16046 26238 16098 26290
rect 16718 26238 16770 26290
rect 18286 26238 18338 26290
rect 18846 26238 18898 26290
rect 19182 26238 19234 26290
rect 25342 26238 25394 26290
rect 30606 26238 30658 26290
rect 36878 26238 36930 26290
rect 37102 26238 37154 26290
rect 37326 26238 37378 26290
rect 39566 26238 39618 26290
rect 40910 26238 40962 26290
rect 41246 26238 41298 26290
rect 41806 26238 41858 26290
rect 4174 26126 4226 26178
rect 6302 26126 6354 26178
rect 6750 26126 6802 26178
rect 9662 26126 9714 26178
rect 13246 26126 13298 26178
rect 16606 26126 16658 26178
rect 18734 26126 18786 26178
rect 20302 26126 20354 26178
rect 24670 26126 24722 26178
rect 28142 26126 28194 26178
rect 30830 26126 30882 26178
rect 31390 26126 31442 26178
rect 31614 26126 31666 26178
rect 32398 26126 32450 26178
rect 7198 26014 7250 26066
rect 14702 26014 14754 26066
rect 15486 26014 15538 26066
rect 17390 26014 17442 26066
rect 17950 26014 18002 26066
rect 18286 26014 18338 26066
rect 19070 26014 19122 26066
rect 31950 26014 32002 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 5630 25678 5682 25730
rect 5966 25678 6018 25730
rect 14926 25678 14978 25730
rect 30718 25678 30770 25730
rect 7198 25566 7250 25618
rect 7646 25566 7698 25618
rect 10334 25566 10386 25618
rect 11230 25566 11282 25618
rect 12350 25566 12402 25618
rect 12798 25566 12850 25618
rect 17278 25566 17330 25618
rect 18622 25566 18674 25618
rect 20750 25566 20802 25618
rect 22094 25566 22146 25618
rect 24222 25566 24274 25618
rect 28590 25566 28642 25618
rect 30494 25566 30546 25618
rect 36542 25566 36594 25618
rect 39454 25566 39506 25618
rect 41582 25566 41634 25618
rect 42814 25566 42866 25618
rect 5630 25454 5682 25506
rect 7310 25454 7362 25506
rect 9550 25454 9602 25506
rect 10782 25454 10834 25506
rect 12238 25454 12290 25506
rect 13022 25454 13074 25506
rect 14478 25454 14530 25506
rect 14702 25454 14754 25506
rect 15150 25454 15202 25506
rect 15934 25454 15986 25506
rect 16606 25454 16658 25506
rect 17390 25454 17442 25506
rect 17838 25454 17890 25506
rect 21310 25454 21362 25506
rect 25790 25454 25842 25506
rect 42366 25454 42418 25506
rect 8766 25342 8818 25394
rect 9326 25342 9378 25394
rect 9662 25342 9714 25394
rect 14142 25342 14194 25394
rect 17502 25342 17554 25394
rect 26462 25342 26514 25394
rect 13806 25230 13858 25282
rect 14590 25230 14642 25282
rect 16046 25230 16098 25282
rect 24670 25230 24722 25282
rect 25342 25230 25394 25282
rect 31054 25230 31106 25282
rect 33630 25230 33682 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 10782 24894 10834 24946
rect 11006 24894 11058 24946
rect 36430 24894 36482 24946
rect 36878 24894 36930 24946
rect 7870 24782 7922 24834
rect 10334 24782 10386 24834
rect 10670 24782 10722 24834
rect 13470 24782 13522 24834
rect 14590 24782 14642 24834
rect 16830 24782 16882 24834
rect 17838 24782 17890 24834
rect 20078 24782 20130 24834
rect 20862 24782 20914 24834
rect 28926 24782 28978 24834
rect 32510 24782 32562 24834
rect 33854 24782 33906 24834
rect 9774 24670 9826 24722
rect 14254 24670 14306 24722
rect 15038 24670 15090 24722
rect 17614 24670 17666 24722
rect 18062 24670 18114 24722
rect 18510 24670 18562 24722
rect 18734 24670 18786 24722
rect 19070 24670 19122 24722
rect 19294 24670 19346 24722
rect 20414 24670 20466 24722
rect 20750 24670 20802 24722
rect 21086 24670 21138 24722
rect 32174 24670 32226 24722
rect 33182 24670 33234 24722
rect 7646 24558 7698 24610
rect 9662 24558 9714 24610
rect 11342 24558 11394 24610
rect 15486 24558 15538 24610
rect 16382 24558 16434 24610
rect 18286 24558 18338 24610
rect 26910 24558 26962 24610
rect 35982 24558 36034 24610
rect 38222 24558 38274 24610
rect 38670 24558 38722 24610
rect 8654 24446 8706 24498
rect 19630 24446 19682 24498
rect 26798 24446 26850 24498
rect 28814 24446 28866 24498
rect 38110 24446 38162 24498
rect 38558 24446 38610 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 9326 24110 9378 24162
rect 14590 24110 14642 24162
rect 32062 24110 32114 24162
rect 8766 23998 8818 24050
rect 12910 23998 12962 24050
rect 14030 23998 14082 24050
rect 18398 23998 18450 24050
rect 26910 23998 26962 24050
rect 29486 23998 29538 24050
rect 35982 23998 36034 24050
rect 39902 23998 39954 24050
rect 5630 23886 5682 23938
rect 7310 23886 7362 23938
rect 8542 23886 8594 23938
rect 10110 23886 10162 23938
rect 13470 23886 13522 23938
rect 14814 23886 14866 23938
rect 15038 23886 15090 23938
rect 15822 23886 15874 23938
rect 15934 23886 15986 23938
rect 16046 23886 16098 23938
rect 16494 23886 16546 23938
rect 18174 23886 18226 23938
rect 19742 23886 19794 23938
rect 20414 23886 20466 23938
rect 20638 23886 20690 23938
rect 23998 23886 24050 23938
rect 32398 23886 32450 23938
rect 33630 23886 33682 23938
rect 36990 23886 37042 23938
rect 5966 23774 6018 23826
rect 6974 23774 7026 23826
rect 7086 23774 7138 23826
rect 7534 23774 7586 23826
rect 7870 23774 7922 23826
rect 9214 23774 9266 23826
rect 10782 23774 10834 23826
rect 14478 23774 14530 23826
rect 16830 23774 16882 23826
rect 17390 23774 17442 23826
rect 18958 23774 19010 23826
rect 20302 23774 20354 23826
rect 21310 23774 21362 23826
rect 23550 23774 23602 23826
rect 24782 23774 24834 23826
rect 27470 23774 27522 23826
rect 27694 23774 27746 23826
rect 28030 23774 28082 23826
rect 29150 23774 29202 23826
rect 32622 23774 32674 23826
rect 33182 23774 33234 23826
rect 37774 23774 37826 23826
rect 5854 23662 5906 23714
rect 7198 23662 7250 23714
rect 15374 23662 15426 23714
rect 19070 23662 19122 23714
rect 21646 23662 21698 23714
rect 22206 23662 22258 23714
rect 23214 23662 23266 23714
rect 23662 23662 23714 23714
rect 27806 23662 27858 23714
rect 29374 23662 29426 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 7310 23326 7362 23378
rect 7534 23326 7586 23378
rect 7646 23326 7698 23378
rect 13582 23326 13634 23378
rect 21422 23326 21474 23378
rect 25566 23326 25618 23378
rect 3950 23214 4002 23266
rect 8318 23214 8370 23266
rect 14254 23214 14306 23266
rect 15150 23214 15202 23266
rect 15374 23214 15426 23266
rect 16494 23214 16546 23266
rect 18398 23214 18450 23266
rect 20750 23214 20802 23266
rect 20862 23214 20914 23266
rect 27246 23214 27298 23266
rect 31726 23214 31778 23266
rect 32062 23214 32114 23266
rect 33182 23214 33234 23266
rect 33742 23214 33794 23266
rect 34078 23214 34130 23266
rect 34862 23214 34914 23266
rect 3278 23102 3330 23154
rect 7422 23102 7474 23154
rect 7870 23102 7922 23154
rect 8206 23102 8258 23154
rect 10110 23102 10162 23154
rect 11454 23102 11506 23154
rect 12910 23102 12962 23154
rect 13470 23102 13522 23154
rect 16718 23102 16770 23154
rect 17390 23102 17442 23154
rect 20974 23102 21026 23154
rect 24670 23102 24722 23154
rect 25230 23102 25282 23154
rect 25566 23102 25618 23154
rect 25902 23102 25954 23154
rect 26126 23102 26178 23154
rect 26462 23102 26514 23154
rect 27694 23102 27746 23154
rect 31054 23102 31106 23154
rect 35870 23102 35922 23154
rect 6078 22990 6130 23042
rect 6526 22990 6578 23042
rect 10334 22990 10386 23042
rect 10782 22990 10834 23042
rect 19182 22990 19234 23042
rect 19742 22990 19794 23042
rect 21758 22990 21810 23042
rect 23886 22990 23938 23042
rect 26238 22990 26290 23042
rect 27358 22990 27410 23042
rect 28478 22990 28530 23042
rect 30606 22990 30658 23042
rect 32510 22990 32562 23042
rect 35310 22990 35362 23042
rect 36542 22990 36594 23042
rect 38670 22990 38722 23042
rect 15486 22878 15538 22930
rect 16718 22878 16770 22930
rect 27022 22878 27074 22930
rect 30942 22878 30994 22930
rect 33518 22878 33570 22930
rect 34750 22878 34802 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 14142 22542 14194 22594
rect 14926 22542 14978 22594
rect 20414 22542 20466 22594
rect 21310 22542 21362 22594
rect 21982 22542 22034 22594
rect 24782 22542 24834 22594
rect 25118 22542 25170 22594
rect 8542 22430 8594 22482
rect 8990 22430 9042 22482
rect 12910 22430 12962 22482
rect 13806 22430 13858 22482
rect 14254 22430 14306 22482
rect 15150 22430 15202 22482
rect 20190 22430 20242 22482
rect 27358 22430 27410 22482
rect 29262 22430 29314 22482
rect 31726 22430 31778 22482
rect 33854 22430 33906 22482
rect 35086 22430 35138 22482
rect 35982 22430 36034 22482
rect 37438 22430 37490 22482
rect 42478 22430 42530 22482
rect 42926 22430 42978 22482
rect 43374 22430 43426 22482
rect 5742 22318 5794 22370
rect 11118 22318 11170 22370
rect 15710 22318 15762 22370
rect 17390 22318 17442 22370
rect 19070 22318 19122 22370
rect 23438 22318 23490 22370
rect 23662 22318 23714 22370
rect 24222 22318 24274 22370
rect 25118 22318 25170 22370
rect 29038 22318 29090 22370
rect 29374 22318 29426 22370
rect 29598 22318 29650 22370
rect 31054 22318 31106 22370
rect 35646 22318 35698 22370
rect 36990 22318 37042 22370
rect 39678 22318 39730 22370
rect 6414 22206 6466 22258
rect 11678 22206 11730 22258
rect 16830 22206 16882 22258
rect 18286 22206 18338 22258
rect 21534 22206 21586 22258
rect 22206 22206 22258 22258
rect 23102 22206 23154 22258
rect 23998 22206 24050 22258
rect 35310 22206 35362 22258
rect 35870 22206 35922 22258
rect 37550 22206 37602 22258
rect 37886 22206 37938 22258
rect 40350 22206 40402 22258
rect 14590 22094 14642 22146
rect 19630 22094 19682 22146
rect 20750 22094 20802 22146
rect 21422 22094 21474 22146
rect 22094 22094 22146 22146
rect 22878 22094 22930 22146
rect 23214 22094 23266 22146
rect 23886 22094 23938 22146
rect 25566 22094 25618 22146
rect 34302 22094 34354 22146
rect 35422 22094 35474 22146
rect 36094 22094 36146 22146
rect 36318 22094 36370 22146
rect 37326 22094 37378 22146
rect 37998 22094 38050 22146
rect 38222 22094 38274 22146
rect 42814 22094 42866 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 5854 21758 5906 21810
rect 6750 21758 6802 21810
rect 7310 21758 7362 21810
rect 21086 21758 21138 21810
rect 21982 21758 22034 21810
rect 28030 21758 28082 21810
rect 28590 21758 28642 21810
rect 35198 21758 35250 21810
rect 40238 21758 40290 21810
rect 6078 21646 6130 21698
rect 6414 21646 6466 21698
rect 6526 21646 6578 21698
rect 7534 21646 7586 21698
rect 11342 21646 11394 21698
rect 17502 21646 17554 21698
rect 20526 21646 20578 21698
rect 21870 21646 21922 21698
rect 29486 21646 29538 21698
rect 33182 21646 33234 21698
rect 33854 21646 33906 21698
rect 39342 21646 39394 21698
rect 5630 21534 5682 21586
rect 5966 21534 6018 21586
rect 10222 21534 10274 21586
rect 12126 21534 12178 21586
rect 15934 21534 15986 21586
rect 16606 21534 16658 21586
rect 17390 21534 17442 21586
rect 19406 21534 19458 21586
rect 21982 21534 22034 21586
rect 22654 21534 22706 21586
rect 23998 21534 24050 21586
rect 24670 21534 24722 21586
rect 27918 21534 27970 21586
rect 29374 21534 29426 21586
rect 29710 21534 29762 21586
rect 32286 21534 32338 21586
rect 33518 21534 33570 21586
rect 34638 21534 34690 21586
rect 35758 21534 35810 21586
rect 39790 21534 39842 21586
rect 40126 21534 40178 21586
rect 40350 21534 40402 21586
rect 40910 21534 40962 21586
rect 7198 21422 7250 21474
rect 12574 21422 12626 21474
rect 13022 21422 13074 21474
rect 15150 21422 15202 21474
rect 16382 21422 16434 21474
rect 22990 21422 23042 21474
rect 23774 21422 23826 21474
rect 25342 21422 25394 21474
rect 30046 21422 30098 21474
rect 34414 21422 34466 21474
rect 36542 21422 36594 21474
rect 38670 21422 38722 21474
rect 39454 21422 39506 21474
rect 41694 21422 41746 21474
rect 43822 21422 43874 21474
rect 44270 21422 44322 21474
rect 6862 21310 6914 21362
rect 16270 21310 16322 21362
rect 16718 21310 16770 21362
rect 23662 21310 23714 21362
rect 24334 21310 24386 21362
rect 24670 21310 24722 21362
rect 28030 21310 28082 21362
rect 33070 21310 33122 21362
rect 34862 21310 34914 21362
rect 39118 21310 39170 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 6302 20974 6354 21026
rect 10782 20862 10834 20914
rect 12462 20862 12514 20914
rect 13582 20862 13634 20914
rect 14926 20862 14978 20914
rect 15598 20862 15650 20914
rect 19182 20862 19234 20914
rect 20526 20862 20578 20914
rect 25342 20862 25394 20914
rect 28590 20862 28642 20914
rect 32062 20862 32114 20914
rect 35646 20862 35698 20914
rect 37102 20862 37154 20914
rect 37998 20862 38050 20914
rect 39678 20862 39730 20914
rect 40574 20862 40626 20914
rect 42366 20862 42418 20914
rect 6638 20750 6690 20802
rect 7982 20750 8034 20802
rect 12574 20750 12626 20802
rect 14030 20750 14082 20802
rect 14366 20750 14418 20802
rect 16606 20750 16658 20802
rect 16942 20750 16994 20802
rect 17502 20750 17554 20802
rect 20414 20750 20466 20802
rect 22430 20750 22482 20802
rect 25678 20750 25730 20802
rect 29262 20750 29314 20802
rect 32622 20750 32674 20802
rect 33294 20750 33346 20802
rect 36430 20750 36482 20802
rect 36878 20750 36930 20802
rect 39006 20750 39058 20802
rect 40126 20750 40178 20802
rect 40462 20750 40514 20802
rect 8654 20638 8706 20690
rect 11454 20638 11506 20690
rect 11790 20638 11842 20690
rect 15374 20638 15426 20690
rect 16718 20638 16770 20690
rect 18398 20638 18450 20690
rect 21870 20638 21922 20690
rect 21982 20638 22034 20690
rect 23214 20638 23266 20690
rect 26462 20638 26514 20690
rect 29934 20638 29986 20690
rect 37326 20638 37378 20690
rect 37550 20638 37602 20690
rect 38334 20638 38386 20690
rect 38446 20638 38498 20690
rect 38670 20638 38722 20690
rect 39790 20638 39842 20690
rect 40686 20638 40738 20690
rect 42254 20638 42306 20690
rect 6414 20526 6466 20578
rect 11230 20526 11282 20578
rect 11342 20526 11394 20578
rect 18958 20526 19010 20578
rect 21534 20526 21586 20578
rect 22206 20526 22258 20578
rect 32398 20526 32450 20578
rect 36094 20526 36146 20578
rect 36318 20526 36370 20578
rect 37886 20526 37938 20578
rect 39566 20526 39618 20578
rect 41246 20526 41298 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 13358 20190 13410 20242
rect 16718 20190 16770 20242
rect 19742 20190 19794 20242
rect 27246 20190 27298 20242
rect 27582 20190 27634 20242
rect 28030 20190 28082 20242
rect 29374 20190 29426 20242
rect 29486 20190 29538 20242
rect 40238 20190 40290 20242
rect 11006 20078 11058 20130
rect 13134 20078 13186 20130
rect 13470 20078 13522 20130
rect 15822 20078 15874 20130
rect 18398 20078 18450 20130
rect 24222 20078 24274 20130
rect 24670 20078 24722 20130
rect 25566 20078 25618 20130
rect 27694 20078 27746 20130
rect 28590 20078 28642 20130
rect 30942 20078 30994 20130
rect 31278 20078 31330 20130
rect 31614 20078 31666 20130
rect 31950 20078 32002 20130
rect 32286 20078 32338 20130
rect 35086 20078 35138 20130
rect 36766 20078 36818 20130
rect 37662 20078 37714 20130
rect 38670 20078 38722 20130
rect 38782 20078 38834 20130
rect 39678 20078 39730 20130
rect 40014 20078 40066 20130
rect 12350 19966 12402 20018
rect 15038 19966 15090 20018
rect 16718 19966 16770 20018
rect 17390 19966 17442 20018
rect 20414 19966 20466 20018
rect 23662 19966 23714 20018
rect 23998 19966 24050 20018
rect 24446 19966 24498 20018
rect 25454 19966 25506 20018
rect 27806 19966 27858 20018
rect 29598 19966 29650 20018
rect 30046 19966 30098 20018
rect 30830 19966 30882 20018
rect 33070 19966 33122 20018
rect 34190 19966 34242 20018
rect 35310 19966 35362 20018
rect 35870 19966 35922 20018
rect 36206 19966 36258 20018
rect 36542 19966 36594 20018
rect 39006 19966 39058 20018
rect 41134 19966 41186 20018
rect 12126 19854 12178 19906
rect 12910 19854 12962 19906
rect 19182 19854 19234 19906
rect 21086 19854 21138 19906
rect 23214 19854 23266 19906
rect 26350 19854 26402 19906
rect 26686 19854 26738 19906
rect 26910 19854 26962 19906
rect 28478 19854 28530 19906
rect 33518 19854 33570 19906
rect 34638 19854 34690 19906
rect 36654 19854 36706 19906
rect 37214 19854 37266 19906
rect 38334 19854 38386 19906
rect 40238 19854 40290 19906
rect 42254 19854 42306 19906
rect 23550 19742 23602 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 12126 19406 12178 19458
rect 12462 19406 12514 19458
rect 32846 19406 32898 19458
rect 33518 19406 33570 19458
rect 8094 19294 8146 19346
rect 10222 19294 10274 19346
rect 10670 19294 10722 19346
rect 16158 19294 16210 19346
rect 19518 19294 19570 19346
rect 20750 19294 20802 19346
rect 22094 19294 22146 19346
rect 23998 19294 24050 19346
rect 33406 19294 33458 19346
rect 35982 19294 36034 19346
rect 37774 19294 37826 19346
rect 39902 19294 39954 19346
rect 42814 19294 42866 19346
rect 7422 19182 7474 19234
rect 12126 19182 12178 19234
rect 14478 19182 14530 19234
rect 15038 19182 15090 19234
rect 17726 19182 17778 19234
rect 21646 19182 21698 19234
rect 21982 19182 22034 19234
rect 22318 19182 22370 19234
rect 22542 19182 22594 19234
rect 22878 19182 22930 19234
rect 27582 19182 27634 19234
rect 29934 19182 29986 19234
rect 33742 19182 33794 19234
rect 35086 19182 35138 19234
rect 35758 19182 35810 19234
rect 37102 19182 37154 19234
rect 41022 19182 41074 19234
rect 15262 19070 15314 19122
rect 18286 19070 18338 19122
rect 22990 19070 23042 19122
rect 24446 19070 24498 19122
rect 32958 19070 33010 19122
rect 34526 19070 34578 19122
rect 34750 19070 34802 19122
rect 35422 19070 35474 19122
rect 36094 19070 36146 19122
rect 43486 19070 43538 19122
rect 14142 18958 14194 19010
rect 19630 18958 19682 19010
rect 21310 18958 21362 19010
rect 23438 18958 23490 19010
rect 26126 18958 26178 19010
rect 27358 18958 27410 19010
rect 29598 18958 29650 19010
rect 29822 18958 29874 19010
rect 34078 18958 34130 19010
rect 34638 18958 34690 19010
rect 43374 18958 43426 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 22542 18622 22594 18674
rect 26350 18622 26402 18674
rect 32398 18622 32450 18674
rect 35422 18622 35474 18674
rect 35870 18622 35922 18674
rect 38782 18622 38834 18674
rect 44270 18622 44322 18674
rect 11790 18510 11842 18562
rect 17502 18510 17554 18562
rect 18510 18510 18562 18562
rect 23326 18510 23378 18562
rect 23662 18510 23714 18562
rect 24670 18510 24722 18562
rect 25230 18510 25282 18562
rect 27358 18510 27410 18562
rect 27470 18510 27522 18562
rect 27806 18510 27858 18562
rect 29262 18510 29314 18562
rect 32510 18510 32562 18562
rect 33294 18510 33346 18562
rect 39118 18510 39170 18562
rect 39790 18510 39842 18562
rect 6078 18398 6130 18450
rect 6750 18398 6802 18450
rect 9662 18398 9714 18450
rect 11902 18398 11954 18450
rect 12350 18398 12402 18450
rect 17838 18398 17890 18450
rect 18286 18398 18338 18450
rect 18846 18398 18898 18450
rect 23102 18398 23154 18450
rect 23998 18398 24050 18450
rect 24334 18398 24386 18450
rect 25566 18398 25618 18450
rect 26014 18398 26066 18450
rect 26574 18398 26626 18450
rect 27022 18398 27074 18450
rect 28030 18398 28082 18450
rect 28366 18398 28418 18450
rect 28814 18398 28866 18450
rect 29038 18398 29090 18450
rect 29710 18398 29762 18450
rect 29822 18398 29874 18450
rect 30270 18398 30322 18450
rect 30494 18398 30546 18450
rect 30718 18398 30770 18450
rect 31166 18398 31218 18450
rect 33070 18398 33122 18450
rect 33630 18398 33682 18450
rect 34414 18398 34466 18450
rect 34638 18398 34690 18450
rect 35086 18398 35138 18450
rect 36094 18398 36146 18450
rect 38110 18398 38162 18450
rect 39454 18398 39506 18450
rect 40014 18398 40066 18450
rect 40350 18398 40402 18450
rect 40910 18398 40962 18450
rect 8878 18286 8930 18338
rect 13134 18286 13186 18338
rect 15262 18286 15314 18338
rect 15710 18286 15762 18338
rect 19630 18286 19682 18338
rect 21758 18286 21810 18338
rect 25342 18286 25394 18338
rect 26462 18286 26514 18338
rect 27918 18286 27970 18338
rect 29150 18286 29202 18338
rect 30046 18286 30098 18338
rect 30942 18286 30994 18338
rect 33518 18286 33570 18338
rect 34862 18286 34914 18338
rect 35982 18286 36034 18338
rect 37998 18286 38050 18338
rect 39902 18286 39954 18338
rect 41694 18286 41746 18338
rect 43822 18286 43874 18338
rect 10782 18174 10834 18226
rect 11118 18174 11170 18226
rect 25678 18174 25730 18226
rect 27358 18174 27410 18226
rect 32398 18174 32450 18226
rect 39454 18174 39506 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 14478 17838 14530 17890
rect 19294 17838 19346 17890
rect 24782 17838 24834 17890
rect 36094 17838 36146 17890
rect 11342 17726 11394 17778
rect 12014 17726 12066 17778
rect 12462 17726 12514 17778
rect 18286 17726 18338 17778
rect 18846 17726 18898 17778
rect 21534 17726 21586 17778
rect 27806 17726 27858 17778
rect 36206 17726 36258 17778
rect 39006 17726 39058 17778
rect 40574 17726 40626 17778
rect 42702 17726 42754 17778
rect 7870 17614 7922 17666
rect 8430 17614 8482 17666
rect 13806 17614 13858 17666
rect 15486 17614 15538 17666
rect 19630 17614 19682 17666
rect 23886 17614 23938 17666
rect 24782 17614 24834 17666
rect 25902 17614 25954 17666
rect 27022 17614 27074 17666
rect 29486 17614 29538 17666
rect 32846 17614 32898 17666
rect 33518 17614 33570 17666
rect 34078 17614 34130 17666
rect 35086 17614 35138 17666
rect 35534 17614 35586 17666
rect 36878 17614 36930 17666
rect 37438 17614 37490 17666
rect 38894 17614 38946 17666
rect 39118 17614 39170 17666
rect 39454 17614 39506 17666
rect 39902 17614 39954 17666
rect 9214 17502 9266 17554
rect 13470 17502 13522 17554
rect 16158 17502 16210 17554
rect 19854 17502 19906 17554
rect 20190 17502 20242 17554
rect 24446 17502 24498 17554
rect 26238 17502 26290 17554
rect 26350 17502 26402 17554
rect 27358 17502 27410 17554
rect 27470 17502 27522 17554
rect 29822 17502 29874 17554
rect 31054 17502 31106 17554
rect 32062 17502 32114 17554
rect 33294 17502 33346 17554
rect 34526 17502 34578 17554
rect 35198 17502 35250 17554
rect 36318 17502 36370 17554
rect 37326 17502 37378 17554
rect 8094 17390 8146 17442
rect 14590 17390 14642 17442
rect 14702 17390 14754 17442
rect 25230 17390 25282 17442
rect 25566 17390 25618 17442
rect 26014 17390 26066 17442
rect 26126 17390 26178 17442
rect 27246 17390 27298 17442
rect 31390 17390 31442 17442
rect 31726 17390 31778 17442
rect 33182 17390 33234 17442
rect 33742 17390 33794 17442
rect 33966 17390 34018 17442
rect 34414 17390 34466 17442
rect 35310 17390 35362 17442
rect 37102 17390 37154 17442
rect 43150 17390 43202 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 9550 17054 9602 17106
rect 16494 17054 16546 17106
rect 20974 17054 21026 17106
rect 22094 17054 22146 17106
rect 22766 17054 22818 17106
rect 26350 17054 26402 17106
rect 28030 17054 28082 17106
rect 29710 17054 29762 17106
rect 30382 17054 30434 17106
rect 39678 17054 39730 17106
rect 16830 16942 16882 16994
rect 17502 16942 17554 16994
rect 18398 16942 18450 16994
rect 19182 16942 19234 16994
rect 19630 16942 19682 16994
rect 21310 16942 21362 16994
rect 22542 16942 22594 16994
rect 26574 16942 26626 16994
rect 27022 16942 27074 16994
rect 27806 16942 27858 16994
rect 28254 16942 28306 16994
rect 30046 16942 30098 16994
rect 31054 16942 31106 16994
rect 31390 16942 31442 16994
rect 32174 16942 32226 16994
rect 33854 16942 33906 16994
rect 37102 16942 37154 16994
rect 42030 16942 42082 16994
rect 9886 16830 9938 16882
rect 13134 16830 13186 16882
rect 16046 16830 16098 16882
rect 17838 16830 17890 16882
rect 18622 16830 18674 16882
rect 19294 16830 19346 16882
rect 21534 16830 21586 16882
rect 22206 16830 22258 16882
rect 22878 16830 22930 16882
rect 23326 16830 23378 16882
rect 23662 16830 23714 16882
rect 24110 16830 24162 16882
rect 24334 16830 24386 16882
rect 24446 16830 24498 16882
rect 25230 16830 25282 16882
rect 25454 16830 25506 16882
rect 25790 16830 25842 16882
rect 26014 16830 26066 16882
rect 26910 16830 26962 16882
rect 27134 16830 27186 16882
rect 27582 16830 27634 16882
rect 30718 16830 30770 16882
rect 31838 16830 31890 16882
rect 33070 16830 33122 16882
rect 36430 16830 36482 16882
rect 41918 16830 41970 16882
rect 12014 16718 12066 16770
rect 14926 16718 14978 16770
rect 22990 16718 23042 16770
rect 25342 16718 25394 16770
rect 35982 16718 36034 16770
rect 39230 16718 39282 16770
rect 22094 16606 22146 16658
rect 23998 16606 24050 16658
rect 26238 16606 26290 16658
rect 27918 16606 27970 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 11230 16270 11282 16322
rect 11566 16270 11618 16322
rect 14702 16270 14754 16322
rect 16270 16270 16322 16322
rect 8654 16158 8706 16210
rect 10782 16158 10834 16210
rect 12910 16158 12962 16210
rect 16718 16158 16770 16210
rect 22766 16158 22818 16210
rect 30718 16158 30770 16210
rect 38222 16158 38274 16210
rect 7982 16046 8034 16098
rect 15150 16046 15202 16098
rect 18958 16046 19010 16098
rect 19294 16046 19346 16098
rect 23886 16046 23938 16098
rect 24446 16046 24498 16098
rect 24558 16046 24610 16098
rect 24782 16046 24834 16098
rect 25006 16046 25058 16098
rect 29598 16046 29650 16098
rect 31838 16046 31890 16098
rect 34302 16046 34354 16098
rect 34526 16046 34578 16098
rect 34862 16046 34914 16098
rect 11902 15934 11954 15986
rect 12126 15934 12178 15986
rect 13918 15934 13970 15986
rect 14366 15934 14418 15986
rect 15486 15934 15538 15986
rect 15934 15934 15986 15986
rect 16158 15934 16210 15986
rect 13582 15822 13634 15874
rect 18734 15822 18786 15874
rect 19182 15822 19234 15874
rect 24558 15822 24610 15874
rect 25902 15822 25954 15874
rect 29934 15822 29986 15874
rect 32062 15822 32114 15874
rect 34638 15822 34690 15874
rect 36206 15822 36258 15874
rect 38110 15822 38162 15874
rect 43822 15822 43874 15874
rect 44270 15822 44322 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 16046 15486 16098 15538
rect 23326 15486 23378 15538
rect 24222 15486 24274 15538
rect 28478 15486 28530 15538
rect 36542 15486 36594 15538
rect 38782 15486 38834 15538
rect 6750 15374 6802 15426
rect 11902 15374 11954 15426
rect 13470 15374 13522 15426
rect 17614 15374 17666 15426
rect 18398 15374 18450 15426
rect 19294 15374 19346 15426
rect 20750 15374 20802 15426
rect 26126 15374 26178 15426
rect 26462 15374 26514 15426
rect 28030 15374 28082 15426
rect 29934 15374 29986 15426
rect 30158 15374 30210 15426
rect 37326 15374 37378 15426
rect 39678 15374 39730 15426
rect 6078 15262 6130 15314
rect 10558 15262 10610 15314
rect 12014 15262 12066 15314
rect 12798 15262 12850 15314
rect 18734 15262 18786 15314
rect 19630 15262 19682 15314
rect 20078 15262 20130 15314
rect 25230 15262 25282 15314
rect 25454 15262 25506 15314
rect 25790 15262 25842 15314
rect 28366 15262 28418 15314
rect 28814 15262 28866 15314
rect 29598 15262 29650 15314
rect 36542 15262 36594 15314
rect 36990 15262 37042 15314
rect 39454 15262 39506 15314
rect 40910 15262 40962 15314
rect 44270 15262 44322 15314
rect 8878 15150 8930 15202
rect 9662 15150 9714 15202
rect 11342 15150 11394 15202
rect 15598 15150 15650 15202
rect 17390 15150 17442 15202
rect 22878 15150 22930 15202
rect 25342 15150 25394 15202
rect 30046 15150 30098 15202
rect 38670 15150 38722 15202
rect 41694 15150 41746 15202
rect 43822 15150 43874 15202
rect 44942 15150 44994 15202
rect 47070 15150 47122 15202
rect 11006 15038 11058 15090
rect 17726 15038 17778 15090
rect 28590 15038 28642 15090
rect 29598 15038 29650 15090
rect 36094 15038 36146 15090
rect 36430 15038 36482 15090
rect 36878 15038 36930 15090
rect 39006 15038 39058 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 21422 14702 21474 14754
rect 21758 14702 21810 14754
rect 24334 14702 24386 14754
rect 35982 14702 36034 14754
rect 42478 14702 42530 14754
rect 11342 14590 11394 14642
rect 11790 14590 11842 14642
rect 18174 14590 18226 14642
rect 20302 14590 20354 14642
rect 20750 14590 20802 14642
rect 27022 14590 27074 14642
rect 28142 14590 28194 14642
rect 31950 14590 32002 14642
rect 37886 14590 37938 14642
rect 40014 14590 40066 14642
rect 8542 14478 8594 14530
rect 16606 14478 16658 14530
rect 17390 14478 17442 14530
rect 24110 14478 24162 14530
rect 24446 14478 24498 14530
rect 25454 14478 25506 14530
rect 25902 14478 25954 14530
rect 26686 14478 26738 14530
rect 27470 14478 27522 14530
rect 28366 14478 28418 14530
rect 29150 14478 29202 14530
rect 30158 14478 30210 14530
rect 31054 14478 31106 14530
rect 35310 14478 35362 14530
rect 35646 14478 35698 14530
rect 36094 14478 36146 14530
rect 40798 14478 40850 14530
rect 41470 14478 41522 14530
rect 43934 14478 43986 14530
rect 9214 14366 9266 14418
rect 16382 14366 16434 14418
rect 16942 14366 16994 14418
rect 21982 14366 22034 14418
rect 22318 14366 22370 14418
rect 23886 14366 23938 14418
rect 26126 14366 26178 14418
rect 26462 14366 26514 14418
rect 26910 14366 26962 14418
rect 27918 14366 27970 14418
rect 30270 14366 30322 14418
rect 31166 14366 31218 14418
rect 32398 14366 32450 14418
rect 33182 14366 33234 14418
rect 34862 14366 34914 14418
rect 35086 14366 35138 14418
rect 36430 14366 36482 14418
rect 41694 14366 41746 14418
rect 42142 14366 42194 14418
rect 42702 14366 42754 14418
rect 43262 14366 43314 14418
rect 44158 14366 44210 14418
rect 23998 14254 24050 14306
rect 25678 14254 25730 14306
rect 25790 14254 25842 14306
rect 27022 14254 27074 14306
rect 29038 14254 29090 14306
rect 31950 14254 32002 14306
rect 32174 14254 32226 14306
rect 32622 14254 32674 14306
rect 32734 14254 32786 14306
rect 32958 14254 33010 14306
rect 35198 14254 35250 14306
rect 35982 14254 36034 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 9550 13918 9602 13970
rect 19742 13918 19794 13970
rect 21310 13918 21362 13970
rect 23326 13918 23378 13970
rect 24110 13918 24162 13970
rect 26014 13918 26066 13970
rect 28814 13918 28866 13970
rect 32062 13918 32114 13970
rect 32174 13918 32226 13970
rect 34302 13918 34354 13970
rect 35310 13918 35362 13970
rect 36430 13918 36482 13970
rect 37662 13918 37714 13970
rect 38222 13918 38274 13970
rect 39902 13918 39954 13970
rect 41022 13918 41074 13970
rect 41918 13918 41970 13970
rect 44718 13918 44770 13970
rect 6414 13806 6466 13858
rect 8990 13806 9042 13858
rect 10222 13806 10274 13858
rect 10558 13806 10610 13858
rect 12014 13806 12066 13858
rect 13694 13806 13746 13858
rect 15486 13806 15538 13858
rect 16494 13806 16546 13858
rect 17614 13806 17666 13858
rect 20638 13806 20690 13858
rect 23886 13806 23938 13858
rect 25342 13806 25394 13858
rect 25566 13806 25618 13858
rect 27918 13806 27970 13858
rect 30270 13806 30322 13858
rect 30830 13806 30882 13858
rect 33294 13806 33346 13858
rect 33406 13806 33458 13858
rect 35870 13806 35922 13858
rect 36990 13806 37042 13858
rect 37214 13806 37266 13858
rect 38110 13806 38162 13858
rect 38446 13806 38498 13858
rect 38894 13806 38946 13858
rect 42590 13806 42642 13858
rect 42814 13806 42866 13858
rect 43598 13806 43650 13858
rect 5742 13694 5794 13746
rect 9886 13694 9938 13746
rect 11118 13694 11170 13746
rect 11454 13694 11506 13746
rect 12238 13694 12290 13746
rect 13582 13694 13634 13746
rect 15822 13694 15874 13746
rect 16606 13694 16658 13746
rect 17726 13694 17778 13746
rect 18622 13694 18674 13746
rect 20078 13694 20130 13746
rect 20862 13694 20914 13746
rect 22542 13694 22594 13746
rect 22766 13694 22818 13746
rect 22990 13694 23042 13746
rect 23326 13694 23378 13746
rect 23662 13694 23714 13746
rect 24446 13694 24498 13746
rect 26574 13694 26626 13746
rect 27470 13694 27522 13746
rect 28366 13694 28418 13746
rect 29262 13694 29314 13746
rect 29934 13694 29986 13746
rect 31054 13694 31106 13746
rect 31950 13694 32002 13746
rect 32510 13694 32562 13746
rect 33070 13694 33122 13746
rect 33854 13694 33906 13746
rect 34190 13694 34242 13746
rect 34414 13694 34466 13746
rect 34750 13694 34802 13746
rect 35422 13694 35474 13746
rect 36094 13694 36146 13746
rect 36542 13694 36594 13746
rect 38782 13694 38834 13746
rect 39566 13694 39618 13746
rect 42254 13694 42306 13746
rect 43822 13694 43874 13746
rect 44382 13694 44434 13746
rect 8542 13582 8594 13634
rect 19182 13582 19234 13634
rect 21758 13582 21810 13634
rect 27246 13582 27298 13634
rect 27806 13582 27858 13634
rect 33294 13582 33346 13634
rect 45278 13582 45330 13634
rect 14366 13470 14418 13522
rect 14702 13470 14754 13522
rect 16718 13470 16770 13522
rect 18286 13470 18338 13522
rect 24222 13470 24274 13522
rect 25678 13470 25730 13522
rect 35646 13470 35698 13522
rect 36766 13470 36818 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 18062 13134 18114 13186
rect 24558 13134 24610 13186
rect 26350 13134 26402 13186
rect 26686 13134 26738 13186
rect 42142 13134 42194 13186
rect 8990 13022 9042 13074
rect 11118 13022 11170 13074
rect 11566 13022 11618 13074
rect 15150 13022 15202 13074
rect 17278 13022 17330 13074
rect 25342 13022 25394 13074
rect 25790 13022 25842 13074
rect 29262 13022 29314 13074
rect 31390 13022 31442 13074
rect 33406 13022 33458 13074
rect 35534 13022 35586 13074
rect 37774 13022 37826 13074
rect 38222 13022 38274 13074
rect 47742 13022 47794 13074
rect 8318 12910 8370 12962
rect 14366 12910 14418 12962
rect 17726 12910 17778 12962
rect 18510 12910 18562 12962
rect 21534 12910 21586 12962
rect 23550 12910 23602 12962
rect 23998 12910 24050 12962
rect 24558 12910 24610 12962
rect 25902 12910 25954 12962
rect 29486 12910 29538 12962
rect 34862 12910 34914 12962
rect 34974 12910 35026 12962
rect 35758 12910 35810 12962
rect 35982 12910 36034 12962
rect 39342 12910 39394 12962
rect 42478 12910 42530 12962
rect 44046 12910 44098 12962
rect 44830 12910 44882 12962
rect 18734 12798 18786 12850
rect 23326 12798 23378 12850
rect 24222 12798 24274 12850
rect 25566 12798 25618 12850
rect 26574 12798 26626 12850
rect 27582 12798 27634 12850
rect 28254 12798 28306 12850
rect 28590 12798 28642 12850
rect 29150 12798 29202 12850
rect 30942 12798 30994 12850
rect 32174 12798 32226 12850
rect 32958 12798 33010 12850
rect 33182 12798 33234 12850
rect 34638 12798 34690 12850
rect 35422 12798 35474 12850
rect 39006 12798 39058 12850
rect 39118 12798 39170 12850
rect 39678 12798 39730 12850
rect 42702 12798 42754 12850
rect 43262 12798 43314 12850
rect 44270 12798 44322 12850
rect 45614 12798 45666 12850
rect 21310 12686 21362 12738
rect 22542 12686 22594 12738
rect 22990 12686 23042 12738
rect 24782 12686 24834 12738
rect 27246 12686 27298 12738
rect 27918 12686 27970 12738
rect 30606 12686 30658 12738
rect 31838 12686 31890 12738
rect 32622 12686 32674 12738
rect 32846 12686 32898 12738
rect 35086 12686 35138 12738
rect 38670 12686 38722 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 17502 12350 17554 12402
rect 23214 12350 23266 12402
rect 23998 12350 24050 12402
rect 25902 12350 25954 12402
rect 27470 12350 27522 12402
rect 27694 12350 27746 12402
rect 28814 12350 28866 12402
rect 31054 12350 31106 12402
rect 32062 12350 32114 12402
rect 34750 12350 34802 12402
rect 35534 12350 35586 12402
rect 36206 12350 36258 12402
rect 37998 12350 38050 12402
rect 38222 12350 38274 12402
rect 44942 12350 44994 12402
rect 15262 12238 15314 12290
rect 20638 12238 20690 12290
rect 24222 12238 24274 12290
rect 25230 12238 25282 12290
rect 30382 12238 30434 12290
rect 33854 12238 33906 12290
rect 34302 12238 34354 12290
rect 35198 12238 35250 12290
rect 35422 12238 35474 12290
rect 37326 12238 37378 12290
rect 39230 12238 39282 12290
rect 39678 12238 39730 12290
rect 42702 12238 42754 12290
rect 43150 12238 43202 12290
rect 43934 12238 43986 12290
rect 11006 12126 11058 12178
rect 14590 12126 14642 12178
rect 15374 12126 15426 12178
rect 19854 12126 19906 12178
rect 23438 12126 23490 12178
rect 23886 12126 23938 12178
rect 24446 12126 24498 12178
rect 25342 12126 25394 12178
rect 27246 12126 27298 12178
rect 28366 12126 28418 12178
rect 28478 12126 28530 12178
rect 28702 12126 28754 12178
rect 28926 12126 28978 12178
rect 29262 12126 29314 12178
rect 29486 12126 29538 12178
rect 30046 12126 30098 12178
rect 30606 12126 30658 12178
rect 31390 12126 31442 12178
rect 31726 12126 31778 12178
rect 33630 12126 33682 12178
rect 34638 12126 34690 12178
rect 34974 12126 35026 12178
rect 35870 12126 35922 12178
rect 35982 12126 36034 12178
rect 36430 12126 36482 12178
rect 36542 12126 36594 12178
rect 37886 12126 37938 12178
rect 43822 12126 43874 12178
rect 44606 12126 44658 12178
rect 11678 12014 11730 12066
rect 13806 12014 13858 12066
rect 22766 12014 22818 12066
rect 27358 12014 27410 12066
rect 29374 12014 29426 12066
rect 37214 12014 37266 12066
rect 14254 11902 14306 11954
rect 29822 11902 29874 11954
rect 37550 11902 37602 11954
rect 38558 11902 38610 11954
rect 38894 11902 38946 11954
rect 42142 11902 42194 11954
rect 42478 11902 42530 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 21422 11566 21474 11618
rect 21758 11566 21810 11618
rect 23102 11566 23154 11618
rect 14030 11454 14082 11506
rect 20190 11454 20242 11506
rect 20638 11454 20690 11506
rect 30270 11454 30322 11506
rect 31054 11454 31106 11506
rect 33854 11454 33906 11506
rect 35982 11454 36034 11506
rect 36430 11454 36482 11506
rect 37662 11454 37714 11506
rect 41022 11454 41074 11506
rect 44270 11454 44322 11506
rect 12462 11342 12514 11394
rect 15710 11342 15762 11394
rect 17278 11342 17330 11394
rect 22990 11342 23042 11394
rect 23886 11342 23938 11394
rect 24334 11342 24386 11394
rect 24446 11342 24498 11394
rect 24782 11342 24834 11394
rect 27470 11342 27522 11394
rect 27806 11342 27858 11394
rect 28142 11342 28194 11394
rect 30718 11342 30770 11394
rect 31838 11342 31890 11394
rect 33182 11342 33234 11394
rect 40574 11342 40626 11394
rect 41358 11342 41410 11394
rect 12126 11230 12178 11282
rect 18062 11230 18114 11282
rect 21982 11230 22034 11282
rect 22318 11230 22370 11282
rect 24222 11230 24274 11282
rect 25118 11230 25170 11282
rect 25454 11230 25506 11282
rect 39790 11230 39842 11282
rect 42142 11230 42194 11282
rect 16270 11118 16322 11170
rect 23102 11118 23154 11170
rect 23550 11118 23602 11170
rect 25902 11118 25954 11170
rect 27022 11118 27074 11170
rect 27694 11118 27746 11170
rect 31502 11118 31554 11170
rect 37326 11118 37378 11170
rect 44942 11118 44994 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 15038 10782 15090 10834
rect 18622 10782 18674 10834
rect 24222 10782 24274 10834
rect 26126 10782 26178 10834
rect 33406 10782 33458 10834
rect 33854 10782 33906 10834
rect 35870 10782 35922 10834
rect 38670 10782 38722 10834
rect 42030 10782 42082 10834
rect 14142 10670 14194 10722
rect 14478 10670 14530 10722
rect 20526 10670 20578 10722
rect 22318 10670 22370 10722
rect 25342 10670 25394 10722
rect 26574 10670 26626 10722
rect 27582 10670 27634 10722
rect 28814 10670 28866 10722
rect 31390 10670 31442 10722
rect 34974 10670 35026 10722
rect 36430 10670 36482 10722
rect 36878 10670 36930 10722
rect 40014 10670 40066 10722
rect 10446 10558 10498 10610
rect 17838 10558 17890 10610
rect 18958 10558 19010 10610
rect 19630 10558 19682 10610
rect 19966 10558 20018 10610
rect 20750 10558 20802 10610
rect 22094 10558 22146 10610
rect 23214 10558 23266 10610
rect 26462 10558 26514 10610
rect 27806 10558 27858 10610
rect 31166 10558 31218 10610
rect 34190 10558 34242 10610
rect 34750 10558 34802 10610
rect 36206 10558 36258 10610
rect 38446 10558 38498 10610
rect 39790 10558 39842 10610
rect 42254 10558 42306 10610
rect 11118 10446 11170 10498
rect 13246 10446 13298 10498
rect 14702 10446 14754 10498
rect 18286 10446 18338 10498
rect 22766 10446 22818 10498
rect 23550 10446 23602 10498
rect 25230 10446 25282 10498
rect 27022 10446 27074 10498
rect 25566 10334 25618 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 14366 9998 14418 10050
rect 25902 9998 25954 10050
rect 27358 9998 27410 10050
rect 29486 9998 29538 10050
rect 31950 9998 32002 10050
rect 33182 9998 33234 10050
rect 13582 9886 13634 9938
rect 17054 9886 17106 9938
rect 22430 9886 22482 9938
rect 23998 9886 24050 9938
rect 27694 9886 27746 9938
rect 31950 9886 32002 9938
rect 39454 9886 39506 9938
rect 41582 9886 41634 9938
rect 42814 9886 42866 9938
rect 14814 9774 14866 9826
rect 17502 9774 17554 9826
rect 18062 9774 18114 9826
rect 18734 9774 18786 9826
rect 19294 9774 19346 9826
rect 22094 9774 22146 9826
rect 22654 9774 22706 9826
rect 24334 9774 24386 9826
rect 32398 9774 32450 9826
rect 33406 9774 33458 9826
rect 33630 9774 33682 9826
rect 42254 9774 42306 9826
rect 11342 9662 11394 9714
rect 11678 9662 11730 9714
rect 14030 9662 14082 9714
rect 14926 9662 14978 9714
rect 17390 9662 17442 9714
rect 17950 9662 18002 9714
rect 19182 9662 19234 9714
rect 19742 9662 19794 9714
rect 22990 9662 23042 9714
rect 25118 9662 25170 9714
rect 25566 9662 25618 9714
rect 26126 9662 26178 9714
rect 26462 9662 26514 9714
rect 27918 9662 27970 9714
rect 28478 9662 28530 9714
rect 29150 9662 29202 9714
rect 38670 9662 38722 9714
rect 17166 9550 17218 9602
rect 17726 9550 17778 9602
rect 18398 9550 18450 9602
rect 18622 9550 18674 9602
rect 18958 9550 19010 9602
rect 20190 9550 20242 9602
rect 21646 9550 21698 9602
rect 24782 9550 24834 9602
rect 29374 9550 29426 9602
rect 32846 9550 32898 9602
rect 33966 9550 34018 9602
rect 35758 9550 35810 9602
rect 36206 9550 36258 9602
rect 37998 9550 38050 9602
rect 38334 9550 38386 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 16718 9214 16770 9266
rect 18622 9214 18674 9266
rect 21198 9214 21250 9266
rect 23662 9214 23714 9266
rect 34302 9214 34354 9266
rect 36430 9214 36482 9266
rect 36990 9214 37042 9266
rect 37998 9214 38050 9266
rect 40238 9214 40290 9266
rect 14926 9102 14978 9154
rect 15598 9102 15650 9154
rect 16046 9102 16098 9154
rect 17614 9102 17666 9154
rect 19630 9102 19682 9154
rect 21870 9102 21922 9154
rect 22654 9102 22706 9154
rect 22766 9102 22818 9154
rect 27134 9102 27186 9154
rect 33182 9102 33234 9154
rect 33294 9102 33346 9154
rect 33742 9102 33794 9154
rect 33854 9102 33906 9154
rect 35310 9102 35362 9154
rect 35870 9102 35922 9154
rect 36542 9102 36594 9154
rect 38446 9102 38498 9154
rect 38558 9102 38610 9154
rect 39342 9102 39394 9154
rect 10558 8990 10610 9042
rect 14254 8990 14306 9042
rect 15038 8990 15090 9042
rect 17950 8990 18002 9042
rect 19406 8990 19458 9042
rect 21534 8990 21586 9042
rect 22206 8990 22258 9042
rect 22430 8990 22482 9042
rect 26350 8990 26402 9042
rect 29710 8990 29762 9042
rect 33518 8990 33570 9042
rect 36206 8990 36258 9042
rect 37438 8990 37490 9042
rect 38782 8990 38834 9042
rect 39118 8990 39170 9042
rect 39902 8990 39954 9042
rect 11342 8878 11394 8930
rect 13470 8878 13522 8930
rect 19070 8878 19122 8930
rect 23214 8878 23266 8930
rect 26014 8878 26066 8930
rect 29262 8878 29314 8930
rect 30382 8878 30434 8930
rect 32510 8878 32562 8930
rect 13918 8766 13970 8818
rect 16382 8766 16434 8818
rect 18734 8766 18786 8818
rect 19070 8766 19122 8818
rect 20190 8766 20242 8818
rect 20526 8766 20578 8818
rect 33182 8766 33234 8818
rect 34750 8766 34802 8818
rect 35086 8766 35138 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 32286 8430 32338 8482
rect 15150 8318 15202 8370
rect 17390 8318 17442 8370
rect 19518 8318 19570 8370
rect 20638 8318 20690 8370
rect 23550 8318 23602 8370
rect 24670 8318 24722 8370
rect 26798 8318 26850 8370
rect 33742 8318 33794 8370
rect 34190 8318 34242 8370
rect 34526 8318 34578 8370
rect 37102 8318 37154 8370
rect 37438 8318 37490 8370
rect 11902 8206 11954 8258
rect 15934 8206 15986 8258
rect 16718 8206 16770 8258
rect 19966 8206 20018 8258
rect 23886 8206 23938 8258
rect 33070 8206 33122 8258
rect 34862 8206 34914 8258
rect 36094 8206 36146 8258
rect 39342 8206 39394 8258
rect 11566 8094 11618 8146
rect 15822 8094 15874 8146
rect 21982 8094 22034 8146
rect 30942 8094 30994 8146
rect 31278 8094 31330 8146
rect 31950 8094 32002 8146
rect 32846 8094 32898 8146
rect 37662 8094 37714 8146
rect 38222 8094 38274 8146
rect 39566 8094 39618 8146
rect 39902 8094 39954 8146
rect 13694 7982 13746 8034
rect 14814 7982 14866 8034
rect 20190 7982 20242 8034
rect 22318 7982 22370 8034
rect 22654 7982 22706 8034
rect 23102 7982 23154 8034
rect 35198 7982 35250 8034
rect 35758 7982 35810 8034
rect 39006 7982 39058 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 17838 7646 17890 7698
rect 24558 7646 24610 7698
rect 28814 7646 28866 7698
rect 33406 7646 33458 7698
rect 33742 7646 33794 7698
rect 37886 7646 37938 7698
rect 18846 7534 18898 7586
rect 20190 7534 20242 7586
rect 22654 7534 22706 7586
rect 23550 7534 23602 7586
rect 27806 7534 27858 7586
rect 28254 7534 28306 7586
rect 35310 7534 35362 7586
rect 38446 7534 38498 7586
rect 39118 7534 39170 7586
rect 39454 7534 39506 7586
rect 39790 7534 39842 7586
rect 12238 7422 12290 7474
rect 18174 7422 18226 7474
rect 18958 7422 19010 7474
rect 19406 7422 19458 7474
rect 22990 7422 23042 7474
rect 23438 7422 23490 7474
rect 29710 7422 29762 7474
rect 34638 7422 34690 7474
rect 38782 7422 38834 7474
rect 12910 7310 12962 7362
rect 15038 7310 15090 7362
rect 15486 7310 15538 7362
rect 22318 7310 22370 7362
rect 30382 7310 30434 7362
rect 32510 7310 32562 7362
rect 37438 7310 37490 7362
rect 24222 7198 24274 7250
rect 28478 7198 28530 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 15486 6862 15538 6914
rect 32398 6862 32450 6914
rect 23998 6750 24050 6802
rect 27246 6750 27298 6802
rect 38222 6750 38274 6802
rect 13806 6638 13858 6690
rect 16270 6638 16322 6690
rect 22542 6638 22594 6690
rect 24334 6638 24386 6690
rect 29374 6638 29426 6690
rect 33070 6638 33122 6690
rect 41134 6638 41186 6690
rect 41582 6638 41634 6690
rect 13470 6526 13522 6578
rect 16046 6526 16098 6578
rect 23214 6526 23266 6578
rect 25118 6526 25170 6578
rect 29934 6526 29986 6578
rect 30942 6526 30994 6578
rect 31278 6526 31330 6578
rect 32062 6526 32114 6578
rect 32958 6526 33010 6578
rect 40350 6526 40402 6578
rect 15150 6414 15202 6466
rect 29150 6414 29202 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 23886 6078 23938 6130
rect 25566 6078 25618 6130
rect 29262 6078 29314 6130
rect 18398 5966 18450 6018
rect 19070 5966 19122 6018
rect 20638 5966 20690 6018
rect 21982 5966 22034 6018
rect 22990 5966 23042 6018
rect 23326 5966 23378 6018
rect 27022 5966 27074 6018
rect 27582 5966 27634 6018
rect 28254 5966 28306 6018
rect 28702 5966 28754 6018
rect 30270 5966 30322 6018
rect 32174 5966 32226 6018
rect 33854 5966 33906 6018
rect 34302 5966 34354 6018
rect 35422 5966 35474 6018
rect 35982 5966 36034 6018
rect 13358 5854 13410 5906
rect 18286 5854 18338 5906
rect 19406 5854 19458 5906
rect 20414 5854 20466 5906
rect 22206 5854 22258 5906
rect 25902 5854 25954 5906
rect 26462 5854 26514 5906
rect 26798 5854 26850 5906
rect 30606 5854 30658 5906
rect 31278 5854 31330 5906
rect 31614 5854 31666 5906
rect 32398 5854 32450 5906
rect 33518 5854 33570 5906
rect 36206 5854 36258 5906
rect 14030 5742 14082 5794
rect 16158 5742 16210 5794
rect 16606 5742 16658 5794
rect 17838 5742 17890 5794
rect 21086 5742 21138 5794
rect 28926 5742 28978 5794
rect 17502 5630 17554 5682
rect 21422 5630 21474 5682
rect 23550 5630 23602 5682
rect 33182 5630 33234 5682
rect 36542 5630 36594 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 34974 5294 35026 5346
rect 18510 5182 18562 5234
rect 20638 5182 20690 5234
rect 22318 5182 22370 5234
rect 26014 5182 26066 5234
rect 31502 5182 31554 5234
rect 33630 5182 33682 5234
rect 34078 5182 34130 5234
rect 36990 5182 37042 5234
rect 40350 5182 40402 5234
rect 14478 5070 14530 5122
rect 17726 5070 17778 5122
rect 23214 5070 23266 5122
rect 27694 5070 27746 5122
rect 30158 5070 30210 5122
rect 30830 5070 30882 5122
rect 35758 5070 35810 5122
rect 39118 5070 39170 5122
rect 39902 5070 39954 5122
rect 14254 4958 14306 5010
rect 21758 4958 21810 5010
rect 22094 4958 22146 5010
rect 23886 4958 23938 5010
rect 27918 4958 27970 5010
rect 28366 4958 28418 5010
rect 30382 4958 30434 5010
rect 35534 4958 35586 5010
rect 22654 4846 22706 4898
rect 27358 4846 27410 4898
rect 34638 4846 34690 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 19630 4510 19682 4562
rect 23886 4510 23938 4562
rect 24334 4510 24386 4562
rect 25566 4510 25618 4562
rect 32510 4510 32562 4562
rect 37326 4510 37378 4562
rect 37774 4510 37826 4562
rect 14702 4398 14754 4450
rect 17390 4398 17442 4450
rect 18734 4398 18786 4450
rect 21086 4398 21138 4450
rect 23550 4398 23602 4450
rect 29934 4398 29986 4450
rect 36990 4398 37042 4450
rect 14030 4286 14082 4338
rect 17614 4286 17666 4338
rect 18510 4286 18562 4338
rect 19294 4286 19346 4338
rect 20414 4286 20466 4338
rect 26014 4286 26066 4338
rect 29262 4286 29314 4338
rect 36654 4286 36706 4338
rect 16830 4174 16882 4226
rect 23214 4174 23266 4226
rect 26686 4174 26738 4226
rect 28814 4174 28866 4226
rect 32062 4174 32114 4226
rect 33742 4174 33794 4226
rect 35870 4174 35922 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 17166 3614 17218 3666
rect 20974 3614 21026 3666
rect 22878 3614 22930 3666
rect 27358 3502 27410 3554
rect 34526 3502 34578 3554
rect 27022 3390 27074 3442
rect 34750 3390 34802 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 4032 59200 4144 60000
rect 4480 59200 4592 60000
rect 4928 59200 5040 60000
rect 5376 59200 5488 60000
rect 5824 59200 5936 60000
rect 6272 59200 6384 60000
rect 6720 59200 6832 60000
rect 7168 59200 7280 60000
rect 7616 59200 7728 60000
rect 8064 59200 8176 60000
rect 8512 59200 8624 60000
rect 8960 59200 9072 60000
rect 9408 59200 9520 60000
rect 9856 59200 9968 60000
rect 10304 59200 10416 60000
rect 10752 59200 10864 60000
rect 11200 59200 11312 60000
rect 11648 59200 11760 60000
rect 12096 59200 12208 60000
rect 12544 59200 12656 60000
rect 12992 59200 13104 60000
rect 13440 59200 13552 60000
rect 13888 59200 14000 60000
rect 14336 59200 14448 60000
rect 14784 59200 14896 60000
rect 15232 59200 15344 60000
rect 15680 59200 15792 60000
rect 16128 59200 16240 60000
rect 16576 59200 16688 60000
rect 17024 59200 17136 60000
rect 17472 59200 17584 60000
rect 17920 59200 18032 60000
rect 18368 59200 18480 60000
rect 18816 59200 18928 60000
rect 19264 59200 19376 60000
rect 19712 59200 19824 60000
rect 20160 59200 20272 60000
rect 20608 59200 20720 60000
rect 21056 59200 21168 60000
rect 21504 59200 21616 60000
rect 21952 59200 22064 60000
rect 22400 59200 22512 60000
rect 22848 59200 22960 60000
rect 23296 59200 23408 60000
rect 23744 59200 23856 60000
rect 24192 59200 24304 60000
rect 24640 59200 24752 60000
rect 25088 59200 25200 60000
rect 25536 59200 25648 60000
rect 25984 59200 26096 60000
rect 26432 59200 26544 60000
rect 26880 59200 26992 60000
rect 27328 59200 27440 60000
rect 27776 59200 27888 60000
rect 28224 59200 28336 60000
rect 28672 59200 28784 60000
rect 29120 59200 29232 60000
rect 29568 59200 29680 60000
rect 30016 59200 30128 60000
rect 30464 59200 30576 60000
rect 30912 59200 31024 60000
rect 31360 59200 31472 60000
rect 31808 59200 31920 60000
rect 32256 59200 32368 60000
rect 32704 59200 32816 60000
rect 33152 59200 33264 60000
rect 33600 59200 33712 60000
rect 34048 59200 34160 60000
rect 34496 59200 34608 60000
rect 34944 59200 35056 60000
rect 35392 59200 35504 60000
rect 35840 59200 35952 60000
rect 36288 59200 36400 60000
rect 36736 59200 36848 60000
rect 37184 59200 37296 60000
rect 37632 59200 37744 60000
rect 38080 59200 38192 60000
rect 38528 59200 38640 60000
rect 38976 59200 39088 60000
rect 39424 59200 39536 60000
rect 39872 59200 39984 60000
rect 40320 59200 40432 60000
rect 40768 59200 40880 60000
rect 41216 59200 41328 60000
rect 41664 59200 41776 60000
rect 42112 59200 42224 60000
rect 42560 59200 42672 60000
rect 43008 59200 43120 60000
rect 43456 59200 43568 60000
rect 43904 59200 44016 60000
rect 44352 59200 44464 60000
rect 44800 59200 44912 60000
rect 45248 59200 45360 60000
rect 45696 59200 45808 60000
rect 46144 59200 46256 60000
rect 46592 59200 46704 60000
rect 47040 59200 47152 60000
rect 47488 59200 47600 60000
rect 47936 59200 48048 60000
rect 48384 59200 48496 60000
rect 48832 59200 48944 60000
rect 49280 59200 49392 60000
rect 49728 59200 49840 60000
rect 50176 59200 50288 60000
rect 50624 59200 50736 60000
rect 51072 59200 51184 60000
rect 51520 59200 51632 60000
rect 51968 59200 52080 60000
rect 52416 59200 52528 60000
rect 52864 59200 52976 60000
rect 53312 59200 53424 60000
rect 53760 59200 53872 60000
rect 54208 59200 54320 60000
rect 54656 59200 54768 60000
rect 55104 59200 55216 60000
rect 55552 59200 55664 60000
rect 2156 55298 2212 55310
rect 2156 55246 2158 55298
rect 2210 55246 2212 55298
rect 1820 54516 1876 54526
rect 2156 54516 2212 55246
rect 2940 55188 2996 55198
rect 2940 55186 3108 55188
rect 2940 55134 2942 55186
rect 2994 55134 3108 55186
rect 2940 55132 3108 55134
rect 2940 55122 2996 55132
rect 1820 54514 2212 54516
rect 1820 54462 1822 54514
rect 1874 54462 2212 54514
rect 1820 54460 2212 54462
rect 1596 53844 1652 53854
rect 1596 29988 1652 53788
rect 1820 52162 1876 54460
rect 2492 54402 2548 54414
rect 2492 54350 2494 54402
rect 2546 54350 2548 54402
rect 2492 53842 2548 54350
rect 2492 53790 2494 53842
rect 2546 53790 2548 53842
rect 2492 53778 2548 53790
rect 2604 53620 2660 53630
rect 2940 53620 2996 53630
rect 2604 53618 2996 53620
rect 2604 53566 2606 53618
rect 2658 53566 2942 53618
rect 2994 53566 2996 53618
rect 2604 53564 2996 53566
rect 2604 53554 2660 53564
rect 2940 53554 2996 53564
rect 2380 53508 2436 53518
rect 1820 52110 1822 52162
rect 1874 52110 1876 52162
rect 1820 50594 1876 52110
rect 1820 50542 1822 50594
rect 1874 50542 1876 50594
rect 1820 48242 1876 50542
rect 2044 53452 2380 53508
rect 2044 50036 2100 53452
rect 2380 53414 2436 53452
rect 3052 52836 3108 55132
rect 3500 54292 3556 54302
rect 3164 53508 3220 53518
rect 3220 53452 3332 53508
rect 3164 53442 3220 53452
rect 3276 53170 3332 53452
rect 3276 53118 3278 53170
rect 3330 53118 3332 53170
rect 3276 53106 3332 53118
rect 3500 53058 3556 54236
rect 3500 53006 3502 53058
rect 3554 53006 3556 53058
rect 3500 52994 3556 53006
rect 3724 53842 3780 53854
rect 3724 53790 3726 53842
rect 3778 53790 3780 53842
rect 3164 52836 3220 52846
rect 3052 52834 3220 52836
rect 3052 52782 3166 52834
rect 3218 52782 3220 52834
rect 3052 52780 3220 52782
rect 3164 52770 3220 52780
rect 2492 52724 2548 52734
rect 2492 52274 2548 52668
rect 3724 52388 3780 53790
rect 4060 53844 4116 59200
rect 4508 56308 4564 59200
rect 5404 56868 5460 59200
rect 5852 57764 5908 59200
rect 5852 57708 6244 57764
rect 4956 56812 5460 56868
rect 4620 56308 4676 56318
rect 4508 56252 4620 56308
rect 4620 56214 4676 56252
rect 4956 55970 5012 56812
rect 5516 56308 5572 56318
rect 5516 56214 5572 56252
rect 6188 56306 6244 57708
rect 6188 56254 6190 56306
rect 6242 56254 6244 56306
rect 6188 56242 6244 56254
rect 5852 56196 5908 56206
rect 5852 56102 5908 56140
rect 4956 55918 4958 55970
rect 5010 55918 5012 55970
rect 4956 55906 5012 55918
rect 6748 55972 6804 59200
rect 7196 56308 7252 59200
rect 7420 56308 7476 56318
rect 7196 56306 7476 56308
rect 7196 56254 7422 56306
rect 7474 56254 7476 56306
rect 7196 56252 7476 56254
rect 7420 56242 7476 56252
rect 6972 55972 7028 55982
rect 6748 55970 7028 55972
rect 6748 55918 6974 55970
rect 7026 55918 7028 55970
rect 6748 55916 7028 55918
rect 8092 55972 8148 59200
rect 8540 56308 8596 59200
rect 8652 56308 8708 56318
rect 8540 56306 8708 56308
rect 8540 56254 8654 56306
rect 8706 56254 8708 56306
rect 8540 56252 8708 56254
rect 8652 56242 8708 56252
rect 9100 56196 9156 56206
rect 8204 55972 8260 55982
rect 8092 55970 8260 55972
rect 8092 55918 8206 55970
rect 8258 55918 8260 55970
rect 8092 55916 8260 55918
rect 6972 55906 7028 55916
rect 8204 55906 8260 55916
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 5068 55410 5124 55422
rect 5068 55358 5070 55410
rect 5122 55358 5124 55410
rect 5068 55076 5124 55358
rect 8764 55298 8820 55310
rect 8764 55246 8766 55298
rect 8818 55246 8820 55298
rect 5964 55076 6020 55086
rect 5068 55074 6020 55076
rect 5068 55022 5966 55074
rect 6018 55022 6020 55074
rect 5068 55020 6020 55022
rect 4620 54402 4676 54414
rect 4620 54350 4622 54402
rect 4674 54350 4676 54402
rect 4620 54292 4676 54350
rect 5516 54292 5572 54302
rect 4620 54236 4900 54292
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4060 53778 4116 53788
rect 3836 53732 3892 53742
rect 3836 53638 3892 53676
rect 4844 53732 4900 54236
rect 5516 54198 5572 54236
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 3724 52322 3780 52332
rect 2492 52222 2494 52274
rect 2546 52222 2548 52274
rect 2492 52210 2548 52222
rect 4620 52274 4676 52286
rect 4620 52222 4622 52274
rect 4674 52222 4676 52274
rect 4620 52164 4676 52222
rect 4620 51490 4676 52108
rect 4620 51438 4622 51490
rect 4674 51438 4676 51490
rect 4620 51426 4676 51438
rect 4844 52276 4900 53676
rect 5852 52946 5908 55020
rect 5964 55010 6020 55020
rect 6300 55074 6356 55086
rect 6300 55022 6302 55074
rect 6354 55022 6356 55074
rect 6300 54514 6356 55022
rect 7308 54740 7364 54750
rect 7308 54738 8148 54740
rect 7308 54686 7310 54738
rect 7362 54686 8148 54738
rect 7308 54684 8148 54686
rect 7308 54674 7364 54684
rect 6300 54462 6302 54514
rect 6354 54462 6356 54514
rect 6188 54402 6244 54414
rect 6188 54350 6190 54402
rect 6242 54350 6244 54402
rect 5964 53842 6020 53854
rect 5964 53790 5966 53842
rect 6018 53790 6020 53842
rect 5964 53060 6020 53790
rect 6076 53060 6132 53070
rect 5964 53004 6076 53060
rect 6076 52966 6132 53004
rect 6188 53058 6244 54350
rect 6188 53006 6190 53058
rect 6242 53006 6244 53058
rect 5852 52894 5854 52946
rect 5906 52894 5908 52946
rect 5852 52882 5908 52894
rect 5180 52836 5236 52846
rect 5180 52742 5236 52780
rect 6188 52836 6244 53006
rect 6300 52948 6356 54462
rect 6972 54292 7028 54302
rect 7196 54292 7252 54302
rect 6972 54198 7028 54236
rect 7084 54290 7252 54292
rect 7084 54238 7198 54290
rect 7250 54238 7252 54290
rect 7084 54236 7252 54238
rect 7084 53956 7140 54236
rect 7196 54226 7252 54236
rect 7308 54290 7364 54302
rect 7308 54238 7310 54290
rect 7362 54238 7364 54290
rect 6636 53900 7140 53956
rect 6636 53172 6692 53900
rect 6300 52882 6356 52892
rect 6524 53170 6692 53172
rect 6524 53118 6638 53170
rect 6690 53118 6692 53170
rect 6524 53116 6692 53118
rect 4844 51378 4900 52220
rect 5068 52722 5124 52734
rect 5068 52670 5070 52722
rect 5122 52670 5124 52722
rect 5068 51602 5124 52670
rect 5404 52722 5460 52734
rect 5404 52670 5406 52722
rect 5458 52670 5460 52722
rect 5068 51550 5070 51602
rect 5122 51550 5124 51602
rect 5068 51538 5124 51550
rect 5180 52388 5236 52398
rect 5180 51490 5236 52332
rect 5180 51438 5182 51490
rect 5234 51438 5236 51490
rect 5180 51426 5236 51438
rect 4844 51326 4846 51378
rect 4898 51326 4900 51378
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4620 50706 4676 50718
rect 4620 50654 4622 50706
rect 4674 50654 4676 50706
rect 2492 50484 2548 50494
rect 2044 49942 2100 49980
rect 2156 50482 2548 50484
rect 2156 50430 2494 50482
rect 2546 50430 2548 50482
rect 2156 50428 2548 50430
rect 2156 50034 2212 50428
rect 2492 50418 2548 50428
rect 2156 49982 2158 50034
rect 2210 49982 2212 50034
rect 2156 49970 2212 49982
rect 2716 50036 2772 50046
rect 2268 49812 2324 49822
rect 2604 49812 2660 49822
rect 2268 49810 2660 49812
rect 2268 49758 2270 49810
rect 2322 49758 2606 49810
rect 2658 49758 2660 49810
rect 2268 49756 2660 49758
rect 2268 49746 2324 49756
rect 2604 49746 2660 49756
rect 2716 49252 2772 49980
rect 3500 49812 3556 49822
rect 3500 49718 3556 49756
rect 4620 49812 4676 50654
rect 4620 49746 4676 49756
rect 4844 49810 4900 51326
rect 5404 51380 5460 52670
rect 5516 52724 5572 52734
rect 5516 52630 5572 52668
rect 5740 52388 5796 52398
rect 6188 52388 6244 52780
rect 6412 52388 6468 52398
rect 6188 52386 6468 52388
rect 6188 52334 6414 52386
rect 6466 52334 6468 52386
rect 6188 52332 6468 52334
rect 5628 52276 5684 52286
rect 5628 52162 5684 52220
rect 5628 52110 5630 52162
rect 5682 52110 5684 52162
rect 5628 52098 5684 52110
rect 5740 51940 5796 52332
rect 6412 52322 6468 52332
rect 5852 52164 5908 52174
rect 5852 52070 5908 52108
rect 5964 52050 6020 52062
rect 5964 51998 5966 52050
rect 6018 51998 6020 52050
rect 5964 51940 6020 51998
rect 5740 51884 6020 51940
rect 5404 51314 5460 51324
rect 5628 51378 5684 51390
rect 5628 51326 5630 51378
rect 5682 51326 5684 51378
rect 4956 49924 5012 49934
rect 4956 49922 5572 49924
rect 4956 49870 4958 49922
rect 5010 49870 5572 49922
rect 4956 49868 5572 49870
rect 4956 49858 5012 49868
rect 4844 49758 4846 49810
rect 4898 49758 4900 49810
rect 4844 49746 4900 49758
rect 2716 49158 2772 49196
rect 3388 49698 3444 49710
rect 3388 49646 3390 49698
rect 3442 49646 3444 49698
rect 2940 48916 2996 48926
rect 2940 48822 2996 48860
rect 3388 48916 3444 49646
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 3388 48850 3444 48860
rect 3500 49252 3556 49262
rect 3500 48914 3556 49196
rect 4732 49028 4788 49038
rect 4620 48972 4732 49028
rect 3500 48862 3502 48914
rect 3554 48862 3556 48914
rect 3500 48850 3556 48862
rect 4396 48916 4452 48926
rect 4396 48822 4452 48860
rect 2828 48802 2884 48814
rect 2828 48750 2830 48802
rect 2882 48750 2884 48802
rect 2828 48468 2884 48750
rect 2492 48412 2884 48468
rect 3836 48802 3892 48814
rect 3836 48750 3838 48802
rect 3890 48750 3892 48802
rect 3836 48468 3892 48750
rect 2492 48354 2548 48412
rect 3836 48402 3892 48412
rect 2492 48302 2494 48354
rect 2546 48302 2548 48354
rect 2492 48290 2548 48302
rect 1820 48190 1822 48242
rect 1874 48190 1876 48242
rect 1820 46676 1876 48190
rect 4620 48130 4676 48972
rect 4732 48934 4788 48972
rect 5516 48244 5572 49868
rect 5628 49140 5684 51326
rect 5740 51380 5796 51884
rect 5852 51380 5908 51390
rect 5740 51378 5908 51380
rect 5740 51326 5854 51378
rect 5906 51326 5908 51378
rect 5740 51324 5908 51326
rect 5740 50594 5796 50606
rect 5740 50542 5742 50594
rect 5794 50542 5796 50594
rect 5740 50484 5796 50542
rect 5740 50418 5796 50428
rect 5852 50148 5908 51324
rect 6076 51380 6132 51390
rect 6076 51286 6132 51324
rect 6188 51156 6244 51166
rect 6188 51154 6468 51156
rect 6188 51102 6190 51154
rect 6242 51102 6468 51154
rect 6188 51100 6468 51102
rect 6188 51090 6244 51100
rect 6412 50706 6468 51100
rect 6412 50654 6414 50706
rect 6466 50654 6468 50706
rect 6412 50642 6468 50654
rect 6524 50428 6580 53116
rect 6636 53106 6692 53116
rect 7196 53172 7252 53182
rect 7308 53172 7364 54238
rect 8092 53842 8148 54684
rect 8092 53790 8094 53842
rect 8146 53790 8148 53842
rect 8092 53778 8148 53790
rect 7196 53170 7364 53172
rect 7196 53118 7198 53170
rect 7250 53118 7364 53170
rect 7196 53116 7364 53118
rect 8764 53730 8820 55246
rect 8764 53678 8766 53730
rect 8818 53678 8820 53730
rect 7196 53106 7252 53116
rect 6972 53060 7028 53070
rect 6860 52946 6916 52958
rect 6860 52894 6862 52946
rect 6914 52894 6916 52946
rect 6860 52836 6916 52894
rect 6860 52770 6916 52780
rect 6972 52388 7028 53004
rect 7420 53060 7476 53070
rect 7308 52948 7364 52958
rect 6860 52386 7028 52388
rect 6860 52334 6974 52386
rect 7026 52334 7028 52386
rect 6860 52332 7028 52334
rect 6748 51492 6804 51502
rect 6860 51492 6916 52332
rect 6972 52322 7028 52332
rect 7084 52892 7308 52948
rect 7084 52386 7140 52892
rect 7308 52854 7364 52892
rect 7420 52946 7476 53004
rect 7420 52894 7422 52946
rect 7474 52894 7476 52946
rect 7420 52882 7476 52894
rect 7084 52334 7086 52386
rect 7138 52334 7140 52386
rect 6972 51604 7028 51614
rect 7084 51604 7140 52334
rect 7420 52388 7476 52398
rect 7420 52386 8036 52388
rect 7420 52334 7422 52386
rect 7474 52334 8036 52386
rect 7420 52332 8036 52334
rect 7420 52322 7476 52332
rect 7308 52164 7364 52174
rect 7756 52164 7812 52174
rect 6972 51602 7140 51604
rect 6972 51550 6974 51602
rect 7026 51550 7140 51602
rect 6972 51548 7140 51550
rect 7196 52162 7812 52164
rect 7196 52110 7310 52162
rect 7362 52110 7758 52162
rect 7810 52110 7812 52162
rect 7196 52108 7812 52110
rect 7196 51602 7252 52108
rect 7308 52098 7364 52108
rect 7756 52098 7812 52108
rect 7868 52164 7924 52174
rect 7868 52070 7924 52108
rect 7196 51550 7198 51602
rect 7250 51550 7252 51602
rect 6972 51538 7028 51548
rect 7196 51538 7252 51550
rect 6748 51490 6916 51492
rect 6748 51438 6750 51490
rect 6802 51438 6916 51490
rect 6748 51436 6916 51438
rect 6748 51426 6804 51436
rect 6972 51156 7028 51166
rect 5852 50082 5908 50092
rect 6076 50372 6580 50428
rect 6860 50484 6916 50494
rect 6972 50484 7028 51100
rect 6916 50428 7028 50484
rect 7308 51154 7364 51166
rect 7308 51102 7310 51154
rect 7362 51102 7364 51154
rect 5852 49810 5908 49822
rect 5852 49758 5854 49810
rect 5906 49758 5908 49810
rect 5740 49140 5796 49150
rect 5628 49138 5796 49140
rect 5628 49086 5742 49138
rect 5794 49086 5796 49138
rect 5628 49084 5796 49086
rect 5740 49074 5796 49084
rect 5628 48916 5684 48926
rect 5852 48916 5908 49758
rect 5964 49812 6020 49822
rect 5964 49026 6020 49756
rect 5964 48974 5966 49026
rect 6018 48974 6020 49026
rect 5964 48962 6020 48974
rect 5684 48860 5908 48916
rect 5628 48822 5684 48860
rect 5628 48244 5684 48254
rect 4620 48078 4622 48130
rect 4674 48078 4676 48130
rect 4620 48066 4676 48078
rect 4844 48242 5684 48244
rect 4844 48190 5630 48242
rect 5682 48190 5684 48242
rect 4844 48188 5684 48190
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4844 47346 4900 48188
rect 5628 48178 5684 48188
rect 5852 48244 5908 48254
rect 6076 48244 6132 50372
rect 6300 50036 6356 50046
rect 6300 49942 6356 49980
rect 6412 49922 6468 49934
rect 6412 49870 6414 49922
rect 6466 49870 6468 49922
rect 6412 49812 6468 49870
rect 6412 49746 6468 49756
rect 6188 49700 6244 49710
rect 6188 49026 6244 49644
rect 6188 48974 6190 49026
rect 6242 48974 6244 49026
rect 6188 48962 6244 48974
rect 5852 48242 6132 48244
rect 5852 48190 5854 48242
rect 5906 48190 6132 48242
rect 5852 48188 6132 48190
rect 6636 48354 6692 48366
rect 6636 48302 6638 48354
rect 6690 48302 6692 48354
rect 5852 47796 5908 48188
rect 6188 48020 6244 48030
rect 5068 47740 5908 47796
rect 6076 48018 6244 48020
rect 6076 47966 6190 48018
rect 6242 47966 6244 48018
rect 6076 47964 6244 47966
rect 5068 47682 5124 47740
rect 5068 47630 5070 47682
rect 5122 47630 5124 47682
rect 5068 47618 5124 47630
rect 5740 47572 5796 47582
rect 4956 47460 5012 47470
rect 4956 47366 5012 47404
rect 4844 47294 4846 47346
rect 4898 47294 4900 47346
rect 4844 47236 4900 47294
rect 5628 47348 5684 47358
rect 5628 47254 5684 47292
rect 4844 47180 5124 47236
rect 2940 47124 2996 47134
rect 2940 46786 2996 47068
rect 2940 46734 2942 46786
rect 2994 46734 2996 46786
rect 2940 46722 2996 46734
rect 2268 46676 2324 46686
rect 1820 46674 2324 46676
rect 1820 46622 2270 46674
rect 2322 46622 2324 46674
rect 1820 46620 2324 46622
rect 2268 46004 2324 46620
rect 4844 46676 4900 46686
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 2268 45938 2324 45948
rect 4396 46004 4452 46014
rect 4396 45106 4452 45948
rect 4844 45778 4900 46620
rect 5068 46562 5124 47180
rect 5516 46676 5572 46686
rect 5740 46676 5796 47516
rect 5964 47460 6020 47470
rect 5964 47366 6020 47404
rect 6076 47458 6132 47964
rect 6188 47954 6244 47964
rect 6636 47572 6692 48302
rect 6636 47506 6692 47516
rect 6076 47406 6078 47458
rect 6130 47406 6132 47458
rect 5516 46674 5796 46676
rect 5516 46622 5518 46674
rect 5570 46622 5796 46674
rect 5516 46620 5796 46622
rect 5964 46788 6020 46798
rect 5964 46674 6020 46732
rect 5964 46622 5966 46674
rect 6018 46622 6020 46674
rect 5516 46610 5572 46620
rect 5964 46610 6020 46622
rect 5068 46510 5070 46562
rect 5122 46510 5124 46562
rect 5068 46498 5124 46510
rect 4956 46452 5012 46462
rect 5404 46452 5460 46462
rect 4956 46002 5012 46396
rect 5180 46450 5460 46452
rect 5180 46398 5406 46450
rect 5458 46398 5460 46450
rect 5180 46396 5460 46398
rect 5068 46116 5124 46126
rect 5068 46022 5124 46060
rect 4956 45950 4958 46002
rect 5010 45950 5012 46002
rect 4956 45938 5012 45950
rect 4844 45726 4846 45778
rect 4898 45726 4900 45778
rect 4844 45714 4900 45726
rect 5068 45220 5124 45230
rect 5180 45220 5236 46396
rect 5404 46386 5460 46396
rect 5740 46452 5796 46462
rect 5740 46358 5796 46396
rect 6076 46116 6132 47406
rect 6860 47460 6916 50428
rect 6972 49812 7028 49822
rect 6972 49718 7028 49756
rect 7084 49810 7140 49822
rect 7084 49758 7086 49810
rect 7138 49758 7140 49810
rect 7084 49028 7140 49758
rect 7196 49812 7252 49822
rect 7196 49718 7252 49756
rect 7084 48962 7140 48972
rect 6972 48468 7028 48478
rect 6972 47908 7028 48412
rect 6972 47842 7028 47852
rect 6972 47460 7028 47470
rect 6860 47458 7028 47460
rect 6860 47406 6974 47458
rect 7026 47406 7028 47458
rect 6860 47404 7028 47406
rect 6860 46788 6916 46798
rect 6860 46694 6916 46732
rect 6300 46676 6356 46686
rect 6300 46582 6356 46620
rect 6524 46450 6580 46462
rect 6524 46398 6526 46450
rect 6578 46398 6580 46450
rect 6076 46050 6132 46060
rect 6412 46116 6468 46126
rect 6524 46116 6580 46398
rect 6468 46060 6580 46116
rect 6412 46050 6468 46060
rect 6972 46004 7028 47404
rect 7308 46786 7364 51102
rect 7644 50148 7700 50158
rect 7644 50034 7700 50092
rect 7644 49982 7646 50034
rect 7698 49982 7700 50034
rect 7644 49970 7700 49982
rect 7980 48354 8036 52332
rect 8428 52164 8484 52174
rect 8764 52164 8820 53678
rect 8428 52162 8820 52164
rect 8428 52110 8430 52162
rect 8482 52110 8820 52162
rect 8428 52108 8820 52110
rect 8876 54292 8932 54302
rect 8428 51156 8484 52108
rect 8876 51380 8932 54236
rect 8876 51314 8932 51324
rect 8428 51090 8484 51100
rect 8652 50372 8708 50382
rect 8204 50370 8708 50372
rect 8204 50318 8654 50370
rect 8706 50318 8708 50370
rect 8204 50316 8708 50318
rect 8204 49812 8260 50316
rect 8652 50306 8708 50316
rect 7980 48302 7982 48354
rect 8034 48302 8036 48354
rect 7980 48290 8036 48302
rect 8092 48354 8148 48366
rect 8092 48302 8094 48354
rect 8146 48302 8148 48354
rect 7756 48020 7812 48030
rect 7756 47570 7812 47964
rect 7756 47518 7758 47570
rect 7810 47518 7812 47570
rect 7756 47506 7812 47518
rect 8092 47012 8148 48302
rect 7308 46734 7310 46786
rect 7362 46734 7364 46786
rect 7308 46722 7364 46734
rect 7644 46956 8148 47012
rect 6972 45910 7028 45948
rect 7196 46676 7252 46686
rect 5068 45218 5236 45220
rect 5068 45166 5070 45218
rect 5122 45166 5236 45218
rect 5068 45164 5236 45166
rect 6972 45444 7028 45454
rect 5068 45154 5124 45164
rect 4396 45054 4398 45106
rect 4450 45054 4452 45106
rect 4396 45042 4452 45054
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 6972 43538 7028 45388
rect 7196 44994 7252 46620
rect 7644 46676 7700 46956
rect 7644 46610 7700 46620
rect 8092 46562 8148 46574
rect 8092 46510 8094 46562
rect 8146 46510 8148 46562
rect 7644 46450 7700 46462
rect 7644 46398 7646 46450
rect 7698 46398 7700 46450
rect 7644 45332 7700 46398
rect 8092 45444 8148 46510
rect 8092 45378 8148 45388
rect 8204 45332 8260 49756
rect 8988 49028 9044 49038
rect 8764 48354 8820 48366
rect 8764 48302 8766 48354
rect 8818 48302 8820 48354
rect 8316 48242 8372 48254
rect 8316 48190 8318 48242
rect 8370 48190 8372 48242
rect 8316 45668 8372 48190
rect 8764 47012 8820 48302
rect 8876 48132 8932 48142
rect 8876 48038 8932 48076
rect 8988 48018 9044 48972
rect 8988 47966 8990 48018
rect 9042 47966 9044 48018
rect 8988 47954 9044 47966
rect 8764 46946 8820 46956
rect 8988 47460 9044 47470
rect 8988 46898 9044 47404
rect 8988 46846 8990 46898
rect 9042 46846 9044 46898
rect 8988 46834 9044 46846
rect 8652 46788 8708 46798
rect 8428 46676 8484 46686
rect 8428 46582 8484 46620
rect 8652 46674 8708 46732
rect 8652 46622 8654 46674
rect 8706 46622 8708 46674
rect 8652 46610 8708 46622
rect 8764 45890 8820 45902
rect 8764 45838 8766 45890
rect 8818 45838 8820 45890
rect 8316 45612 8596 45668
rect 8204 45276 8484 45332
rect 7644 45266 7700 45276
rect 8092 45220 8148 45230
rect 8092 45106 8148 45164
rect 8092 45054 8094 45106
rect 8146 45054 8148 45106
rect 8092 45042 8148 45054
rect 8428 45106 8484 45276
rect 8428 45054 8430 45106
rect 8482 45054 8484 45106
rect 7196 44942 7198 44994
rect 7250 44942 7252 44994
rect 7196 44930 7252 44942
rect 7420 44436 7476 44446
rect 7420 44342 7476 44380
rect 7980 44436 8036 44446
rect 7308 44324 7364 44334
rect 7308 44230 7364 44268
rect 7868 44322 7924 44334
rect 7868 44270 7870 44322
rect 7922 44270 7924 44322
rect 7196 44212 7252 44222
rect 7196 44118 7252 44156
rect 7868 43988 7924 44270
rect 7868 43922 7924 43932
rect 6972 43486 6974 43538
rect 7026 43486 7028 43538
rect 6972 43474 7028 43486
rect 7644 43764 7700 43774
rect 7532 43426 7588 43438
rect 7532 43374 7534 43426
rect 7586 43374 7588 43426
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 6748 42756 6804 42766
rect 6076 41972 6132 41982
rect 6748 41972 6804 42700
rect 7532 42756 7588 43374
rect 7532 42690 7588 42700
rect 6076 41970 6804 41972
rect 6076 41918 6078 41970
rect 6130 41918 6804 41970
rect 6076 41916 6804 41918
rect 7420 42642 7476 42654
rect 7420 42590 7422 42642
rect 7474 42590 7476 42642
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 5068 40964 5124 40974
rect 1820 40404 1876 40414
rect 1820 39618 1876 40348
rect 4060 40404 4116 40414
rect 4060 40310 4116 40348
rect 4844 40402 4900 40414
rect 4844 40350 4846 40402
rect 4898 40350 4900 40402
rect 3276 40292 3332 40302
rect 3276 40198 3332 40236
rect 2940 40180 2996 40190
rect 2492 40178 2996 40180
rect 2492 40126 2942 40178
rect 2994 40126 2996 40178
rect 2492 40124 2996 40126
rect 2492 39730 2548 40124
rect 2940 40114 2996 40124
rect 3052 40180 3108 40190
rect 3052 40086 3108 40124
rect 3388 40180 3444 40190
rect 3948 40180 4004 40190
rect 3388 40178 3556 40180
rect 3388 40126 3390 40178
rect 3442 40126 3556 40178
rect 3388 40124 3556 40126
rect 3388 40114 3444 40124
rect 2492 39678 2494 39730
rect 2546 39678 2548 39730
rect 2492 39666 2548 39678
rect 1820 39566 1822 39618
rect 1874 39566 1876 39618
rect 1820 36482 1876 39566
rect 3500 39058 3556 40124
rect 3500 39006 3502 39058
rect 3554 39006 3556 39058
rect 3500 38994 3556 39006
rect 3612 39284 3668 39294
rect 2940 38948 2996 38958
rect 2940 38854 2996 38892
rect 2716 38834 2772 38846
rect 2716 38782 2718 38834
rect 2770 38782 2772 38834
rect 2716 37940 2772 38782
rect 3052 38836 3108 38846
rect 3052 38742 3108 38780
rect 3388 38836 3444 38846
rect 3388 38668 3444 38780
rect 3388 38612 3556 38668
rect 2380 37492 2436 37502
rect 2380 37398 2436 37436
rect 2716 37378 2772 37884
rect 2716 37326 2718 37378
rect 2770 37326 2772 37378
rect 1820 36430 1822 36482
rect 1874 36430 1876 36482
rect 1820 35028 1876 36430
rect 2156 37266 2212 37278
rect 2156 37214 2158 37266
rect 2210 37214 2212 37266
rect 2156 36036 2212 37214
rect 2492 37044 2548 37054
rect 2492 36594 2548 36988
rect 2492 36542 2494 36594
rect 2546 36542 2548 36594
rect 2492 36530 2548 36542
rect 2156 35970 2212 35980
rect 2716 35698 2772 37326
rect 3500 37938 3556 38612
rect 3500 37886 3502 37938
rect 3554 37886 3556 37938
rect 3500 37492 3556 37886
rect 3612 37604 3668 39228
rect 3948 39058 4004 40124
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4844 39732 4900 40350
rect 5068 40404 5124 40908
rect 6076 40964 6132 41916
rect 6860 41860 6916 41870
rect 6860 41766 6916 41804
rect 6076 40898 6132 40908
rect 5068 40338 5124 40348
rect 7308 40402 7364 40414
rect 7308 40350 7310 40402
rect 7362 40350 7364 40402
rect 6972 40292 7028 40302
rect 7308 40292 7364 40350
rect 7420 40404 7476 42590
rect 7644 40740 7700 43708
rect 7868 40852 7924 40862
rect 7420 40338 7476 40348
rect 7532 40684 7700 40740
rect 7756 40796 7868 40852
rect 6972 40290 7364 40292
rect 6972 40238 6974 40290
rect 7026 40238 7364 40290
rect 6972 40236 7364 40238
rect 4844 39666 4900 39676
rect 5740 39732 5796 39742
rect 5740 39638 5796 39676
rect 6076 39620 6132 39630
rect 6076 39526 6132 39564
rect 6412 39618 6468 39630
rect 6412 39566 6414 39618
rect 6466 39566 6468 39618
rect 3948 39006 3950 39058
rect 4002 39006 4004 39058
rect 3948 38994 4004 39006
rect 4060 39508 4116 39518
rect 3836 38948 3892 38958
rect 3724 38836 3780 38846
rect 3724 38742 3780 38780
rect 3836 38668 3892 38892
rect 3724 38612 3892 38668
rect 3724 37828 3780 38612
rect 4060 38274 4116 39452
rect 5628 39508 5684 39518
rect 5852 39508 5908 39518
rect 5628 39414 5684 39452
rect 5740 39506 5908 39508
rect 5740 39454 5854 39506
rect 5906 39454 5908 39506
rect 5740 39452 5908 39454
rect 4732 39396 4788 39406
rect 4620 39394 4788 39396
rect 4620 39342 4734 39394
rect 4786 39342 4788 39394
rect 4620 39340 4788 39342
rect 4284 38948 4340 38958
rect 4060 38222 4062 38274
rect 4114 38222 4116 38274
rect 4060 38210 4116 38222
rect 4172 38834 4228 38846
rect 4172 38782 4174 38834
rect 4226 38782 4228 38834
rect 3948 37940 4004 37950
rect 4172 37940 4228 38782
rect 4284 38834 4340 38892
rect 4284 38782 4286 38834
rect 4338 38782 4340 38834
rect 4284 38770 4340 38782
rect 4620 38612 4676 39340
rect 4732 39330 4788 39340
rect 5740 39060 5796 39452
rect 5852 39442 5908 39452
rect 6412 39284 6468 39566
rect 6412 39218 6468 39228
rect 5292 39004 5796 39060
rect 5180 38948 5236 38958
rect 4732 38836 4788 38874
rect 4732 38770 4788 38780
rect 5180 38834 5236 38892
rect 5180 38782 5182 38834
rect 5234 38782 5236 38834
rect 5180 38770 5236 38782
rect 4844 38722 4900 38734
rect 4844 38670 4846 38722
rect 4898 38670 4900 38722
rect 4844 38668 4900 38670
rect 4844 38612 5012 38668
rect 5292 38612 5348 39004
rect 6076 38834 6132 38846
rect 6076 38782 6078 38834
rect 6130 38782 6132 38834
rect 4956 38556 5348 38612
rect 4620 38546 4676 38556
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4844 38388 4900 38398
rect 4004 37884 4228 37940
rect 4844 38050 4900 38332
rect 4844 37998 4846 38050
rect 4898 37998 4900 38050
rect 3948 37846 4004 37884
rect 3724 37734 3780 37772
rect 4508 37826 4564 37838
rect 4508 37774 4510 37826
rect 4562 37774 4564 37826
rect 3612 37548 3892 37604
rect 3052 37266 3108 37278
rect 3052 37214 3054 37266
rect 3106 37214 3108 37266
rect 3052 37156 3108 37214
rect 3500 37266 3556 37436
rect 3724 37268 3780 37278
rect 3500 37214 3502 37266
rect 3554 37214 3556 37266
rect 3500 37202 3556 37214
rect 3612 37212 3724 37268
rect 3052 37090 3108 37100
rect 3612 37154 3668 37212
rect 3724 37202 3780 37212
rect 3612 37102 3614 37154
rect 3666 37102 3668 37154
rect 3612 37090 3668 37102
rect 3836 37042 3892 37548
rect 4508 37378 4564 37774
rect 4508 37326 4510 37378
rect 4562 37326 4564 37378
rect 3836 36990 3838 37042
rect 3890 36990 3892 37042
rect 3836 36978 3892 36990
rect 3948 37044 4004 37054
rect 4508 37044 4564 37326
rect 4620 37268 4676 37278
rect 4844 37268 4900 37998
rect 5068 37828 5124 37838
rect 5068 37734 5124 37772
rect 5292 37378 5348 38556
rect 5404 38612 5460 38622
rect 5404 38518 5460 38556
rect 5740 38612 5796 38622
rect 5740 38518 5796 38556
rect 5292 37326 5294 37378
rect 5346 37326 5348 37378
rect 5292 37314 5348 37326
rect 5852 38050 5908 38062
rect 5852 37998 5854 38050
rect 5906 37998 5908 38050
rect 5180 37268 5236 37278
rect 4844 37212 5180 37268
rect 4620 37174 4676 37212
rect 5180 37174 5236 37212
rect 5852 37268 5908 37998
rect 5852 37202 5908 37212
rect 6076 37156 6132 38782
rect 6300 38834 6356 38846
rect 6300 38782 6302 38834
rect 6354 38782 6356 38834
rect 6300 38612 6356 38782
rect 3948 36950 4004 36988
rect 4284 36988 4564 37044
rect 4732 37044 4788 37054
rect 5068 37044 5124 37054
rect 4732 37042 4900 37044
rect 4732 36990 4734 37042
rect 4786 36990 4900 37042
rect 4732 36988 4900 36990
rect 2716 35646 2718 35698
rect 2770 35646 2772 35698
rect 2716 35634 2772 35646
rect 3052 36036 3108 36046
rect 3052 35698 3108 35980
rect 3052 35646 3054 35698
rect 3106 35646 3108 35698
rect 3052 35634 3108 35646
rect 3948 35588 4004 35598
rect 3948 35494 4004 35532
rect 4284 35588 4340 36988
rect 4732 36978 4788 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4620 36594 4676 36606
rect 4620 36542 4622 36594
rect 4674 36542 4676 36594
rect 4620 36372 4676 36542
rect 4844 36484 4900 36988
rect 5068 36706 5124 36988
rect 5068 36654 5070 36706
rect 5122 36654 5124 36706
rect 5068 36642 5124 36654
rect 5292 36708 5348 36718
rect 4396 35700 4452 35710
rect 4620 35700 4676 36316
rect 4732 36428 4900 36484
rect 4732 35924 4788 36428
rect 4956 36372 5012 36382
rect 4956 36278 5012 36316
rect 5292 36036 5348 36652
rect 4732 35868 5012 35924
rect 4732 35700 4788 35710
rect 4396 35698 4788 35700
rect 4396 35646 4398 35698
rect 4450 35646 4734 35698
rect 4786 35646 4788 35698
rect 4396 35644 4788 35646
rect 4396 35634 4452 35644
rect 4732 35634 4788 35644
rect 4956 35700 5012 35868
rect 5292 35922 5348 35980
rect 5292 35870 5294 35922
rect 5346 35870 5348 35922
rect 5292 35858 5348 35870
rect 5740 36484 5796 36494
rect 4956 35698 5460 35700
rect 4956 35646 4958 35698
rect 5010 35646 5460 35698
rect 4956 35644 5460 35646
rect 4956 35634 5012 35644
rect 4284 35522 4340 35532
rect 3164 35474 3220 35486
rect 3164 35422 3166 35474
rect 3218 35422 3220 35474
rect 3164 35138 3220 35422
rect 5404 35476 5460 35644
rect 5740 35586 5796 36428
rect 6076 36484 6132 37100
rect 6076 36418 6132 36428
rect 6188 37380 6244 37390
rect 6188 37044 6244 37324
rect 6300 37156 6356 38556
rect 6300 37090 6356 37100
rect 6412 38834 6468 38846
rect 6412 38782 6414 38834
rect 6466 38782 6468 38834
rect 6188 36482 6244 36988
rect 6412 36708 6468 38782
rect 6860 38722 6916 38734
rect 6860 38670 6862 38722
rect 6914 38670 6916 38722
rect 6860 38612 6916 38670
rect 6860 38546 6916 38556
rect 6860 37940 6916 37950
rect 6972 37940 7028 40236
rect 6860 37938 7028 37940
rect 6860 37886 6862 37938
rect 6914 37886 7028 37938
rect 6860 37884 7028 37886
rect 7084 39732 7140 39742
rect 7084 39506 7140 39676
rect 7084 39454 7086 39506
rect 7138 39454 7140 39506
rect 6860 37874 6916 37884
rect 6412 36642 6468 36652
rect 6188 36430 6190 36482
rect 6242 36430 6244 36482
rect 6188 36418 6244 36430
rect 5740 35534 5742 35586
rect 5794 35534 5796 35586
rect 5740 35522 5796 35534
rect 5964 36370 6020 36382
rect 5964 36318 5966 36370
rect 6018 36318 6020 36370
rect 5964 36260 6020 36318
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 3164 35086 3166 35138
rect 3218 35086 3220 35138
rect 3164 35074 3220 35086
rect 4620 35140 4676 35150
rect 2828 35028 2884 35038
rect 1820 34130 1876 34972
rect 2492 35026 2884 35028
rect 2492 34974 2830 35026
rect 2882 34974 2884 35026
rect 2492 34972 2884 34974
rect 2492 34242 2548 34972
rect 2828 34962 2884 34972
rect 3276 35028 3332 35038
rect 2492 34190 2494 34242
rect 2546 34190 2548 34242
rect 2492 34178 2548 34190
rect 2940 34690 2996 34702
rect 2940 34638 2942 34690
rect 2994 34638 2996 34690
rect 1820 34078 1822 34130
rect 1874 34078 1876 34130
rect 1820 34066 1876 34078
rect 2940 33908 2996 34638
rect 2940 33842 2996 33852
rect 3276 32562 3332 34972
rect 4620 34018 4676 35084
rect 4620 33966 4622 34018
rect 4674 33966 4676 34018
rect 4620 33954 4676 33966
rect 4844 35028 4900 35038
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4732 33572 4788 33582
rect 3948 33570 4788 33572
rect 3948 33518 4734 33570
rect 4786 33518 4788 33570
rect 3948 33516 4788 33518
rect 3948 32674 4004 33516
rect 4732 33506 4788 33516
rect 4844 33458 4900 34972
rect 5292 34692 5348 34702
rect 5068 34580 5124 34590
rect 5068 34130 5124 34524
rect 5068 34078 5070 34130
rect 5122 34078 5124 34130
rect 4956 33906 5012 33918
rect 4956 33854 4958 33906
rect 5010 33854 5012 33906
rect 4956 33570 5012 33854
rect 5068 33908 5124 34078
rect 5292 34130 5348 34636
rect 5292 34078 5294 34130
rect 5346 34078 5348 34130
rect 5292 34066 5348 34078
rect 5404 34130 5460 35420
rect 5964 34916 6020 36204
rect 6412 36370 6468 36382
rect 6412 36318 6414 36370
rect 6466 36318 6468 36370
rect 6076 35700 6132 35710
rect 6412 35700 6468 36318
rect 6076 35698 6468 35700
rect 6076 35646 6078 35698
rect 6130 35646 6468 35698
rect 6076 35644 6468 35646
rect 6748 36258 6804 36270
rect 6748 36206 6750 36258
rect 6802 36206 6804 36258
rect 6748 35700 6804 36206
rect 6076 35364 6132 35644
rect 6748 35634 6804 35644
rect 6076 35298 6132 35308
rect 6076 34916 6132 34926
rect 5964 34860 6076 34916
rect 5404 34078 5406 34130
rect 5458 34078 5460 34130
rect 5404 34066 5460 34078
rect 5964 34132 6020 34142
rect 5068 33842 5124 33852
rect 4956 33518 4958 33570
rect 5010 33518 5012 33570
rect 4956 33506 5012 33518
rect 4844 33406 4846 33458
rect 4898 33406 4900 33458
rect 4844 32788 4900 33406
rect 5964 33458 6020 34076
rect 5964 33406 5966 33458
rect 6018 33406 6020 33458
rect 5964 33394 6020 33406
rect 4900 32732 5124 32788
rect 4844 32722 4900 32732
rect 3948 32622 3950 32674
rect 4002 32622 4004 32674
rect 3948 32610 4004 32622
rect 3276 32510 3278 32562
rect 3330 32510 3332 32562
rect 3276 32498 3332 32510
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 5068 30994 5124 32732
rect 6076 32450 6132 34860
rect 6748 34916 6804 34926
rect 7084 34916 7140 39454
rect 7196 39620 7252 39630
rect 7196 39058 7252 39564
rect 7196 39006 7198 39058
rect 7250 39006 7252 39058
rect 7196 38994 7252 39006
rect 7420 39620 7476 39630
rect 7532 39620 7588 40684
rect 7420 39618 7588 39620
rect 7420 39566 7422 39618
rect 7474 39566 7588 39618
rect 7420 39564 7588 39566
rect 7644 40516 7700 40526
rect 7756 40516 7812 40796
rect 7868 40786 7924 40796
rect 7644 40514 7812 40516
rect 7644 40462 7646 40514
rect 7698 40462 7812 40514
rect 7644 40460 7812 40462
rect 7308 36372 7364 36382
rect 7196 34916 7252 34926
rect 7084 34860 7196 34916
rect 6748 34822 6804 34860
rect 7196 34822 7252 34860
rect 6972 34804 7028 34814
rect 6972 34710 7028 34748
rect 7196 34132 7252 34142
rect 7308 34132 7364 36316
rect 7420 35812 7476 39564
rect 7532 38834 7588 38846
rect 7532 38782 7534 38834
rect 7586 38782 7588 38834
rect 7532 38612 7588 38782
rect 7644 38724 7700 40460
rect 7980 39844 8036 44380
rect 8316 44324 8372 44334
rect 8428 44324 8484 45054
rect 8540 44994 8596 45612
rect 8764 45444 8820 45838
rect 8988 45780 9044 45790
rect 8764 45378 8820 45388
rect 8876 45724 8988 45780
rect 8876 45330 8932 45724
rect 8988 45714 9044 45724
rect 9100 45668 9156 56140
rect 9436 55972 9492 59200
rect 9884 56308 9940 59200
rect 10108 56308 10164 56318
rect 9884 56306 10164 56308
rect 9884 56254 10110 56306
rect 10162 56254 10164 56306
rect 9884 56252 10164 56254
rect 10108 56242 10164 56252
rect 9660 55972 9716 55982
rect 9436 55970 9716 55972
rect 9436 55918 9662 55970
rect 9714 55918 9716 55970
rect 9436 55916 9716 55918
rect 9660 55906 9716 55916
rect 10780 55970 10836 59200
rect 11228 56306 11284 59200
rect 12124 57876 12180 59200
rect 11228 56254 11230 56306
rect 11282 56254 11284 56306
rect 11228 56242 11284 56254
rect 11788 57820 12180 57876
rect 10780 55918 10782 55970
rect 10834 55918 10836 55970
rect 10780 55906 10836 55918
rect 11676 55972 11732 55982
rect 11788 55972 11844 57820
rect 12572 57764 12628 59200
rect 12124 57708 12628 57764
rect 12124 56306 12180 57708
rect 12124 56254 12126 56306
rect 12178 56254 12180 56306
rect 12124 56242 12180 56254
rect 12572 56866 12628 56878
rect 12572 56814 12574 56866
rect 12626 56814 12628 56866
rect 11676 55970 11844 55972
rect 11676 55918 11678 55970
rect 11730 55918 11844 55970
rect 11676 55916 11844 55918
rect 12572 55970 12628 56814
rect 13356 56868 13412 56878
rect 13468 56868 13524 59200
rect 13916 57428 13972 59200
rect 13356 56866 13524 56868
rect 13356 56814 13358 56866
rect 13410 56814 13524 56866
rect 13356 56812 13524 56814
rect 13692 57372 13972 57428
rect 13356 56802 13412 56812
rect 12572 55918 12574 55970
rect 12626 55918 12628 55970
rect 11676 55906 11732 55916
rect 12572 55906 12628 55918
rect 13468 56642 13524 56654
rect 13468 56590 13470 56642
rect 13522 56590 13524 56642
rect 13468 55970 13524 56590
rect 13468 55918 13470 55970
rect 13522 55918 13524 55970
rect 13468 55906 13524 55918
rect 11676 55412 11732 55422
rect 10556 55410 11732 55412
rect 10556 55358 11678 55410
rect 11730 55358 11732 55410
rect 10556 55356 11732 55358
rect 9548 55188 9604 55198
rect 9548 55186 9828 55188
rect 9548 55134 9550 55186
rect 9602 55134 9828 55186
rect 9548 55132 9828 55134
rect 9548 55122 9604 55132
rect 9772 54402 9828 55132
rect 9772 54350 9774 54402
rect 9826 54350 9828 54402
rect 9772 54338 9828 54350
rect 9884 54626 9940 54638
rect 9884 54574 9886 54626
rect 9938 54574 9940 54626
rect 9884 54292 9940 54574
rect 9884 54226 9940 54236
rect 9996 54628 10052 54638
rect 9996 53842 10052 54572
rect 10444 54514 10500 54526
rect 10444 54462 10446 54514
rect 10498 54462 10500 54514
rect 9996 53790 9998 53842
rect 10050 53790 10052 53842
rect 9996 53778 10052 53790
rect 10108 54290 10164 54302
rect 10108 54238 10110 54290
rect 10162 54238 10164 54290
rect 10108 53058 10164 54238
rect 10108 53006 10110 53058
rect 10162 53006 10164 53058
rect 10108 52994 10164 53006
rect 10444 52834 10500 54462
rect 10556 52948 10612 55356
rect 11676 55346 11732 55356
rect 13692 55186 13748 57372
rect 14812 56642 14868 59200
rect 14812 56590 14814 56642
rect 14866 56590 14868 56642
rect 14812 56578 14868 56590
rect 14364 56308 14420 56318
rect 14364 56214 14420 56252
rect 15036 56196 15092 56206
rect 15036 56102 15092 56140
rect 14812 56082 14868 56094
rect 14812 56030 14814 56082
rect 14866 56030 14868 56082
rect 13916 55972 13972 55982
rect 13916 55878 13972 55916
rect 14700 55412 14756 55422
rect 14812 55412 14868 56030
rect 15260 55468 15316 59200
rect 15708 56644 15764 59200
rect 15484 56588 15764 56644
rect 14700 55410 14812 55412
rect 14700 55358 14702 55410
rect 14754 55358 14812 55410
rect 14700 55356 14812 55358
rect 14700 55346 14756 55356
rect 14812 55346 14868 55356
rect 15036 55412 15316 55468
rect 15372 56196 15428 56206
rect 15372 55524 15428 56140
rect 13692 55134 13694 55186
rect 13746 55134 13748 55186
rect 13692 55122 13748 55134
rect 15036 55186 15092 55412
rect 15372 55298 15428 55468
rect 15372 55246 15374 55298
rect 15426 55246 15428 55298
rect 15372 55234 15428 55246
rect 15484 56082 15540 56588
rect 15484 56030 15486 56082
rect 15538 56030 15540 56082
rect 15036 55134 15038 55186
rect 15090 55134 15092 55186
rect 15036 55122 15092 55134
rect 15484 54738 15540 56030
rect 15932 56084 15988 56094
rect 15932 55990 15988 56028
rect 16156 55972 16212 59200
rect 16604 56308 16660 59200
rect 16604 56242 16660 56252
rect 16156 55906 16212 55916
rect 16492 55970 16548 55982
rect 16716 55972 16772 55982
rect 16492 55918 16494 55970
rect 16546 55918 16548 55970
rect 16492 55636 16548 55918
rect 16492 55570 16548 55580
rect 16604 55916 16716 55972
rect 16380 55524 16436 55534
rect 15484 54686 15486 54738
rect 15538 54686 15540 54738
rect 15484 54674 15540 54686
rect 15596 55298 15652 55310
rect 15596 55246 15598 55298
rect 15650 55246 15652 55298
rect 15596 54740 15652 55246
rect 15932 55300 15988 55310
rect 15932 55206 15988 55244
rect 16380 55076 16436 55468
rect 16492 55412 16548 55422
rect 16604 55412 16660 55916
rect 16716 55906 16772 55916
rect 17052 55860 17108 59200
rect 17500 56532 17556 59200
rect 17500 56476 17780 56532
rect 16940 55804 17108 55860
rect 16828 55524 16884 55534
rect 16492 55410 16660 55412
rect 16492 55358 16494 55410
rect 16546 55358 16660 55410
rect 16492 55356 16660 55358
rect 16716 55412 16772 55422
rect 16828 55412 16884 55468
rect 16716 55410 16884 55412
rect 16716 55358 16718 55410
rect 16770 55358 16884 55410
rect 16716 55356 16884 55358
rect 16940 55412 16996 55804
rect 17052 55524 17108 55534
rect 17612 55524 17668 55534
rect 17052 55522 17668 55524
rect 17052 55470 17054 55522
rect 17106 55470 17614 55522
rect 17666 55470 17668 55522
rect 17052 55468 17668 55470
rect 17052 55458 17108 55468
rect 17612 55458 17668 55468
rect 16492 55346 16548 55356
rect 16716 55346 16772 55356
rect 16940 55346 16996 55356
rect 17500 55300 17556 55310
rect 17500 55186 17556 55244
rect 17500 55134 17502 55186
rect 17554 55134 17556 55186
rect 17500 55122 17556 55134
rect 17612 55076 17668 55086
rect 16380 55020 16772 55076
rect 15596 54674 15652 54684
rect 16604 54740 16660 54750
rect 10668 54628 10724 54638
rect 10668 54534 10724 54572
rect 11452 54628 11508 54638
rect 11508 54572 11620 54628
rect 11452 54562 11508 54572
rect 10780 54516 10836 54526
rect 10780 54514 10948 54516
rect 10780 54462 10782 54514
rect 10834 54462 10948 54514
rect 10780 54460 10948 54462
rect 10780 54450 10836 54460
rect 10892 52948 10948 54460
rect 11452 52948 11508 52958
rect 10556 52946 10836 52948
rect 10556 52894 10558 52946
rect 10610 52894 10836 52946
rect 10556 52892 10836 52894
rect 10892 52946 11508 52948
rect 10892 52894 11454 52946
rect 11506 52894 11508 52946
rect 10892 52892 11508 52894
rect 11564 52948 11620 54572
rect 16604 54626 16660 54684
rect 16716 54738 16772 55020
rect 16716 54686 16718 54738
rect 16770 54686 16772 54738
rect 16716 54674 16772 54686
rect 17612 54738 17668 55020
rect 17612 54686 17614 54738
rect 17666 54686 17668 54738
rect 17612 54674 17668 54686
rect 16604 54574 16606 54626
rect 16658 54574 16660 54626
rect 16604 54562 16660 54574
rect 16940 54628 16996 54638
rect 16940 54626 17444 54628
rect 16940 54574 16942 54626
rect 16994 54574 17444 54626
rect 16940 54572 17444 54574
rect 16940 54562 16996 54572
rect 16380 54516 16436 54526
rect 16380 54422 16436 54460
rect 17388 54514 17444 54572
rect 17388 54462 17390 54514
rect 17442 54462 17444 54514
rect 17388 54450 17444 54462
rect 15820 54402 15876 54414
rect 15820 54350 15822 54402
rect 15874 54350 15876 54402
rect 12796 53730 12852 53742
rect 12796 53678 12798 53730
rect 12850 53678 12852 53730
rect 12124 53620 12180 53630
rect 11676 53618 12180 53620
rect 11676 53566 12126 53618
rect 12178 53566 12180 53618
rect 11676 53564 12180 53566
rect 11676 53170 11732 53564
rect 12124 53554 12180 53564
rect 12796 53620 12852 53678
rect 12796 53554 12852 53564
rect 13580 53730 13636 53742
rect 13580 53678 13582 53730
rect 13634 53678 13636 53730
rect 13580 53620 13636 53678
rect 13580 53554 13636 53564
rect 14252 53618 14308 53630
rect 14252 53566 14254 53618
rect 14306 53566 14308 53618
rect 11676 53118 11678 53170
rect 11730 53118 11732 53170
rect 11676 53106 11732 53118
rect 14252 53172 14308 53566
rect 14252 53106 14308 53116
rect 15148 53620 15204 53630
rect 11676 52948 11732 52958
rect 11564 52946 11732 52948
rect 11564 52894 11678 52946
rect 11730 52894 11732 52946
rect 11564 52892 11732 52894
rect 10556 52882 10612 52892
rect 10444 52782 10446 52834
rect 10498 52782 10500 52834
rect 10444 52770 10500 52782
rect 9212 52052 9268 52062
rect 9212 52050 10052 52052
rect 9212 51998 9214 52050
rect 9266 51998 10052 52050
rect 9212 51996 10052 51998
rect 9212 51986 9268 51996
rect 9660 51604 9716 51614
rect 9548 50036 9604 50046
rect 9548 49922 9604 49980
rect 9660 50034 9716 51548
rect 9996 51602 10052 51996
rect 9996 51550 9998 51602
rect 10050 51550 10052 51602
rect 9996 51538 10052 51550
rect 10780 51490 10836 52892
rect 11340 52274 11396 52286
rect 11340 52222 11342 52274
rect 11394 52222 11396 52274
rect 11004 51604 11060 51614
rect 11004 51510 11060 51548
rect 11340 51604 11396 52222
rect 11452 52276 11508 52892
rect 11676 52388 11732 52892
rect 11676 52322 11732 52332
rect 11900 52946 11956 52958
rect 11900 52894 11902 52946
rect 11954 52894 11956 52946
rect 11788 52276 11844 52286
rect 11900 52276 11956 52894
rect 11452 52220 11620 52276
rect 11340 51538 11396 51548
rect 11452 52052 11508 52062
rect 10780 51438 10782 51490
rect 10834 51438 10836 51490
rect 10780 51426 10836 51438
rect 9772 51380 9828 51390
rect 9772 50482 9828 51324
rect 9884 51378 9940 51390
rect 9884 51326 9886 51378
rect 9938 51326 9940 51378
rect 9884 50708 9940 51326
rect 10220 51380 10276 51390
rect 10220 51286 10276 51324
rect 10444 51378 10500 51390
rect 10444 51326 10446 51378
rect 10498 51326 10500 51378
rect 10444 50820 10500 51326
rect 11340 51380 11396 51390
rect 11340 51044 11396 51324
rect 11452 51378 11508 51996
rect 11564 51940 11620 52220
rect 11788 52274 11956 52276
rect 11788 52222 11790 52274
rect 11842 52222 11956 52274
rect 11788 52220 11956 52222
rect 13132 52834 13188 52846
rect 13132 52782 13134 52834
rect 13186 52782 13188 52834
rect 11788 52210 11844 52220
rect 11900 52052 11956 52062
rect 11900 51958 11956 51996
rect 11676 51940 11732 51950
rect 12124 51940 12180 51950
rect 11564 51938 11732 51940
rect 11564 51886 11678 51938
rect 11730 51886 11732 51938
rect 11564 51884 11732 51886
rect 11452 51326 11454 51378
rect 11506 51326 11508 51378
rect 11452 51314 11508 51326
rect 11340 50988 11508 51044
rect 10444 50754 10500 50764
rect 11340 50820 11396 50830
rect 9884 50642 9940 50652
rect 11228 50708 11284 50718
rect 10892 50596 10948 50606
rect 10892 50502 10948 50540
rect 11228 50594 11284 50652
rect 11340 50706 11396 50764
rect 11340 50654 11342 50706
rect 11394 50654 11396 50706
rect 11340 50642 11396 50654
rect 11228 50542 11230 50594
rect 11282 50542 11284 50594
rect 11228 50530 11284 50542
rect 11452 50594 11508 50988
rect 11452 50542 11454 50594
rect 11506 50542 11508 50594
rect 9772 50430 9774 50482
rect 9826 50430 9828 50482
rect 9772 50418 9828 50430
rect 10108 50484 10164 50494
rect 10108 50390 10164 50428
rect 10780 50484 10836 50494
rect 11452 50484 11508 50542
rect 10780 50372 11060 50428
rect 11452 50418 11508 50428
rect 9660 49982 9662 50034
rect 9714 49982 9716 50034
rect 9660 49970 9716 49982
rect 10668 49924 10724 49934
rect 9548 49870 9550 49922
rect 9602 49870 9604 49922
rect 9548 49858 9604 49870
rect 10220 49922 10724 49924
rect 10220 49870 10670 49922
rect 10722 49870 10724 49922
rect 10220 49868 10724 49870
rect 9660 49586 9716 49598
rect 9660 49534 9662 49586
rect 9714 49534 9716 49586
rect 9660 48356 9716 49534
rect 10108 49140 10164 49150
rect 9100 45602 9156 45612
rect 9436 48300 9716 48356
rect 9772 49026 9828 49038
rect 9772 48974 9774 49026
rect 9826 48974 9828 49026
rect 8876 45278 8878 45330
rect 8930 45278 8932 45330
rect 8876 45266 8932 45278
rect 8540 44942 8542 44994
rect 8594 44942 8596 44994
rect 8540 44930 8596 44942
rect 8316 44322 8484 44324
rect 8316 44270 8318 44322
rect 8370 44270 8484 44322
rect 8316 44268 8484 44270
rect 8316 44258 8372 44268
rect 9436 43988 9492 48300
rect 9548 48020 9604 48030
rect 9548 47926 9604 47964
rect 9660 48018 9716 48030
rect 9660 47966 9662 48018
rect 9714 47966 9716 48018
rect 9660 47908 9716 47966
rect 9660 47842 9716 47852
rect 9772 47572 9828 48974
rect 9996 49028 10052 49038
rect 9996 48934 10052 48972
rect 10108 48804 10164 49084
rect 9996 48748 10164 48804
rect 9996 48242 10052 48748
rect 9996 48190 9998 48242
rect 10050 48190 10052 48242
rect 9996 48178 10052 48190
rect 9884 48132 9940 48142
rect 9884 48038 9940 48076
rect 10108 47908 10164 47918
rect 10220 47908 10276 49868
rect 10668 49812 10724 49868
rect 10668 49746 10724 49756
rect 11004 49810 11060 50372
rect 11004 49758 11006 49810
rect 11058 49758 11060 49810
rect 10332 49140 10388 49150
rect 10332 49046 10388 49084
rect 10444 49084 10948 49140
rect 10164 47852 10276 47908
rect 10108 47842 10164 47852
rect 9884 47572 9940 47582
rect 9772 47570 9940 47572
rect 9772 47518 9886 47570
rect 9938 47518 9940 47570
rect 9772 47516 9940 47518
rect 9884 47012 9940 47516
rect 9772 46564 9828 46574
rect 9884 46564 9940 46956
rect 10220 46676 10276 46686
rect 10444 46676 10500 49084
rect 10668 48914 10724 48926
rect 10668 48862 10670 48914
rect 10722 48862 10724 48914
rect 10276 46620 10500 46676
rect 10220 46582 10276 46620
rect 9772 46562 9940 46564
rect 9772 46510 9774 46562
rect 9826 46510 9940 46562
rect 9772 46508 9940 46510
rect 9772 45890 9828 46508
rect 10332 46450 10388 46462
rect 10332 46398 10334 46450
rect 10386 46398 10388 46450
rect 9772 45838 9774 45890
rect 9826 45838 9828 45890
rect 9772 45826 9828 45838
rect 10108 46002 10164 46014
rect 10108 45950 10110 46002
rect 10162 45950 10164 46002
rect 9660 45780 9716 45790
rect 9660 45686 9716 45724
rect 9660 45444 9716 45454
rect 9660 45330 9716 45388
rect 10108 45332 10164 45950
rect 9660 45278 9662 45330
rect 9714 45278 9716 45330
rect 9660 45266 9716 45278
rect 9772 45276 10164 45332
rect 9436 43922 9492 43932
rect 9548 44434 9604 44446
rect 9548 44382 9550 44434
rect 9602 44382 9604 44434
rect 9548 44324 9604 44382
rect 9548 43538 9604 44268
rect 9772 44212 9828 45276
rect 10220 45220 10276 45230
rect 9772 43650 9828 44156
rect 9884 44212 9940 44222
rect 10220 44212 10276 45164
rect 10332 44322 10388 46398
rect 10444 45780 10500 46620
rect 10556 48130 10612 48142
rect 10556 48078 10558 48130
rect 10610 48078 10612 48130
rect 10556 46900 10612 48078
rect 10556 46674 10612 46844
rect 10668 46788 10724 48862
rect 10892 48914 10948 49084
rect 10892 48862 10894 48914
rect 10946 48862 10948 48914
rect 10892 48850 10948 48862
rect 10780 48802 10836 48814
rect 10780 48750 10782 48802
rect 10834 48750 10836 48802
rect 10780 48244 10836 48750
rect 10780 48188 10948 48244
rect 10780 48018 10836 48030
rect 10780 47966 10782 48018
rect 10834 47966 10836 48018
rect 10780 47460 10836 47966
rect 10892 47682 10948 48188
rect 11004 48132 11060 49758
rect 11564 49812 11620 49822
rect 11564 49718 11620 49756
rect 11228 49588 11284 49598
rect 11228 49028 11284 49532
rect 11452 49586 11508 49598
rect 11452 49534 11454 49586
rect 11506 49534 11508 49586
rect 11452 49028 11508 49534
rect 11676 49252 11732 51884
rect 12012 51938 12180 51940
rect 12012 51886 12126 51938
rect 12178 51886 12180 51938
rect 12012 51884 12180 51886
rect 11900 50596 11956 50606
rect 12012 50596 12068 51884
rect 12124 51874 12180 51884
rect 12348 51604 12404 51614
rect 12348 51492 12404 51548
rect 11956 50540 12068 50596
rect 12236 51490 12404 51492
rect 12236 51438 12350 51490
rect 12402 51438 12404 51490
rect 12236 51436 12404 51438
rect 12236 50594 12292 51436
rect 12348 51426 12404 51436
rect 12460 51380 12516 51390
rect 13132 51380 13188 52782
rect 12460 51378 12852 51380
rect 12460 51326 12462 51378
rect 12514 51326 12852 51378
rect 12460 51324 12852 51326
rect 12460 51314 12516 51324
rect 12572 50708 12628 50718
rect 12628 50652 12740 50708
rect 12572 50642 12628 50652
rect 12236 50542 12238 50594
rect 12290 50542 12292 50594
rect 11900 50502 11956 50540
rect 12236 50530 12292 50542
rect 12460 50484 12516 50494
rect 12516 50428 12628 50484
rect 12460 50390 12516 50428
rect 11900 49812 11956 49822
rect 11900 49718 11956 49756
rect 12348 49810 12404 49822
rect 12348 49758 12350 49810
rect 12402 49758 12404 49810
rect 12348 49700 12404 49758
rect 12460 49812 12516 49822
rect 12460 49718 12516 49756
rect 12572 49810 12628 50428
rect 12572 49758 12574 49810
rect 12626 49758 12628 49810
rect 12348 49634 12404 49644
rect 11788 49588 11844 49598
rect 11788 49494 11844 49532
rect 11676 49186 11732 49196
rect 12012 49364 12068 49374
rect 12012 49140 12068 49308
rect 11788 49084 12068 49140
rect 11788 49028 11844 49084
rect 11452 48972 11620 49028
rect 11116 48916 11172 48926
rect 11116 48466 11172 48860
rect 11228 48804 11284 48972
rect 11452 48804 11508 48814
rect 11228 48802 11508 48804
rect 11228 48750 11454 48802
rect 11506 48750 11508 48802
rect 11228 48748 11508 48750
rect 11452 48738 11508 48748
rect 11116 48414 11118 48466
rect 11170 48414 11172 48466
rect 11116 48402 11172 48414
rect 11564 48356 11620 48972
rect 11564 48290 11620 48300
rect 11676 48972 11844 49028
rect 12012 49026 12068 49084
rect 12012 48974 12014 49026
rect 12066 48974 12068 49026
rect 11452 48132 11508 48142
rect 11676 48132 11732 48972
rect 12012 48962 12068 48974
rect 12236 49028 12292 49038
rect 12572 49028 12628 49758
rect 12236 49026 12628 49028
rect 12236 48974 12238 49026
rect 12290 48974 12628 49026
rect 12236 48972 12628 48974
rect 12684 49700 12740 50652
rect 12236 48962 12292 48972
rect 11900 48916 11956 48926
rect 11900 48822 11956 48860
rect 12572 48804 12628 48814
rect 12684 48804 12740 49644
rect 12796 49810 12852 51324
rect 13132 51286 13188 51324
rect 15148 51380 15204 53564
rect 15820 53620 15876 54350
rect 17724 53954 17780 56476
rect 17836 56194 17892 56206
rect 17836 56142 17838 56194
rect 17890 56142 17892 56194
rect 17836 55300 17892 56142
rect 17836 54626 17892 55244
rect 17836 54574 17838 54626
rect 17890 54574 17892 54626
rect 17836 54562 17892 54574
rect 17724 53902 17726 53954
rect 17778 53902 17780 53954
rect 17724 53890 17780 53902
rect 15820 53554 15876 53564
rect 16380 53842 16436 53854
rect 16380 53790 16382 53842
rect 16434 53790 16436 53842
rect 16380 53508 16436 53790
rect 17948 53620 18004 59200
rect 18396 56420 18452 59200
rect 18172 56364 18452 56420
rect 18060 55636 18116 55646
rect 18060 55076 18116 55580
rect 18060 55010 18116 55020
rect 18172 53844 18228 56364
rect 18732 56308 18788 56318
rect 18172 53778 18228 53788
rect 18284 56306 18788 56308
rect 18284 56254 18734 56306
rect 18786 56254 18788 56306
rect 18284 56252 18788 56254
rect 18172 53620 18228 53630
rect 17948 53618 18228 53620
rect 17948 53566 18174 53618
rect 18226 53566 18228 53618
rect 17948 53564 18228 53566
rect 18172 53554 18228 53564
rect 16380 53442 16436 53452
rect 16716 53506 16772 53518
rect 16716 53454 16718 53506
rect 16770 53454 16772 53506
rect 16044 53172 16100 53210
rect 16044 53106 16100 53116
rect 15820 52946 15876 52958
rect 15820 52894 15822 52946
rect 15874 52894 15876 52946
rect 15820 52388 15876 52894
rect 16156 52948 16212 52958
rect 16604 52948 16660 52958
rect 16156 52946 16436 52948
rect 16156 52894 16158 52946
rect 16210 52894 16436 52946
rect 16156 52892 16436 52894
rect 16156 52882 16212 52892
rect 16268 52724 16324 52734
rect 15820 52322 15876 52332
rect 16156 52722 16324 52724
rect 16156 52670 16270 52722
rect 16322 52670 16324 52722
rect 16156 52668 16324 52670
rect 16380 52724 16436 52892
rect 16604 52854 16660 52892
rect 16716 52724 16772 53454
rect 17052 53508 17108 53518
rect 17108 53452 17332 53508
rect 17052 53414 17108 53452
rect 16380 52668 16772 52724
rect 16156 52274 16212 52668
rect 16268 52658 16324 52668
rect 16156 52222 16158 52274
rect 16210 52222 16212 52274
rect 16156 52210 16212 52222
rect 16268 52388 16324 52398
rect 15708 52164 15764 52174
rect 16268 52164 16324 52332
rect 15708 52162 16100 52164
rect 15708 52110 15710 52162
rect 15762 52110 16100 52162
rect 15708 52108 16100 52110
rect 15708 52098 15764 52108
rect 15484 52052 15540 52062
rect 15484 51958 15540 51996
rect 16044 52052 16100 52108
rect 16268 52162 16548 52164
rect 16268 52110 16270 52162
rect 16322 52110 16548 52162
rect 16268 52108 16548 52110
rect 16268 52098 16324 52108
rect 16044 52050 16212 52052
rect 16044 51998 16046 52050
rect 16098 51998 16212 52050
rect 16044 51996 16212 51998
rect 16044 51986 16100 51996
rect 15148 51314 15204 51324
rect 15596 51938 15652 51950
rect 15596 51886 15598 51938
rect 15650 51886 15652 51938
rect 13916 51266 13972 51278
rect 13916 51214 13918 51266
rect 13970 51214 13972 51266
rect 13916 50372 13972 51214
rect 15596 50818 15652 51886
rect 16156 51604 16212 51996
rect 16492 51828 16548 52108
rect 16604 52162 16660 52668
rect 16604 52110 16606 52162
rect 16658 52110 16660 52162
rect 16604 52052 16660 52110
rect 17052 52164 17108 52174
rect 17052 52070 17108 52108
rect 16604 51986 16660 51996
rect 16940 51940 16996 51950
rect 16828 51884 16940 51940
rect 16492 51772 16660 51828
rect 16492 51604 16548 51614
rect 16156 51602 16548 51604
rect 16156 51550 16494 51602
rect 16546 51550 16548 51602
rect 16156 51548 16548 51550
rect 16492 51538 16548 51548
rect 15596 50766 15598 50818
rect 15650 50766 15652 50818
rect 15596 50754 15652 50766
rect 15932 51380 15988 51390
rect 16156 51380 16212 51390
rect 15932 50708 15988 51324
rect 16044 51324 16156 51380
rect 16044 51266 16100 51324
rect 16156 51314 16212 51324
rect 16044 51214 16046 51266
rect 16098 51214 16100 51266
rect 16044 51202 16100 51214
rect 16044 50820 16100 50830
rect 16044 50818 16324 50820
rect 16044 50766 16046 50818
rect 16098 50766 16324 50818
rect 16044 50764 16324 50766
rect 16044 50754 16100 50764
rect 15932 50614 15988 50652
rect 16268 50594 16324 50764
rect 16268 50542 16270 50594
rect 16322 50542 16324 50594
rect 16268 50530 16324 50542
rect 16604 50594 16660 51772
rect 16716 51492 16772 51502
rect 16716 51398 16772 51436
rect 16828 51490 16884 51884
rect 16940 51874 16996 51884
rect 17276 51938 17332 53452
rect 18284 53172 18340 56252
rect 18732 56242 18788 56252
rect 18732 56082 18788 56094
rect 18732 56030 18734 56082
rect 18786 56030 18788 56082
rect 18732 55636 18788 56030
rect 18844 55748 18900 59200
rect 19068 55972 19124 55982
rect 19068 55878 19124 55916
rect 19292 55748 19348 59200
rect 19740 56644 19796 59200
rect 19628 56588 19796 56644
rect 20188 56642 20244 59200
rect 20188 56590 20190 56642
rect 20242 56590 20244 56642
rect 19628 56196 19684 56588
rect 20188 56578 20244 56590
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19628 56140 20020 56196
rect 19852 55972 19908 55982
rect 18844 55692 19124 55748
rect 19292 55692 19572 55748
rect 18732 55580 18900 55636
rect 18844 55412 18900 55580
rect 18844 55346 18900 55356
rect 18396 55300 18452 55310
rect 18396 54626 18452 55244
rect 18956 55298 19012 55310
rect 18956 55246 18958 55298
rect 19010 55246 19012 55298
rect 18844 55188 18900 55198
rect 18844 55094 18900 55132
rect 18956 55076 19012 55246
rect 18956 55010 19012 55020
rect 18396 54574 18398 54626
rect 18450 54574 18452 54626
rect 18396 54562 18452 54574
rect 18732 54516 18788 54526
rect 18956 54516 19012 54526
rect 18788 54514 19012 54516
rect 18788 54462 18958 54514
rect 19010 54462 19012 54514
rect 18788 54460 19012 54462
rect 18732 54450 18788 54460
rect 18956 54450 19012 54460
rect 19068 53954 19124 55692
rect 19292 55412 19348 55422
rect 19292 54516 19348 55356
rect 19516 54740 19572 55692
rect 19628 55522 19684 55534
rect 19628 55470 19630 55522
rect 19682 55470 19684 55522
rect 19628 55300 19684 55470
rect 19628 55234 19684 55244
rect 19852 55298 19908 55916
rect 19964 55412 20020 56140
rect 19964 55346 20020 55356
rect 20524 55412 20580 55422
rect 19852 55246 19854 55298
rect 19906 55246 19908 55298
rect 19852 55234 19908 55246
rect 20300 55298 20356 55310
rect 20300 55246 20302 55298
rect 20354 55246 20356 55298
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19516 54684 19796 54740
rect 19404 54628 19460 54638
rect 19460 54572 19572 54628
rect 19404 54562 19460 54572
rect 19292 54422 19348 54460
rect 19516 54514 19572 54572
rect 19516 54462 19518 54514
rect 19570 54462 19572 54514
rect 19516 54450 19572 54462
rect 19404 54404 19460 54414
rect 19404 54310 19460 54348
rect 19068 53902 19070 53954
rect 19122 53902 19124 53954
rect 19068 53890 19124 53902
rect 18844 53844 18900 53854
rect 18844 53750 18900 53788
rect 19740 53620 19796 54684
rect 19852 54514 19908 54526
rect 19852 54462 19854 54514
rect 19906 54462 19908 54514
rect 19852 53844 19908 54462
rect 20300 54516 20356 55246
rect 20300 54402 20356 54460
rect 20300 54350 20302 54402
rect 20354 54350 20356 54402
rect 20300 54338 20356 54350
rect 19852 53778 19908 53788
rect 20524 53842 20580 55356
rect 20636 55186 20692 59200
rect 20748 56642 20804 56654
rect 20748 56590 20750 56642
rect 20802 56590 20804 56642
rect 20748 55970 20804 56590
rect 21196 56084 21252 56094
rect 20748 55918 20750 55970
rect 20802 55918 20804 55970
rect 20748 55906 20804 55918
rect 20972 56082 21252 56084
rect 20972 56030 21198 56082
rect 21250 56030 21252 56082
rect 20972 56028 21252 56030
rect 20636 55134 20638 55186
rect 20690 55134 20692 55186
rect 20636 55122 20692 55134
rect 20748 54628 20804 54638
rect 20748 54534 20804 54572
rect 20524 53790 20526 53842
rect 20578 53790 20580 53842
rect 20524 53778 20580 53790
rect 19852 53620 19908 53630
rect 19740 53618 19908 53620
rect 19740 53566 19854 53618
rect 19906 53566 19908 53618
rect 19740 53564 19908 53566
rect 19852 53554 19908 53564
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 18172 53116 18340 53172
rect 17948 52834 18004 52846
rect 17948 52782 17950 52834
rect 18002 52782 18004 52834
rect 17276 51886 17278 51938
rect 17330 51886 17332 51938
rect 17276 51874 17332 51886
rect 17500 52388 17556 52398
rect 17500 51938 17556 52332
rect 17948 52386 18004 52782
rect 17948 52334 17950 52386
rect 18002 52334 18004 52386
rect 17948 52322 18004 52334
rect 17612 52164 17668 52174
rect 17836 52164 17892 52174
rect 17668 52162 17892 52164
rect 17668 52110 17838 52162
rect 17890 52110 17892 52162
rect 17668 52108 17892 52110
rect 17612 52098 17668 52108
rect 17500 51886 17502 51938
rect 17554 51886 17556 51938
rect 17500 51874 17556 51886
rect 17612 51938 17668 51950
rect 17612 51886 17614 51938
rect 17666 51886 17668 51938
rect 16828 51438 16830 51490
rect 16882 51438 16884 51490
rect 16828 51426 16884 51438
rect 17612 51378 17668 51886
rect 17612 51326 17614 51378
rect 17666 51326 17668 51378
rect 17612 51314 17668 51326
rect 17388 51268 17444 51278
rect 16940 51266 17444 51268
rect 16940 51214 17390 51266
rect 17442 51214 17444 51266
rect 16940 51212 17444 51214
rect 16828 50820 16884 50830
rect 16940 50820 16996 51212
rect 17388 51202 17444 51212
rect 16828 50818 16996 50820
rect 16828 50766 16830 50818
rect 16882 50766 16996 50818
rect 16828 50764 16996 50766
rect 16828 50754 16884 50764
rect 16604 50542 16606 50594
rect 16658 50542 16660 50594
rect 16604 50428 16660 50542
rect 17052 50594 17108 50606
rect 17052 50542 17054 50594
rect 17106 50542 17108 50594
rect 16716 50484 16772 50494
rect 13916 50306 13972 50316
rect 16380 50372 16436 50382
rect 16604 50372 16772 50428
rect 16380 50278 16436 50316
rect 12796 49758 12798 49810
rect 12850 49758 12852 49810
rect 12796 49364 12852 49758
rect 16604 49922 16660 49934
rect 16604 49870 16606 49922
rect 16658 49870 16660 49922
rect 12796 49298 12852 49308
rect 16492 49586 16548 49598
rect 16492 49534 16494 49586
rect 16546 49534 16548 49586
rect 12796 49026 12852 49038
rect 12796 48974 12798 49026
rect 12850 48974 12852 49026
rect 12796 48916 12852 48974
rect 12796 48850 12852 48860
rect 14364 49026 14420 49038
rect 14364 48974 14366 49026
rect 14418 48974 14420 49026
rect 11004 48076 11172 48132
rect 10892 47630 10894 47682
rect 10946 47630 10948 47682
rect 10892 47618 10948 47630
rect 11004 47460 11060 47470
rect 10780 47404 11004 47460
rect 11004 47366 11060 47404
rect 11116 47236 11172 48076
rect 11452 48130 11732 48132
rect 11452 48078 11454 48130
rect 11506 48078 11732 48130
rect 11452 48076 11732 48078
rect 12236 48802 12740 48804
rect 12236 48750 12574 48802
rect 12626 48750 12740 48802
rect 12236 48748 12740 48750
rect 11452 48066 11508 48076
rect 11228 47572 11284 47582
rect 11788 47572 11844 47582
rect 11284 47570 11844 47572
rect 11284 47518 11790 47570
rect 11842 47518 11844 47570
rect 11284 47516 11844 47518
rect 11228 47478 11284 47516
rect 11788 47506 11844 47516
rect 12012 47458 12068 47470
rect 12012 47406 12014 47458
rect 12066 47406 12068 47458
rect 11340 47346 11396 47358
rect 11340 47294 11342 47346
rect 11394 47294 11396 47346
rect 11228 47236 11284 47246
rect 11116 47180 11228 47236
rect 11228 47170 11284 47180
rect 10668 46722 10724 46732
rect 10556 46622 10558 46674
rect 10610 46622 10612 46674
rect 10556 46610 10612 46622
rect 11340 46116 11396 47294
rect 11676 47346 11732 47358
rect 11676 47294 11678 47346
rect 11730 47294 11732 47346
rect 11676 46788 11732 47294
rect 11676 46722 11732 46732
rect 11788 47236 11844 47246
rect 12012 47236 12068 47406
rect 12236 47458 12292 48748
rect 12572 48738 12628 48748
rect 13580 48356 13636 48366
rect 13580 48262 13636 48300
rect 14364 48244 14420 48974
rect 15036 48914 15092 48926
rect 15036 48862 15038 48914
rect 15090 48862 15092 48914
rect 15036 48356 15092 48862
rect 15036 48290 15092 48300
rect 16044 48356 16100 48366
rect 16044 48262 16100 48300
rect 14812 48244 14868 48254
rect 14364 48242 14868 48244
rect 14364 48190 14366 48242
rect 14418 48190 14814 48242
rect 14866 48190 14868 48242
rect 14364 48188 14868 48190
rect 14364 48178 14420 48188
rect 14812 47572 14868 48188
rect 16156 48244 16212 48254
rect 12236 47406 12238 47458
rect 12290 47406 12292 47458
rect 12236 47394 12292 47406
rect 12572 47460 12628 47470
rect 12572 47366 12628 47404
rect 12684 47236 12740 47246
rect 12012 47234 12740 47236
rect 12012 47182 12686 47234
rect 12738 47182 12740 47234
rect 12012 47180 12740 47182
rect 11340 46050 11396 46060
rect 10668 45780 10724 45790
rect 10444 45778 11172 45780
rect 10444 45726 10670 45778
rect 10722 45726 11172 45778
rect 10444 45724 11172 45726
rect 10668 45714 10724 45724
rect 10332 44270 10334 44322
rect 10386 44270 10388 44322
rect 10332 44258 10388 44270
rect 10556 45332 10612 45342
rect 9884 44210 10276 44212
rect 9884 44158 9886 44210
rect 9938 44158 10276 44210
rect 9884 44156 10276 44158
rect 10556 44210 10612 45276
rect 11116 45330 11172 45724
rect 11116 45278 11118 45330
rect 11170 45278 11172 45330
rect 11116 45266 11172 45278
rect 11788 44546 11844 47180
rect 12684 47170 12740 47180
rect 12796 47234 12852 47246
rect 12796 47182 12798 47234
rect 12850 47182 12852 47234
rect 11900 46900 11956 46910
rect 11900 46564 11956 46844
rect 12796 46900 12852 47182
rect 12796 46834 12852 46844
rect 14028 46788 14084 46798
rect 14028 46694 14084 46732
rect 14812 46674 14868 47516
rect 15260 47572 15316 47582
rect 16156 47572 16212 48188
rect 16380 48244 16436 48254
rect 16492 48244 16548 49534
rect 16604 49476 16660 49870
rect 16604 49410 16660 49420
rect 16380 48242 16548 48244
rect 16380 48190 16382 48242
rect 16434 48190 16548 48242
rect 16380 48188 16548 48190
rect 16604 48244 16660 48254
rect 16716 48244 16772 50372
rect 16828 49812 16884 49822
rect 16828 49718 16884 49756
rect 17052 49588 17108 50542
rect 17724 50594 17780 52108
rect 17836 52098 17892 52108
rect 17948 52052 18004 52062
rect 17948 51958 18004 51996
rect 18060 51492 18116 51502
rect 18060 51378 18116 51436
rect 18060 51326 18062 51378
rect 18114 51326 18116 51378
rect 18060 51314 18116 51326
rect 18172 50932 18228 53116
rect 18284 52946 18340 52958
rect 18284 52894 18286 52946
rect 18338 52894 18340 52946
rect 18284 52388 18340 52894
rect 19180 52946 19236 52958
rect 19180 52894 19182 52946
rect 19234 52894 19236 52946
rect 18732 52836 18788 52846
rect 18732 52742 18788 52780
rect 18284 52276 18340 52332
rect 18508 52276 18564 52286
rect 18284 52220 18508 52276
rect 18508 52182 18564 52220
rect 18396 51940 18452 51950
rect 18396 51846 18452 51884
rect 17724 50542 17726 50594
rect 17778 50542 17780 50594
rect 17388 50484 17444 50522
rect 17724 50428 17780 50542
rect 17388 50418 17444 50428
rect 17500 50372 17780 50428
rect 18060 50876 18228 50932
rect 18284 51604 18340 51614
rect 19180 51604 19236 52894
rect 19628 52948 19684 52958
rect 19404 52836 19460 52846
rect 19404 52386 19460 52780
rect 19404 52334 19406 52386
rect 19458 52334 19460 52386
rect 19404 52322 19460 52334
rect 19628 52164 19684 52892
rect 19852 52834 19908 52846
rect 19852 52782 19854 52834
rect 19906 52782 19908 52834
rect 19740 52388 19796 52398
rect 19852 52388 19908 52782
rect 19740 52386 19908 52388
rect 19740 52334 19742 52386
rect 19794 52334 19908 52386
rect 19740 52332 19908 52334
rect 19740 52322 19796 52332
rect 19740 52164 19796 52174
rect 19628 52108 19740 52164
rect 19292 51604 19348 51614
rect 19180 51548 19292 51604
rect 18060 50428 18116 50876
rect 18172 50708 18228 50718
rect 18284 50708 18340 51548
rect 19292 51378 19348 51548
rect 19292 51326 19294 51378
rect 19346 51326 19348 51378
rect 19292 51314 19348 51326
rect 19180 51268 19236 51278
rect 18228 50652 18340 50708
rect 19068 51212 19180 51268
rect 18172 50614 18228 50652
rect 18956 50596 19012 50606
rect 18956 50502 19012 50540
rect 18844 50484 18900 50494
rect 18060 50372 18452 50428
rect 18844 50390 18900 50428
rect 17388 50036 17444 50046
rect 17500 50036 17556 50372
rect 17388 50034 17556 50036
rect 17388 49982 17390 50034
rect 17442 49982 17556 50034
rect 17388 49980 17556 49982
rect 17388 49970 17444 49980
rect 17724 49812 17780 49822
rect 17724 49718 17780 49756
rect 17052 49522 17108 49532
rect 17948 49698 18004 49710
rect 17948 49646 17950 49698
rect 18002 49646 18004 49698
rect 17164 49476 17220 49486
rect 17164 49138 17220 49420
rect 17948 49476 18004 49646
rect 17948 49410 18004 49420
rect 17164 49086 17166 49138
rect 17218 49086 17220 49138
rect 17164 49074 17220 49086
rect 16604 48242 16772 48244
rect 16604 48190 16606 48242
rect 16658 48190 16772 48242
rect 16604 48188 16772 48190
rect 17276 48916 17332 48926
rect 16380 48178 16436 48188
rect 16604 48178 16660 48188
rect 15260 46898 15316 47516
rect 15932 47516 16212 47572
rect 16604 47572 16660 47582
rect 15932 47458 15988 47516
rect 16268 47460 16324 47470
rect 15932 47406 15934 47458
rect 15986 47406 15988 47458
rect 15932 47394 15988 47406
rect 16156 47404 16268 47460
rect 16156 47346 16212 47404
rect 16268 47394 16324 47404
rect 16604 47458 16660 47516
rect 17276 47570 17332 48860
rect 17500 48802 17556 48814
rect 17500 48750 17502 48802
rect 17554 48750 17556 48802
rect 17500 48244 17556 48750
rect 17836 48804 17892 48814
rect 17836 48710 17892 48748
rect 17276 47518 17278 47570
rect 17330 47518 17332 47570
rect 17276 47506 17332 47518
rect 17388 48188 17500 48244
rect 16604 47406 16606 47458
rect 16658 47406 16660 47458
rect 16604 47394 16660 47406
rect 16156 47294 16158 47346
rect 16210 47294 16212 47346
rect 16156 47282 16212 47294
rect 15260 46846 15262 46898
rect 15314 46846 15316 46898
rect 15260 46834 15316 46846
rect 14812 46622 14814 46674
rect 14866 46622 14868 46674
rect 14812 46610 14868 46622
rect 11900 46562 12292 46564
rect 11900 46510 11902 46562
rect 11954 46510 12292 46562
rect 11900 46508 12292 46510
rect 11900 46498 11956 46508
rect 12236 45890 12292 46508
rect 12236 45838 12238 45890
rect 12290 45838 12292 45890
rect 12236 45826 12292 45838
rect 13356 46116 13412 46126
rect 13244 45668 13300 45678
rect 11788 44494 11790 44546
rect 11842 44494 11844 44546
rect 11788 44482 11844 44494
rect 12796 45332 12852 45342
rect 12124 44436 12180 44446
rect 12124 44342 12180 44380
rect 12796 44434 12852 45276
rect 12796 44382 12798 44434
rect 12850 44382 12852 44434
rect 12796 44370 12852 44382
rect 13244 44436 13300 45612
rect 13356 45218 13412 46060
rect 17276 46116 17332 46126
rect 17388 46116 17444 48188
rect 17500 48178 17556 48188
rect 17948 48242 18004 48254
rect 17948 48190 17950 48242
rect 18002 48190 18004 48242
rect 17276 46114 17444 46116
rect 17276 46062 17278 46114
rect 17330 46062 17444 46114
rect 17276 46060 17444 46062
rect 17948 46676 18004 48190
rect 17276 46050 17332 46060
rect 16940 46004 16996 46014
rect 16940 45910 16996 45948
rect 17612 46004 17668 46014
rect 17612 45910 17668 45948
rect 17836 46004 17892 46014
rect 13356 45166 13358 45218
rect 13410 45166 13412 45218
rect 13356 45154 13412 45166
rect 14140 45890 14196 45902
rect 14140 45838 14142 45890
rect 14194 45838 14196 45890
rect 14140 45108 14196 45838
rect 14812 45780 14868 45790
rect 14812 45686 14868 45724
rect 15372 45780 15428 45790
rect 14140 45014 14196 45052
rect 14588 45108 14644 45118
rect 14588 45014 14644 45052
rect 10556 44158 10558 44210
rect 10610 44158 10612 44210
rect 9884 44146 9940 44156
rect 10556 44146 10612 44158
rect 12348 44210 12404 44222
rect 12348 44158 12350 44210
rect 12402 44158 12404 44210
rect 11676 44100 11732 44110
rect 10556 43988 10612 43998
rect 10108 43764 10164 43774
rect 10108 43670 10164 43708
rect 9772 43598 9774 43650
rect 9826 43598 9828 43650
rect 9772 43586 9828 43598
rect 9548 43486 9550 43538
rect 9602 43486 9604 43538
rect 9548 43474 9604 43486
rect 10556 43538 10612 43932
rect 11452 43652 11508 43662
rect 11452 43558 11508 43596
rect 10556 43486 10558 43538
rect 10610 43486 10612 43538
rect 10556 43474 10612 43486
rect 11004 43538 11060 43550
rect 11004 43486 11006 43538
rect 11058 43486 11060 43538
rect 9548 42868 9604 42878
rect 9548 42866 9940 42868
rect 9548 42814 9550 42866
rect 9602 42814 9940 42866
rect 9548 42812 9940 42814
rect 9548 42802 9604 42812
rect 9884 42194 9940 42812
rect 9884 42142 9886 42194
rect 9938 42142 9940 42194
rect 8988 41972 9044 41982
rect 8876 41860 8932 41870
rect 8092 40964 8148 40974
rect 8092 40626 8148 40908
rect 8092 40574 8094 40626
rect 8146 40574 8148 40626
rect 8092 40562 8148 40574
rect 8876 40626 8932 41804
rect 8988 41858 9044 41916
rect 8988 41806 8990 41858
rect 9042 41806 9044 41858
rect 8988 41794 9044 41806
rect 9884 41298 9940 42142
rect 9884 41246 9886 41298
rect 9938 41246 9940 41298
rect 9884 41234 9940 41246
rect 9996 42532 10052 42542
rect 9212 40964 9268 40974
rect 9212 40870 9268 40908
rect 9996 40964 10052 42476
rect 10780 42532 10836 42542
rect 10780 42438 10836 42476
rect 10668 42196 10724 42206
rect 10332 42194 10724 42196
rect 10332 42142 10670 42194
rect 10722 42142 10724 42194
rect 10332 42140 10724 42142
rect 10220 42084 10276 42094
rect 10332 42084 10388 42140
rect 10668 42130 10724 42140
rect 10892 42196 10948 42206
rect 11004 42196 11060 43486
rect 11676 43538 11732 44044
rect 12348 44100 12404 44158
rect 12348 44034 12404 44044
rect 11676 43486 11678 43538
rect 11730 43486 11732 43538
rect 11676 43474 11732 43486
rect 12236 43538 12292 43550
rect 12236 43486 12238 43538
rect 12290 43486 12292 43538
rect 10892 42194 11060 42196
rect 10892 42142 10894 42194
rect 10946 42142 11060 42194
rect 10892 42140 11060 42142
rect 10892 42130 10948 42140
rect 10220 42082 10388 42084
rect 10220 42030 10222 42082
rect 10274 42030 10388 42082
rect 10220 42028 10388 42030
rect 10220 42018 10276 42028
rect 9996 40898 10052 40908
rect 10108 41972 10164 41982
rect 10108 41186 10164 41916
rect 10108 41134 10110 41186
rect 10162 41134 10164 41186
rect 10108 40740 10164 41134
rect 8876 40574 8878 40626
rect 8930 40574 8932 40626
rect 8876 40562 8932 40574
rect 9996 40684 10164 40740
rect 9884 40516 9940 40526
rect 9660 40514 9940 40516
rect 9660 40462 9886 40514
rect 9938 40462 9940 40514
rect 9660 40460 9940 40462
rect 8316 40404 8372 40414
rect 8540 40404 8596 40414
rect 9660 40404 9716 40460
rect 9884 40450 9940 40460
rect 8372 40348 8484 40404
rect 8316 40338 8372 40348
rect 7980 39730 8036 39788
rect 7980 39678 7982 39730
rect 8034 39678 8036 39730
rect 7980 39666 8036 39678
rect 8316 39620 8372 39630
rect 8316 39526 8372 39564
rect 8428 39060 8484 40348
rect 8540 40402 9716 40404
rect 8540 40350 8542 40402
rect 8594 40350 9716 40402
rect 8540 40348 9716 40350
rect 8540 40338 8596 40348
rect 9772 40292 9828 40302
rect 9772 40198 9828 40236
rect 8764 40178 8820 40190
rect 8764 40126 8766 40178
rect 8818 40126 8820 40178
rect 8764 39732 8820 40126
rect 8876 40180 8932 40190
rect 8876 40178 9380 40180
rect 8876 40126 8878 40178
rect 8930 40126 9380 40178
rect 8876 40124 9380 40126
rect 8876 40114 8932 40124
rect 8764 39666 8820 39676
rect 9324 39730 9380 40124
rect 9324 39678 9326 39730
rect 9378 39678 9380 39730
rect 9324 39666 9380 39678
rect 9660 39620 9716 39630
rect 9660 39526 9716 39564
rect 9884 39620 9940 39630
rect 9996 39620 10052 40684
rect 10108 40516 10164 40526
rect 10108 40422 10164 40460
rect 10220 40404 10276 40414
rect 10220 40310 10276 40348
rect 10332 40180 10388 42028
rect 10556 41972 10612 41982
rect 10556 41878 10612 41916
rect 11004 41748 11060 42140
rect 11116 42532 11172 42542
rect 11116 41970 11172 42476
rect 11788 42532 11844 42542
rect 11788 42438 11844 42476
rect 12236 42532 12292 43486
rect 12236 42466 12292 42476
rect 12908 43426 12964 43438
rect 12908 43374 12910 43426
rect 12962 43374 12964 43426
rect 11116 41918 11118 41970
rect 11170 41918 11172 41970
rect 11116 41906 11172 41918
rect 11900 41860 11956 41870
rect 11900 41858 12068 41860
rect 11900 41806 11902 41858
rect 11954 41806 12068 41858
rect 11900 41804 12068 41806
rect 11900 41794 11956 41804
rect 11004 41692 11284 41748
rect 10444 40964 10500 40974
rect 10444 40962 10612 40964
rect 10444 40910 10446 40962
rect 10498 40910 10612 40962
rect 10444 40908 10612 40910
rect 10444 40898 10500 40908
rect 10556 40516 10612 40908
rect 10668 40628 10724 40638
rect 10668 40516 10724 40572
rect 11228 40570 11284 41692
rect 10556 40514 10724 40516
rect 10556 40462 10558 40514
rect 10610 40462 10724 40514
rect 10556 40460 10724 40462
rect 10892 40514 10948 40526
rect 10892 40462 10894 40514
rect 10946 40462 10948 40514
rect 11228 40518 11230 40570
rect 11282 40518 11284 40570
rect 11452 40628 11508 40638
rect 11228 40506 11284 40518
rect 11340 40514 11396 40526
rect 10556 40450 10612 40460
rect 10332 40114 10388 40124
rect 10892 40404 10948 40462
rect 11340 40462 11342 40514
rect 11394 40462 11396 40514
rect 11340 40404 11396 40462
rect 10948 40348 11396 40404
rect 10108 39844 10164 39854
rect 10108 39750 10164 39788
rect 9884 39618 10052 39620
rect 9884 39566 9886 39618
rect 9938 39566 10052 39618
rect 9884 39564 10052 39566
rect 9884 39554 9940 39564
rect 8764 39508 8820 39518
rect 8652 39506 8820 39508
rect 8652 39454 8766 39506
rect 8818 39454 8820 39506
rect 8652 39452 8820 39454
rect 8540 39060 8596 39070
rect 8428 39058 8596 39060
rect 8428 39006 8542 39058
rect 8594 39006 8596 39058
rect 8428 39004 8596 39006
rect 8540 38994 8596 39004
rect 7644 38658 7700 38668
rect 8316 38834 8372 38846
rect 8316 38782 8318 38834
rect 8370 38782 8372 38834
rect 8316 38668 8372 38782
rect 8540 38836 8596 38846
rect 8652 38836 8708 39452
rect 8764 39442 8820 39452
rect 9212 39396 9268 39406
rect 9212 39302 9268 39340
rect 9436 39396 9492 39406
rect 9884 39396 9940 39406
rect 9436 39394 9828 39396
rect 9436 39342 9438 39394
rect 9490 39342 9828 39394
rect 9436 39340 9828 39342
rect 9436 39330 9492 39340
rect 8540 38834 8708 38836
rect 8540 38782 8542 38834
rect 8594 38782 8708 38834
rect 8540 38780 8708 38782
rect 8764 38836 8820 38846
rect 8540 38770 8596 38780
rect 8764 38742 8820 38780
rect 8988 38834 9044 38846
rect 8988 38782 8990 38834
rect 9042 38782 9044 38834
rect 8988 38668 9044 38782
rect 9660 38834 9716 38846
rect 9660 38782 9662 38834
rect 9714 38782 9716 38834
rect 8316 38612 8484 38668
rect 8988 38612 9604 38668
rect 7532 38052 7588 38556
rect 8316 38388 8372 38398
rect 7532 37986 7588 37996
rect 7644 38050 7700 38062
rect 7644 37998 7646 38050
rect 7698 37998 7700 38050
rect 7644 36708 7700 37998
rect 8204 37826 8260 37838
rect 8204 37774 8206 37826
rect 8258 37774 8260 37826
rect 7756 37380 7812 37390
rect 7756 37286 7812 37324
rect 7980 36708 8036 36718
rect 7644 36706 8036 36708
rect 7644 36654 7646 36706
rect 7698 36654 7982 36706
rect 8034 36654 8036 36706
rect 7644 36652 8036 36654
rect 7644 36642 7700 36652
rect 7980 36642 8036 36652
rect 8204 36596 8260 37774
rect 8316 37154 8372 38332
rect 8428 37828 8484 38612
rect 8428 37762 8484 37772
rect 9212 37828 9268 37838
rect 8316 37102 8318 37154
rect 8370 37102 8372 37154
rect 8316 37090 8372 37102
rect 8876 37266 8932 37278
rect 8876 37214 8878 37266
rect 8930 37214 8932 37266
rect 8316 36708 8372 36718
rect 8316 36614 8372 36652
rect 8204 36530 8260 36540
rect 8652 36482 8708 36494
rect 8652 36430 8654 36482
rect 8706 36430 8708 36482
rect 7532 36372 7588 36382
rect 7532 36278 7588 36316
rect 8204 36260 8260 36270
rect 8204 36166 8260 36204
rect 7868 35812 7924 35822
rect 7420 35810 7924 35812
rect 7420 35758 7870 35810
rect 7922 35758 7924 35810
rect 7420 35756 7924 35758
rect 7868 35746 7924 35756
rect 7980 35698 8036 35710
rect 7980 35646 7982 35698
rect 8034 35646 8036 35698
rect 7420 35476 7476 35486
rect 7420 35382 7476 35420
rect 7980 35140 8036 35646
rect 8204 35700 8260 35710
rect 8204 35698 8372 35700
rect 8204 35646 8206 35698
rect 8258 35646 8372 35698
rect 8204 35644 8372 35646
rect 8204 35634 8260 35644
rect 8204 35140 8260 35150
rect 7644 35138 8260 35140
rect 7644 35086 8206 35138
rect 8258 35086 8260 35138
rect 7644 35084 8260 35086
rect 7644 34916 7700 35084
rect 7532 34914 7700 34916
rect 7532 34862 7646 34914
rect 7698 34862 7700 34914
rect 7532 34860 7700 34862
rect 7420 34692 7476 34702
rect 7420 34598 7476 34636
rect 7420 34356 7476 34366
rect 7532 34356 7588 34860
rect 7644 34850 7700 34860
rect 7756 34916 7812 34926
rect 7420 34354 7588 34356
rect 7420 34302 7422 34354
rect 7474 34302 7588 34354
rect 7420 34300 7588 34302
rect 7420 34290 7476 34300
rect 7756 34242 7812 34860
rect 7868 34804 7924 34814
rect 7868 34710 7924 34748
rect 7756 34190 7758 34242
rect 7810 34190 7812 34242
rect 7756 34178 7812 34190
rect 7980 34242 8036 35084
rect 8204 35074 8260 35084
rect 8204 34804 8260 34814
rect 8316 34804 8372 35644
rect 8652 35588 8708 36430
rect 8876 36484 8932 37214
rect 9100 36820 9156 36830
rect 8876 36418 8932 36428
rect 8988 36764 9100 36820
rect 8652 35494 8708 35532
rect 8652 35252 8708 35262
rect 8428 34916 8484 34926
rect 8428 34822 8484 34860
rect 8652 34914 8708 35196
rect 8652 34862 8654 34914
rect 8706 34862 8708 34914
rect 8652 34850 8708 34862
rect 8876 34916 8932 34926
rect 8988 34916 9044 36764
rect 9100 36754 9156 36764
rect 8876 34914 9044 34916
rect 8876 34862 8878 34914
rect 8930 34862 9044 34914
rect 8876 34860 9044 34862
rect 8876 34850 8932 34860
rect 9212 34804 9268 37772
rect 9548 37490 9604 38612
rect 9660 38164 9716 38782
rect 9772 38276 9828 39340
rect 9772 38210 9828 38220
rect 9996 39396 10052 39564
rect 10444 39508 10500 39518
rect 10332 39506 10500 39508
rect 10332 39454 10446 39506
rect 10498 39454 10500 39506
rect 10332 39452 10500 39454
rect 9996 39340 10164 39396
rect 9884 39060 9940 39340
rect 9660 38098 9716 38108
rect 9548 37438 9550 37490
rect 9602 37438 9604 37490
rect 9548 37426 9604 37438
rect 9884 37380 9940 39004
rect 9772 37324 9940 37380
rect 9996 38836 10052 38846
rect 9660 37154 9716 37166
rect 9660 37102 9662 37154
rect 9714 37102 9716 37154
rect 9660 36820 9716 37102
rect 9660 36754 9716 36764
rect 9436 36484 9492 36494
rect 9436 36390 9492 36428
rect 8260 34748 8372 34804
rect 8988 34748 9268 34804
rect 9324 35588 9380 35598
rect 8204 34738 8260 34748
rect 8764 34690 8820 34702
rect 8764 34638 8766 34690
rect 8818 34638 8820 34690
rect 7980 34190 7982 34242
rect 8034 34190 8036 34242
rect 7980 34178 8036 34190
rect 8092 34354 8148 34366
rect 8092 34302 8094 34354
rect 8146 34302 8148 34354
rect 7252 34076 7364 34132
rect 7196 34038 7252 34076
rect 8092 33458 8148 34302
rect 8652 34354 8708 34366
rect 8652 34302 8654 34354
rect 8706 34302 8708 34354
rect 8540 34132 8596 34142
rect 8652 34132 8708 34302
rect 8540 34130 8708 34132
rect 8540 34078 8542 34130
rect 8594 34078 8708 34130
rect 8540 34076 8708 34078
rect 8540 34066 8596 34076
rect 8316 33908 8372 33918
rect 8764 33908 8820 34638
rect 8876 34356 8932 34366
rect 8988 34356 9044 34748
rect 8876 34354 9044 34356
rect 8876 34302 8878 34354
rect 8930 34302 8990 34354
rect 9042 34302 9044 34354
rect 8876 34300 9044 34302
rect 8876 34290 8932 34300
rect 8988 34290 9044 34300
rect 8316 33906 8820 33908
rect 8316 33854 8318 33906
rect 8370 33854 8820 33906
rect 8316 33852 8820 33854
rect 8316 33842 8372 33852
rect 9324 33572 9380 35532
rect 9772 35364 9828 37324
rect 9884 37156 9940 37166
rect 9884 36370 9940 37100
rect 9884 36318 9886 36370
rect 9938 36318 9940 36370
rect 9884 36306 9940 36318
rect 9660 35308 9828 35364
rect 9660 35252 9716 35308
rect 9996 35252 10052 38780
rect 10108 38724 10164 39340
rect 10332 39058 10388 39452
rect 10444 39442 10500 39452
rect 10556 39396 10612 39406
rect 10556 39302 10612 39340
rect 10780 39394 10836 39406
rect 10780 39342 10782 39394
rect 10834 39342 10836 39394
rect 10780 39284 10836 39342
rect 10780 39218 10836 39228
rect 10332 39006 10334 39058
rect 10386 39006 10388 39058
rect 10332 38994 10388 39006
rect 10892 39060 10948 40348
rect 11340 40178 11396 40190
rect 11340 40126 11342 40178
rect 11394 40126 11396 40178
rect 11116 39844 11172 39854
rect 11116 39730 11172 39788
rect 11116 39678 11118 39730
rect 11170 39678 11172 39730
rect 11116 39666 11172 39678
rect 11004 39620 11060 39630
rect 11004 39526 11060 39564
rect 11340 39172 11396 40126
rect 11340 39106 11396 39116
rect 10892 39004 11060 39060
rect 10220 38948 10276 38958
rect 10220 38854 10276 38892
rect 10668 38946 10724 38958
rect 10668 38894 10670 38946
rect 10722 38894 10724 38946
rect 10556 38724 10612 38734
rect 10108 38722 10612 38724
rect 10108 38670 10558 38722
rect 10610 38670 10612 38722
rect 10108 38668 10612 38670
rect 10556 38658 10612 38668
rect 10444 38500 10500 38510
rect 10332 38388 10388 38398
rect 10220 38276 10276 38286
rect 10220 38050 10276 38220
rect 10220 37998 10222 38050
rect 10274 37998 10276 38050
rect 10220 37986 10276 37998
rect 10332 37380 10388 38332
rect 10444 37940 10500 38444
rect 10668 38388 10724 38894
rect 10892 38836 10948 38846
rect 10668 38322 10724 38332
rect 10780 38834 10948 38836
rect 10780 38782 10894 38834
rect 10946 38782 10948 38834
rect 10780 38780 10948 38782
rect 10668 38164 10724 38174
rect 10556 38108 10668 38164
rect 10556 38050 10612 38108
rect 10668 38098 10724 38108
rect 10556 37998 10558 38050
rect 10610 37998 10612 38050
rect 10556 37986 10612 37998
rect 10444 37846 10500 37884
rect 10556 37716 10612 37726
rect 10332 37324 10500 37380
rect 10332 37156 10388 37166
rect 10220 37154 10388 37156
rect 10220 37102 10334 37154
rect 10386 37102 10388 37154
rect 10220 37100 10388 37102
rect 10108 36708 10164 36718
rect 10108 36484 10164 36652
rect 10220 36706 10276 37100
rect 10332 37090 10388 37100
rect 10220 36654 10222 36706
rect 10274 36654 10276 36706
rect 10220 36642 10276 36654
rect 10108 36390 10164 36428
rect 9660 35186 9716 35196
rect 9772 35196 10052 35252
rect 9772 34356 9828 35196
rect 10108 35140 10164 35150
rect 10332 35140 10388 35150
rect 10108 35138 10332 35140
rect 10108 35086 10110 35138
rect 10162 35086 10332 35138
rect 10108 35084 10332 35086
rect 10108 35074 10164 35084
rect 10332 35074 10388 35084
rect 9884 35028 9940 35038
rect 9884 34802 9940 34972
rect 9884 34750 9886 34802
rect 9938 34750 9940 34802
rect 9884 34738 9940 34750
rect 9996 34804 10052 34814
rect 9996 34710 10052 34748
rect 10444 34802 10500 37324
rect 10556 36370 10612 37660
rect 10556 36318 10558 36370
rect 10610 36318 10612 36370
rect 10556 36306 10612 36318
rect 10668 36482 10724 36494
rect 10668 36430 10670 36482
rect 10722 36430 10724 36482
rect 10668 36372 10724 36430
rect 10780 36484 10836 38780
rect 10892 38770 10948 38780
rect 10892 37268 10948 37278
rect 11004 37268 11060 39004
rect 11340 38836 11396 38846
rect 11452 38836 11508 40572
rect 12012 40626 12068 41804
rect 12012 40574 12014 40626
rect 12066 40574 12068 40626
rect 12012 40562 12068 40574
rect 12460 40740 12516 40750
rect 11564 40516 11620 40526
rect 11564 39396 11620 40460
rect 12012 40402 12068 40414
rect 12460 40404 12516 40684
rect 12908 40516 12964 43374
rect 12908 40450 12964 40460
rect 12012 40350 12014 40402
rect 12066 40350 12068 40402
rect 12012 40292 12068 40350
rect 11900 39396 11956 39406
rect 11564 39394 11900 39396
rect 11564 39342 11566 39394
rect 11618 39342 11900 39394
rect 11564 39340 11900 39342
rect 11564 39330 11620 39340
rect 11564 39060 11620 39070
rect 11564 38966 11620 39004
rect 11900 39058 11956 39340
rect 11900 39006 11902 39058
rect 11954 39006 11956 39058
rect 11900 38994 11956 39006
rect 12012 38948 12068 40236
rect 12012 38882 12068 38892
rect 12236 40402 12516 40404
rect 12236 40350 12462 40402
rect 12514 40350 12516 40402
rect 12236 40348 12516 40350
rect 11340 38834 11508 38836
rect 11340 38782 11342 38834
rect 11394 38782 11508 38834
rect 11340 38780 11508 38782
rect 11340 38770 11396 38780
rect 12236 38668 12292 40348
rect 12460 40338 12516 40348
rect 12796 40402 12852 40414
rect 12796 40350 12798 40402
rect 12850 40350 12852 40402
rect 12348 40178 12404 40190
rect 12348 40126 12350 40178
rect 12402 40126 12404 40178
rect 12348 39732 12404 40126
rect 12348 39666 12404 39676
rect 12796 39620 12852 40350
rect 12796 39554 12852 39564
rect 12908 39506 12964 39518
rect 12908 39454 12910 39506
rect 12962 39454 12964 39506
rect 12796 39396 12852 39406
rect 12348 39394 12852 39396
rect 12348 39342 12798 39394
rect 12850 39342 12852 39394
rect 12348 39340 12852 39342
rect 12348 38834 12404 39340
rect 12796 39330 12852 39340
rect 12684 39172 12740 39182
rect 12348 38782 12350 38834
rect 12402 38782 12404 38834
rect 12348 38770 12404 38782
rect 12460 38836 12516 38846
rect 12236 38612 12404 38668
rect 11564 38500 11620 38510
rect 11116 38050 11172 38062
rect 11564 38052 11620 38444
rect 11116 37998 11118 38050
rect 11170 37998 11172 38050
rect 11116 37716 11172 37998
rect 11116 37650 11172 37660
rect 11228 38050 11620 38052
rect 11228 37998 11566 38050
rect 11618 37998 11620 38050
rect 11228 37996 11620 37998
rect 10892 37266 11060 37268
rect 10892 37214 10894 37266
rect 10946 37214 11060 37266
rect 10892 37212 11060 37214
rect 10892 37202 10948 37212
rect 10780 36418 10836 36428
rect 10668 35698 10724 36316
rect 10892 35924 10948 35934
rect 10668 35646 10670 35698
rect 10722 35646 10724 35698
rect 10668 35634 10724 35646
rect 10780 35868 10892 35924
rect 10668 34916 10724 34926
rect 10780 34916 10836 35868
rect 10892 35858 10948 35868
rect 10892 35700 10948 35710
rect 11004 35700 11060 37212
rect 11228 37266 11284 37996
rect 11564 37986 11620 37996
rect 11228 37214 11230 37266
rect 11282 37214 11284 37266
rect 11228 36372 11284 37214
rect 11676 37938 11732 37950
rect 11676 37886 11678 37938
rect 11730 37886 11732 37938
rect 11340 37044 11396 37054
rect 11340 36950 11396 36988
rect 10892 35698 11060 35700
rect 10892 35646 10894 35698
rect 10946 35646 11060 35698
rect 10892 35644 11060 35646
rect 11116 36316 11284 36372
rect 11564 36708 11620 36718
rect 11564 36594 11620 36652
rect 11564 36542 11566 36594
rect 11618 36542 11620 36594
rect 10892 35634 10948 35644
rect 11116 35140 11172 36316
rect 11228 36148 11284 36158
rect 11228 35922 11284 36092
rect 11228 35870 11230 35922
rect 11282 35870 11284 35922
rect 11228 35858 11284 35870
rect 11564 35924 11620 36542
rect 11564 35858 11620 35868
rect 11676 36484 11732 37886
rect 12348 37378 12404 38612
rect 12348 37326 12350 37378
rect 12402 37326 12404 37378
rect 12348 37314 12404 37326
rect 11788 37266 11844 37278
rect 11788 37214 11790 37266
rect 11842 37214 11844 37266
rect 11788 37156 11844 37214
rect 11788 37090 11844 37100
rect 11676 35700 11732 36428
rect 12124 36596 12180 36606
rect 12124 36260 12180 36540
rect 12124 35810 12180 36204
rect 12124 35758 12126 35810
rect 12178 35758 12180 35810
rect 12124 35746 12180 35758
rect 11788 35700 11844 35710
rect 11676 35698 11844 35700
rect 11676 35646 11790 35698
rect 11842 35646 11844 35698
rect 11676 35644 11844 35646
rect 11788 35634 11844 35644
rect 11116 35074 11172 35084
rect 11452 35252 11508 35262
rect 10668 34914 10836 34916
rect 10668 34862 10670 34914
rect 10722 34862 10836 34914
rect 10668 34860 10836 34862
rect 10668 34850 10724 34860
rect 10444 34750 10446 34802
rect 10498 34750 10500 34802
rect 10332 34692 10388 34702
rect 10220 34690 10388 34692
rect 10220 34638 10334 34690
rect 10386 34638 10388 34690
rect 10220 34636 10388 34638
rect 9996 34356 10052 34366
rect 9772 34354 10052 34356
rect 9772 34302 9998 34354
rect 10050 34302 10052 34354
rect 9772 34300 10052 34302
rect 9996 34290 10052 34300
rect 10108 34356 10164 34366
rect 10220 34356 10276 34636
rect 10108 34354 10276 34356
rect 10108 34302 10110 34354
rect 10162 34302 10276 34354
rect 10108 34300 10276 34302
rect 10108 34290 10164 34300
rect 9884 34130 9940 34142
rect 9884 34078 9886 34130
rect 9938 34078 9940 34130
rect 9884 34020 9940 34078
rect 9884 33954 9940 33964
rect 10332 33684 10388 34636
rect 10444 34468 10500 34750
rect 10444 34402 10500 34412
rect 10780 34242 10836 34860
rect 10892 34804 10948 34814
rect 10892 34710 10948 34748
rect 11452 34802 11508 35196
rect 12460 35140 12516 38780
rect 12572 38612 12628 38622
rect 12572 38518 12628 38556
rect 12684 38050 12740 39116
rect 12796 38948 12852 38958
rect 12796 38854 12852 38892
rect 12684 37998 12686 38050
rect 12738 37998 12740 38050
rect 12684 37986 12740 37998
rect 12796 38276 12852 38286
rect 12796 37938 12852 38220
rect 12908 38164 12964 39454
rect 13132 39396 13188 39406
rect 13020 38834 13076 38846
rect 13020 38782 13022 38834
rect 13074 38782 13076 38834
rect 13020 38724 13076 38782
rect 13020 38658 13076 38668
rect 13132 38722 13188 39340
rect 13132 38670 13134 38722
rect 13186 38670 13188 38722
rect 13132 38658 13188 38670
rect 12908 38098 12964 38108
rect 12796 37886 12798 37938
rect 12850 37886 12852 37938
rect 12796 37874 12852 37886
rect 13020 37826 13076 37838
rect 13020 37774 13022 37826
rect 13074 37774 13076 37826
rect 13020 37380 13076 37774
rect 13020 37314 13076 37324
rect 13244 36484 13300 44380
rect 14812 44436 14868 44446
rect 14812 44342 14868 44380
rect 15148 44436 15204 44446
rect 15148 44322 15204 44380
rect 15148 44270 15150 44322
rect 15202 44270 15204 44322
rect 15148 44258 15204 44270
rect 15036 43426 15092 43438
rect 15036 43374 15038 43426
rect 15090 43374 15092 43426
rect 14924 42756 14980 42766
rect 15036 42756 15092 43374
rect 14924 42754 15092 42756
rect 14924 42702 14926 42754
rect 14978 42702 15092 42754
rect 14924 42700 15092 42702
rect 14924 42690 14980 42700
rect 15036 42644 15092 42700
rect 15036 42588 15316 42644
rect 14588 42532 14644 42542
rect 14588 42530 15092 42532
rect 14588 42478 14590 42530
rect 14642 42478 15092 42530
rect 14588 42476 15092 42478
rect 14588 42466 14644 42476
rect 14476 42084 14532 42094
rect 14812 42084 14868 42094
rect 14476 42082 14868 42084
rect 14476 42030 14478 42082
rect 14530 42030 14814 42082
rect 14866 42030 14868 42082
rect 14476 42028 14868 42030
rect 14364 41972 14420 41982
rect 14028 41916 14364 41972
rect 14028 41858 14084 41916
rect 14364 41878 14420 41916
rect 14028 41806 14030 41858
rect 14082 41806 14084 41858
rect 14028 41794 14084 41806
rect 14252 41748 14308 41758
rect 14252 41298 14308 41692
rect 14252 41246 14254 41298
rect 14306 41246 14308 41298
rect 14252 41234 14308 41246
rect 13580 41186 13636 41198
rect 13580 41134 13582 41186
rect 13634 41134 13636 41186
rect 13468 40628 13524 40638
rect 13468 40534 13524 40572
rect 13580 40404 13636 41134
rect 14364 41188 14420 41198
rect 14476 41188 14532 42028
rect 14812 42018 14868 42028
rect 14364 41186 14532 41188
rect 14364 41134 14366 41186
rect 14418 41134 14532 41186
rect 14364 41132 14532 41134
rect 14812 41186 14868 41198
rect 15036 41188 15092 42476
rect 15260 41970 15316 42588
rect 15260 41918 15262 41970
rect 15314 41918 15316 41970
rect 15260 41906 15316 41918
rect 14812 41134 14814 41186
rect 14866 41134 14868 41186
rect 14364 41122 14420 41132
rect 14812 41076 14868 41134
rect 14812 41010 14868 41020
rect 14924 41186 15092 41188
rect 14924 41134 15038 41186
rect 15090 41134 15092 41186
rect 14924 41132 15092 41134
rect 13804 40964 13860 40974
rect 14140 40964 14196 40974
rect 13580 40310 13636 40348
rect 13692 40962 14196 40964
rect 13692 40910 13806 40962
rect 13858 40910 14142 40962
rect 14194 40910 14196 40962
rect 13692 40908 14196 40910
rect 13468 40180 13524 40190
rect 13468 39844 13524 40124
rect 13468 39778 13524 39788
rect 13580 39732 13636 39742
rect 13580 39638 13636 39676
rect 13468 39620 13524 39630
rect 13468 39058 13524 39564
rect 13468 39006 13470 39058
rect 13522 39006 13524 39058
rect 13468 38994 13524 39006
rect 13692 39618 13748 40908
rect 13804 40898 13860 40908
rect 14140 40898 14196 40908
rect 14252 40964 14308 40974
rect 13804 40404 13860 40414
rect 14252 40404 14308 40908
rect 14924 40852 14980 41132
rect 15036 41122 15092 41132
rect 15260 41188 15316 41198
rect 13804 40402 14308 40404
rect 13804 40350 13806 40402
rect 13858 40350 14254 40402
rect 14306 40350 14308 40402
rect 13804 40348 14308 40350
rect 13804 40338 13860 40348
rect 13692 39566 13694 39618
rect 13746 39566 13748 39618
rect 13580 38948 13636 38958
rect 13580 38854 13636 38892
rect 13692 38834 13748 39566
rect 14028 39618 14084 40348
rect 14252 40338 14308 40348
rect 14476 40796 14980 40852
rect 15148 40962 15204 40974
rect 15148 40910 15150 40962
rect 15202 40910 15204 40962
rect 15148 40852 15204 40910
rect 15260 40964 15316 41132
rect 15260 40898 15316 40908
rect 14476 40404 14532 40796
rect 15148 40786 15204 40796
rect 14812 40628 14868 40638
rect 14812 40534 14868 40572
rect 14588 40516 14644 40526
rect 14644 40460 14756 40516
rect 14588 40450 14644 40460
rect 14476 40310 14532 40348
rect 14028 39566 14030 39618
rect 14082 39566 14084 39618
rect 14028 39554 14084 39566
rect 14364 38948 14420 38958
rect 14420 38892 14644 38948
rect 14364 38882 14420 38892
rect 13692 38782 13694 38834
rect 13746 38782 13748 38834
rect 13356 38724 13412 38734
rect 13692 38668 13748 38782
rect 14140 38834 14196 38846
rect 14140 38782 14142 38834
rect 14194 38782 14196 38834
rect 13356 38612 13524 38668
rect 13692 38612 14084 38668
rect 13468 38500 13524 38612
rect 13468 38434 13524 38444
rect 13804 38052 13860 38062
rect 13804 37958 13860 37996
rect 14028 38050 14084 38612
rect 14140 38162 14196 38782
rect 14252 38836 14308 38846
rect 14252 38742 14308 38780
rect 14588 38834 14644 38892
rect 14588 38782 14590 38834
rect 14642 38782 14644 38834
rect 14588 38770 14644 38782
rect 14476 38722 14532 38734
rect 14476 38670 14478 38722
rect 14530 38670 14532 38722
rect 14476 38668 14532 38670
rect 14700 38668 14756 40460
rect 15148 40292 15204 40302
rect 14924 39508 14980 39518
rect 14924 38946 14980 39452
rect 14924 38894 14926 38946
rect 14978 38894 14980 38946
rect 14924 38882 14980 38894
rect 14476 38612 14756 38668
rect 15148 38724 15204 40236
rect 15372 40068 15428 45724
rect 16268 45220 16324 45230
rect 16044 44322 16100 44334
rect 16044 44270 16046 44322
rect 16098 44270 16100 44322
rect 15484 44100 15540 44110
rect 16044 44100 16100 44270
rect 16268 44210 16324 45164
rect 17836 45220 17892 45948
rect 17948 45444 18004 46620
rect 17948 45378 18004 45388
rect 17836 45154 17892 45164
rect 16268 44158 16270 44210
rect 16322 44158 16324 44210
rect 16268 44146 16324 44158
rect 16716 45108 16772 45118
rect 16716 44322 16772 45052
rect 18060 45106 18116 45118
rect 18060 45054 18062 45106
rect 18114 45054 18116 45106
rect 17500 44996 17556 45006
rect 18060 44996 18116 45054
rect 17500 44994 18116 44996
rect 17500 44942 17502 44994
rect 17554 44942 18116 44994
rect 17500 44940 18116 44942
rect 17500 44930 17556 44940
rect 16716 44270 16718 44322
rect 16770 44270 16772 44322
rect 15540 44044 16100 44100
rect 15484 44006 15540 44044
rect 16044 42756 16100 44044
rect 16716 43988 16772 44270
rect 16716 43922 16772 43932
rect 17388 44210 17444 44222
rect 17388 44158 17390 44210
rect 17442 44158 17444 44210
rect 17052 43652 17108 43662
rect 16716 42980 16772 42990
rect 16268 42756 16324 42766
rect 16044 42754 16324 42756
rect 16044 42702 16270 42754
rect 16322 42702 16324 42754
rect 16044 42700 16324 42702
rect 16268 42690 16324 42700
rect 16380 42532 16436 42542
rect 16380 42530 16660 42532
rect 16380 42478 16382 42530
rect 16434 42478 16660 42530
rect 16380 42476 16660 42478
rect 16380 42466 16436 42476
rect 15820 42082 15876 42094
rect 15820 42030 15822 42082
rect 15874 42030 15876 42082
rect 15484 41860 15540 41870
rect 15484 41858 15764 41860
rect 15484 41806 15486 41858
rect 15538 41806 15764 41858
rect 15484 41804 15764 41806
rect 15484 41794 15540 41804
rect 15484 40962 15540 40974
rect 15484 40910 15486 40962
rect 15538 40910 15540 40962
rect 15484 40404 15540 40910
rect 15708 40964 15764 41804
rect 15820 41188 15876 42030
rect 16044 41972 16100 41982
rect 16044 41878 16100 41916
rect 15820 41122 15876 41132
rect 16268 41188 16324 41198
rect 16268 41094 16324 41132
rect 15932 41074 15988 41086
rect 15932 41022 15934 41074
rect 15986 41022 15988 41074
rect 15708 40908 15876 40964
rect 15820 40740 15876 40908
rect 15932 40740 15988 41022
rect 15820 40684 15988 40740
rect 16044 41076 16100 41086
rect 16044 40962 16100 41020
rect 16044 40910 16046 40962
rect 16098 40910 16100 40962
rect 15708 40404 15764 40414
rect 15484 40402 15764 40404
rect 15484 40350 15710 40402
rect 15762 40350 15764 40402
rect 15484 40348 15764 40350
rect 15372 40002 15428 40012
rect 15708 39956 15764 40348
rect 15820 40292 15876 40684
rect 15932 40516 15988 40526
rect 16044 40516 16100 40910
rect 16380 41076 16436 41086
rect 16156 40852 16212 40862
rect 16212 40796 16324 40852
rect 16156 40786 16212 40796
rect 15932 40514 16044 40516
rect 15932 40462 15934 40514
rect 15986 40462 16044 40514
rect 15932 40460 16044 40462
rect 15932 40450 15988 40460
rect 16044 40450 16100 40460
rect 16268 40514 16324 40796
rect 16380 40626 16436 41020
rect 16380 40574 16382 40626
rect 16434 40574 16436 40626
rect 16380 40562 16436 40574
rect 16268 40462 16270 40514
rect 16322 40462 16324 40514
rect 16268 40450 16324 40462
rect 15820 40226 15876 40236
rect 16268 40068 16324 40078
rect 15708 39900 15988 39956
rect 15932 39732 15988 39900
rect 16156 39732 16212 39742
rect 15932 39730 16212 39732
rect 15932 39678 16158 39730
rect 16210 39678 16212 39730
rect 15932 39676 16212 39678
rect 15484 39620 15540 39630
rect 15820 39620 15876 39630
rect 15484 39618 15820 39620
rect 15484 39566 15486 39618
rect 15538 39566 15820 39618
rect 15484 39564 15820 39566
rect 15484 39554 15540 39564
rect 15820 39526 15876 39564
rect 15932 39508 15988 39518
rect 15932 39058 15988 39452
rect 15932 39006 15934 39058
rect 15986 39006 15988 39058
rect 15932 38994 15988 39006
rect 15372 38948 15428 38958
rect 15148 38658 15204 38668
rect 15260 38946 15428 38948
rect 15260 38894 15374 38946
rect 15426 38894 15428 38946
rect 15260 38892 15428 38894
rect 14476 38500 14532 38510
rect 14532 38444 14644 38500
rect 14476 38434 14532 38444
rect 14140 38110 14142 38162
rect 14194 38110 14196 38162
rect 14140 38098 14196 38110
rect 14028 37998 14030 38050
rect 14082 37998 14084 38050
rect 14028 37986 14084 37998
rect 14364 38050 14420 38062
rect 14364 37998 14366 38050
rect 14418 37998 14420 38050
rect 13468 37940 13524 37950
rect 13468 36596 13524 37884
rect 14252 37826 14308 37838
rect 14252 37774 14254 37826
rect 14306 37774 14308 37826
rect 13580 37380 13636 37390
rect 13580 37378 13860 37380
rect 13580 37326 13582 37378
rect 13634 37326 13860 37378
rect 13580 37324 13860 37326
rect 13580 37314 13636 37324
rect 13468 36530 13524 36540
rect 13804 36708 13860 37324
rect 13804 36652 14196 36708
rect 12908 36428 13300 36484
rect 12684 36370 12740 36382
rect 12684 36318 12686 36370
rect 12738 36318 12740 36370
rect 12684 36036 12740 36318
rect 12796 36372 12852 36382
rect 12796 36278 12852 36316
rect 12684 35970 12740 35980
rect 12796 35140 12852 35150
rect 12460 35138 12852 35140
rect 12460 35086 12798 35138
rect 12850 35086 12852 35138
rect 12460 35084 12852 35086
rect 12796 35074 12852 35084
rect 11452 34750 11454 34802
rect 11506 34750 11508 34802
rect 11452 34738 11508 34750
rect 11564 34804 11620 34814
rect 11620 34748 11732 34804
rect 11564 34738 11620 34748
rect 10780 34190 10782 34242
rect 10834 34190 10836 34242
rect 10780 34178 10836 34190
rect 11004 34692 11060 34702
rect 10444 34132 10500 34142
rect 10444 34038 10500 34076
rect 11004 34132 11060 34636
rect 11564 34468 11620 34478
rect 11060 34076 11508 34132
rect 11004 34038 11060 34076
rect 10332 33628 10836 33684
rect 9324 33506 9380 33516
rect 10780 33570 10836 33628
rect 10780 33518 10782 33570
rect 10834 33518 10836 33570
rect 10780 33506 10836 33518
rect 8092 33406 8094 33458
rect 8146 33406 8148 33458
rect 8092 33394 8148 33406
rect 8764 33346 8820 33358
rect 8764 33294 8766 33346
rect 8818 33294 8820 33346
rect 8540 33124 8596 33134
rect 6076 32398 6078 32450
rect 6130 32398 6132 32450
rect 6076 32386 6132 32398
rect 6524 32788 6580 32798
rect 6524 31892 6580 32732
rect 6524 31826 6580 31836
rect 6748 32452 6804 32462
rect 6300 31668 6356 31678
rect 6748 31668 6804 32396
rect 7756 31892 7812 31902
rect 7756 31778 7812 31836
rect 8204 31892 8260 31902
rect 8260 31836 8372 31892
rect 8204 31826 8260 31836
rect 7756 31726 7758 31778
rect 7810 31726 7812 31778
rect 7756 31714 7812 31726
rect 6300 31666 6804 31668
rect 6300 31614 6302 31666
rect 6354 31614 6804 31666
rect 6300 31612 6804 31614
rect 6300 31602 6356 31612
rect 6188 31556 6244 31566
rect 5740 31554 6244 31556
rect 5740 31502 6190 31554
rect 6242 31502 6244 31554
rect 5740 31500 6244 31502
rect 5740 31106 5796 31500
rect 6188 31490 6244 31500
rect 5740 31054 5742 31106
rect 5794 31054 5796 31106
rect 5740 31042 5796 31054
rect 7868 31332 7924 31342
rect 5068 30942 5070 30994
rect 5122 30942 5124 30994
rect 5068 30930 5124 30942
rect 7868 30882 7924 31276
rect 7868 30830 7870 30882
rect 7922 30830 7924 30882
rect 7868 30818 7924 30830
rect 8204 31106 8260 31118
rect 8204 31054 8206 31106
rect 8258 31054 8260 31106
rect 7308 30772 7364 30782
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 7308 30434 7364 30716
rect 7308 30382 7310 30434
rect 7362 30382 7364 30434
rect 7308 30370 7364 30382
rect 6972 30324 7028 30334
rect 1596 29922 1652 29932
rect 6860 30322 7028 30324
rect 6860 30270 6974 30322
rect 7026 30270 7028 30322
rect 6860 30268 7028 30270
rect 6860 29538 6916 30268
rect 6972 30258 7028 30268
rect 6860 29486 6862 29538
rect 6914 29486 6916 29538
rect 6860 29474 6916 29486
rect 7084 29988 7140 29998
rect 8204 29988 8260 31054
rect 8316 30210 8372 31836
rect 8540 31890 8596 33068
rect 8764 33124 8820 33294
rect 10556 33346 10612 33358
rect 10556 33294 10558 33346
rect 10610 33294 10612 33346
rect 9324 33124 9380 33134
rect 8764 33122 9380 33124
rect 8764 33070 9326 33122
rect 9378 33070 9380 33122
rect 8764 33068 9380 33070
rect 8764 32004 8820 33068
rect 9324 33058 9380 33068
rect 8764 31938 8820 31948
rect 9100 32788 9156 32798
rect 8540 31838 8542 31890
rect 8594 31838 8596 31890
rect 8540 31826 8596 31838
rect 8540 31220 8596 31230
rect 9100 31220 9156 32732
rect 8540 31218 9156 31220
rect 8540 31166 8542 31218
rect 8594 31166 9102 31218
rect 9154 31166 9156 31218
rect 8540 31164 9156 31166
rect 8540 31154 8596 31164
rect 9100 31154 9156 31164
rect 9660 32004 9716 32014
rect 9660 31218 9716 31948
rect 10556 31892 10612 33294
rect 11452 33234 11508 34076
rect 11564 34130 11620 34412
rect 11564 34078 11566 34130
rect 11618 34078 11620 34130
rect 11564 34066 11620 34078
rect 11676 34132 11732 34748
rect 12684 34802 12740 34814
rect 12684 34750 12686 34802
rect 12738 34750 12740 34802
rect 11788 34692 11844 34702
rect 11788 34598 11844 34636
rect 12012 34132 12068 34142
rect 11676 34130 12068 34132
rect 11676 34078 12014 34130
rect 12066 34078 12068 34130
rect 11676 34076 12068 34078
rect 12012 34066 12068 34076
rect 12012 33908 12068 33918
rect 12012 33906 12180 33908
rect 12012 33854 12014 33906
rect 12066 33854 12180 33906
rect 12012 33852 12180 33854
rect 12012 33842 12068 33852
rect 12124 33460 12180 33852
rect 12684 33570 12740 34750
rect 12796 34690 12852 34702
rect 12796 34638 12798 34690
rect 12850 34638 12852 34690
rect 12796 34132 12852 34638
rect 12796 34066 12852 34076
rect 12684 33518 12686 33570
rect 12738 33518 12740 33570
rect 12684 33506 12740 33518
rect 12124 33458 12628 33460
rect 12124 33406 12126 33458
rect 12178 33406 12628 33458
rect 12124 33404 12628 33406
rect 12124 33394 12180 33404
rect 11452 33182 11454 33234
rect 11506 33182 11508 33234
rect 11452 33170 11508 33182
rect 11676 33346 11732 33358
rect 11676 33294 11678 33346
rect 11730 33294 11732 33346
rect 11116 33122 11172 33134
rect 11116 33070 11118 33122
rect 11170 33070 11172 33122
rect 10892 32450 10948 32462
rect 10892 32398 10894 32450
rect 10946 32398 10948 32450
rect 10892 32004 10948 32398
rect 10892 31938 10948 31948
rect 10556 31826 10612 31836
rect 10668 31892 10724 31902
rect 10668 31890 10836 31892
rect 10668 31838 10670 31890
rect 10722 31838 10836 31890
rect 10668 31836 10836 31838
rect 10668 31826 10724 31836
rect 10780 31780 10836 31836
rect 11004 31780 11060 31790
rect 10780 31778 11060 31780
rect 10780 31726 11006 31778
rect 11058 31726 11060 31778
rect 10780 31724 11060 31726
rect 10556 31444 10612 31454
rect 9660 31166 9662 31218
rect 9714 31166 9716 31218
rect 9660 31154 9716 31166
rect 10332 31220 10388 31230
rect 10332 31126 10388 31164
rect 10556 31106 10612 31388
rect 10556 31054 10558 31106
rect 10610 31054 10612 31106
rect 10556 31042 10612 31054
rect 10892 30994 10948 31724
rect 11004 31714 11060 31724
rect 11116 31444 11172 33070
rect 11116 31378 11172 31388
rect 11228 32004 11284 32014
rect 11676 31948 11732 33294
rect 12572 33236 12628 33404
rect 12684 33236 12740 33246
rect 12572 33234 12740 33236
rect 12572 33182 12686 33234
rect 12738 33182 12740 33234
rect 12572 33180 12740 33182
rect 12684 33170 12740 33180
rect 12796 33234 12852 33246
rect 12796 33182 12798 33234
rect 12850 33182 12852 33234
rect 12236 33122 12292 33134
rect 12236 33070 12238 33122
rect 12290 33070 12292 33122
rect 10892 30942 10894 30994
rect 10946 30942 10948 30994
rect 10892 30930 10948 30942
rect 11116 30996 11172 31006
rect 8316 30158 8318 30210
rect 8370 30158 8372 30210
rect 8316 30146 8372 30158
rect 8988 30884 9044 30894
rect 8988 30210 9044 30828
rect 10220 30772 10276 30782
rect 10220 30678 10276 30716
rect 9212 30324 9268 30334
rect 8988 30158 8990 30210
rect 9042 30158 9044 30210
rect 8988 30146 9044 30158
rect 9100 30268 9212 30324
rect 7084 29986 8260 29988
rect 7084 29934 7086 29986
rect 7138 29934 8260 29986
rect 7084 29932 8260 29934
rect 6188 29426 6244 29438
rect 6188 29374 6190 29426
rect 6242 29374 6244 29426
rect 5180 29316 5236 29326
rect 5068 29260 5180 29316
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 5068 28532 5124 29260
rect 5180 29250 5236 29260
rect 6188 29316 6244 29374
rect 6188 29250 6244 29260
rect 6748 29316 6804 29326
rect 6524 29092 6580 29102
rect 6524 28642 6580 29036
rect 6524 28590 6526 28642
rect 6578 28590 6580 28642
rect 6524 28578 6580 28590
rect 4956 28476 5124 28532
rect 4956 27858 5012 28476
rect 6188 28420 6244 28430
rect 4956 27806 4958 27858
rect 5010 27806 5012 27858
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 3500 26292 3556 26302
rect 3500 26198 3556 26236
rect 4956 26292 5012 27806
rect 5852 28418 6244 28420
rect 5852 28366 6190 28418
rect 6242 28366 6244 28418
rect 5852 28364 6244 28366
rect 5628 27748 5684 27758
rect 5628 27746 5796 27748
rect 5628 27694 5630 27746
rect 5682 27694 5796 27746
rect 5628 27692 5796 27694
rect 5628 27682 5684 27692
rect 5740 27298 5796 27692
rect 5740 27246 5742 27298
rect 5794 27246 5796 27298
rect 5740 27234 5796 27246
rect 5852 26962 5908 28364
rect 6188 28354 6244 28364
rect 6524 27412 6580 27422
rect 6076 27188 6132 27198
rect 6524 27188 6580 27356
rect 6076 27186 6580 27188
rect 6076 27134 6078 27186
rect 6130 27134 6526 27186
rect 6578 27134 6580 27186
rect 6076 27132 6580 27134
rect 6076 27122 6132 27132
rect 6524 27122 6580 27132
rect 5852 26910 5854 26962
rect 5906 26910 5908 26962
rect 5852 26908 5908 26910
rect 4956 26226 5012 26236
rect 5740 26852 5908 26908
rect 4172 26180 4228 26190
rect 4172 26086 4228 26124
rect 5628 26180 5684 26190
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 5628 25730 5684 26124
rect 5628 25678 5630 25730
rect 5682 25678 5684 25730
rect 5628 25666 5684 25678
rect 5628 25508 5684 25518
rect 5740 25508 5796 26852
rect 5964 26180 6020 26190
rect 5964 25732 6020 26124
rect 5628 25506 5796 25508
rect 5628 25454 5630 25506
rect 5682 25454 5796 25506
rect 5628 25452 5796 25454
rect 5852 25730 6020 25732
rect 5852 25678 5966 25730
rect 6018 25678 6020 25730
rect 5852 25676 6020 25678
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 5628 23938 5684 25452
rect 5852 23940 5908 25676
rect 5964 25666 6020 25676
rect 6300 26178 6356 26190
rect 6300 26126 6302 26178
rect 6354 26126 6356 26178
rect 6300 25508 6356 26126
rect 6300 25442 6356 25452
rect 6748 26178 6804 29260
rect 6972 29092 7028 29102
rect 6972 28754 7028 29036
rect 6972 28702 6974 28754
rect 7026 28702 7028 28754
rect 6972 28690 7028 28702
rect 7084 26908 7140 29932
rect 8204 29316 8260 29326
rect 8204 28082 8260 29260
rect 8988 29316 9044 29326
rect 9100 29316 9156 30268
rect 9212 30258 9268 30268
rect 11116 30322 11172 30940
rect 11116 30270 11118 30322
rect 11170 30270 11172 30322
rect 11116 30258 11172 30270
rect 11228 29650 11284 31948
rect 11452 31892 11732 31948
rect 12012 32004 12068 32014
rect 11340 31332 11396 31342
rect 11340 30994 11396 31276
rect 11340 30942 11342 30994
rect 11394 30942 11396 30994
rect 11340 30930 11396 30942
rect 11452 30324 11508 31836
rect 11564 31780 11620 31790
rect 12012 31780 12068 31948
rect 11564 31778 12068 31780
rect 11564 31726 11566 31778
rect 11618 31726 12014 31778
rect 12066 31726 12068 31778
rect 11564 31724 12068 31726
rect 11564 31714 11620 31724
rect 12012 31714 12068 31724
rect 12236 31780 12292 33070
rect 12236 31714 12292 31724
rect 12460 31778 12516 31790
rect 12460 31726 12462 31778
rect 12514 31726 12516 31778
rect 12460 31220 12516 31726
rect 12460 31154 12516 31164
rect 12012 30996 12068 31006
rect 12012 30902 12068 30940
rect 12572 30996 12628 31006
rect 12572 30902 12628 30940
rect 11788 30772 11844 30782
rect 12348 30772 12404 30782
rect 11788 30770 12292 30772
rect 11788 30718 11790 30770
rect 11842 30718 12292 30770
rect 11788 30716 12292 30718
rect 11788 30706 11844 30716
rect 12236 30434 12292 30716
rect 12236 30382 12238 30434
rect 12290 30382 12292 30434
rect 12236 30370 12292 30382
rect 12348 30434 12404 30716
rect 12796 30660 12852 33182
rect 12796 30594 12852 30604
rect 12572 30436 12628 30446
rect 12908 30436 12964 36428
rect 13020 36260 13076 36270
rect 13468 36260 13524 36270
rect 13020 36258 13412 36260
rect 13020 36206 13022 36258
rect 13074 36206 13412 36258
rect 13020 36204 13412 36206
rect 13020 36194 13076 36204
rect 13356 35140 13412 36204
rect 13468 36258 13748 36260
rect 13468 36206 13470 36258
rect 13522 36206 13748 36258
rect 13468 36204 13748 36206
rect 13468 36194 13524 36204
rect 13468 35700 13524 35710
rect 13468 35606 13524 35644
rect 13580 35140 13636 35150
rect 13356 35138 13636 35140
rect 13356 35086 13582 35138
rect 13634 35086 13636 35138
rect 13356 35084 13636 35086
rect 13580 35074 13636 35084
rect 13468 34690 13524 34702
rect 13468 34638 13470 34690
rect 13522 34638 13524 34690
rect 13468 34580 13524 34638
rect 13468 34514 13524 34524
rect 13580 34468 13636 34478
rect 13468 34356 13524 34366
rect 13468 34262 13524 34300
rect 13020 34130 13076 34142
rect 13020 34078 13022 34130
rect 13074 34078 13076 34130
rect 13020 31780 13076 34078
rect 13020 31714 13076 31724
rect 13244 34132 13300 34142
rect 12348 30382 12350 30434
rect 12402 30382 12404 30434
rect 12348 30370 12404 30382
rect 12460 30434 12964 30436
rect 12460 30382 12574 30434
rect 12626 30382 12964 30434
rect 12460 30380 12964 30382
rect 11452 30258 11508 30268
rect 11788 30212 11844 30222
rect 12460 30212 12516 30380
rect 12572 30370 12628 30380
rect 11788 30210 12516 30212
rect 11788 30158 11790 30210
rect 11842 30158 12516 30210
rect 11788 30156 12516 30158
rect 12796 30212 12852 30222
rect 11788 30146 11844 30156
rect 11228 29598 11230 29650
rect 11282 29598 11284 29650
rect 11228 29586 11284 29598
rect 11564 30100 11620 30110
rect 8988 29314 9156 29316
rect 8988 29262 8990 29314
rect 9042 29262 9156 29314
rect 8988 29260 9156 29262
rect 9772 29316 9828 29326
rect 8988 29250 9044 29260
rect 9772 29222 9828 29260
rect 11564 29314 11620 30044
rect 12684 29986 12740 29998
rect 12684 29934 12686 29986
rect 12738 29934 12740 29986
rect 12012 29652 12068 29662
rect 12012 29558 12068 29596
rect 12684 29426 12740 29934
rect 12684 29374 12686 29426
rect 12738 29374 12740 29426
rect 12684 29362 12740 29374
rect 12796 29428 12852 30156
rect 12796 29362 12852 29372
rect 11564 29262 11566 29314
rect 11618 29262 11620 29314
rect 11564 29250 11620 29262
rect 12460 29204 12516 29214
rect 12460 29110 12516 29148
rect 8204 28030 8206 28082
rect 8258 28030 8260 28082
rect 8204 28018 8260 28030
rect 12908 28084 12964 30380
rect 12908 28018 12964 28028
rect 13132 30548 13188 30558
rect 13132 29538 13188 30492
rect 13132 29486 13134 29538
rect 13186 29486 13188 29538
rect 9660 27972 9716 27982
rect 7756 27860 7812 27870
rect 7756 27746 7812 27804
rect 7756 27694 7758 27746
rect 7810 27694 7812 27746
rect 7756 27682 7812 27694
rect 8428 27860 8484 27870
rect 7980 27636 8036 27646
rect 7980 27074 8036 27580
rect 7980 27022 7982 27074
rect 8034 27022 8036 27074
rect 7980 27010 8036 27022
rect 7644 26964 7700 27002
rect 6748 26126 6750 26178
rect 6802 26126 6804 26178
rect 5628 23886 5630 23938
rect 5682 23886 5684 23938
rect 3948 23716 4004 23726
rect 3948 23266 4004 23660
rect 3948 23214 3950 23266
rect 4002 23214 4004 23266
rect 3948 23202 4004 23214
rect 3276 23156 3332 23166
rect 3276 23062 3332 23100
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 5628 21586 5684 23886
rect 5740 23884 5908 23940
rect 5740 23380 5796 23884
rect 5964 23826 6020 23838
rect 5964 23774 5966 23826
rect 6018 23774 6020 23826
rect 5852 23716 5908 23726
rect 5852 23622 5908 23660
rect 5964 23380 6020 23774
rect 6524 23492 6580 23502
rect 5740 23324 5908 23380
rect 5740 23156 5796 23166
rect 5740 22484 5796 23100
rect 5740 22370 5796 22428
rect 5740 22318 5742 22370
rect 5794 22318 5796 22370
rect 5740 22306 5796 22318
rect 5852 22148 5908 23324
rect 5964 23314 6020 23324
rect 6412 23436 6524 23492
rect 6076 23044 6132 23054
rect 6076 22950 6132 22988
rect 6412 22484 6468 23436
rect 6524 23426 6580 23436
rect 6524 23044 6580 23054
rect 6748 23044 6804 26126
rect 6524 23042 6804 23044
rect 6524 22990 6526 23042
rect 6578 22990 6804 23042
rect 6524 22988 6804 22990
rect 6524 22978 6580 22988
rect 6748 22484 6804 22988
rect 6412 22428 6580 22484
rect 5628 21534 5630 21586
rect 5682 21534 5684 21586
rect 5628 21522 5684 21534
rect 5740 22092 5908 22148
rect 6412 22258 6468 22270
rect 6412 22206 6414 22258
rect 6466 22206 6468 22258
rect 5740 21364 5796 22092
rect 6412 22036 6468 22206
rect 5852 21980 6468 22036
rect 5852 21810 5908 21980
rect 5852 21758 5854 21810
rect 5906 21758 5908 21810
rect 5852 21746 5908 21758
rect 6076 21698 6132 21710
rect 6076 21646 6078 21698
rect 6130 21646 6132 21698
rect 5964 21588 6020 21598
rect 6076 21588 6132 21646
rect 6412 21700 6468 21710
rect 6524 21700 6580 22428
rect 6748 22418 6804 22428
rect 6860 26852 7140 26908
rect 7532 26852 7700 26908
rect 6748 21812 6804 21822
rect 6860 21812 6916 26852
rect 7196 26516 7252 26526
rect 7196 26514 7476 26516
rect 7196 26462 7198 26514
rect 7250 26462 7476 26514
rect 7196 26460 7476 26462
rect 7196 26450 7252 26460
rect 7308 26292 7364 26302
rect 7308 26198 7364 26236
rect 6972 26068 7028 26078
rect 6972 23826 7028 26012
rect 7196 26066 7252 26078
rect 7196 26014 7198 26066
rect 7250 26014 7252 26066
rect 7196 25618 7252 26014
rect 7196 25566 7198 25618
rect 7250 25566 7252 25618
rect 7196 25554 7252 25566
rect 7308 25508 7364 25518
rect 7308 25414 7364 25452
rect 7420 25396 7476 26460
rect 7420 25330 7476 25340
rect 7532 24388 7588 26852
rect 7756 26292 7812 26302
rect 7644 25620 7700 25630
rect 7644 25526 7700 25564
rect 7644 25060 7700 25070
rect 7756 25060 7812 26236
rect 8428 26290 8484 27804
rect 9548 27636 9604 27646
rect 9436 27634 9604 27636
rect 9436 27582 9550 27634
rect 9602 27582 9604 27634
rect 9436 27580 9604 27582
rect 8876 27074 8932 27086
rect 8876 27022 8878 27074
rect 8930 27022 8932 27074
rect 8540 26964 8596 27002
rect 8540 26898 8596 26908
rect 8876 26402 8932 27022
rect 9324 26962 9380 26974
rect 9324 26910 9326 26962
rect 9378 26910 9380 26962
rect 9324 26908 9380 26910
rect 8876 26350 8878 26402
rect 8930 26350 8932 26402
rect 8876 26338 8932 26350
rect 9212 26852 9380 26908
rect 8428 26238 8430 26290
rect 8482 26238 8484 26290
rect 7700 25004 7812 25060
rect 7980 25396 8036 25406
rect 7644 24610 7700 25004
rect 7868 24836 7924 24846
rect 7980 24836 8036 25340
rect 8428 24948 8484 26238
rect 8764 26292 8820 26302
rect 8764 26198 8820 26236
rect 8764 25396 8820 25406
rect 8764 25302 8820 25340
rect 8428 24882 8484 24892
rect 9212 24948 9268 26852
rect 9436 26292 9492 27580
rect 9548 27570 9604 27580
rect 9548 27412 9604 27422
rect 9548 27186 9604 27356
rect 9548 27134 9550 27186
rect 9602 27134 9604 27186
rect 9548 27122 9604 27134
rect 9660 27074 9716 27916
rect 10220 27972 10276 27982
rect 9884 27860 9940 27898
rect 10220 27878 10276 27916
rect 9884 27794 9940 27804
rect 10556 27860 10612 27870
rect 13132 27860 13188 29486
rect 10556 27766 10612 27804
rect 12460 27858 13188 27860
rect 12460 27806 13134 27858
rect 13186 27806 13188 27858
rect 12460 27804 13188 27806
rect 9884 27636 9940 27646
rect 9884 27634 10276 27636
rect 9884 27582 9886 27634
rect 9938 27582 10276 27634
rect 9884 27580 10276 27582
rect 9884 27570 9940 27580
rect 10220 27186 10276 27580
rect 11228 27244 11620 27300
rect 11228 27188 11284 27244
rect 10220 27134 10222 27186
rect 10274 27134 10276 27186
rect 10220 27122 10276 27134
rect 10892 27132 11284 27188
rect 9660 27022 9662 27074
rect 9714 27022 9716 27074
rect 9660 26908 9716 27022
rect 10444 27074 10500 27086
rect 10444 27022 10446 27074
rect 10498 27022 10500 27074
rect 9436 26226 9492 26236
rect 9548 26852 9716 26908
rect 9996 26964 10052 26974
rect 9548 26290 9604 26852
rect 9996 26514 10052 26908
rect 9996 26462 9998 26514
rect 10050 26462 10052 26514
rect 9996 26450 10052 26462
rect 9548 26238 9550 26290
rect 9602 26238 9604 26290
rect 9548 26068 9604 26238
rect 9772 26290 9828 26302
rect 9772 26238 9774 26290
rect 9826 26238 9828 26290
rect 9660 26180 9716 26190
rect 9660 26086 9716 26124
rect 9548 26002 9604 26012
rect 9772 25844 9828 26238
rect 9324 25788 9828 25844
rect 10108 26292 10164 26302
rect 9324 25508 9380 25788
rect 9324 25394 9380 25452
rect 9324 25342 9326 25394
rect 9378 25342 9380 25394
rect 9324 25330 9380 25342
rect 9548 25506 9604 25518
rect 9548 25454 9550 25506
rect 9602 25454 9604 25506
rect 9548 25060 9604 25454
rect 9548 24994 9604 25004
rect 9660 25394 9716 25406
rect 9660 25342 9662 25394
rect 9714 25342 9716 25394
rect 9212 24882 9268 24892
rect 7868 24834 8036 24836
rect 7868 24782 7870 24834
rect 7922 24782 8036 24834
rect 7868 24780 8036 24782
rect 7868 24770 7924 24780
rect 7644 24558 7646 24610
rect 7698 24558 7700 24610
rect 7644 24546 7700 24558
rect 7308 24332 7588 24388
rect 7308 23940 7364 24332
rect 7308 23938 7476 23940
rect 7308 23886 7310 23938
rect 7362 23886 7476 23938
rect 7308 23884 7476 23886
rect 7308 23874 7364 23884
rect 6972 23774 6974 23826
rect 7026 23774 7028 23826
rect 6972 23380 7028 23774
rect 7084 23828 7140 23838
rect 7084 23734 7140 23772
rect 7196 23716 7252 23726
rect 7196 23714 7364 23716
rect 7196 23662 7198 23714
rect 7250 23662 7364 23714
rect 7196 23660 7364 23662
rect 7196 23650 7252 23660
rect 7308 23604 7364 23660
rect 7420 23604 7476 23884
rect 7532 23828 7588 23838
rect 7868 23828 7924 23838
rect 7532 23826 7924 23828
rect 7532 23774 7534 23826
rect 7586 23774 7870 23826
rect 7922 23774 7924 23826
rect 7532 23772 7924 23774
rect 7532 23762 7588 23772
rect 7420 23548 7700 23604
rect 7308 23538 7364 23548
rect 7308 23380 7364 23390
rect 6972 23378 7364 23380
rect 6972 23326 7310 23378
rect 7362 23326 7364 23378
rect 6972 23324 7364 23326
rect 7308 23314 7364 23324
rect 7532 23380 7588 23390
rect 7420 23268 7476 23278
rect 7420 23154 7476 23212
rect 7420 23102 7422 23154
rect 7474 23102 7476 23154
rect 7420 23044 7476 23102
rect 7420 22978 7476 22988
rect 7308 21812 7364 21822
rect 6412 21698 6580 21700
rect 6412 21646 6414 21698
rect 6466 21646 6526 21698
rect 6578 21646 6580 21698
rect 6412 21644 6580 21646
rect 6412 21634 6468 21644
rect 6524 21634 6580 21644
rect 6636 21810 7364 21812
rect 6636 21758 6750 21810
rect 6802 21758 7310 21810
rect 7362 21758 7364 21810
rect 6636 21756 7364 21758
rect 5964 21586 6132 21588
rect 5964 21534 5966 21586
rect 6018 21534 6132 21586
rect 5964 21532 6132 21534
rect 5964 21522 6020 21532
rect 5740 21308 6356 21364
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 6300 21026 6356 21308
rect 6300 20974 6302 21026
rect 6354 20974 6356 21026
rect 6300 20962 6356 20974
rect 6636 20802 6692 21756
rect 6748 21746 6804 21756
rect 7308 21746 7364 21756
rect 7532 21698 7588 23324
rect 7644 23378 7700 23548
rect 7868 23492 7924 23772
rect 7868 23426 7924 23436
rect 7644 23326 7646 23378
rect 7698 23326 7700 23378
rect 7644 23314 7700 23326
rect 7980 23380 8036 24780
rect 9660 24612 9716 25342
rect 10108 24836 10164 26236
rect 10220 26290 10276 26302
rect 10220 26238 10222 26290
rect 10274 26238 10276 26290
rect 10220 25620 10276 26238
rect 10332 25620 10388 25630
rect 10220 25564 10332 25620
rect 10332 25526 10388 25564
rect 10332 24836 10388 24846
rect 10108 24780 10332 24836
rect 10332 24742 10388 24780
rect 8764 24610 9716 24612
rect 8764 24558 9662 24610
rect 9714 24558 9716 24610
rect 8764 24556 9716 24558
rect 8652 24500 8708 24510
rect 7980 23314 8036 23324
rect 8316 24444 8652 24500
rect 8316 23266 8372 24444
rect 8652 24406 8708 24444
rect 8540 24164 8596 24174
rect 8540 23938 8596 24108
rect 8764 24050 8820 24556
rect 9660 24546 9716 24556
rect 9772 24722 9828 24734
rect 9772 24670 9774 24722
rect 9826 24670 9828 24722
rect 9772 24276 9828 24670
rect 9324 24220 9828 24276
rect 9324 24164 9380 24220
rect 9324 24070 9380 24108
rect 8764 23998 8766 24050
rect 8818 23998 8820 24050
rect 8764 23986 8820 23998
rect 8540 23886 8542 23938
rect 8594 23886 8596 23938
rect 8540 23874 8596 23886
rect 10108 23940 10164 23950
rect 10108 23938 10276 23940
rect 10108 23886 10110 23938
rect 10162 23886 10276 23938
rect 10108 23884 10276 23886
rect 10108 23874 10164 23884
rect 8316 23214 8318 23266
rect 8370 23214 8372 23266
rect 8316 23202 8372 23214
rect 8428 23828 8484 23838
rect 7868 23156 7924 23166
rect 8204 23156 8260 23166
rect 7868 23154 8260 23156
rect 7868 23102 7870 23154
rect 7922 23102 8206 23154
rect 8258 23102 8260 23154
rect 7868 23100 8260 23102
rect 7868 23090 7924 23100
rect 8204 23090 8260 23100
rect 7532 21646 7534 21698
rect 7586 21646 7588 21698
rect 7532 21634 7588 21646
rect 7980 22484 8036 22494
rect 8428 22484 8484 23772
rect 9212 23828 9268 23838
rect 9212 23734 9268 23772
rect 10108 23154 10164 23166
rect 10108 23102 10110 23154
rect 10162 23102 10164 23154
rect 8540 22484 8596 22494
rect 8428 22482 8596 22484
rect 8428 22430 8542 22482
rect 8594 22430 8596 22482
rect 8428 22428 8596 22430
rect 6636 20750 6638 20802
rect 6690 20750 6692 20802
rect 6636 20738 6692 20750
rect 6748 21532 7252 21588
rect 6412 20578 6468 20590
rect 6412 20526 6414 20578
rect 6466 20526 6468 20578
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 6076 18452 6132 18462
rect 6076 18358 6132 18396
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 6076 15314 6132 15326
rect 6076 15262 6078 15314
rect 6130 15262 6132 15314
rect 6076 15204 6132 15262
rect 5964 15148 6076 15204
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 5740 13748 5796 13758
rect 5964 13748 6020 15148
rect 6076 15138 6132 15148
rect 6412 13858 6468 20526
rect 6748 18450 6804 21532
rect 7196 21474 7252 21532
rect 7196 21422 7198 21474
rect 7250 21422 7252 21474
rect 7196 21410 7252 21422
rect 6748 18398 6750 18450
rect 6802 18398 6804 18450
rect 6748 18386 6804 18398
rect 6860 21362 6916 21374
rect 6860 21310 6862 21362
rect 6914 21310 6916 21362
rect 6748 15428 6804 15438
rect 6860 15428 6916 21310
rect 7980 20804 8036 22428
rect 8540 22418 8596 22428
rect 8988 22484 9044 22494
rect 8988 22390 9044 22428
rect 10108 21588 10164 23102
rect 10220 22484 10276 23884
rect 10332 23492 10388 23502
rect 10332 23042 10388 23436
rect 10444 23380 10500 27022
rect 10892 26290 10948 27132
rect 11116 26964 11172 27002
rect 11116 26898 11172 26908
rect 10892 26238 10894 26290
rect 10946 26238 10948 26290
rect 10892 26226 10948 26238
rect 11228 25618 11284 27132
rect 11452 27074 11508 27086
rect 11452 27022 11454 27074
rect 11506 27022 11508 27074
rect 11452 26908 11508 27022
rect 11228 25566 11230 25618
rect 11282 25566 11284 25618
rect 11228 25554 11284 25566
rect 11340 26852 11508 26908
rect 11564 26962 11620 27244
rect 12460 27298 12516 27804
rect 13132 27794 13188 27804
rect 13244 28644 13300 34076
rect 13580 34130 13636 34412
rect 13580 34078 13582 34130
rect 13634 34078 13636 34130
rect 13580 34066 13636 34078
rect 13356 34018 13412 34030
rect 13356 33966 13358 34018
rect 13410 33966 13412 34018
rect 13356 33348 13412 33966
rect 13692 33572 13748 36204
rect 13804 35700 13860 36652
rect 14028 36484 14084 36494
rect 14028 36390 14084 36428
rect 14140 36482 14196 36652
rect 14140 36430 14142 36482
rect 14194 36430 14196 36482
rect 14140 36418 14196 36430
rect 13916 36370 13972 36382
rect 13916 36318 13918 36370
rect 13970 36318 13972 36370
rect 13916 36260 13972 36318
rect 13916 36194 13972 36204
rect 14140 36260 14196 36270
rect 13804 35634 13860 35644
rect 13916 35588 13972 35598
rect 13804 35252 13860 35262
rect 13804 35138 13860 35196
rect 13804 35086 13806 35138
rect 13858 35086 13860 35138
rect 13804 35074 13860 35086
rect 13916 33908 13972 35532
rect 14028 34692 14084 34702
rect 14028 34130 14084 34636
rect 14028 34078 14030 34130
rect 14082 34078 14084 34130
rect 14028 34066 14084 34078
rect 14140 34132 14196 36204
rect 14252 35252 14308 37774
rect 14364 36372 14420 37998
rect 14476 36820 14532 36830
rect 14476 36706 14532 36764
rect 14476 36654 14478 36706
rect 14530 36654 14532 36706
rect 14476 36642 14532 36654
rect 14588 36484 14644 38444
rect 15036 38276 15092 38286
rect 14924 37828 14980 37838
rect 14812 37826 14980 37828
rect 14812 37774 14926 37826
rect 14978 37774 14980 37826
rect 14812 37772 14980 37774
rect 14812 37268 14868 37772
rect 14924 37762 14980 37772
rect 14812 37202 14868 37212
rect 14924 37266 14980 37278
rect 14924 37214 14926 37266
rect 14978 37214 14980 37266
rect 14364 36306 14420 36316
rect 14476 36428 14644 36484
rect 14700 37044 14756 37054
rect 14252 35186 14308 35196
rect 14476 35140 14532 36428
rect 14588 36260 14644 36270
rect 14588 36166 14644 36204
rect 14700 35924 14756 36988
rect 14924 36708 14980 37214
rect 15036 37154 15092 38220
rect 15036 37102 15038 37154
rect 15090 37102 15092 37154
rect 15036 37090 15092 37102
rect 15260 37826 15316 38892
rect 15372 38882 15428 38892
rect 15484 38834 15540 38846
rect 15484 38782 15486 38834
rect 15538 38782 15540 38834
rect 15260 37774 15262 37826
rect 15314 37774 15316 37826
rect 15036 36708 15092 36718
rect 14924 36652 15036 36708
rect 15036 36642 15092 36652
rect 14812 36484 14868 36494
rect 14812 36390 14868 36428
rect 15036 36370 15092 36382
rect 15036 36318 15038 36370
rect 15090 36318 15092 36370
rect 14700 35810 14756 35868
rect 14924 36036 14980 36046
rect 14924 35924 14980 35980
rect 15036 35924 15092 36318
rect 14924 35868 15092 35924
rect 15148 36372 15204 36382
rect 14700 35758 14702 35810
rect 14754 35758 14756 35810
rect 14700 35746 14756 35758
rect 14812 35812 14868 35822
rect 14812 35718 14868 35756
rect 14364 35084 14532 35140
rect 14364 35028 14420 35084
rect 14252 34972 14420 35028
rect 14252 34914 14308 34972
rect 14252 34862 14254 34914
rect 14306 34862 14308 34914
rect 14252 34468 14308 34862
rect 14364 34802 14420 34814
rect 14364 34750 14366 34802
rect 14418 34750 14420 34802
rect 14364 34692 14420 34750
rect 14812 34692 14868 34702
rect 14364 34690 14868 34692
rect 14364 34638 14814 34690
rect 14866 34638 14868 34690
rect 14364 34636 14868 34638
rect 14252 34402 14308 34412
rect 14588 34468 14644 34478
rect 14588 34354 14644 34412
rect 14588 34302 14590 34354
rect 14642 34302 14644 34354
rect 14588 34290 14644 34302
rect 14700 34132 14756 34142
rect 14140 34076 14420 34132
rect 14252 33908 14308 33918
rect 13916 33906 14308 33908
rect 13916 33854 14254 33906
rect 14306 33854 14308 33906
rect 13916 33852 14308 33854
rect 13692 33516 13860 33572
rect 13692 33348 13748 33358
rect 13356 33346 13748 33348
rect 13356 33294 13694 33346
rect 13746 33294 13748 33346
rect 13356 33292 13748 33294
rect 13692 33282 13748 33292
rect 13804 32676 13860 33516
rect 13916 33124 13972 33134
rect 13916 33030 13972 33068
rect 13580 32620 13860 32676
rect 13916 32788 13972 32798
rect 13468 31780 13524 31790
rect 13468 31686 13524 31724
rect 13580 30436 13636 32620
rect 13804 32452 13860 32462
rect 13916 32452 13972 32732
rect 13804 32450 13972 32452
rect 13804 32398 13806 32450
rect 13858 32398 13972 32450
rect 13804 32396 13972 32398
rect 13804 32386 13860 32396
rect 14028 31668 14084 33852
rect 14252 33842 14308 33852
rect 14364 33460 14420 34076
rect 14700 33460 14756 34076
rect 14812 33908 14868 34636
rect 14812 33842 14868 33852
rect 14812 33460 14868 33470
rect 14252 33404 14420 33460
rect 14476 33458 14868 33460
rect 14476 33406 14814 33458
rect 14866 33406 14868 33458
rect 14476 33404 14868 33406
rect 14140 33348 14196 33358
rect 14140 33254 14196 33292
rect 14140 32338 14196 32350
rect 14140 32286 14142 32338
rect 14194 32286 14196 32338
rect 14140 31778 14196 32286
rect 14140 31726 14142 31778
rect 14194 31726 14196 31778
rect 14140 31714 14196 31726
rect 14028 31602 14084 31612
rect 13692 31554 13748 31566
rect 13692 31502 13694 31554
rect 13746 31502 13748 31554
rect 13692 30548 13748 31502
rect 13804 31554 13860 31566
rect 13804 31502 13806 31554
rect 13858 31502 13860 31554
rect 13804 30994 13860 31502
rect 13804 30942 13806 30994
rect 13858 30942 13860 30994
rect 13804 30930 13860 30942
rect 13916 31556 13972 31566
rect 13916 30996 13972 31500
rect 14252 31220 14308 33404
rect 14364 33236 14420 33246
rect 14476 33236 14532 33404
rect 14812 33394 14868 33404
rect 14364 33234 14532 33236
rect 14364 33182 14366 33234
rect 14418 33182 14532 33234
rect 14364 33180 14532 33182
rect 14364 33170 14420 33180
rect 14700 33012 14756 33022
rect 14364 32788 14420 32798
rect 14700 32788 14756 32956
rect 14364 32786 14756 32788
rect 14364 32734 14366 32786
rect 14418 32734 14756 32786
rect 14364 32732 14756 32734
rect 14364 32722 14420 32732
rect 14700 32674 14756 32732
rect 14700 32622 14702 32674
rect 14754 32622 14756 32674
rect 14700 32610 14756 32622
rect 14924 32452 14980 35868
rect 15036 35698 15092 35710
rect 15036 35646 15038 35698
rect 15090 35646 15092 35698
rect 15036 34242 15092 35646
rect 15148 34354 15204 36316
rect 15260 35140 15316 37774
rect 15372 38610 15428 38622
rect 15372 38558 15374 38610
rect 15426 38558 15428 38610
rect 15372 36932 15428 38558
rect 15484 38388 15540 38782
rect 16156 38668 16212 39676
rect 15484 38322 15540 38332
rect 16044 38612 16212 38668
rect 15708 38164 15764 38174
rect 15708 38070 15764 38108
rect 15820 38050 15876 38062
rect 15820 37998 15822 38050
rect 15874 37998 15876 38050
rect 15820 37604 15876 37998
rect 15372 36866 15428 36876
rect 15484 37548 15876 37604
rect 16044 37938 16100 38612
rect 16044 37886 16046 37938
rect 16098 37886 16100 37938
rect 15484 36706 15540 37548
rect 15932 37492 15988 37502
rect 15932 37266 15988 37436
rect 15932 37214 15934 37266
rect 15986 37214 15988 37266
rect 15932 37202 15988 37214
rect 15708 37154 15764 37166
rect 15708 37102 15710 37154
rect 15762 37102 15764 37154
rect 15596 37044 15652 37054
rect 15596 36950 15652 36988
rect 15484 36654 15486 36706
rect 15538 36654 15540 36706
rect 15484 36642 15540 36654
rect 15372 36484 15428 36494
rect 15708 36484 15764 37102
rect 15372 36482 15764 36484
rect 15372 36430 15374 36482
rect 15426 36430 15764 36482
rect 15372 36428 15764 36430
rect 15372 36418 15428 36428
rect 15708 36036 15764 36428
rect 16044 36482 16100 37886
rect 16268 37380 16324 40012
rect 16604 39732 16660 42476
rect 16716 41300 16772 42924
rect 17052 42868 17108 43596
rect 17388 43204 17444 44158
rect 18060 43988 18116 44940
rect 18060 43922 18116 43932
rect 18172 44212 18228 44222
rect 17836 43652 17892 43662
rect 17836 43540 17892 43596
rect 18060 43652 18116 43662
rect 18172 43652 18228 44156
rect 18060 43650 18228 43652
rect 18060 43598 18062 43650
rect 18114 43598 18228 43650
rect 18060 43596 18228 43598
rect 18396 43652 18452 50372
rect 19068 50034 19124 51212
rect 19180 51202 19236 51212
rect 19292 50482 19348 50494
rect 19292 50430 19294 50482
rect 19346 50430 19348 50482
rect 19292 50428 19348 50430
rect 19068 49982 19070 50034
rect 19122 49982 19124 50034
rect 19068 49970 19124 49982
rect 19180 50372 19348 50428
rect 19516 50484 19572 50494
rect 18732 49810 18788 49822
rect 18732 49758 18734 49810
rect 18786 49758 18788 49810
rect 18732 49588 18788 49758
rect 18956 49812 19012 49822
rect 18956 49718 19012 49756
rect 19180 49810 19236 50372
rect 19180 49758 19182 49810
rect 19234 49758 19236 49810
rect 19180 49746 19236 49758
rect 19516 49922 19572 50428
rect 19628 50372 19684 52108
rect 19740 52070 19796 52108
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19964 51268 20020 51278
rect 19964 51174 20020 51212
rect 19964 50932 20020 50942
rect 19964 50594 20020 50876
rect 19964 50542 19966 50594
rect 20018 50542 20020 50594
rect 19964 50530 20020 50542
rect 20076 50706 20132 50718
rect 20076 50654 20078 50706
rect 20130 50654 20132 50706
rect 20076 50428 20132 50654
rect 20972 50428 21028 56028
rect 21196 56018 21252 56028
rect 21084 55412 21140 55422
rect 21084 54626 21140 55356
rect 21420 55298 21476 55310
rect 21420 55246 21422 55298
rect 21474 55246 21476 55298
rect 21420 54740 21476 55246
rect 21420 54674 21476 54684
rect 21532 54738 21588 59200
rect 21980 55970 22036 59200
rect 21980 55918 21982 55970
rect 22034 55918 22036 55970
rect 21980 55906 22036 55918
rect 22764 56082 22820 56094
rect 22764 56030 22766 56082
rect 22818 56030 22820 56082
rect 22092 55188 22148 55198
rect 21532 54686 21534 54738
rect 21586 54686 21588 54738
rect 21532 54674 21588 54686
rect 21868 55186 22148 55188
rect 21868 55134 22094 55186
rect 22146 55134 22148 55186
rect 21868 55132 22148 55134
rect 21084 54574 21086 54626
rect 21138 54574 21140 54626
rect 21084 54562 21140 54574
rect 21868 53954 21924 55132
rect 22092 55122 22148 55132
rect 21980 54740 22036 54750
rect 22652 54740 22708 54750
rect 21980 54646 22036 54684
rect 22428 54684 22652 54740
rect 21868 53902 21870 53954
rect 21922 53902 21924 53954
rect 21868 53890 21924 53902
rect 21868 53730 21924 53742
rect 21868 53678 21870 53730
rect 21922 53678 21924 53730
rect 21532 53618 21588 53630
rect 21532 53566 21534 53618
rect 21586 53566 21588 53618
rect 21532 52164 21588 53566
rect 21532 52098 21588 52108
rect 21868 52612 21924 53678
rect 22428 53172 22484 54684
rect 22652 54646 22708 54684
rect 22428 53170 22596 53172
rect 22428 53118 22430 53170
rect 22482 53118 22596 53170
rect 22428 53116 22596 53118
rect 22428 53106 22484 53116
rect 21868 52162 21924 52556
rect 21868 52110 21870 52162
rect 21922 52110 21924 52162
rect 21868 52098 21924 52110
rect 21980 52834 22036 52846
rect 21980 52782 21982 52834
rect 22034 52782 22036 52834
rect 21980 52276 22036 52782
rect 21980 52050 22036 52220
rect 21980 51998 21982 52050
rect 22034 51998 22036 52050
rect 21980 51986 22036 51998
rect 21756 51604 21812 51614
rect 21532 50708 21588 50718
rect 21532 50596 21588 50652
rect 20076 50372 20244 50428
rect 19628 50306 19684 50316
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19516 49870 19518 49922
rect 19570 49870 19572 49922
rect 19068 49588 19124 49598
rect 18732 49522 18788 49532
rect 18956 49532 19068 49588
rect 18732 49364 18788 49374
rect 18620 49028 18676 49038
rect 18508 48916 18564 48926
rect 18508 48822 18564 48860
rect 18620 47460 18676 48972
rect 18620 47394 18676 47404
rect 18620 46004 18676 46014
rect 18732 46004 18788 49308
rect 18844 49252 18900 49262
rect 18956 49252 19012 49532
rect 19068 49522 19124 49532
rect 18844 49250 19012 49252
rect 18844 49198 18846 49250
rect 18898 49198 19012 49250
rect 18844 49196 19012 49198
rect 19180 49364 19236 49374
rect 18844 49186 18900 49196
rect 19068 49140 19124 49150
rect 19068 49026 19124 49084
rect 19068 48974 19070 49026
rect 19122 48974 19124 49026
rect 19068 48962 19124 48974
rect 19180 46004 19236 49308
rect 19516 49026 19572 49870
rect 19740 49812 19796 49822
rect 19516 48974 19518 49026
rect 19570 48974 19572 49026
rect 19404 47572 19460 47582
rect 19516 47572 19572 48974
rect 19628 49810 19796 49812
rect 19628 49758 19742 49810
rect 19794 49758 19796 49810
rect 19628 49756 19796 49758
rect 19628 49028 19684 49756
rect 19740 49746 19796 49756
rect 20076 49810 20132 49822
rect 20076 49758 20078 49810
rect 20130 49758 20132 49810
rect 19964 49698 20020 49710
rect 19964 49646 19966 49698
rect 20018 49646 20020 49698
rect 19964 49588 20020 49646
rect 19964 49522 20020 49532
rect 20076 49364 20132 49758
rect 20076 49298 20132 49308
rect 20188 49252 20244 50372
rect 20188 49158 20244 49196
rect 20412 50372 20468 50382
rect 19628 48934 19684 48972
rect 19740 49028 19796 49038
rect 19740 49026 20356 49028
rect 19740 48974 19742 49026
rect 19794 48974 20356 49026
rect 19740 48972 20356 48974
rect 19740 48962 19796 48972
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19740 48468 19796 48478
rect 19740 48132 19796 48412
rect 19740 48130 19908 48132
rect 19740 48078 19742 48130
rect 19794 48078 19908 48130
rect 19740 48076 19908 48078
rect 19740 48066 19796 48076
rect 19404 47570 19572 47572
rect 19404 47518 19406 47570
rect 19458 47518 19572 47570
rect 19404 47516 19572 47518
rect 19852 47572 19908 48076
rect 20188 47684 20244 47694
rect 20300 47684 20356 48972
rect 20412 48804 20468 50316
rect 20748 50372 21028 50428
rect 21196 50594 21588 50596
rect 21196 50542 21534 50594
rect 21586 50542 21588 50594
rect 21196 50540 21588 50542
rect 20636 49812 20692 49822
rect 20636 49718 20692 49756
rect 20412 48738 20468 48748
rect 20524 49364 20580 49374
rect 20524 48916 20580 49308
rect 20748 49028 20804 50372
rect 21196 49812 21252 50540
rect 21532 50530 21588 50540
rect 21308 50372 21364 50382
rect 21308 50370 21476 50372
rect 21308 50318 21310 50370
rect 21362 50318 21476 50370
rect 21308 50316 21476 50318
rect 21308 50306 21364 50316
rect 21308 49812 21364 49822
rect 21196 49810 21364 49812
rect 21196 49758 21310 49810
rect 21362 49758 21364 49810
rect 21196 49756 21364 49758
rect 21308 49746 21364 49756
rect 21308 49364 21364 49374
rect 20524 48356 20580 48860
rect 20636 48972 20804 49028
rect 20860 49028 20916 49038
rect 20636 48468 20692 48972
rect 20748 48802 20804 48814
rect 20748 48750 20750 48802
rect 20802 48750 20804 48802
rect 20748 48692 20804 48750
rect 20748 48626 20804 48636
rect 20636 48412 20804 48468
rect 20524 48354 20692 48356
rect 20524 48302 20526 48354
rect 20578 48302 20692 48354
rect 20524 48300 20692 48302
rect 20524 48290 20580 48300
rect 20188 47682 20356 47684
rect 20188 47630 20190 47682
rect 20242 47630 20356 47682
rect 20188 47628 20356 47630
rect 20188 47618 20244 47628
rect 19404 47506 19460 47516
rect 19852 47478 19908 47516
rect 19404 47348 19460 47358
rect 19404 47068 19460 47292
rect 19836 47068 20100 47078
rect 19404 47012 19572 47068
rect 18620 46002 19012 46004
rect 18620 45950 18622 46002
rect 18674 45950 19012 46002
rect 18620 45948 19012 45950
rect 19180 45948 19460 46004
rect 18620 45938 18676 45948
rect 18956 45892 19012 45948
rect 18956 45890 19348 45892
rect 18956 45838 18958 45890
rect 19010 45838 19348 45890
rect 18956 45836 19348 45838
rect 18956 45826 19012 45836
rect 19068 45666 19124 45678
rect 19068 45614 19070 45666
rect 19122 45614 19124 45666
rect 19068 45332 19124 45614
rect 19180 45668 19236 45678
rect 19180 45574 19236 45612
rect 18732 45276 19124 45332
rect 18732 45218 18788 45276
rect 18732 45166 18734 45218
rect 18786 45166 18788 45218
rect 18732 45154 18788 45166
rect 18956 44436 19012 44446
rect 18508 43652 18564 43662
rect 18452 43650 18564 43652
rect 18452 43598 18510 43650
rect 18562 43598 18564 43650
rect 18452 43596 18564 43598
rect 17836 43538 18004 43540
rect 17836 43486 17838 43538
rect 17890 43486 18004 43538
rect 17836 43484 18004 43486
rect 17836 43474 17892 43484
rect 17388 43148 17780 43204
rect 17052 42774 17108 42812
rect 17276 42756 17332 42766
rect 17164 42700 17276 42756
rect 16716 41298 16884 41300
rect 16716 41246 16718 41298
rect 16770 41246 16884 41298
rect 16716 41244 16884 41246
rect 16716 41234 16772 41244
rect 16828 40404 16884 41244
rect 16940 41186 16996 41198
rect 16940 41134 16942 41186
rect 16994 41134 16996 41186
rect 16940 40628 16996 41134
rect 16940 40562 16996 40572
rect 16828 40338 16884 40348
rect 17164 40292 17220 42700
rect 17276 42690 17332 42700
rect 17388 42642 17444 42654
rect 17388 42590 17390 42642
rect 17442 42590 17444 42642
rect 17388 41748 17444 42590
rect 17388 41682 17444 41692
rect 17612 42642 17668 42654
rect 17612 42590 17614 42642
rect 17666 42590 17668 42642
rect 17276 41412 17332 41422
rect 17276 41318 17332 41356
rect 17612 41300 17668 42590
rect 17724 42530 17780 43148
rect 17836 42868 17892 42878
rect 17836 42774 17892 42812
rect 17948 42644 18004 43484
rect 18060 42980 18116 43596
rect 18396 43558 18452 43596
rect 18508 43586 18564 43596
rect 18956 43650 19012 44380
rect 18956 43598 18958 43650
rect 19010 43598 19012 43650
rect 18956 43586 19012 43598
rect 18844 43316 18900 43326
rect 18060 42914 18116 42924
rect 18620 43314 18900 43316
rect 18620 43262 18846 43314
rect 18898 43262 18900 43314
rect 18620 43260 18900 43262
rect 17724 42478 17726 42530
rect 17778 42478 17780 42530
rect 17724 42466 17780 42478
rect 17836 42588 18004 42644
rect 18060 42754 18116 42766
rect 18060 42702 18062 42754
rect 18114 42702 18116 42754
rect 17724 41972 17780 41982
rect 17724 41878 17780 41916
rect 17836 41300 17892 42588
rect 17948 42420 18004 42430
rect 17948 41970 18004 42364
rect 17948 41918 17950 41970
rect 18002 41918 18004 41970
rect 17948 41906 18004 41918
rect 16940 40236 17220 40292
rect 17388 41244 17668 41300
rect 17724 41244 17892 41300
rect 17948 41748 18004 41758
rect 16604 39620 16660 39676
rect 16380 39618 16660 39620
rect 16380 39566 16606 39618
rect 16658 39566 16660 39618
rect 16380 39564 16660 39566
rect 16380 38834 16436 39564
rect 16604 39554 16660 39564
rect 16828 39956 16884 39966
rect 16828 39060 16884 39900
rect 16828 38994 16884 39004
rect 16380 38782 16382 38834
rect 16434 38782 16436 38834
rect 16380 38770 16436 38782
rect 16828 38836 16884 38846
rect 16828 38742 16884 38780
rect 16044 36430 16046 36482
rect 16098 36430 16100 36482
rect 16044 36418 16100 36430
rect 16156 37324 16324 37380
rect 16604 38164 16660 38174
rect 16156 36372 16212 37324
rect 16156 36306 16212 36316
rect 16268 37154 16324 37166
rect 16268 37102 16270 37154
rect 16322 37102 16324 37154
rect 16044 36260 16100 36270
rect 16044 36166 16100 36204
rect 16268 36260 16324 37102
rect 16268 36194 16324 36204
rect 15708 35980 16324 36036
rect 15372 35924 15428 35934
rect 15372 35830 15428 35868
rect 15596 35700 15652 35710
rect 15596 35606 15652 35644
rect 15484 35588 15540 35598
rect 15260 35074 15316 35084
rect 15372 35586 15540 35588
rect 15372 35534 15486 35586
rect 15538 35534 15540 35586
rect 15372 35532 15540 35534
rect 15372 35028 15428 35532
rect 15484 35522 15540 35532
rect 15820 35586 15876 35598
rect 15820 35534 15822 35586
rect 15874 35534 15876 35586
rect 15820 35364 15876 35534
rect 16268 35586 16324 35980
rect 16492 35700 16548 35710
rect 16492 35606 16548 35644
rect 16268 35534 16270 35586
rect 16322 35534 16324 35586
rect 16268 35522 16324 35534
rect 16044 35476 16100 35486
rect 15932 35364 15988 35374
rect 15820 35308 15932 35364
rect 15484 35028 15540 35038
rect 15372 34972 15484 35028
rect 15932 35028 15988 35308
rect 16044 35308 16100 35420
rect 16044 35252 16436 35308
rect 15932 34972 16212 35028
rect 15484 34962 15540 34972
rect 15260 34902 15316 34914
rect 15260 34850 15262 34902
rect 15314 34850 15316 34902
rect 15260 34468 15316 34850
rect 15932 34804 15988 34814
rect 15932 34802 16100 34804
rect 15932 34750 15934 34802
rect 15986 34750 16100 34802
rect 15932 34748 16100 34750
rect 15932 34738 15988 34748
rect 15596 34580 15652 34590
rect 15260 34412 15540 34468
rect 15148 34302 15150 34354
rect 15202 34302 15204 34354
rect 15148 34290 15204 34302
rect 15036 34190 15038 34242
rect 15090 34190 15092 34242
rect 15036 33348 15092 34190
rect 15260 34242 15316 34254
rect 15260 34190 15262 34242
rect 15314 34190 15316 34242
rect 15036 33282 15092 33292
rect 15148 34132 15204 34142
rect 14700 32396 14980 32452
rect 14364 32340 14420 32350
rect 14588 32340 14644 32350
rect 14364 32338 14644 32340
rect 14364 32286 14366 32338
rect 14418 32286 14590 32338
rect 14642 32286 14644 32338
rect 14364 32284 14644 32286
rect 14364 32274 14420 32284
rect 14588 32274 14644 32284
rect 14700 31890 14756 32396
rect 15148 31948 15204 34076
rect 15260 33124 15316 34190
rect 15484 34020 15540 34412
rect 15484 33954 15540 33964
rect 15596 33796 15652 34524
rect 16044 34354 16100 34748
rect 16044 34302 16046 34354
rect 16098 34302 16100 34354
rect 16044 34290 16100 34302
rect 15260 33058 15316 33068
rect 15484 33740 15652 33796
rect 15932 34130 15988 34142
rect 15932 34078 15934 34130
rect 15986 34078 15988 34130
rect 15260 32676 15316 32686
rect 15484 32676 15540 33740
rect 15596 33124 15652 33134
rect 15652 33068 15764 33124
rect 15596 33030 15652 33068
rect 15260 32674 15540 32676
rect 15260 32622 15262 32674
rect 15314 32622 15540 32674
rect 15260 32620 15540 32622
rect 15596 32676 15652 32686
rect 15260 32610 15316 32620
rect 15596 32582 15652 32620
rect 15372 32452 15428 32462
rect 15708 32452 15764 33068
rect 15820 32788 15876 32798
rect 15820 32674 15876 32732
rect 15820 32622 15822 32674
rect 15874 32622 15876 32674
rect 15820 32610 15876 32622
rect 15820 32452 15876 32462
rect 15708 32396 15820 32452
rect 15372 32358 15428 32396
rect 15820 32386 15876 32396
rect 14700 31838 14702 31890
rect 14754 31838 14756 31890
rect 14700 31826 14756 31838
rect 14924 31892 15204 31948
rect 15372 32116 15428 32126
rect 14812 31668 14868 31678
rect 14812 31574 14868 31612
rect 14588 31556 14644 31566
rect 13916 30930 13972 30940
rect 14140 31164 14308 31220
rect 14364 31554 14644 31556
rect 14364 31502 14590 31554
rect 14642 31502 14644 31554
rect 14364 31500 14644 31502
rect 14028 30884 14084 30894
rect 14028 30790 14084 30828
rect 13692 30482 13748 30492
rect 13804 30660 13860 30670
rect 13468 30380 13636 30436
rect 13468 30324 13524 30380
rect 13804 30324 13860 30604
rect 13356 30268 13524 30324
rect 13580 30322 13860 30324
rect 13580 30270 13806 30322
rect 13858 30270 13860 30322
rect 13580 30268 13860 30270
rect 13356 29652 13412 30268
rect 13468 30100 13524 30110
rect 13468 30006 13524 30044
rect 13356 29538 13412 29596
rect 13356 29486 13358 29538
rect 13410 29486 13412 29538
rect 13356 29474 13412 29486
rect 13468 29314 13524 29326
rect 13468 29262 13470 29314
rect 13522 29262 13524 29314
rect 13468 28980 13524 29262
rect 13468 28914 13524 28924
rect 13020 27636 13076 27646
rect 13020 27542 13076 27580
rect 12460 27246 12462 27298
rect 12514 27246 12516 27298
rect 12460 27234 12516 27246
rect 12236 27076 12292 27086
rect 12236 26982 12292 27020
rect 13132 27076 13188 27086
rect 11564 26910 11566 26962
rect 11618 26910 11620 26962
rect 11564 26898 11620 26910
rect 11900 26962 11956 26974
rect 11900 26910 11902 26962
rect 11954 26910 11956 26962
rect 11340 26404 11396 26852
rect 10780 25508 10836 25518
rect 10780 25506 10948 25508
rect 10780 25454 10782 25506
rect 10834 25454 10948 25506
rect 10780 25452 10948 25454
rect 10780 25442 10836 25452
rect 10780 24948 10836 24958
rect 10780 24854 10836 24892
rect 10668 24836 10724 24846
rect 10668 24742 10724 24780
rect 10780 23828 10836 23838
rect 10780 23734 10836 23772
rect 10892 23380 10948 25452
rect 11004 24948 11060 24958
rect 11340 24948 11396 26348
rect 11900 25172 11956 26910
rect 12236 26404 12292 26414
rect 12236 26310 12292 26348
rect 13132 26402 13188 27020
rect 13132 26350 13134 26402
rect 13186 26350 13188 26402
rect 13132 26338 13188 26350
rect 13244 26178 13300 28588
rect 13356 28868 13412 28878
rect 13580 28868 13636 30268
rect 13804 30258 13860 30268
rect 14140 30212 14196 31164
rect 14252 30994 14308 31006
rect 14252 30942 14254 30994
rect 14306 30942 14308 30994
rect 14252 30436 14308 30942
rect 14252 30370 14308 30380
rect 14364 30212 14420 31500
rect 14588 31490 14644 31500
rect 14924 31220 14980 31892
rect 14476 31218 14980 31220
rect 14476 31166 14926 31218
rect 14978 31166 14980 31218
rect 14476 31164 14980 31166
rect 14476 31106 14532 31164
rect 14924 31154 14980 31164
rect 15036 31780 15092 31790
rect 14476 31054 14478 31106
rect 14530 31054 14532 31106
rect 14476 31042 14532 31054
rect 15036 30660 15092 31724
rect 15260 31778 15316 31790
rect 15260 31726 15262 31778
rect 15314 31726 15316 31778
rect 15260 31556 15316 31726
rect 15260 31490 15316 31500
rect 15036 30594 15092 30604
rect 15148 31108 15204 31118
rect 14924 30436 14980 30446
rect 14924 30342 14980 30380
rect 15036 30324 15092 30334
rect 14476 30212 14532 30222
rect 14700 30212 14756 30222
rect 14196 30156 14308 30212
rect 14364 30210 14756 30212
rect 14364 30158 14478 30210
rect 14530 30158 14702 30210
rect 14754 30158 14756 30210
rect 14364 30156 14756 30158
rect 14140 30146 14196 30156
rect 14252 30100 14308 30156
rect 14476 30146 14532 30156
rect 14700 30100 14756 30156
rect 15036 30210 15092 30268
rect 15036 30158 15038 30210
rect 15090 30158 15092 30210
rect 15036 30146 15092 30158
rect 14252 30044 14420 30100
rect 13692 29986 13748 29998
rect 13692 29934 13694 29986
rect 13746 29934 13748 29986
rect 13692 29204 13748 29934
rect 13916 29986 13972 29998
rect 13916 29934 13918 29986
rect 13970 29934 13972 29986
rect 13804 29428 13860 29438
rect 13916 29428 13972 29934
rect 14140 29988 14196 29998
rect 14140 29986 14308 29988
rect 14140 29934 14142 29986
rect 14194 29934 14308 29986
rect 14140 29932 14308 29934
rect 14140 29922 14196 29932
rect 14252 29652 14308 29932
rect 14364 29986 14420 30044
rect 15148 30100 15204 31052
rect 15260 31108 15316 31118
rect 15372 31108 15428 32060
rect 15820 31220 15876 31230
rect 15932 31220 15988 34078
rect 16156 33572 16212 34972
rect 16268 34916 16324 34926
rect 16268 34244 16324 34860
rect 16380 34580 16436 35252
rect 16380 34514 16436 34524
rect 16268 34150 16324 34188
rect 16492 34132 16548 34142
rect 16492 34038 16548 34076
rect 16604 33908 16660 38108
rect 16716 37266 16772 37278
rect 16716 37214 16718 37266
rect 16770 37214 16772 37266
rect 16716 37156 16772 37214
rect 16828 37156 16884 37166
rect 16716 37100 16828 37156
rect 16828 37090 16884 37100
rect 16940 37044 16996 40236
rect 17164 40068 17220 40078
rect 17388 40068 17444 41244
rect 17612 41076 17668 41086
rect 17612 40982 17668 41020
rect 17164 39730 17220 40012
rect 17164 39678 17166 39730
rect 17218 39678 17220 39730
rect 17164 38164 17220 39678
rect 17164 38098 17220 38108
rect 17276 40012 17444 40068
rect 17164 37940 17220 37950
rect 16716 36372 16772 36382
rect 16940 36372 16996 36988
rect 16716 36370 16996 36372
rect 16716 36318 16718 36370
rect 16770 36318 16996 36370
rect 16716 36316 16996 36318
rect 16716 36306 16772 36316
rect 16828 35924 16884 35934
rect 16716 35810 16772 35822
rect 16716 35758 16718 35810
rect 16770 35758 16772 35810
rect 16716 35588 16772 35758
rect 16828 35810 16884 35868
rect 16828 35758 16830 35810
rect 16882 35758 16884 35810
rect 16828 35746 16884 35758
rect 16716 35308 16772 35532
rect 16716 35252 16884 35308
rect 16268 33572 16324 33582
rect 16156 33570 16324 33572
rect 16156 33518 16270 33570
rect 16322 33518 16324 33570
rect 16156 33516 16324 33518
rect 16156 32676 16212 32686
rect 16156 32562 16212 32620
rect 16156 32510 16158 32562
rect 16210 32510 16212 32562
rect 16156 32498 16212 32510
rect 16044 31780 16100 31790
rect 16268 31780 16324 33516
rect 16492 33570 16548 33582
rect 16492 33518 16494 33570
rect 16546 33518 16548 33570
rect 16492 33458 16548 33518
rect 16492 33406 16494 33458
rect 16546 33406 16548 33458
rect 16492 33394 16548 33406
rect 16604 32788 16660 33852
rect 16604 32732 16772 32788
rect 16044 31332 16100 31724
rect 16044 31266 16100 31276
rect 16156 31724 16324 31780
rect 16604 32562 16660 32574
rect 16604 32510 16606 32562
rect 16658 32510 16660 32562
rect 16604 31780 16660 32510
rect 15820 31218 15988 31220
rect 15820 31166 15822 31218
rect 15874 31166 15988 31218
rect 15820 31164 15988 31166
rect 15820 31154 15876 31164
rect 15260 31106 15428 31108
rect 15260 31054 15262 31106
rect 15314 31054 15428 31106
rect 15260 31052 15428 31054
rect 15708 31108 15764 31118
rect 15260 30324 15316 31052
rect 15708 31014 15764 31052
rect 15484 30994 15540 31006
rect 15484 30942 15486 30994
rect 15538 30942 15540 30994
rect 15484 30772 15540 30942
rect 15484 30716 15876 30772
rect 15596 30548 15652 30558
rect 15596 30434 15652 30492
rect 15596 30382 15598 30434
rect 15650 30382 15652 30434
rect 15596 30370 15652 30382
rect 15260 30258 15316 30268
rect 15708 30324 15764 30334
rect 15708 30230 15764 30268
rect 15820 30212 15876 30716
rect 15932 30212 15988 30222
rect 15820 30210 15988 30212
rect 15820 30158 15934 30210
rect 15986 30158 15988 30210
rect 15820 30156 15988 30158
rect 15260 30100 15316 30110
rect 15148 30098 15316 30100
rect 15148 30046 15262 30098
rect 15314 30046 15316 30098
rect 15148 30044 15316 30046
rect 14700 30034 14756 30044
rect 15260 30034 15316 30044
rect 14364 29934 14366 29986
rect 14418 29934 14420 29986
rect 14364 29922 14420 29934
rect 14476 29876 14532 29886
rect 14252 29596 14420 29652
rect 14252 29428 14308 29438
rect 13916 29426 14308 29428
rect 13916 29374 14254 29426
rect 14306 29374 14308 29426
rect 13916 29372 14308 29374
rect 13804 29334 13860 29372
rect 14252 29316 14308 29372
rect 14252 29250 14308 29260
rect 13692 29148 13860 29204
rect 13804 28980 13860 29148
rect 13804 28914 13860 28924
rect 13692 28868 13748 28878
rect 13580 28866 13748 28868
rect 13580 28814 13694 28866
rect 13746 28814 13748 28866
rect 13580 28812 13748 28814
rect 13356 27858 13412 28812
rect 13692 28802 13748 28812
rect 13468 28644 13524 28654
rect 13468 28550 13524 28588
rect 14364 28532 14420 29596
rect 14476 29202 14532 29820
rect 14476 29150 14478 29202
rect 14530 29150 14532 29202
rect 14476 28868 14532 29150
rect 14812 29764 14868 29774
rect 14476 28802 14532 28812
rect 14700 28868 14756 28878
rect 14700 28754 14756 28812
rect 14812 28866 14868 29708
rect 15932 29764 15988 30156
rect 16156 29764 16212 31724
rect 16604 31714 16660 31724
rect 16268 31556 16324 31566
rect 16268 30996 16324 31500
rect 16268 30902 16324 30940
rect 16604 31108 16660 31118
rect 16156 29708 16324 29764
rect 15932 29698 15988 29708
rect 15148 29652 15204 29662
rect 15036 29540 15092 29550
rect 15036 29446 15092 29484
rect 15148 29538 15204 29596
rect 15148 29486 15150 29538
rect 15202 29486 15204 29538
rect 15148 29474 15204 29486
rect 16156 29540 16212 29550
rect 15820 29428 15876 29438
rect 15820 29334 15876 29372
rect 15036 29204 15092 29214
rect 15596 29204 15652 29214
rect 14812 28814 14814 28866
rect 14866 28814 14868 28866
rect 14812 28802 14868 28814
rect 14924 29202 15092 29204
rect 14924 29150 15038 29202
rect 15090 29150 15092 29202
rect 14924 29148 15092 29150
rect 14700 28702 14702 28754
rect 14754 28702 14756 28754
rect 14700 28690 14756 28702
rect 14364 28466 14420 28476
rect 14028 28420 14084 28430
rect 14028 28326 14084 28364
rect 13356 27806 13358 27858
rect 13410 27806 13412 27858
rect 13356 27794 13412 27806
rect 13580 27860 13636 27870
rect 13580 27766 13636 27804
rect 14700 27860 14756 27870
rect 14924 27860 14980 29148
rect 15036 29138 15092 29148
rect 15372 29202 15652 29204
rect 15372 29150 15598 29202
rect 15650 29150 15652 29202
rect 15372 29148 15652 29150
rect 14756 27804 14980 27860
rect 14364 27636 14420 27646
rect 14252 27076 14308 27086
rect 14252 26962 14308 27020
rect 14252 26910 14254 26962
rect 14306 26910 14308 26962
rect 13244 26126 13246 26178
rect 13298 26126 13300 26178
rect 13244 26114 13300 26126
rect 13356 26290 13412 26302
rect 13356 26238 13358 26290
rect 13410 26238 13412 26290
rect 12348 25618 12404 25630
rect 12348 25566 12350 25618
rect 12402 25566 12404 25618
rect 11900 25106 11956 25116
rect 12236 25506 12292 25518
rect 12236 25454 12238 25506
rect 12290 25454 12292 25506
rect 11004 24946 11396 24948
rect 11004 24894 11006 24946
rect 11058 24894 11396 24946
rect 11004 24892 11396 24894
rect 11452 25060 11508 25070
rect 11004 24882 11060 24892
rect 11340 24612 11396 24622
rect 11452 24612 11508 25004
rect 11340 24610 11508 24612
rect 11340 24558 11342 24610
rect 11394 24558 11508 24610
rect 11340 24556 11508 24558
rect 11340 24546 11396 24556
rect 12236 24388 12292 25454
rect 12236 24322 12292 24332
rect 12348 24500 12404 25566
rect 12348 23716 12404 24444
rect 12348 23650 12404 23660
rect 12796 25618 12852 25630
rect 12796 25566 12798 25618
rect 12850 25566 12852 25618
rect 10444 23324 10724 23380
rect 10332 22990 10334 23042
rect 10386 22990 10388 23042
rect 10332 22978 10388 22990
rect 10668 22820 10724 23324
rect 10892 23314 10948 23324
rect 11452 23154 11508 23166
rect 11452 23102 11454 23154
rect 11506 23102 11508 23154
rect 10780 23042 10836 23054
rect 10780 22990 10782 23042
rect 10834 22990 10836 23042
rect 10780 22932 10836 22990
rect 11452 22932 11508 23102
rect 12796 23156 12852 25566
rect 13020 25506 13076 25518
rect 13020 25454 13022 25506
rect 13074 25454 13076 25506
rect 13020 24836 13076 25454
rect 13020 24770 13076 24780
rect 13356 25172 13412 26238
rect 14140 26292 14196 26302
rect 14140 25508 14196 26236
rect 14140 25394 14196 25452
rect 14140 25342 14142 25394
rect 14194 25342 14196 25394
rect 14140 25330 14196 25342
rect 13692 25284 13748 25294
rect 13356 24612 13412 25116
rect 13468 25228 13692 25284
rect 13468 24834 13524 25228
rect 13692 25218 13748 25228
rect 13804 25282 13860 25294
rect 13804 25230 13806 25282
rect 13858 25230 13860 25282
rect 13804 25060 13860 25230
rect 13804 24994 13860 25004
rect 13468 24782 13470 24834
rect 13522 24782 13524 24834
rect 13468 24770 13524 24782
rect 14252 24724 14308 26910
rect 14364 26402 14420 27580
rect 14700 27186 14756 27804
rect 14700 27134 14702 27186
rect 14754 27134 14756 27186
rect 14700 27122 14756 27134
rect 15148 27746 15204 27758
rect 15148 27694 15150 27746
rect 15202 27694 15204 27746
rect 15148 27634 15204 27694
rect 15148 27582 15150 27634
rect 15202 27582 15204 27634
rect 15036 27076 15092 27086
rect 15036 26982 15092 27020
rect 14588 26852 14644 26862
rect 14588 26850 14756 26852
rect 14588 26798 14590 26850
rect 14642 26798 14756 26850
rect 14588 26796 14756 26798
rect 14588 26786 14644 26796
rect 14588 26516 14644 26526
rect 14364 26350 14366 26402
rect 14418 26350 14420 26402
rect 14364 26338 14420 26350
rect 14476 26514 14644 26516
rect 14476 26462 14590 26514
rect 14642 26462 14644 26514
rect 14476 26460 14644 26462
rect 14476 26292 14532 26460
rect 14588 26450 14644 26460
rect 14700 26292 14756 26796
rect 15148 26404 15204 27582
rect 15036 26292 15092 26302
rect 14476 26226 14532 26236
rect 14588 26290 15092 26292
rect 14588 26238 15038 26290
rect 15090 26238 15092 26290
rect 14588 26236 15092 26238
rect 14476 25508 14532 25518
rect 14588 25508 14644 26236
rect 15036 26226 15092 26236
rect 14700 26068 14756 26078
rect 14924 26068 14980 26078
rect 14700 26066 14924 26068
rect 14700 26014 14702 26066
rect 14754 26014 14924 26066
rect 14700 26012 14924 26014
rect 14700 26002 14756 26012
rect 14924 25730 14980 26012
rect 14924 25678 14926 25730
rect 14978 25678 14980 25730
rect 14924 25666 14980 25678
rect 14476 25506 14644 25508
rect 14476 25454 14478 25506
rect 14530 25454 14644 25506
rect 14476 25452 14644 25454
rect 14700 25508 14756 25518
rect 14756 25452 15092 25508
rect 14476 25442 14532 25452
rect 14700 25414 14756 25452
rect 14588 25284 14644 25294
rect 14588 25190 14644 25228
rect 14588 24836 14644 24846
rect 14588 24742 14644 24780
rect 13804 24722 14308 24724
rect 13804 24670 14254 24722
rect 14306 24670 14308 24722
rect 13804 24668 14308 24670
rect 13356 24556 13636 24612
rect 12908 24388 12964 24398
rect 12908 24052 12964 24332
rect 12908 24050 13524 24052
rect 12908 23998 12910 24050
rect 12962 23998 13524 24050
rect 12908 23996 13524 23998
rect 12908 23986 12964 23996
rect 13468 23938 13524 23996
rect 13468 23886 13470 23938
rect 13522 23886 13524 23938
rect 13468 23874 13524 23886
rect 13468 23716 13524 23726
rect 12908 23156 12964 23166
rect 12796 23154 12964 23156
rect 12796 23102 12910 23154
rect 12962 23102 12964 23154
rect 12796 23100 12964 23102
rect 12908 23090 12964 23100
rect 13468 23154 13524 23660
rect 13580 23378 13636 24556
rect 13580 23326 13582 23378
rect 13634 23326 13636 23378
rect 13580 23314 13636 23326
rect 13468 23102 13470 23154
rect 13522 23102 13524 23154
rect 13468 23090 13524 23102
rect 10780 22876 11508 22932
rect 10668 22764 11172 22820
rect 10220 22418 10276 22428
rect 10220 21588 10276 21598
rect 10108 21586 10276 21588
rect 10108 21534 10222 21586
rect 10274 21534 10276 21586
rect 10108 21532 10276 21534
rect 7420 20802 8036 20804
rect 7420 20750 7982 20802
rect 8034 20750 8036 20802
rect 7420 20748 8036 20750
rect 7420 19234 7476 20748
rect 7980 20738 8036 20748
rect 8652 20690 8708 20702
rect 8652 20638 8654 20690
rect 8706 20638 8708 20690
rect 8092 20580 8148 20590
rect 8092 19346 8148 20524
rect 8652 19460 8708 20638
rect 8652 19394 8708 19404
rect 8092 19294 8094 19346
rect 8146 19294 8148 19346
rect 8092 19282 8148 19294
rect 10220 19346 10276 21532
rect 10780 20914 10836 22764
rect 10780 20862 10782 20914
rect 10834 20862 10836 20914
rect 10780 20850 10836 20862
rect 11004 22484 11060 22494
rect 11004 20132 11060 22428
rect 11116 22370 11172 22764
rect 12908 22484 12964 22494
rect 12908 22390 12964 22428
rect 13804 22484 13860 24668
rect 14252 24658 14308 24668
rect 15036 24722 15092 25452
rect 15148 25506 15204 26348
rect 15260 26292 15316 26302
rect 15260 26198 15316 26236
rect 15148 25454 15150 25506
rect 15202 25454 15204 25506
rect 15148 25442 15204 25454
rect 15372 25284 15428 29148
rect 15596 29138 15652 29148
rect 15708 29204 15764 29214
rect 15596 27748 15652 27758
rect 15596 27654 15652 27692
rect 15484 26068 15540 26078
rect 15484 25974 15540 26012
rect 15708 25508 15764 29148
rect 16156 28866 16212 29484
rect 16156 28814 16158 28866
rect 16210 28814 16212 28866
rect 16156 28802 16212 28814
rect 16044 28532 16100 28542
rect 16044 28438 16100 28476
rect 16156 28418 16212 28430
rect 16156 28366 16158 28418
rect 16210 28366 16212 28418
rect 16044 28308 16100 28318
rect 16044 28084 16100 28252
rect 16156 28196 16212 28366
rect 16156 28130 16212 28140
rect 15932 28082 16100 28084
rect 15932 28030 16046 28082
rect 16098 28030 16100 28082
rect 15932 28028 16100 28030
rect 15820 27188 15876 27198
rect 15820 27094 15876 27132
rect 15820 26516 15876 26554
rect 15820 26450 15876 26460
rect 15820 26292 15876 26302
rect 15932 26292 15988 28028
rect 16044 28018 16100 28028
rect 16268 27634 16324 29708
rect 16492 29426 16548 29438
rect 16492 29374 16494 29426
rect 16546 29374 16548 29426
rect 16492 28420 16548 29374
rect 16604 29314 16660 31052
rect 16716 29428 16772 32732
rect 16716 29362 16772 29372
rect 16604 29262 16606 29314
rect 16658 29262 16660 29314
rect 16604 29250 16660 29262
rect 16492 28084 16548 28364
rect 16716 28532 16772 28542
rect 16828 28532 16884 35252
rect 16940 32676 16996 36316
rect 17052 37884 17164 37940
rect 17052 33458 17108 37884
rect 17164 37874 17220 37884
rect 17052 33406 17054 33458
rect 17106 33406 17108 33458
rect 17052 32788 17108 33406
rect 17164 37604 17220 37614
rect 17164 33348 17220 37548
rect 17276 33796 17332 40012
rect 17500 39732 17556 39742
rect 17724 39732 17780 41244
rect 17836 41074 17892 41086
rect 17836 41022 17838 41074
rect 17890 41022 17892 41074
rect 17836 40964 17892 41022
rect 17836 40898 17892 40908
rect 17948 40962 18004 41692
rect 18060 41636 18116 42702
rect 18284 42756 18340 42766
rect 18620 42756 18676 43260
rect 18844 43250 18900 43260
rect 18284 42754 18676 42756
rect 18284 42702 18286 42754
rect 18338 42702 18676 42754
rect 18284 42700 18676 42702
rect 18844 42754 18900 42766
rect 18844 42702 18846 42754
rect 18898 42702 18900 42754
rect 18284 42690 18340 42700
rect 18620 42532 18676 42542
rect 18508 42530 18676 42532
rect 18508 42478 18622 42530
rect 18674 42478 18676 42530
rect 18508 42476 18676 42478
rect 18172 41970 18228 41982
rect 18172 41918 18174 41970
rect 18226 41918 18228 41970
rect 18172 41748 18228 41918
rect 18396 41972 18452 41982
rect 18508 41972 18564 42476
rect 18620 42466 18676 42476
rect 18844 42532 18900 42702
rect 18844 42466 18900 42476
rect 18396 41970 18564 41972
rect 18396 41918 18398 41970
rect 18450 41918 18564 41970
rect 18396 41916 18564 41918
rect 18620 42308 18676 42318
rect 18396 41860 18452 41916
rect 18172 41682 18228 41692
rect 18284 41804 18396 41860
rect 18060 41570 18116 41580
rect 18060 41412 18116 41422
rect 18284 41412 18340 41804
rect 18396 41794 18452 41804
rect 18060 41410 18340 41412
rect 18060 41358 18062 41410
rect 18114 41358 18340 41410
rect 18060 41356 18340 41358
rect 18060 41346 18116 41356
rect 18396 41300 18452 41310
rect 18284 41188 18340 41198
rect 18396 41188 18452 41244
rect 18284 41186 18452 41188
rect 18284 41134 18286 41186
rect 18338 41134 18452 41186
rect 18284 41132 18452 41134
rect 18284 41122 18340 41132
rect 17948 40910 17950 40962
rect 18002 40910 18004 40962
rect 17948 40898 18004 40910
rect 18508 41074 18564 41086
rect 18508 41022 18510 41074
rect 18562 41022 18564 41074
rect 18508 40740 18564 41022
rect 18508 40514 18564 40684
rect 18508 40462 18510 40514
rect 18562 40462 18564 40514
rect 18508 40450 18564 40462
rect 17500 38724 17556 39676
rect 17612 39676 17724 39732
rect 17612 39284 17668 39676
rect 17724 39666 17780 39676
rect 17836 40404 17892 40414
rect 17836 39618 17892 40348
rect 18284 40404 18340 40414
rect 18340 40348 18452 40404
rect 18284 40338 18340 40348
rect 17836 39566 17838 39618
rect 17890 39566 17892 39618
rect 17836 39554 17892 39566
rect 18284 39956 18340 39966
rect 18284 39618 18340 39900
rect 18284 39566 18286 39618
rect 18338 39566 18340 39618
rect 18284 39554 18340 39566
rect 17724 39506 17780 39518
rect 17724 39454 17726 39506
rect 17778 39454 17780 39506
rect 17724 39396 17780 39454
rect 17724 39340 17892 39396
rect 17612 39228 17780 39284
rect 17724 39002 17780 39228
rect 17612 38946 17668 38958
rect 17612 38894 17614 38946
rect 17666 38894 17668 38946
rect 17724 38950 17726 39002
rect 17778 38950 17780 39002
rect 17724 38938 17780 38950
rect 17836 39004 17892 39340
rect 17836 38948 18004 39004
rect 17612 38836 17668 38894
rect 17836 38836 17892 38846
rect 17612 38780 17780 38836
rect 17500 38658 17556 38668
rect 17612 38610 17668 38622
rect 17612 38558 17614 38610
rect 17666 38558 17668 38610
rect 17500 38050 17556 38062
rect 17500 37998 17502 38050
rect 17554 37998 17556 38050
rect 17388 37828 17444 37838
rect 17388 37492 17444 37772
rect 17388 37398 17444 37436
rect 17500 36484 17556 37998
rect 17612 37156 17668 38558
rect 17612 37090 17668 37100
rect 17724 37490 17780 38780
rect 17836 37604 17892 38780
rect 17836 37538 17892 37548
rect 17724 37438 17726 37490
rect 17778 37438 17780 37490
rect 17724 36820 17780 37438
rect 17948 37492 18004 38948
rect 18284 38946 18340 38958
rect 18284 38894 18286 38946
rect 18338 38894 18340 38946
rect 18284 38836 18340 38894
rect 18284 38770 18340 38780
rect 18172 38724 18228 38762
rect 18172 38658 18228 38668
rect 17948 37426 18004 37436
rect 18284 37380 18340 37390
rect 18396 37380 18452 40348
rect 18508 39620 18564 39630
rect 18508 39526 18564 39564
rect 18508 38834 18564 38846
rect 18508 38782 18510 38834
rect 18562 38782 18564 38834
rect 18508 38164 18564 38782
rect 18508 38098 18564 38108
rect 18284 37378 18452 37380
rect 18284 37326 18286 37378
rect 18338 37326 18452 37378
rect 18284 37324 18452 37326
rect 18284 37314 18340 37324
rect 18508 37268 18564 37278
rect 18396 37266 18564 37268
rect 18396 37214 18510 37266
rect 18562 37214 18564 37266
rect 18396 37212 18564 37214
rect 17724 36764 18340 36820
rect 17612 36484 17668 36494
rect 17500 36482 17892 36484
rect 17500 36430 17614 36482
rect 17666 36430 17892 36482
rect 17500 36428 17892 36430
rect 17612 36418 17668 36428
rect 17388 35588 17444 35598
rect 17388 35494 17444 35532
rect 17612 35474 17668 35486
rect 17612 35422 17614 35474
rect 17666 35422 17668 35474
rect 17500 34916 17556 34926
rect 17500 34354 17556 34860
rect 17500 34302 17502 34354
rect 17554 34302 17556 34354
rect 17500 34132 17556 34302
rect 17500 34066 17556 34076
rect 17612 34468 17668 35422
rect 17612 33908 17668 34412
rect 17612 33842 17668 33852
rect 17724 35476 17780 35486
rect 17276 33740 17556 33796
rect 17164 33292 17332 33348
rect 17052 32722 17108 32732
rect 17164 33124 17220 33134
rect 16940 32610 16996 32620
rect 17164 31666 17220 33068
rect 17164 31614 17166 31666
rect 17218 31614 17220 31666
rect 17164 31602 17220 31614
rect 17276 31444 17332 33292
rect 17388 32788 17444 32798
rect 17388 32694 17444 32732
rect 17164 31388 17332 31444
rect 17388 31556 17444 31566
rect 17164 30772 17220 31388
rect 17388 31220 17444 31500
rect 17388 31126 17444 31164
rect 17500 31218 17556 33740
rect 17500 31166 17502 31218
rect 17554 31166 17556 31218
rect 17500 31154 17556 31166
rect 17612 31108 17668 31118
rect 17612 31014 17668 31052
rect 17724 30884 17780 35420
rect 17164 30210 17220 30716
rect 17164 30158 17166 30210
rect 17218 30158 17220 30210
rect 17164 30146 17220 30158
rect 17388 30828 17780 30884
rect 17836 31890 17892 36428
rect 17948 36372 18004 36382
rect 17948 35922 18004 36316
rect 17948 35870 17950 35922
rect 18002 35870 18004 35922
rect 17948 35858 18004 35870
rect 18284 35812 18340 36764
rect 18172 35810 18340 35812
rect 18172 35758 18286 35810
rect 18338 35758 18340 35810
rect 18172 35756 18340 35758
rect 18060 35028 18116 35038
rect 18172 35028 18228 35756
rect 18284 35746 18340 35756
rect 18396 35586 18452 37212
rect 18508 37202 18564 37212
rect 18396 35534 18398 35586
rect 18450 35534 18452 35586
rect 18284 35476 18340 35486
rect 18396 35476 18452 35534
rect 18340 35420 18452 35476
rect 18284 35410 18340 35420
rect 18060 35026 18228 35028
rect 18060 34974 18062 35026
rect 18114 34974 18228 35026
rect 18060 34972 18228 34974
rect 18060 34962 18116 34972
rect 17948 33124 18004 33134
rect 17948 33030 18004 33068
rect 18172 32676 18228 34972
rect 18620 34916 18676 42252
rect 19292 42196 19348 45836
rect 19180 42140 19348 42196
rect 18732 41970 18788 41982
rect 18732 41918 18734 41970
rect 18786 41918 18788 41970
rect 18732 41412 18788 41918
rect 18844 41972 18900 41982
rect 18844 41878 18900 41916
rect 19068 41970 19124 41982
rect 19068 41918 19070 41970
rect 19122 41918 19124 41970
rect 18732 41346 18788 41356
rect 19068 41748 19124 41918
rect 19068 41074 19124 41692
rect 19068 41022 19070 41074
rect 19122 41022 19124 41074
rect 19068 40964 19124 41022
rect 19068 40898 19124 40908
rect 18844 40404 18900 40414
rect 18844 40310 18900 40348
rect 19068 40404 19124 40414
rect 18844 39732 18900 39742
rect 18844 39638 18900 39676
rect 18844 39172 18900 39182
rect 18732 38834 18788 38846
rect 18732 38782 18734 38834
rect 18786 38782 18788 38834
rect 18732 36484 18788 38782
rect 18844 38276 18900 39116
rect 19068 38668 19124 40348
rect 19180 39620 19236 42140
rect 19292 41970 19348 41982
rect 19292 41918 19294 41970
rect 19346 41918 19348 41970
rect 19292 41860 19348 41918
rect 19292 41524 19348 41804
rect 19404 41636 19460 45948
rect 19516 45890 19572 47012
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20300 46898 20356 47628
rect 20524 47684 20580 47694
rect 20524 47590 20580 47628
rect 20300 46846 20302 46898
rect 20354 46846 20356 46898
rect 20300 46834 20356 46846
rect 20412 47012 20468 47022
rect 20412 46676 20468 46956
rect 20636 46898 20692 48300
rect 20748 47684 20804 48412
rect 20860 48242 20916 48972
rect 21308 49026 21364 49308
rect 21308 48974 21310 49026
rect 21362 48974 21364 49026
rect 21308 48962 21364 48974
rect 21420 49028 21476 50316
rect 21644 49810 21700 49822
rect 21644 49758 21646 49810
rect 21698 49758 21700 49810
rect 21644 49252 21700 49758
rect 21644 49186 21700 49196
rect 21420 48962 21476 48972
rect 21532 49026 21588 49038
rect 21532 48974 21534 49026
rect 21586 48974 21588 49026
rect 21532 48916 21588 48974
rect 21084 48804 21140 48814
rect 20972 48468 21028 48478
rect 20972 48374 21028 48412
rect 20860 48190 20862 48242
rect 20914 48190 20916 48242
rect 20860 48178 20916 48190
rect 21084 48242 21140 48748
rect 21420 48802 21476 48814
rect 21420 48750 21422 48802
rect 21474 48750 21476 48802
rect 21420 48356 21476 48750
rect 21084 48190 21086 48242
rect 21138 48190 21140 48242
rect 21084 48178 21140 48190
rect 21196 48300 21476 48356
rect 21084 48020 21140 48030
rect 21196 48020 21252 48300
rect 21084 48018 21252 48020
rect 21084 47966 21086 48018
rect 21138 47966 21252 48018
rect 21084 47964 21252 47966
rect 21084 47954 21140 47964
rect 21420 47684 21476 47694
rect 20748 47628 20916 47684
rect 20748 47458 20804 47470
rect 20748 47406 20750 47458
rect 20802 47406 20804 47458
rect 20748 47348 20804 47406
rect 20748 47282 20804 47292
rect 20636 46846 20638 46898
rect 20690 46846 20692 46898
rect 20636 46834 20692 46846
rect 19516 45838 19518 45890
rect 19570 45838 19572 45890
rect 19516 45826 19572 45838
rect 19628 46562 19684 46574
rect 19628 46510 19630 46562
rect 19682 46510 19684 46562
rect 19628 45668 19684 46510
rect 20412 46002 20468 46620
rect 20412 45950 20414 46002
rect 20466 45950 20468 46002
rect 20412 45938 20468 45950
rect 19516 45220 19572 45230
rect 19516 44436 19572 45164
rect 19516 44342 19572 44380
rect 19628 43988 19684 45612
rect 20076 45780 20132 45790
rect 20076 45668 20132 45724
rect 20076 45666 20244 45668
rect 20076 45614 20078 45666
rect 20130 45614 20244 45666
rect 20076 45612 20244 45614
rect 20076 45602 20132 45612
rect 20188 45556 20244 45612
rect 19836 45500 20100 45510
rect 20188 45500 20356 45556
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20076 44884 20132 44894
rect 19852 44212 19908 44222
rect 19852 44118 19908 44156
rect 20076 44098 20132 44828
rect 20076 44046 20078 44098
rect 20130 44046 20132 44098
rect 20076 44034 20132 44046
rect 20188 44210 20244 44222
rect 20188 44158 20190 44210
rect 20242 44158 20244 44210
rect 19628 43428 19684 43932
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19740 43428 19796 43438
rect 19628 43426 19796 43428
rect 19628 43374 19742 43426
rect 19794 43374 19796 43426
rect 19628 43372 19796 43374
rect 19516 42532 19572 42542
rect 19516 42084 19572 42476
rect 19628 42308 19684 43372
rect 19740 43362 19796 43372
rect 20188 42756 20244 44158
rect 20300 43316 20356 45500
rect 20860 45220 20916 47628
rect 21308 47628 21420 47684
rect 21308 47236 21364 47628
rect 21420 47618 21476 47628
rect 21420 47460 21476 47470
rect 21532 47460 21588 48860
rect 21756 48692 21812 51548
rect 22540 51604 22596 53116
rect 22764 52388 22820 56030
rect 22876 54740 22932 59200
rect 22988 54740 23044 54750
rect 22876 54738 23044 54740
rect 22876 54686 22990 54738
rect 23042 54686 23044 54738
rect 22876 54684 23044 54686
rect 23324 54740 23380 59200
rect 24220 57204 24276 59200
rect 24220 57148 24612 57204
rect 23660 56642 23716 56654
rect 23660 56590 23662 56642
rect 23714 56590 23716 56642
rect 23660 56194 23716 56590
rect 23660 56142 23662 56194
rect 23714 56142 23716 56194
rect 23660 56130 23716 56142
rect 24220 55412 24276 55422
rect 24220 55410 24388 55412
rect 24220 55358 24222 55410
rect 24274 55358 24388 55410
rect 24220 55356 24388 55358
rect 24220 55346 24276 55356
rect 23548 55076 23604 55086
rect 23436 54740 23492 54750
rect 23324 54738 23492 54740
rect 23324 54686 23438 54738
rect 23490 54686 23492 54738
rect 23324 54684 23492 54686
rect 22988 54674 23044 54684
rect 23436 54674 23492 54684
rect 23324 53844 23380 53854
rect 22876 53732 22932 53742
rect 22876 52946 22932 53676
rect 23100 53508 23156 53518
rect 23324 53508 23380 53788
rect 23100 53506 23380 53508
rect 23100 53454 23102 53506
rect 23154 53454 23380 53506
rect 23100 53452 23380 53454
rect 23100 53442 23156 53452
rect 22876 52894 22878 52946
rect 22930 52894 22932 52946
rect 22876 52882 22932 52894
rect 22988 52722 23044 52734
rect 22988 52670 22990 52722
rect 23042 52670 23044 52722
rect 22988 52500 23044 52670
rect 22988 52444 23268 52500
rect 22764 52332 23156 52388
rect 22764 52162 22820 52174
rect 22764 52110 22766 52162
rect 22818 52110 22820 52162
rect 22540 51510 22596 51548
rect 22652 51938 22708 51950
rect 22652 51886 22654 51938
rect 22706 51886 22708 51938
rect 22652 51380 22708 51886
rect 22652 51314 22708 51324
rect 22092 51266 22148 51278
rect 22092 51214 22094 51266
rect 22146 51214 22148 51266
rect 22092 50932 22148 51214
rect 22092 50428 22148 50876
rect 22764 50706 22820 52110
rect 22764 50654 22766 50706
rect 22818 50654 22820 50706
rect 22764 50642 22820 50654
rect 22988 51268 23044 51278
rect 22652 50596 22708 50606
rect 22428 50484 22484 50522
rect 22652 50428 22708 50540
rect 22092 50372 22372 50428
rect 22428 50418 22484 50428
rect 22316 50036 22372 50372
rect 22540 50372 22708 50428
rect 22876 50372 22932 50382
rect 22988 50372 23044 51212
rect 22428 50036 22484 50046
rect 22316 50034 22484 50036
rect 22316 49982 22430 50034
rect 22482 49982 22484 50034
rect 22316 49980 22484 49982
rect 22428 49970 22484 49980
rect 22540 49922 22596 50372
rect 22876 50370 23044 50372
rect 22876 50318 22878 50370
rect 22930 50318 23044 50370
rect 22876 50316 23044 50318
rect 22876 50306 22932 50316
rect 22540 49870 22542 49922
rect 22594 49870 22596 49922
rect 22540 49858 22596 49870
rect 21868 49812 21924 49822
rect 22204 49812 22260 49822
rect 21868 49810 22260 49812
rect 21868 49758 21870 49810
rect 21922 49758 22206 49810
rect 22258 49758 22260 49810
rect 21868 49756 22260 49758
rect 21868 49364 21924 49756
rect 22204 49746 22260 49756
rect 21868 49298 21924 49308
rect 22092 49252 22148 49262
rect 21868 49028 21924 49038
rect 21868 48934 21924 48972
rect 22092 49026 22148 49196
rect 22092 48974 22094 49026
rect 22146 48974 22148 49026
rect 22092 48962 22148 48974
rect 22988 49026 23044 50316
rect 22988 48974 22990 49026
rect 23042 48974 23044 49026
rect 22988 48962 23044 48974
rect 22428 48916 22484 48926
rect 22876 48916 22932 48926
rect 22428 48914 22932 48916
rect 22428 48862 22430 48914
rect 22482 48862 22878 48914
rect 22930 48862 22932 48914
rect 22428 48860 22932 48862
rect 22428 48850 22484 48860
rect 21756 48244 21812 48636
rect 22316 48802 22372 48814
rect 22316 48750 22318 48802
rect 22370 48750 22372 48802
rect 21868 48244 21924 48254
rect 21756 48242 21924 48244
rect 21756 48190 21870 48242
rect 21922 48190 21924 48242
rect 21756 48188 21924 48190
rect 21868 48178 21924 48188
rect 21644 47684 21700 47694
rect 22204 47684 22260 47694
rect 21644 47682 22260 47684
rect 21644 47630 21646 47682
rect 21698 47630 22206 47682
rect 22258 47630 22260 47682
rect 21644 47628 22260 47630
rect 21644 47618 21700 47628
rect 22204 47618 22260 47628
rect 21756 47460 21812 47470
rect 21532 47458 21812 47460
rect 21532 47406 21758 47458
rect 21810 47406 21812 47458
rect 21532 47404 21812 47406
rect 21420 47366 21476 47404
rect 21756 47394 21812 47404
rect 22316 47348 22372 48750
rect 22540 48468 22596 48478
rect 22540 48354 22596 48412
rect 22540 48302 22542 48354
rect 22594 48302 22596 48354
rect 22540 48290 22596 48302
rect 22540 47684 22596 47694
rect 22652 47684 22708 48860
rect 22876 48850 22932 48860
rect 22596 47628 22708 47684
rect 22540 47590 22596 47628
rect 22316 47254 22372 47292
rect 21308 47180 21588 47236
rect 21308 46564 21364 46574
rect 20860 45154 20916 45164
rect 21196 46508 21308 46564
rect 21196 45668 21252 46508
rect 21308 46470 21364 46508
rect 21532 46562 21588 47180
rect 21756 47234 21812 47246
rect 21756 47182 21758 47234
rect 21810 47182 21812 47234
rect 21756 46788 21812 47182
rect 22988 47236 23044 47246
rect 22988 47142 23044 47180
rect 21756 46722 21812 46732
rect 21532 46510 21534 46562
rect 21586 46510 21588 46562
rect 21532 46498 21588 46510
rect 21196 45108 21252 45612
rect 21420 45668 21476 45678
rect 21868 45668 21924 45678
rect 21420 45666 21924 45668
rect 21420 45614 21422 45666
rect 21474 45614 21870 45666
rect 21922 45614 21924 45666
rect 21420 45612 21924 45614
rect 21420 45108 21476 45612
rect 21868 45602 21924 45612
rect 21196 45106 21476 45108
rect 21196 45054 21198 45106
rect 21250 45054 21476 45106
rect 21196 45052 21476 45054
rect 21196 45042 21252 45052
rect 20860 44996 20916 45006
rect 20748 44994 20916 44996
rect 20748 44942 20862 44994
rect 20914 44942 20916 44994
rect 20748 44940 20916 44942
rect 20412 44324 20468 44334
rect 20412 44230 20468 44268
rect 20412 43316 20468 43326
rect 20300 43260 20412 43316
rect 20412 43250 20468 43260
rect 20188 42690 20244 42700
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19628 42242 19684 42252
rect 19628 42084 19684 42094
rect 19516 42082 19684 42084
rect 19516 42030 19630 42082
rect 19682 42030 19684 42082
rect 19516 42028 19684 42030
rect 19628 42018 19684 42028
rect 19852 42084 19908 42094
rect 19404 41580 19684 41636
rect 19292 41468 19572 41524
rect 19516 41410 19572 41468
rect 19516 41358 19518 41410
rect 19570 41358 19572 41410
rect 19516 41346 19572 41358
rect 19292 41188 19348 41198
rect 19292 41094 19348 41132
rect 19516 41076 19572 41086
rect 19292 40628 19348 40666
rect 19292 40562 19348 40572
rect 19516 40402 19572 41020
rect 19516 40350 19518 40402
rect 19570 40350 19572 40402
rect 19292 39956 19348 39966
rect 19292 39730 19348 39900
rect 19292 39678 19294 39730
rect 19346 39678 19348 39730
rect 19292 39666 19348 39678
rect 19180 39508 19236 39564
rect 19180 39452 19348 39508
rect 19180 38948 19236 38958
rect 19180 38854 19236 38892
rect 19068 38612 19236 38668
rect 18844 38220 19124 38276
rect 18732 35922 18788 36428
rect 18732 35870 18734 35922
rect 18786 35870 18788 35922
rect 18732 35858 18788 35870
rect 18844 38050 18900 38062
rect 18844 37998 18846 38050
rect 18898 37998 18900 38050
rect 18844 35252 18900 37998
rect 18956 37492 19012 37502
rect 18956 36820 19012 37436
rect 19068 36932 19124 38220
rect 19180 37492 19236 38612
rect 19180 37426 19236 37436
rect 19068 36876 19236 36932
rect 18956 36764 19124 36820
rect 18284 34914 18676 34916
rect 18284 34862 18622 34914
rect 18674 34862 18676 34914
rect 18284 34860 18676 34862
rect 18284 34020 18340 34860
rect 18620 34850 18676 34860
rect 18732 35196 18900 35252
rect 18956 35698 19012 35710
rect 18956 35646 18958 35698
rect 19010 35646 19012 35698
rect 18396 34692 18452 34702
rect 18396 34132 18452 34636
rect 18396 34066 18452 34076
rect 18620 34130 18676 34142
rect 18620 34078 18622 34130
rect 18674 34078 18676 34130
rect 18284 33954 18340 33964
rect 18508 34018 18564 34030
rect 18508 33966 18510 34018
rect 18562 33966 18564 34018
rect 18284 33124 18340 33134
rect 18508 33124 18564 33966
rect 18620 33236 18676 34078
rect 18620 33170 18676 33180
rect 18284 33122 18564 33124
rect 18284 33070 18286 33122
rect 18338 33070 18564 33122
rect 18284 33068 18564 33070
rect 18284 33012 18340 33068
rect 18732 33012 18788 35196
rect 18956 35140 19012 35646
rect 18844 35138 19012 35140
rect 18844 35086 18958 35138
rect 19010 35086 19012 35138
rect 18844 35084 19012 35086
rect 18844 33234 18900 35084
rect 18956 35074 19012 35084
rect 18956 34132 19012 34142
rect 19068 34132 19124 36764
rect 19180 35140 19236 36876
rect 19292 35364 19348 39452
rect 19404 38834 19460 38846
rect 19404 38782 19406 38834
rect 19458 38782 19460 38834
rect 19404 38724 19460 38782
rect 19404 38658 19460 38668
rect 19516 36260 19572 40350
rect 19628 39956 19684 41580
rect 19852 41298 19908 42028
rect 19964 42082 20020 42094
rect 19964 42030 19966 42082
rect 20018 42030 20020 42082
rect 19964 41860 20020 42030
rect 19964 41636 20020 41804
rect 19964 41570 20020 41580
rect 19852 41246 19854 41298
rect 19906 41246 19908 41298
rect 19852 41234 19908 41246
rect 19740 41188 19796 41198
rect 19740 41094 19796 41132
rect 19964 41074 20020 41086
rect 19964 41022 19966 41074
rect 20018 41022 20020 41074
rect 19964 40964 20020 41022
rect 20636 41076 20692 41086
rect 20636 40982 20692 41020
rect 20300 40964 20356 40974
rect 19964 40908 20244 40964
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20188 40628 20244 40908
rect 20300 40870 20356 40908
rect 20636 40628 20692 40638
rect 20188 40572 20636 40628
rect 20636 40534 20692 40572
rect 19628 39890 19684 39900
rect 20076 39508 20132 39518
rect 19628 39452 20076 39508
rect 19628 39060 19684 39452
rect 20076 39414 20132 39452
rect 20188 39394 20244 39406
rect 20188 39342 20190 39394
rect 20242 39342 20244 39394
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19740 39060 19796 39070
rect 19628 39058 19796 39060
rect 19628 39006 19742 39058
rect 19794 39006 19796 39058
rect 19628 39004 19796 39006
rect 19628 38164 19684 38174
rect 19628 38070 19684 38108
rect 19740 38050 19796 39004
rect 20076 38724 20132 38762
rect 20076 38658 20132 38668
rect 20188 38500 20244 39342
rect 20748 39396 20804 44940
rect 20860 44930 20916 44940
rect 21420 44434 21476 45052
rect 21420 44382 21422 44434
rect 21474 44382 21476 44434
rect 21420 44370 21476 44382
rect 21756 45220 21812 45230
rect 21308 44212 21364 44222
rect 21196 43652 21252 43662
rect 20860 43538 20916 43550
rect 20860 43486 20862 43538
rect 20914 43486 20916 43538
rect 20860 42084 20916 43486
rect 21196 43538 21252 43596
rect 21308 43650 21364 44156
rect 21308 43598 21310 43650
rect 21362 43598 21364 43650
rect 21308 43586 21364 43598
rect 21532 43764 21588 43774
rect 21196 43486 21198 43538
rect 21250 43486 21252 43538
rect 21196 43474 21252 43486
rect 21420 43538 21476 43550
rect 21420 43486 21422 43538
rect 21474 43486 21476 43538
rect 21420 43092 21476 43486
rect 21196 43036 21476 43092
rect 21196 42532 21252 43036
rect 21532 42980 21588 43708
rect 21756 43428 21812 45164
rect 23100 45220 23156 52332
rect 23212 52164 23268 52444
rect 23212 51490 23268 52108
rect 23324 51940 23380 53452
rect 23436 53730 23492 53742
rect 23436 53678 23438 53730
rect 23490 53678 23492 53730
rect 23436 53508 23492 53678
rect 23436 52724 23492 53452
rect 23436 52658 23492 52668
rect 23324 51874 23380 51884
rect 23548 51604 23604 55020
rect 24220 54514 24276 54526
rect 24220 54462 24222 54514
rect 24274 54462 24276 54514
rect 23660 53844 23716 53854
rect 23660 53750 23716 53788
rect 23996 53506 24052 53518
rect 23996 53454 23998 53506
rect 24050 53454 24052 53506
rect 23660 53058 23716 53070
rect 23660 53006 23662 53058
rect 23714 53006 23716 53058
rect 23660 52052 23716 53006
rect 23884 53058 23940 53070
rect 23884 53006 23886 53058
rect 23938 53006 23940 53058
rect 23884 52612 23940 53006
rect 23884 52546 23940 52556
rect 23996 52162 24052 53454
rect 24220 52948 24276 54462
rect 24332 53732 24388 55356
rect 24556 55186 24612 57148
rect 24668 56642 24724 59200
rect 24668 56590 24670 56642
rect 24722 56590 24724 56642
rect 24668 56578 24724 56590
rect 24556 55134 24558 55186
rect 24610 55134 24612 55186
rect 24556 55122 24612 55134
rect 24668 56082 24724 56094
rect 24668 56030 24670 56082
rect 24722 56030 24724 56082
rect 24668 55300 24724 56030
rect 25340 55972 25396 55982
rect 24668 54740 24724 55244
rect 24668 54646 24724 54684
rect 25228 55970 25396 55972
rect 25228 55918 25342 55970
rect 25394 55918 25396 55970
rect 25228 55916 25396 55918
rect 25228 54738 25284 55916
rect 25340 55906 25396 55916
rect 25564 55524 25620 59200
rect 26012 56980 26068 59200
rect 26012 56924 26740 56980
rect 25340 55468 25620 55524
rect 25340 55186 25396 55468
rect 25676 55300 25732 55310
rect 25676 55206 25732 55244
rect 25340 55134 25342 55186
rect 25394 55134 25396 55186
rect 25340 55122 25396 55134
rect 26460 55188 26516 55198
rect 26460 55094 26516 55132
rect 25228 54686 25230 54738
rect 25282 54686 25284 54738
rect 25228 54674 25284 54686
rect 25564 54514 25620 54526
rect 26348 54516 26404 54526
rect 25564 54462 25566 54514
rect 25618 54462 25620 54514
rect 24332 53638 24388 53676
rect 24892 53730 24948 53742
rect 24892 53678 24894 53730
rect 24946 53678 24948 53730
rect 24220 52892 24388 52948
rect 24220 52724 24276 52734
rect 24220 52630 24276 52668
rect 23996 52110 23998 52162
rect 24050 52110 24052 52162
rect 23996 52098 24052 52110
rect 23660 51986 23716 51996
rect 23436 51548 23604 51604
rect 23772 51940 23828 51950
rect 23212 51438 23214 51490
rect 23266 51438 23268 51490
rect 23212 51426 23268 51438
rect 23324 51490 23380 51502
rect 23324 51438 23326 51490
rect 23378 51438 23380 51490
rect 23324 50932 23380 51438
rect 23436 51156 23492 51548
rect 23548 51380 23604 51390
rect 23548 51378 23716 51380
rect 23548 51326 23550 51378
rect 23602 51326 23716 51378
rect 23548 51324 23716 51326
rect 23548 51314 23604 51324
rect 23436 51100 23604 51156
rect 23324 50866 23380 50876
rect 23100 45154 23156 45164
rect 21980 44996 22036 45006
rect 21980 44994 22260 44996
rect 21980 44942 21982 44994
rect 22034 44942 22260 44994
rect 21980 44940 22260 44942
rect 21980 44930 22036 44940
rect 22204 44434 22260 44940
rect 23548 44548 23604 51100
rect 23660 50596 23716 51324
rect 23772 51378 23828 51884
rect 23884 51492 23940 51502
rect 23884 51398 23940 51436
rect 23772 51326 23774 51378
rect 23826 51326 23828 51378
rect 23772 51268 23828 51326
rect 23772 51202 23828 51212
rect 23884 51156 23940 51166
rect 23884 51154 24052 51156
rect 23884 51102 23886 51154
rect 23938 51102 24052 51154
rect 23884 51100 24052 51102
rect 23884 51090 23940 51100
rect 23660 49810 23716 50540
rect 23772 50594 23828 50606
rect 23772 50542 23774 50594
rect 23826 50542 23828 50594
rect 23772 50484 23828 50542
rect 23996 50594 24052 51100
rect 23996 50542 23998 50594
rect 24050 50542 24052 50594
rect 23996 50428 24052 50542
rect 24108 50596 24164 50606
rect 24108 50502 24164 50540
rect 24332 50428 24388 52892
rect 24556 52724 24612 52734
rect 24556 52630 24612 52668
rect 24892 52612 24948 53678
rect 25564 53732 25620 54462
rect 25564 53666 25620 53676
rect 26236 54514 26404 54516
rect 26236 54462 26350 54514
rect 26402 54462 26404 54514
rect 26236 54460 26404 54462
rect 24892 52546 24948 52556
rect 24892 52274 24948 52286
rect 24892 52222 24894 52274
rect 24946 52222 24948 52274
rect 24444 52164 24500 52174
rect 24444 52070 24500 52108
rect 24668 52052 24724 52062
rect 24668 50708 24724 51996
rect 24892 51604 24948 52222
rect 26124 52164 26180 52174
rect 25900 51938 25956 51950
rect 25900 51886 25902 51938
rect 25954 51886 25956 51938
rect 25900 51716 25956 51886
rect 25452 51660 25956 51716
rect 25452 51604 25508 51660
rect 24892 51548 25508 51604
rect 23772 50418 23828 50428
rect 23884 50372 24052 50428
rect 24220 50372 24388 50428
rect 24444 50596 24500 50606
rect 23884 49922 23940 50372
rect 23884 49870 23886 49922
rect 23938 49870 23940 49922
rect 23884 49858 23940 49870
rect 23660 49758 23662 49810
rect 23714 49758 23716 49810
rect 23660 49746 23716 49758
rect 23660 49476 23716 49486
rect 23660 49250 23716 49420
rect 23660 49198 23662 49250
rect 23714 49198 23716 49250
rect 23660 49186 23716 49198
rect 23996 48916 24052 48926
rect 23996 48822 24052 48860
rect 23660 46788 23716 46798
rect 23660 46694 23716 46732
rect 24108 44996 24164 45006
rect 24220 44996 24276 50372
rect 24444 49922 24500 50540
rect 24556 50484 24612 50522
rect 24556 50418 24612 50428
rect 24444 49870 24446 49922
rect 24498 49870 24500 49922
rect 24332 46674 24388 46686
rect 24332 46622 24334 46674
rect 24386 46622 24388 46674
rect 24332 46564 24388 46622
rect 24332 46498 24388 46508
rect 24108 44994 24276 44996
rect 24108 44942 24110 44994
rect 24162 44942 24276 44994
rect 24108 44940 24276 44942
rect 23548 44492 24052 44548
rect 22204 44382 22206 44434
rect 22258 44382 22260 44434
rect 22204 44370 22260 44382
rect 22428 44322 22484 44334
rect 22428 44270 22430 44322
rect 22482 44270 22484 44322
rect 22092 44212 22148 44222
rect 22092 44118 22148 44156
rect 22428 43540 22484 44270
rect 23324 44322 23380 44334
rect 23324 44270 23326 44322
rect 23378 44270 23380 44322
rect 22988 44210 23044 44222
rect 22988 44158 22990 44210
rect 23042 44158 23044 44210
rect 22988 43764 23044 44158
rect 22988 43698 23044 43708
rect 23100 44098 23156 44110
rect 23100 44046 23102 44098
rect 23154 44046 23156 44098
rect 22484 43484 22596 43540
rect 22428 43474 22484 43484
rect 21420 42924 21588 42980
rect 21644 43426 21812 43428
rect 21644 43374 21758 43426
rect 21810 43374 21812 43426
rect 21644 43372 21812 43374
rect 21308 42644 21364 42654
rect 21308 42550 21364 42588
rect 21196 42466 21252 42476
rect 21420 42420 21476 42924
rect 21644 42644 21700 43372
rect 21756 43362 21812 43372
rect 21756 42868 21812 42878
rect 22316 42868 22372 42878
rect 21756 42866 22372 42868
rect 21756 42814 21758 42866
rect 21810 42814 22318 42866
rect 22370 42814 22372 42866
rect 21756 42812 22372 42814
rect 21756 42802 21812 42812
rect 22316 42802 22372 42812
rect 21644 42588 21812 42644
rect 21532 42532 21588 42542
rect 21532 42530 21700 42532
rect 21532 42478 21534 42530
rect 21586 42478 21700 42530
rect 21532 42476 21700 42478
rect 21532 42466 21588 42476
rect 20860 42018 20916 42028
rect 21308 42364 21476 42420
rect 20972 41972 21028 41982
rect 21196 41972 21252 41982
rect 20972 41878 21028 41916
rect 21084 41970 21252 41972
rect 21084 41918 21198 41970
rect 21250 41918 21252 41970
rect 21084 41916 21252 41918
rect 21084 40628 21140 41916
rect 21196 41906 21252 41916
rect 21308 41970 21364 42364
rect 21532 42308 21588 42318
rect 21420 42252 21532 42308
rect 21420 42194 21476 42252
rect 21532 42242 21588 42252
rect 21420 42142 21422 42194
rect 21474 42142 21476 42194
rect 21420 42130 21476 42142
rect 21308 41918 21310 41970
rect 21362 41918 21364 41970
rect 21308 41906 21364 41918
rect 21532 41972 21588 41982
rect 21532 41878 21588 41916
rect 21644 41748 21700 42476
rect 21756 42530 21812 42588
rect 22540 42642 22596 43484
rect 22652 43428 22708 43438
rect 22652 42978 22708 43372
rect 22652 42926 22654 42978
rect 22706 42926 22708 42978
rect 22652 42914 22708 42926
rect 23100 42868 23156 44046
rect 23324 43540 23380 44270
rect 23324 43474 23380 43484
rect 23884 43428 23940 43438
rect 23884 43334 23940 43372
rect 23100 42802 23156 42812
rect 22540 42590 22542 42642
rect 22594 42590 22596 42642
rect 22540 42578 22596 42590
rect 23548 42756 23604 42766
rect 21756 42478 21758 42530
rect 21810 42478 21812 42530
rect 21756 42466 21812 42478
rect 21868 42532 21924 42542
rect 21868 42308 21924 42476
rect 21756 42252 21924 42308
rect 23212 42532 23268 42542
rect 23548 42532 23604 42700
rect 23212 42530 23604 42532
rect 23212 42478 23214 42530
rect 23266 42478 23604 42530
rect 23212 42476 23604 42478
rect 21756 41972 21812 42252
rect 22092 42196 22148 42206
rect 22092 42102 22148 42140
rect 23212 42196 23268 42476
rect 23212 42130 23268 42140
rect 21756 41906 21812 41916
rect 21420 41692 21700 41748
rect 21420 41298 21476 41692
rect 21420 41246 21422 41298
rect 21474 41246 21476 41298
rect 21420 41234 21476 41246
rect 22092 41300 22148 41310
rect 22428 41300 22484 41310
rect 22148 41244 22372 41300
rect 22092 41234 22148 41244
rect 21980 41188 22036 41198
rect 20972 40572 21140 40628
rect 21308 40962 21364 40974
rect 21532 40964 21588 40974
rect 21308 40910 21310 40962
rect 21362 40910 21364 40962
rect 20860 40402 20916 40414
rect 20860 40350 20862 40402
rect 20914 40350 20916 40402
rect 20860 39508 20916 40350
rect 20972 40290 21028 40572
rect 20972 40238 20974 40290
rect 21026 40238 21028 40290
rect 20972 40226 21028 40238
rect 21084 40404 21140 40414
rect 21308 40404 21364 40910
rect 21084 40402 21364 40404
rect 21084 40350 21086 40402
rect 21138 40350 21364 40402
rect 21084 40348 21364 40350
rect 21420 40962 21588 40964
rect 21420 40910 21534 40962
rect 21586 40910 21588 40962
rect 21420 40908 21588 40910
rect 21084 39844 21140 40348
rect 21084 39778 21140 39788
rect 20860 39452 21364 39508
rect 20748 39340 21252 39396
rect 21084 39060 21140 39070
rect 20300 38836 20356 38846
rect 20860 38836 20916 38846
rect 20300 38742 20356 38780
rect 20412 38834 20916 38836
rect 20412 38782 20862 38834
rect 20914 38782 20916 38834
rect 20412 38780 20916 38782
rect 20188 38434 20244 38444
rect 20412 38500 20468 38780
rect 20860 38770 20916 38780
rect 21084 38834 21140 39004
rect 21084 38782 21086 38834
rect 21138 38782 21140 38834
rect 21084 38770 21140 38782
rect 20636 38612 20692 38622
rect 20636 38518 20692 38556
rect 20412 38434 20468 38444
rect 21196 38500 21252 39340
rect 21196 38434 21252 38444
rect 19740 37998 19742 38050
rect 19794 37998 19796 38050
rect 19740 37986 19796 37998
rect 20524 38388 20580 38398
rect 20524 38274 20580 38332
rect 20524 38222 20526 38274
rect 20578 38222 20580 38274
rect 19964 37938 20020 37950
rect 19964 37886 19966 37938
rect 20018 37886 20020 37938
rect 19964 37828 20020 37886
rect 20524 37940 20580 38222
rect 20636 38276 20692 38286
rect 20636 38182 20692 38220
rect 21308 38052 21364 39452
rect 21420 38276 21476 40908
rect 21532 40898 21588 40908
rect 21756 40962 21812 40974
rect 21756 40910 21758 40962
rect 21810 40910 21812 40962
rect 21756 40628 21812 40910
rect 21756 40562 21812 40572
rect 21644 40516 21700 40526
rect 21532 39508 21588 39518
rect 21532 39414 21588 39452
rect 21532 38948 21588 38958
rect 21644 38948 21700 40460
rect 21532 38946 21700 38948
rect 21532 38894 21534 38946
rect 21586 38894 21700 38946
rect 21532 38892 21700 38894
rect 21756 39844 21812 39854
rect 21756 38946 21812 39788
rect 21756 38894 21758 38946
rect 21810 38894 21812 38946
rect 21532 38724 21588 38892
rect 21756 38882 21812 38894
rect 21868 39508 21924 39518
rect 21868 38834 21924 39452
rect 21868 38782 21870 38834
rect 21922 38782 21924 38834
rect 21868 38770 21924 38782
rect 21980 38668 22036 41132
rect 22316 40740 22372 41244
rect 22428 41206 22484 41244
rect 23212 41300 23268 41310
rect 22316 40626 22372 40684
rect 22316 40574 22318 40626
rect 22370 40574 22372 40626
rect 22316 40562 22372 40574
rect 23212 40628 23268 41244
rect 23212 40534 23268 40572
rect 23324 40740 23380 40750
rect 22540 40404 22596 40414
rect 22540 40310 22596 40348
rect 23212 40290 23268 40302
rect 23212 40238 23214 40290
rect 23266 40238 23268 40290
rect 22988 40178 23044 40190
rect 22988 40126 22990 40178
rect 23042 40126 23044 40178
rect 22988 39844 23044 40126
rect 22988 39778 23044 39788
rect 22092 39620 22148 39630
rect 22148 39564 22372 39620
rect 22092 39526 22148 39564
rect 22092 38948 22148 38958
rect 22092 38834 22148 38892
rect 22092 38782 22094 38834
rect 22146 38782 22148 38834
rect 22092 38770 22148 38782
rect 22316 38668 22372 39564
rect 22876 38834 22932 38846
rect 22876 38782 22878 38834
rect 22930 38782 22932 38834
rect 21532 38658 21588 38668
rect 21868 38612 22036 38668
rect 22092 38612 22372 38668
rect 22764 38722 22820 38734
rect 22764 38670 22766 38722
rect 22818 38670 22820 38722
rect 21532 38500 21588 38510
rect 21588 38444 21812 38500
rect 21532 38434 21588 38444
rect 21420 38220 21588 38276
rect 21084 37996 21364 38052
rect 20636 37940 20692 37950
rect 20524 37884 20636 37940
rect 20692 37884 20916 37940
rect 20636 37846 20692 37884
rect 19628 37772 20020 37828
rect 20188 37828 20244 37838
rect 19628 37156 19684 37772
rect 20188 37734 20244 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20524 37604 20580 37614
rect 19852 37492 19908 37502
rect 19852 37268 19908 37436
rect 20524 37378 20580 37548
rect 20524 37326 20526 37378
rect 20578 37326 20580 37378
rect 20524 37314 20580 37326
rect 20748 37492 20804 37502
rect 20300 37268 20356 37278
rect 19852 37266 20020 37268
rect 19852 37214 19854 37266
rect 19906 37214 20020 37266
rect 19852 37212 20020 37214
rect 19852 37202 19908 37212
rect 19628 37100 19796 37156
rect 19628 36932 19684 36942
rect 19628 36482 19684 36876
rect 19628 36430 19630 36482
rect 19682 36430 19684 36482
rect 19628 36418 19684 36430
rect 19740 36260 19796 37100
rect 19964 36820 20020 37212
rect 20300 37174 20356 37212
rect 19964 36370 20020 36764
rect 19964 36318 19966 36370
rect 20018 36318 20020 36370
rect 19964 36306 20020 36318
rect 20188 37154 20244 37166
rect 20188 37102 20190 37154
rect 20242 37102 20244 37154
rect 19292 35298 19348 35308
rect 19404 36204 19572 36260
rect 19628 36204 19796 36260
rect 19292 35140 19348 35150
rect 19180 35138 19348 35140
rect 19180 35086 19294 35138
rect 19346 35086 19348 35138
rect 19180 35084 19348 35086
rect 19292 35074 19348 35084
rect 19292 34356 19348 34366
rect 19404 34356 19460 36204
rect 19628 36036 19684 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19628 35970 19684 35980
rect 19516 35924 19572 35934
rect 19516 35830 19572 35868
rect 19852 35028 19908 35038
rect 19628 35026 19908 35028
rect 19628 34974 19854 35026
rect 19906 34974 19908 35026
rect 19628 34972 19908 34974
rect 20188 35028 20244 37102
rect 20412 37044 20468 37054
rect 20412 36482 20468 36988
rect 20412 36430 20414 36482
rect 20466 36430 20468 36482
rect 20412 36418 20468 36430
rect 20748 36482 20804 37436
rect 20860 37044 20916 37884
rect 20860 36978 20916 36988
rect 20748 36430 20750 36482
rect 20802 36430 20804 36482
rect 20748 36418 20804 36430
rect 20636 36372 20692 36382
rect 20636 36278 20692 36316
rect 20636 35700 20692 35710
rect 20636 35140 20692 35644
rect 20860 35588 20916 35598
rect 20412 35084 20692 35140
rect 20748 35364 20804 35374
rect 20188 34972 20356 35028
rect 19516 34916 19572 34926
rect 19516 34822 19572 34860
rect 19292 34354 19460 34356
rect 19292 34302 19294 34354
rect 19346 34302 19460 34354
rect 19292 34300 19460 34302
rect 19292 34290 19348 34300
rect 18956 34130 19572 34132
rect 18956 34078 18958 34130
rect 19010 34078 19572 34130
rect 18956 34076 19572 34078
rect 18956 34066 19012 34076
rect 19404 33908 19460 33918
rect 18844 33182 18846 33234
rect 18898 33182 18900 33234
rect 18844 33170 18900 33182
rect 18956 33906 19460 33908
rect 18956 33854 19406 33906
rect 19458 33854 19460 33906
rect 18956 33852 19460 33854
rect 18284 32946 18340 32956
rect 18508 32956 18788 33012
rect 18172 32610 18228 32620
rect 17948 32452 18004 32462
rect 17948 32358 18004 32396
rect 17836 31838 17838 31890
rect 17890 31838 17892 31890
rect 17388 30098 17444 30828
rect 17836 30324 17892 31838
rect 18396 31780 18452 31790
rect 18284 31444 18340 31454
rect 18060 31220 18116 31230
rect 18060 30994 18116 31164
rect 18060 30942 18062 30994
rect 18114 30942 18116 30994
rect 18060 30930 18116 30942
rect 18284 30548 18340 31388
rect 18396 31218 18452 31724
rect 18396 31166 18398 31218
rect 18450 31166 18452 31218
rect 18396 30996 18452 31166
rect 18396 30930 18452 30940
rect 18396 30548 18452 30558
rect 18284 30492 18396 30548
rect 18396 30434 18452 30492
rect 18396 30382 18398 30434
rect 18450 30382 18452 30434
rect 18396 30370 18452 30382
rect 17612 30268 17892 30324
rect 18508 30324 18564 32956
rect 18956 32900 19012 33852
rect 19404 33842 19460 33852
rect 19516 33684 19572 34076
rect 19628 33906 19684 34972
rect 19852 34962 19908 34972
rect 19964 34916 20020 34926
rect 19964 34802 20020 34860
rect 19964 34750 19966 34802
rect 20018 34750 20020 34802
rect 19964 34738 20020 34750
rect 20188 34802 20244 34814
rect 20188 34750 20190 34802
rect 20242 34750 20244 34802
rect 20188 34692 20244 34750
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20188 34356 20244 34636
rect 20188 34290 20244 34300
rect 19852 34132 19908 34142
rect 20300 34132 20356 34972
rect 19852 34130 20356 34132
rect 19852 34078 19854 34130
rect 19906 34078 20356 34130
rect 19852 34076 20356 34078
rect 19852 34066 19908 34076
rect 19628 33854 19630 33906
rect 19682 33854 19684 33906
rect 19628 33842 19684 33854
rect 19740 33908 19796 33918
rect 20076 33908 20132 33918
rect 19516 33628 19684 33684
rect 19292 33460 19348 33470
rect 19180 33404 19292 33460
rect 19180 33346 19236 33404
rect 19292 33394 19348 33404
rect 19180 33294 19182 33346
rect 19234 33294 19236 33346
rect 19180 33282 19236 33294
rect 18732 32844 19012 32900
rect 19068 33236 19124 33246
rect 19068 33122 19124 33180
rect 19068 33070 19070 33122
rect 19122 33070 19124 33122
rect 18620 32676 18676 32714
rect 18620 32610 18676 32620
rect 18620 32452 18676 32462
rect 18620 32004 18676 32396
rect 18620 31666 18676 31948
rect 18620 31614 18622 31666
rect 18674 31614 18676 31666
rect 18620 31602 18676 31614
rect 18732 31444 18788 32844
rect 17500 30212 17556 30222
rect 17500 30118 17556 30156
rect 17388 30046 17390 30098
rect 17442 30046 17444 30098
rect 17388 30034 17444 30046
rect 17500 29428 17556 29438
rect 17500 29334 17556 29372
rect 17276 29202 17332 29214
rect 17612 29204 17668 30268
rect 18508 30258 18564 30268
rect 18620 31388 18788 31444
rect 18844 32674 18900 32686
rect 18844 32622 18846 32674
rect 18898 32622 18900 32674
rect 18844 32340 18900 32622
rect 19068 32676 19124 33070
rect 19180 33124 19236 33134
rect 19180 32786 19236 33068
rect 19292 33122 19348 33134
rect 19292 33070 19294 33122
rect 19346 33070 19348 33122
rect 19292 33012 19348 33070
rect 19292 32900 19348 32956
rect 19292 32844 19572 32900
rect 19180 32734 19182 32786
rect 19234 32734 19236 32786
rect 19180 32722 19236 32734
rect 19516 32788 19572 32844
rect 19516 32722 19572 32732
rect 19404 32676 19460 32686
rect 19068 32610 19124 32620
rect 19292 32674 19460 32676
rect 19292 32622 19406 32674
rect 19458 32622 19460 32674
rect 19292 32620 19460 32622
rect 18956 32452 19012 32462
rect 19292 32452 19348 32620
rect 19404 32610 19460 32620
rect 18956 32450 19348 32452
rect 18956 32398 18958 32450
rect 19010 32398 19348 32450
rect 18956 32396 19348 32398
rect 19516 32562 19572 32574
rect 19516 32510 19518 32562
rect 19570 32510 19572 32562
rect 18956 32386 19012 32396
rect 18172 30212 18228 30222
rect 18620 30212 18676 31388
rect 18228 30156 18452 30212
rect 18172 30118 18228 30156
rect 17836 30098 17892 30110
rect 17836 30046 17838 30098
rect 17890 30046 17892 30098
rect 17836 29876 17892 30046
rect 17836 29810 17892 29820
rect 17948 29986 18004 29998
rect 17948 29934 17950 29986
rect 18002 29934 18004 29986
rect 17948 29652 18004 29934
rect 18284 29652 18340 29662
rect 17948 29586 18004 29596
rect 18060 29596 18284 29652
rect 17276 29150 17278 29202
rect 17330 29150 17332 29202
rect 17052 28644 17108 28654
rect 17052 28550 17108 28588
rect 17276 28642 17332 29150
rect 17276 28590 17278 28642
rect 17330 28590 17332 28642
rect 16716 28530 16884 28532
rect 16716 28478 16718 28530
rect 16770 28478 16884 28530
rect 16716 28476 16884 28478
rect 17276 28532 17332 28590
rect 16604 28084 16660 28094
rect 16492 28082 16660 28084
rect 16492 28030 16606 28082
rect 16658 28030 16660 28082
rect 16492 28028 16660 28030
rect 16604 28018 16660 28028
rect 16716 27970 16772 28476
rect 17276 28466 17332 28476
rect 17388 29148 17668 29204
rect 17948 29428 18004 29438
rect 18060 29428 18116 29596
rect 18284 29586 18340 29596
rect 17948 29426 18116 29428
rect 17948 29374 17950 29426
rect 18002 29374 18116 29426
rect 17948 29372 18116 29374
rect 17948 29202 18004 29372
rect 17948 29150 17950 29202
rect 18002 29150 18004 29202
rect 16716 27918 16718 27970
rect 16770 27918 16772 27970
rect 16716 27906 16772 27918
rect 16268 27582 16270 27634
rect 16322 27582 16324 27634
rect 16268 27570 16324 27582
rect 16380 27748 16436 27758
rect 16380 26516 16436 27692
rect 17388 26908 17444 29148
rect 17948 29138 18004 29150
rect 18060 28812 18340 28868
rect 17724 28644 17780 28654
rect 18060 28644 18116 28812
rect 17780 28588 18116 28644
rect 17724 28578 17780 28588
rect 17724 28420 17780 28430
rect 17724 28326 17780 28364
rect 17836 28418 17892 28430
rect 17836 28366 17838 28418
rect 17890 28366 17892 28418
rect 17500 27860 17556 27870
rect 17500 27858 17780 27860
rect 17500 27806 17502 27858
rect 17554 27806 17780 27858
rect 17500 27804 17780 27806
rect 17500 27794 17556 27804
rect 17724 26908 17780 27804
rect 17836 27076 17892 28366
rect 17948 28420 18004 28430
rect 17948 28326 18004 28364
rect 17948 27188 18004 27198
rect 18060 27188 18116 28588
rect 18172 28644 18228 28654
rect 18172 27970 18228 28588
rect 18284 28642 18340 28812
rect 18396 28754 18452 30156
rect 18620 30118 18676 30156
rect 18732 30994 18788 31006
rect 18732 30942 18734 30994
rect 18786 30942 18788 30994
rect 18620 29652 18676 29662
rect 18620 29558 18676 29596
rect 18396 28702 18398 28754
rect 18450 28702 18452 28754
rect 18396 28690 18452 28702
rect 18732 28756 18788 30942
rect 18732 28690 18788 28700
rect 18284 28590 18286 28642
rect 18338 28590 18340 28642
rect 18284 28578 18340 28590
rect 18620 28532 18676 28542
rect 18844 28532 18900 32284
rect 19068 31218 19124 32396
rect 19516 31668 19572 32510
rect 19068 31166 19070 31218
rect 19122 31166 19124 31218
rect 19068 31154 19124 31166
rect 19292 31612 19572 31668
rect 19628 31780 19684 33628
rect 19740 33346 19796 33852
rect 19964 33906 20132 33908
rect 19964 33854 20078 33906
rect 20130 33854 20132 33906
rect 19964 33852 20132 33854
rect 19964 33570 20020 33852
rect 20076 33842 20132 33852
rect 19964 33518 19966 33570
rect 20018 33518 20020 33570
rect 19964 33460 20020 33518
rect 20188 33570 20244 34076
rect 20300 33908 20356 33918
rect 20300 33814 20356 33852
rect 20188 33518 20190 33570
rect 20242 33518 20244 33570
rect 20188 33506 20244 33518
rect 19964 33394 20020 33404
rect 20300 33460 20356 33470
rect 20300 33366 20356 33404
rect 19740 33294 19742 33346
rect 19794 33294 19796 33346
rect 19740 33282 19796 33294
rect 20412 33236 20468 35084
rect 20748 34916 20804 35308
rect 20300 33180 20468 33236
rect 20524 34860 20804 34916
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20300 31890 20356 33180
rect 20524 32676 20580 34860
rect 20636 34692 20692 34702
rect 20636 33570 20692 34636
rect 20748 34020 20804 34030
rect 20748 33926 20804 33964
rect 20636 33518 20638 33570
rect 20690 33518 20692 33570
rect 20636 33506 20692 33518
rect 20748 33572 20804 33582
rect 20860 33572 20916 35532
rect 21084 35028 21140 37996
rect 21308 37828 21364 37838
rect 21364 37772 21476 37828
rect 21308 37734 21364 37772
rect 21308 37268 21364 37278
rect 21420 37268 21476 37772
rect 21532 37492 21588 38220
rect 21644 37828 21700 37838
rect 21644 37734 21700 37772
rect 21532 37436 21700 37492
rect 21532 37268 21588 37278
rect 21420 37266 21588 37268
rect 21420 37214 21534 37266
rect 21586 37214 21588 37266
rect 21420 37212 21588 37214
rect 21308 37174 21364 37212
rect 21532 37202 21588 37212
rect 21532 36708 21588 36718
rect 21420 36596 21476 36606
rect 21420 36502 21476 36540
rect 21532 36482 21588 36652
rect 21532 36430 21534 36482
rect 21586 36430 21588 36482
rect 21532 36418 21588 36430
rect 21308 36260 21364 36270
rect 21196 35588 21252 35598
rect 21196 35494 21252 35532
rect 20804 33516 20916 33572
rect 20972 34972 21140 35028
rect 20748 33506 20804 33516
rect 20748 33234 20804 33246
rect 20748 33182 20750 33234
rect 20802 33182 20804 33234
rect 20748 33124 20804 33182
rect 20524 32620 20692 32676
rect 20300 31838 20302 31890
rect 20354 31838 20356 31890
rect 20300 31826 20356 31838
rect 20412 32562 20468 32574
rect 20412 32510 20414 32562
rect 20466 32510 20468 32562
rect 19740 31780 19796 31790
rect 19628 31778 19796 31780
rect 19628 31726 19742 31778
rect 19794 31726 19796 31778
rect 19628 31724 19796 31726
rect 19628 31668 19684 31724
rect 19740 31714 19796 31724
rect 20412 31780 20468 32510
rect 20412 31686 20468 31724
rect 20524 32450 20580 32462
rect 20524 32398 20526 32450
rect 20578 32398 20580 32450
rect 19292 30994 19348 31612
rect 19628 31602 19684 31612
rect 20188 31556 20244 31566
rect 20524 31556 20580 32398
rect 20244 31500 20580 31556
rect 20188 31462 20244 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19852 31106 19908 31118
rect 19852 31054 19854 31106
rect 19906 31054 19908 31106
rect 19292 30942 19294 30994
rect 19346 30942 19348 30994
rect 18956 30324 19012 30334
rect 18956 30210 19012 30268
rect 18956 30158 18958 30210
rect 19010 30158 19012 30210
rect 18956 30146 19012 30158
rect 19068 30212 19124 30222
rect 18676 28476 18900 28532
rect 18956 29652 19012 29662
rect 18956 28642 19012 29596
rect 19068 29538 19124 30156
rect 19292 29876 19348 30942
rect 19628 30996 19684 31006
rect 19628 30902 19684 30940
rect 19404 30884 19460 30894
rect 19404 30790 19460 30828
rect 19852 30100 19908 31054
rect 20188 30994 20244 31006
rect 20188 30942 20190 30994
rect 20242 30942 20244 30994
rect 20188 30660 20244 30942
rect 20524 30882 20580 30894
rect 20524 30830 20526 30882
rect 20578 30830 20580 30882
rect 20524 30772 20580 30830
rect 20524 30706 20580 30716
rect 20188 30594 20244 30604
rect 20636 30548 20692 32620
rect 20748 32340 20804 33068
rect 20860 32676 20916 32686
rect 20972 32676 21028 34972
rect 21308 34914 21364 36204
rect 21644 35812 21700 37436
rect 21308 34862 21310 34914
rect 21362 34862 21364 34914
rect 21084 34804 21140 34814
rect 21084 34242 21140 34748
rect 21084 34190 21086 34242
rect 21138 34190 21140 34242
rect 21084 34178 21140 34190
rect 21308 34130 21364 34862
rect 21532 35756 21700 35812
rect 21420 34804 21476 34814
rect 21420 34710 21476 34748
rect 21308 34078 21310 34130
rect 21362 34078 21364 34130
rect 21308 34066 21364 34078
rect 21532 33684 21588 35756
rect 21644 35588 21700 35598
rect 21644 35494 21700 35532
rect 21644 34690 21700 34702
rect 21644 34638 21646 34690
rect 21698 34638 21700 34690
rect 21644 34580 21700 34638
rect 21644 34514 21700 34524
rect 21644 34356 21700 34366
rect 21644 34262 21700 34300
rect 21308 33628 21588 33684
rect 20860 32674 21028 32676
rect 20860 32622 20862 32674
rect 20914 32622 21028 32674
rect 20860 32620 21028 32622
rect 20860 32610 20916 32620
rect 20972 32564 21028 32620
rect 20972 32498 21028 32508
rect 21196 33572 21252 33582
rect 21196 32450 21252 33516
rect 21196 32398 21198 32450
rect 21250 32398 21252 32450
rect 21196 32386 21252 32398
rect 21308 32562 21364 33628
rect 21756 33460 21812 38444
rect 21868 34804 21924 38612
rect 21980 37268 22036 37278
rect 21980 37174 22036 37212
rect 21980 36484 22036 36494
rect 22092 36484 22148 38612
rect 22204 37940 22260 37950
rect 22204 37846 22260 37884
rect 22540 37940 22596 37950
rect 22540 37846 22596 37884
rect 22316 37828 22372 37838
rect 21980 36482 22148 36484
rect 21980 36430 21982 36482
rect 22034 36430 22148 36482
rect 21980 36428 22148 36430
rect 22204 37268 22260 37278
rect 22316 37268 22372 37772
rect 22764 37716 22820 38670
rect 22764 37650 22820 37660
rect 22540 37380 22596 37390
rect 22540 37286 22596 37324
rect 22204 37266 22372 37268
rect 22204 37214 22206 37266
rect 22258 37214 22372 37266
rect 22204 37212 22372 37214
rect 22764 37266 22820 37278
rect 22764 37214 22766 37266
rect 22818 37214 22820 37266
rect 21980 36418 22036 36428
rect 22204 35588 22260 37212
rect 22428 37154 22484 37166
rect 22428 37102 22430 37154
rect 22482 37102 22484 37154
rect 22428 35812 22484 37102
rect 22764 36596 22820 37214
rect 22876 37268 22932 38782
rect 23212 38836 23268 40238
rect 23100 37492 23156 37502
rect 23212 37492 23268 38780
rect 23100 37490 23268 37492
rect 23100 37438 23102 37490
rect 23154 37438 23268 37490
rect 23100 37436 23268 37438
rect 23100 37426 23156 37436
rect 23324 37378 23380 40684
rect 23436 40180 23492 40190
rect 23436 39618 23492 40124
rect 23436 39566 23438 39618
rect 23490 39566 23492 39618
rect 23436 39554 23492 39566
rect 23772 39506 23828 39518
rect 23772 39454 23774 39506
rect 23826 39454 23828 39506
rect 23660 39394 23716 39406
rect 23660 39342 23662 39394
rect 23714 39342 23716 39394
rect 23548 38948 23604 38958
rect 23548 38854 23604 38892
rect 23660 38612 23716 39342
rect 23660 38546 23716 38556
rect 23324 37326 23326 37378
rect 23378 37326 23380 37378
rect 22876 37212 23156 37268
rect 22988 37044 23044 37054
rect 22764 36530 22820 36540
rect 22876 37042 23044 37044
rect 22876 36990 22990 37042
rect 23042 36990 23044 37042
rect 22876 36988 23044 36990
rect 22652 36370 22708 36382
rect 22652 36318 22654 36370
rect 22706 36318 22708 36370
rect 22540 35924 22596 35934
rect 22540 35830 22596 35868
rect 22428 35746 22484 35756
rect 22652 35700 22708 36318
rect 22764 36372 22820 36382
rect 22764 36278 22820 36316
rect 22204 35522 22260 35532
rect 22540 35588 22596 35598
rect 22316 35474 22372 35486
rect 22316 35422 22318 35474
rect 22370 35422 22372 35474
rect 22204 35028 22260 35038
rect 22316 35028 22372 35422
rect 22204 35026 22372 35028
rect 22204 34974 22206 35026
rect 22258 34974 22372 35026
rect 22204 34972 22372 34974
rect 22428 35364 22484 35374
rect 21868 34748 22148 34804
rect 21532 33404 21812 33460
rect 21980 34580 22036 34590
rect 21420 33124 21476 33134
rect 21420 33030 21476 33068
rect 21308 32510 21310 32562
rect 21362 32510 21364 32562
rect 21308 32452 21364 32510
rect 21308 32386 21364 32396
rect 20748 32274 20804 32284
rect 21196 31892 21252 31902
rect 20748 31780 20804 31790
rect 20748 31686 20804 31724
rect 21084 31668 21140 31678
rect 21084 31220 21140 31612
rect 21084 31126 21140 31164
rect 21196 31108 21252 31836
rect 21420 31778 21476 31790
rect 21420 31726 21422 31778
rect 21474 31726 21476 31778
rect 20972 30996 21028 31006
rect 20972 30902 21028 30940
rect 21196 30994 21252 31052
rect 21196 30942 21198 30994
rect 21250 30942 21252 30994
rect 19292 29810 19348 29820
rect 19516 29986 19572 29998
rect 19852 29988 19908 30044
rect 19516 29934 19518 29986
rect 19570 29934 19572 29986
rect 19068 29486 19070 29538
rect 19122 29486 19124 29538
rect 19068 29474 19124 29486
rect 19180 29202 19236 29214
rect 19180 29150 19182 29202
rect 19234 29150 19236 29202
rect 18956 28590 18958 28642
rect 19010 28590 19012 28642
rect 18620 28438 18676 28476
rect 18172 27918 18174 27970
rect 18226 27918 18228 27970
rect 18172 27906 18228 27918
rect 17948 27186 18116 27188
rect 17948 27134 17950 27186
rect 18002 27134 18116 27186
rect 17948 27132 18116 27134
rect 18732 27188 18788 27198
rect 18956 27188 19012 28590
rect 19068 28644 19124 28654
rect 19068 28550 19124 28588
rect 19180 28642 19236 29150
rect 19516 28756 19572 29934
rect 19516 28690 19572 28700
rect 19628 29932 19908 29988
rect 20524 30492 20692 30548
rect 19180 28590 19182 28642
rect 19234 28590 19236 28642
rect 19180 28578 19236 28590
rect 19404 28644 19460 28654
rect 19404 28550 19460 28588
rect 19628 28196 19684 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20524 29650 20580 30492
rect 21196 30324 21252 30942
rect 21196 30258 21252 30268
rect 21308 31220 21364 31230
rect 20524 29598 20526 29650
rect 20578 29598 20580 29650
rect 19964 29540 20020 29550
rect 19964 28754 20020 29484
rect 20524 29540 20580 29598
rect 21308 29652 21364 31164
rect 21420 30994 21476 31726
rect 21420 30942 21422 30994
rect 21474 30942 21476 30994
rect 21420 30434 21476 30942
rect 21532 30996 21588 33404
rect 21644 33348 21700 33404
rect 21644 33282 21700 33292
rect 21980 33346 22036 34524
rect 22092 33572 22148 34748
rect 22204 34356 22260 34972
rect 22428 34914 22484 35308
rect 22428 34862 22430 34914
rect 22482 34862 22484 34914
rect 22428 34850 22484 34862
rect 22260 34300 22372 34356
rect 22204 34290 22260 34300
rect 22092 33506 22148 33516
rect 21980 33294 21982 33346
rect 22034 33294 22036 33346
rect 21980 33282 22036 33294
rect 22316 33346 22372 34300
rect 22316 33294 22318 33346
rect 22370 33294 22372 33346
rect 22316 33282 22372 33294
rect 21756 33236 21812 33246
rect 21756 33142 21812 33180
rect 22540 33234 22596 35532
rect 22652 35586 22708 35644
rect 22652 35534 22654 35586
rect 22706 35534 22708 35586
rect 22652 35522 22708 35534
rect 22652 35252 22708 35262
rect 22652 34132 22708 35196
rect 22652 34038 22708 34076
rect 22652 33796 22708 33806
rect 22652 33570 22708 33740
rect 22652 33518 22654 33570
rect 22706 33518 22708 33570
rect 22652 33506 22708 33518
rect 22540 33182 22542 33234
rect 22594 33182 22596 33234
rect 22540 33170 22596 33182
rect 22092 33124 22148 33134
rect 21868 32674 21924 32686
rect 21868 32622 21870 32674
rect 21922 32622 21924 32674
rect 21644 32116 21700 32126
rect 21644 31778 21700 32060
rect 21868 31892 21924 32622
rect 21980 32452 22036 32462
rect 21980 32358 22036 32396
rect 21868 31826 21924 31836
rect 21980 32116 22036 32126
rect 21644 31726 21646 31778
rect 21698 31726 21700 31778
rect 21644 31714 21700 31726
rect 21980 31780 22036 32060
rect 22092 32002 22148 33068
rect 22092 31950 22094 32002
rect 22146 31950 22148 32002
rect 22092 31938 22148 31950
rect 22204 32564 22260 32574
rect 21980 31724 22148 31780
rect 21644 30996 21700 31006
rect 21532 30994 22036 30996
rect 21532 30942 21646 30994
rect 21698 30942 22036 30994
rect 21532 30940 22036 30942
rect 21644 30930 21700 30940
rect 21420 30382 21422 30434
rect 21474 30382 21476 30434
rect 21420 30370 21476 30382
rect 21868 30772 21924 30782
rect 21532 30212 21588 30222
rect 21532 30118 21588 30156
rect 21420 29988 21476 29998
rect 21420 29986 21588 29988
rect 21420 29934 21422 29986
rect 21474 29934 21588 29986
rect 21420 29932 21588 29934
rect 21420 29922 21476 29932
rect 21308 29586 21364 29596
rect 20524 29474 20580 29484
rect 20860 29540 20916 29550
rect 20860 29446 20916 29484
rect 19964 28702 19966 28754
rect 20018 28702 20020 28754
rect 19964 28644 20020 28702
rect 19964 28578 20020 28588
rect 20300 29316 20356 29326
rect 20300 28644 20356 29260
rect 20972 29316 21028 29326
rect 20972 29314 21476 29316
rect 20972 29262 20974 29314
rect 21026 29262 21476 29314
rect 20972 29260 21476 29262
rect 20972 29250 21028 29260
rect 20636 28756 20692 28766
rect 20300 28642 20580 28644
rect 20300 28590 20302 28642
rect 20354 28590 20580 28642
rect 20300 28588 20580 28590
rect 20300 28578 20356 28588
rect 20188 28532 20244 28542
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 28130 19684 28140
rect 20188 27748 20244 28476
rect 20300 27748 20356 27758
rect 20188 27746 20356 27748
rect 20188 27694 20302 27746
rect 20354 27694 20356 27746
rect 20188 27692 20356 27694
rect 20524 27748 20580 28588
rect 20636 28530 20692 28700
rect 20636 28478 20638 28530
rect 20690 28478 20692 28530
rect 20636 28466 20692 28478
rect 21420 28642 21476 29260
rect 21532 28756 21588 29932
rect 21532 28690 21588 28700
rect 21420 28590 21422 28642
rect 21474 28590 21476 28642
rect 21420 28532 21476 28590
rect 21868 28644 21924 30716
rect 21980 30210 22036 30940
rect 21980 30158 21982 30210
rect 22034 30158 22036 30210
rect 21980 30146 22036 30158
rect 22092 29652 22148 31724
rect 22204 30882 22260 32508
rect 22428 32562 22484 32574
rect 22428 32510 22430 32562
rect 22482 32510 22484 32562
rect 22428 31892 22484 32510
rect 22428 31826 22484 31836
rect 22540 31780 22596 31790
rect 22540 31686 22596 31724
rect 22652 31668 22708 31678
rect 22652 31574 22708 31612
rect 22876 31668 22932 36988
rect 22988 36978 23044 36988
rect 22988 36820 23044 36830
rect 22988 36482 23044 36764
rect 22988 36430 22990 36482
rect 23042 36430 23044 36482
rect 22988 36418 23044 36430
rect 22988 35252 23044 35262
rect 23100 35252 23156 37212
rect 23324 35924 23380 37326
rect 23436 37940 23492 37950
rect 23436 36484 23492 37884
rect 23660 37938 23716 37950
rect 23660 37886 23662 37938
rect 23714 37886 23716 37938
rect 23660 36484 23716 37886
rect 23772 37940 23828 39454
rect 23996 38668 24052 44492
rect 24108 43652 24164 44940
rect 24444 44324 24500 49870
rect 24668 48130 24724 50652
rect 25452 51490 25508 51548
rect 25452 51438 25454 51490
rect 25506 51438 25508 51490
rect 25340 50482 25396 50494
rect 25340 50430 25342 50482
rect 25394 50430 25396 50482
rect 25340 50428 25396 50430
rect 24780 50372 25396 50428
rect 24780 49922 24836 50372
rect 24780 49870 24782 49922
rect 24834 49870 24836 49922
rect 24780 49858 24836 49870
rect 25340 49588 25396 50372
rect 25452 49924 25508 51438
rect 25564 51490 25620 51502
rect 25564 51438 25566 51490
rect 25618 51438 25620 51490
rect 25564 51380 25620 51438
rect 25620 51324 25732 51380
rect 25564 51314 25620 51324
rect 25564 51156 25620 51166
rect 25564 51062 25620 51100
rect 25564 50820 25620 50830
rect 25676 50820 25732 51324
rect 25564 50818 25732 50820
rect 25564 50766 25566 50818
rect 25618 50766 25732 50818
rect 25564 50764 25732 50766
rect 25564 50754 25620 50764
rect 25452 49858 25508 49868
rect 25340 49522 25396 49532
rect 25676 49026 25732 50764
rect 25900 50820 25956 50830
rect 26124 50820 26180 52108
rect 26236 50932 26292 54460
rect 26348 54450 26404 54460
rect 26684 54402 26740 56924
rect 26908 55468 26964 59200
rect 26908 55412 27188 55468
rect 26684 54350 26686 54402
rect 26738 54350 26740 54402
rect 26684 54338 26740 54350
rect 27132 53618 27188 55412
rect 27356 55412 27412 59200
rect 27468 56084 27524 56094
rect 27468 55970 27524 56028
rect 27468 55918 27470 55970
rect 27522 55918 27524 55970
rect 27468 55906 27524 55918
rect 28252 55468 28308 59200
rect 28700 56642 28756 59200
rect 28700 56590 28702 56642
rect 28754 56590 28756 56642
rect 28700 56578 28756 56590
rect 29372 56642 29428 56654
rect 29372 56590 29374 56642
rect 29426 56590 29428 56642
rect 28700 56084 28756 56094
rect 28700 55990 28756 56028
rect 29372 55970 29428 56590
rect 29372 55918 29374 55970
rect 29426 55918 29428 55970
rect 29372 55906 29428 55918
rect 28588 55748 28644 55758
rect 29596 55748 29652 59200
rect 30044 56308 30100 59200
rect 30044 56242 30100 56252
rect 28252 55412 28532 55468
rect 27356 55346 27412 55356
rect 27804 55188 27860 55198
rect 27804 54738 27860 55132
rect 27804 54686 27806 54738
rect 27858 54686 27860 54738
rect 27804 54674 27860 54686
rect 27132 53566 27134 53618
rect 27186 53566 27188 53618
rect 27132 53554 27188 53566
rect 28140 54514 28196 54526
rect 28140 54462 28142 54514
rect 28194 54462 28196 54514
rect 28028 52948 28084 52958
rect 28028 52854 28084 52892
rect 27804 52834 27860 52846
rect 27804 52782 27806 52834
rect 27858 52782 27860 52834
rect 26908 52724 26964 52734
rect 26908 52276 26964 52668
rect 27468 52500 27524 52510
rect 27356 52444 27468 52500
rect 27524 52444 27636 52500
rect 26908 52274 27076 52276
rect 26908 52222 26910 52274
rect 26962 52222 27076 52274
rect 26908 52220 27076 52222
rect 26908 52210 26964 52220
rect 26460 52162 26516 52174
rect 26460 52110 26462 52162
rect 26514 52110 26516 52162
rect 26348 51828 26404 51838
rect 26348 51266 26404 51772
rect 26460 51716 26516 52110
rect 26460 51650 26516 51660
rect 26460 51492 26516 51502
rect 26460 51490 26628 51492
rect 26460 51438 26462 51490
rect 26514 51438 26628 51490
rect 26460 51436 26628 51438
rect 26460 51426 26516 51436
rect 26348 51214 26350 51266
rect 26402 51214 26404 51266
rect 26348 51202 26404 51214
rect 26236 50876 26516 50932
rect 25900 50818 26180 50820
rect 25900 50766 25902 50818
rect 25954 50766 26180 50818
rect 25900 50764 26180 50766
rect 25900 50754 25956 50764
rect 26124 50148 26180 50764
rect 26236 50484 26292 50522
rect 26236 50418 26292 50428
rect 26124 50092 26292 50148
rect 25676 48974 25678 49026
rect 25730 48974 25732 49026
rect 25676 48962 25732 48974
rect 26124 49810 26180 49822
rect 26124 49758 26126 49810
rect 26178 49758 26180 49810
rect 26124 48916 26180 49758
rect 26236 49810 26292 50092
rect 26236 49758 26238 49810
rect 26290 49758 26292 49810
rect 26236 49746 26292 49758
rect 26236 49028 26292 49038
rect 26236 48934 26292 48972
rect 26124 48468 26180 48860
rect 26236 48468 26292 48478
rect 26124 48466 26292 48468
rect 26124 48414 26238 48466
rect 26290 48414 26292 48466
rect 26124 48412 26292 48414
rect 26236 48402 26292 48412
rect 24668 48078 24670 48130
rect 24722 48078 24724 48130
rect 24668 48066 24724 48078
rect 25228 47348 25284 47358
rect 25228 46562 25284 47292
rect 25228 46510 25230 46562
rect 25282 46510 25284 46562
rect 25228 46498 25284 46510
rect 25788 46564 25844 46574
rect 25788 46114 25844 46508
rect 25788 46062 25790 46114
rect 25842 46062 25844 46114
rect 25788 46050 25844 46062
rect 25788 45890 25844 45902
rect 25788 45838 25790 45890
rect 25842 45838 25844 45890
rect 25452 45778 25508 45790
rect 25452 45726 25454 45778
rect 25506 45726 25508 45778
rect 24444 44258 24500 44268
rect 25116 45668 25172 45678
rect 25452 45668 25508 45726
rect 25116 45666 25508 45668
rect 25116 45614 25118 45666
rect 25170 45614 25508 45666
rect 25116 45612 25508 45614
rect 25788 45668 25844 45838
rect 26236 45668 26292 45678
rect 25844 45612 25956 45668
rect 24108 43586 24164 43596
rect 24556 43538 24612 43550
rect 24556 43486 24558 43538
rect 24610 43486 24612 43538
rect 24332 42868 24388 42878
rect 24332 42774 24388 42812
rect 24556 42756 24612 43486
rect 24556 42690 24612 42700
rect 24780 43316 24836 43326
rect 24556 41076 24612 41086
rect 24444 41074 24612 41076
rect 24444 41022 24558 41074
rect 24610 41022 24612 41074
rect 24444 41020 24612 41022
rect 24220 40514 24276 40526
rect 24220 40462 24222 40514
rect 24274 40462 24276 40514
rect 24220 39508 24276 40462
rect 24220 39442 24276 39452
rect 24444 39058 24500 41020
rect 24556 41010 24612 41020
rect 24556 40628 24612 40638
rect 24556 40514 24612 40572
rect 24556 40462 24558 40514
rect 24610 40462 24612 40514
rect 24556 40450 24612 40462
rect 24444 39006 24446 39058
rect 24498 39006 24500 39058
rect 24444 38994 24500 39006
rect 24556 39060 24612 39070
rect 24556 38966 24612 39004
rect 24108 38948 24164 38958
rect 24108 38834 24164 38892
rect 24108 38782 24110 38834
rect 24162 38782 24164 38834
rect 24108 38770 24164 38782
rect 24332 38836 24388 38874
rect 24332 38770 24388 38780
rect 23772 37874 23828 37884
rect 23884 38610 23940 38622
rect 23996 38612 24164 38668
rect 23884 38558 23886 38610
rect 23938 38558 23940 38610
rect 23884 37826 23940 38558
rect 23884 37774 23886 37826
rect 23938 37774 23940 37826
rect 23884 37762 23940 37774
rect 23996 37938 24052 37950
rect 23996 37886 23998 37938
rect 24050 37886 24052 37938
rect 23996 37716 24052 37886
rect 23996 37650 24052 37660
rect 24108 36708 24164 38612
rect 24332 38612 24388 38622
rect 24388 38556 24612 38612
rect 24332 38546 24388 38556
rect 24220 38276 24276 38286
rect 24276 38220 24388 38276
rect 24220 38210 24276 38220
rect 24220 37938 24276 37950
rect 24220 37886 24222 37938
rect 24274 37886 24276 37938
rect 24220 37156 24276 37886
rect 24220 37090 24276 37100
rect 24108 36652 24276 36708
rect 24108 36484 24164 36494
rect 23660 36428 23828 36484
rect 23436 36390 23492 36428
rect 23548 36258 23604 36270
rect 23548 36206 23550 36258
rect 23602 36206 23604 36258
rect 23548 36036 23604 36206
rect 23324 35858 23380 35868
rect 23436 35980 23604 36036
rect 23660 36258 23716 36270
rect 23660 36206 23662 36258
rect 23714 36206 23716 36258
rect 23044 35196 23156 35252
rect 23436 35252 23492 35980
rect 23548 35700 23604 35710
rect 23660 35700 23716 36206
rect 23604 35644 23716 35700
rect 23772 35700 23828 36428
rect 23548 35606 23604 35644
rect 23772 35606 23828 35644
rect 23884 36428 24108 36484
rect 23884 35476 23940 36428
rect 24108 36390 24164 36428
rect 23996 35924 24052 35934
rect 23996 35830 24052 35868
rect 24220 35700 24276 36652
rect 24332 36482 24388 38220
rect 24556 38050 24612 38556
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24556 37986 24612 37998
rect 24332 36430 24334 36482
rect 24386 36430 24388 36482
rect 24332 36418 24388 36430
rect 24556 36372 24612 36382
rect 24556 36278 24612 36316
rect 24444 36260 24500 36270
rect 24444 36166 24500 36204
rect 22988 35186 23044 35196
rect 23436 35186 23492 35196
rect 23660 35420 23940 35476
rect 23996 35644 24276 35700
rect 23660 35138 23716 35420
rect 23996 35252 24052 35644
rect 23660 35086 23662 35138
rect 23714 35086 23716 35138
rect 23660 35074 23716 35086
rect 23772 35196 24052 35252
rect 24108 35474 24164 35486
rect 24108 35422 24110 35474
rect 24162 35422 24164 35474
rect 22988 34916 23044 34926
rect 23436 34916 23492 34926
rect 22988 34914 23492 34916
rect 22988 34862 22990 34914
rect 23042 34862 23438 34914
rect 23490 34862 23492 34914
rect 22988 34860 23492 34862
rect 22988 34850 23044 34860
rect 23436 34850 23492 34860
rect 23100 34130 23156 34142
rect 23100 34078 23102 34130
rect 23154 34078 23156 34130
rect 23100 33236 23156 34078
rect 23100 33170 23156 33180
rect 22876 31602 22932 31612
rect 22988 32562 23044 32574
rect 22988 32510 22990 32562
rect 23042 32510 23044 32562
rect 22764 31108 22820 31118
rect 22204 30830 22206 30882
rect 22258 30830 22260 30882
rect 22204 30818 22260 30830
rect 22316 30994 22372 31006
rect 22316 30942 22318 30994
rect 22370 30942 22372 30994
rect 22316 30210 22372 30942
rect 22764 30994 22820 31052
rect 22764 30942 22766 30994
rect 22818 30942 22820 30994
rect 22764 30930 22820 30942
rect 22988 30434 23044 32510
rect 23772 32116 23828 35196
rect 23884 34914 23940 34926
rect 24108 34916 24164 35422
rect 24332 35140 24388 35150
rect 24668 35140 24724 35150
rect 24388 35084 24612 35140
rect 24332 35074 24388 35084
rect 23884 34862 23886 34914
rect 23938 34862 23940 34914
rect 23884 34804 23940 34862
rect 23884 34244 23940 34748
rect 23884 34178 23940 34188
rect 23996 34860 24164 34916
rect 24332 34916 24388 34926
rect 23996 33684 24052 34860
rect 24332 34822 24388 34860
rect 24108 34692 24164 34702
rect 24108 34598 24164 34636
rect 24220 34690 24276 34702
rect 24220 34638 24222 34690
rect 24274 34638 24276 34690
rect 24220 34468 24276 34638
rect 24220 34402 24276 34412
rect 24556 34354 24612 35084
rect 24556 34302 24558 34354
rect 24610 34302 24612 34354
rect 24556 34290 24612 34302
rect 24668 34130 24724 35084
rect 24668 34078 24670 34130
rect 24722 34078 24724 34130
rect 24220 33908 24276 33918
rect 24220 33814 24276 33852
rect 24444 33906 24500 33918
rect 24444 33854 24446 33906
rect 24498 33854 24500 33906
rect 23996 33618 24052 33628
rect 23772 32050 23828 32060
rect 24220 32788 24276 32798
rect 23548 31892 23604 31902
rect 23212 31780 23268 31790
rect 23100 31724 23212 31780
rect 23100 30772 23156 31724
rect 23212 31686 23268 31724
rect 23548 31780 23604 31836
rect 23660 31780 23716 31790
rect 23548 31778 23716 31780
rect 23548 31726 23662 31778
rect 23714 31726 23716 31778
rect 23548 31724 23716 31726
rect 23324 31332 23380 31342
rect 23324 30994 23380 31276
rect 23324 30942 23326 30994
rect 23378 30942 23380 30994
rect 23324 30930 23380 30942
rect 23100 30706 23156 30716
rect 23324 30772 23380 30782
rect 22988 30382 22990 30434
rect 23042 30382 23044 30434
rect 22988 30370 23044 30382
rect 23324 30434 23380 30716
rect 23324 30382 23326 30434
rect 23378 30382 23380 30434
rect 23324 30370 23380 30382
rect 22988 30212 23044 30222
rect 22316 30158 22318 30210
rect 22370 30158 22372 30210
rect 22316 30146 22372 30158
rect 22876 30210 23044 30212
rect 22876 30158 22990 30210
rect 23042 30158 23044 30210
rect 22876 30156 23044 30158
rect 22428 30100 22484 30110
rect 22652 30100 22708 30110
rect 22484 30044 22596 30100
rect 22428 30034 22484 30044
rect 22540 29986 22596 30044
rect 22652 30006 22708 30044
rect 22540 29934 22542 29986
rect 22594 29934 22596 29986
rect 22540 29764 22596 29934
rect 22876 29764 22932 30156
rect 22988 30146 23044 30156
rect 23548 30212 23604 31724
rect 23660 31714 23716 31724
rect 24220 31778 24276 32732
rect 24332 32564 24388 32574
rect 24332 32470 24388 32508
rect 24220 31726 24222 31778
rect 24274 31726 24276 31778
rect 24220 31714 24276 31726
rect 24444 31668 24500 33854
rect 24556 33012 24612 33022
rect 24556 32674 24612 32956
rect 24668 32900 24724 34078
rect 24668 32834 24724 32844
rect 24780 32788 24836 43260
rect 25116 38668 25172 45612
rect 25788 45602 25844 45612
rect 25340 45444 25396 45454
rect 25340 44994 25396 45388
rect 25900 45330 25956 45612
rect 26236 45574 26292 45612
rect 25900 45278 25902 45330
rect 25954 45278 25956 45330
rect 25900 45266 25956 45278
rect 26348 45444 26404 45454
rect 26348 45106 26404 45388
rect 26348 45054 26350 45106
rect 26402 45054 26404 45106
rect 26348 45042 26404 45054
rect 25340 44942 25342 44994
rect 25394 44942 25396 44994
rect 25340 42756 25396 44942
rect 25676 44884 25732 44894
rect 25676 44790 25732 44828
rect 26012 44884 26068 44894
rect 26012 44790 26068 44828
rect 25452 44434 25508 44446
rect 25452 44382 25454 44434
rect 25506 44382 25508 44434
rect 25452 44324 25508 44382
rect 25452 44258 25508 44268
rect 25340 41972 25396 42700
rect 26460 42866 26516 50876
rect 26572 50034 26628 51436
rect 26684 51156 26740 51166
rect 26684 51154 26964 51156
rect 26684 51102 26686 51154
rect 26738 51102 26964 51154
rect 26684 51100 26964 51102
rect 26684 51090 26740 51100
rect 26908 50820 26964 51100
rect 27020 51044 27076 52220
rect 27132 52164 27188 52174
rect 27132 52070 27188 52108
rect 27356 52162 27412 52444
rect 27468 52434 27524 52444
rect 27356 52110 27358 52162
rect 27410 52110 27412 52162
rect 27356 52098 27412 52110
rect 27468 52276 27524 52286
rect 27244 51604 27300 51614
rect 27468 51604 27524 52220
rect 27244 51602 27524 51604
rect 27244 51550 27246 51602
rect 27298 51550 27524 51602
rect 27244 51548 27524 51550
rect 27244 51538 27300 51548
rect 27132 51490 27188 51502
rect 27132 51438 27134 51490
rect 27186 51438 27188 51490
rect 27132 51380 27188 51438
rect 27132 51314 27188 51324
rect 27580 51268 27636 52444
rect 27804 52164 27860 52782
rect 27916 52724 27972 52734
rect 27916 52386 27972 52668
rect 27916 52334 27918 52386
rect 27970 52334 27972 52386
rect 27916 52322 27972 52334
rect 28140 52388 28196 54462
rect 28476 53618 28532 55412
rect 28588 55410 28644 55692
rect 28588 55358 28590 55410
rect 28642 55358 28644 55410
rect 28588 55346 28644 55358
rect 28700 55692 29652 55748
rect 30268 56082 30324 56094
rect 30268 56030 30270 56082
rect 30322 56030 30324 56082
rect 30268 55748 30324 56030
rect 28588 54740 28644 54750
rect 28700 54740 28756 55692
rect 30268 55682 30324 55692
rect 29596 55412 29652 55422
rect 29596 55318 29652 55356
rect 30940 55186 30996 59200
rect 31052 56308 31108 56318
rect 31052 56214 31108 56252
rect 31388 56308 31444 59200
rect 32284 57428 32340 59200
rect 32732 57652 32788 59200
rect 32732 57596 33236 57652
rect 32284 57372 33124 57428
rect 31388 56242 31444 56252
rect 32620 56308 32676 56318
rect 32284 56082 32340 56094
rect 32284 56030 32286 56082
rect 32338 56030 32340 56082
rect 30940 55134 30942 55186
rect 30994 55134 30996 55186
rect 30940 55122 30996 55134
rect 31500 55298 31556 55310
rect 31500 55246 31502 55298
rect 31554 55246 31556 55298
rect 30380 55076 30436 55086
rect 30380 54982 30436 55020
rect 28588 54738 28756 54740
rect 28588 54686 28590 54738
rect 28642 54686 28756 54738
rect 28588 54684 28756 54686
rect 28588 54674 28644 54684
rect 31276 54516 31332 54526
rect 31500 54516 31556 55246
rect 32172 55186 32228 55198
rect 32172 55134 32174 55186
rect 32226 55134 32228 55186
rect 32172 54738 32228 55134
rect 32172 54686 32174 54738
rect 32226 54686 32228 54738
rect 32172 54674 32228 54686
rect 31836 54516 31892 54526
rect 31500 54514 31892 54516
rect 31500 54462 31838 54514
rect 31890 54462 31892 54514
rect 31500 54460 31892 54462
rect 28924 54404 28980 54414
rect 31052 54404 31108 54414
rect 28924 54310 28980 54348
rect 30604 54402 31108 54404
rect 30604 54350 31054 54402
rect 31106 54350 31108 54402
rect 30604 54348 31108 54350
rect 28476 53566 28478 53618
rect 28530 53566 28532 53618
rect 28476 53554 28532 53566
rect 29372 53732 29428 53742
rect 29708 53732 29764 53742
rect 29372 53506 29428 53676
rect 29372 53454 29374 53506
rect 29426 53454 29428 53506
rect 29372 53442 29428 53454
rect 29596 53730 29764 53732
rect 29596 53678 29710 53730
rect 29762 53678 29764 53730
rect 29596 53676 29764 53678
rect 28364 53170 28420 53182
rect 28364 53118 28366 53170
rect 28418 53118 28420 53170
rect 28364 53060 28420 53118
rect 28364 52994 28420 53004
rect 29596 53060 29652 53676
rect 29708 53666 29764 53676
rect 30380 53732 30436 53742
rect 30380 53730 30548 53732
rect 30380 53678 30382 53730
rect 30434 53678 30548 53730
rect 30380 53676 30548 53678
rect 30380 53666 30436 53676
rect 28140 52322 28196 52332
rect 28588 52946 28644 52958
rect 28588 52894 28590 52946
rect 28642 52894 28644 52946
rect 28588 52276 28644 52894
rect 28924 52946 28980 52958
rect 28924 52894 28926 52946
rect 28978 52894 28980 52946
rect 28812 52836 28868 52846
rect 28812 52742 28868 52780
rect 28588 52210 28644 52220
rect 28924 52500 28980 52894
rect 28924 52276 28980 52444
rect 29148 52948 29204 52958
rect 29148 52388 29204 52892
rect 29596 52946 29652 53004
rect 29932 53618 29988 53630
rect 29932 53566 29934 53618
rect 29986 53566 29988 53618
rect 29932 53060 29988 53566
rect 30492 53170 30548 53676
rect 30604 53618 30660 54348
rect 31052 54338 31108 54348
rect 30604 53566 30606 53618
rect 30658 53566 30660 53618
rect 30604 53554 30660 53566
rect 30492 53118 30494 53170
rect 30546 53118 30548 53170
rect 30492 53106 30548 53118
rect 31276 53170 31332 54460
rect 31836 53732 31892 54460
rect 32284 54404 32340 56030
rect 32620 55970 32676 56252
rect 32620 55918 32622 55970
rect 32674 55918 32676 55970
rect 32620 55906 32676 55918
rect 33068 54738 33124 57372
rect 33180 57092 33236 57596
rect 33180 57026 33236 57036
rect 33628 56308 33684 59200
rect 33628 56242 33684 56252
rect 34076 55636 34132 59200
rect 34636 57092 34692 57102
rect 34076 55570 34132 55580
rect 34300 56082 34356 56094
rect 34300 56030 34302 56082
rect 34354 56030 34356 56082
rect 34300 55410 34356 56030
rect 34636 55970 34692 57036
rect 34972 56084 35028 59200
rect 35420 56642 35476 59200
rect 35420 56590 35422 56642
rect 35474 56590 35476 56642
rect 35420 56578 35476 56590
rect 35308 56308 35364 56318
rect 35308 56214 35364 56252
rect 36316 56308 36372 59200
rect 36764 57092 36820 59200
rect 36764 57026 36820 57036
rect 36316 56242 36372 56252
rect 36764 56642 36820 56654
rect 36764 56590 36766 56642
rect 36818 56590 36820 56642
rect 36764 56306 36820 56590
rect 36764 56254 36766 56306
rect 36818 56254 36820 56306
rect 36764 56242 36820 56254
rect 37436 56196 37492 56206
rect 34636 55918 34638 55970
rect 34690 55918 34692 55970
rect 34636 55906 34692 55918
rect 34860 56028 35028 56084
rect 36092 56082 36148 56094
rect 36092 56030 36094 56082
rect 36146 56030 36148 56082
rect 34300 55358 34302 55410
rect 34354 55358 34356 55410
rect 34300 55346 34356 55358
rect 33068 54686 33070 54738
rect 33122 54686 33124 54738
rect 33068 54674 33124 54686
rect 34748 55298 34804 55310
rect 34748 55246 34750 55298
rect 34802 55246 34804 55298
rect 32396 54516 32452 54526
rect 32396 54422 32452 54460
rect 32284 54338 32340 54348
rect 34188 53956 34244 53966
rect 31948 53732 32004 53742
rect 31836 53676 31948 53732
rect 31948 53638 32004 53676
rect 33180 53732 33236 53742
rect 32620 53620 32676 53630
rect 31276 53118 31278 53170
rect 31330 53118 31332 53170
rect 31276 53106 31332 53118
rect 32172 53618 32676 53620
rect 32172 53566 32622 53618
rect 32674 53566 32676 53618
rect 32172 53564 32676 53566
rect 29932 52994 29988 53004
rect 30716 53060 30772 53070
rect 30716 52966 30772 53004
rect 29596 52894 29598 52946
rect 29650 52894 29652 52946
rect 29596 52882 29652 52894
rect 30268 52836 30324 52846
rect 29820 52724 29876 52734
rect 30044 52724 30100 52734
rect 29820 52630 29876 52668
rect 29932 52722 30100 52724
rect 29932 52670 30046 52722
rect 30098 52670 30100 52722
rect 29932 52668 30100 52670
rect 29932 52388 29988 52668
rect 30044 52658 30100 52668
rect 28924 52210 28980 52220
rect 29036 52332 29204 52388
rect 29484 52332 29988 52388
rect 30044 52388 30100 52398
rect 27692 51492 27748 51502
rect 27804 51492 27860 52108
rect 28924 51604 28980 51614
rect 28924 51510 28980 51548
rect 27692 51490 27860 51492
rect 27692 51438 27694 51490
rect 27746 51438 27860 51490
rect 27692 51436 27860 51438
rect 28700 51492 28756 51502
rect 27692 51426 27748 51436
rect 28700 51398 28756 51436
rect 27916 51380 27972 51390
rect 27804 51268 27860 51278
rect 27580 51266 27860 51268
rect 27580 51214 27806 51266
rect 27858 51214 27860 51266
rect 27580 51212 27860 51214
rect 27804 51202 27860 51212
rect 27356 51154 27412 51166
rect 27356 51102 27358 51154
rect 27410 51102 27412 51154
rect 27020 50988 27300 51044
rect 27132 50820 27188 50830
rect 26908 50818 27188 50820
rect 26908 50766 27134 50818
rect 27186 50766 27188 50818
rect 26908 50764 27188 50766
rect 27132 50754 27188 50764
rect 26796 50596 26852 50606
rect 26796 50502 26852 50540
rect 27132 50594 27188 50606
rect 27132 50542 27134 50594
rect 27186 50542 27188 50594
rect 27132 50484 27188 50542
rect 27132 50418 27188 50428
rect 26572 49982 26574 50034
rect 26626 49982 26628 50034
rect 26572 49476 26628 49982
rect 26684 49924 26740 49934
rect 26684 49698 26740 49868
rect 26684 49646 26686 49698
rect 26738 49646 26740 49698
rect 26684 49634 26740 49646
rect 26796 49812 26852 49822
rect 26572 49410 26628 49420
rect 26572 49252 26628 49262
rect 26572 49158 26628 49196
rect 26796 49138 26852 49756
rect 26796 49086 26798 49138
rect 26850 49086 26852 49138
rect 26796 49074 26852 49086
rect 27132 49252 27188 49262
rect 27244 49252 27300 50988
rect 27356 50372 27412 51102
rect 27468 51156 27524 51166
rect 27468 50820 27524 51100
rect 27468 50726 27524 50764
rect 27916 51156 27972 51324
rect 28252 51380 28308 51390
rect 28252 51378 28420 51380
rect 28252 51326 28254 51378
rect 28306 51326 28420 51378
rect 28252 51324 28420 51326
rect 28252 51314 28308 51324
rect 28028 51156 28084 51166
rect 27916 51154 28084 51156
rect 27916 51102 28030 51154
rect 28082 51102 28084 51154
rect 27916 51100 28084 51102
rect 27356 50306 27412 50316
rect 27692 50596 27748 50606
rect 27692 50148 27748 50540
rect 27356 50092 27748 50148
rect 27356 49922 27412 50092
rect 27356 49870 27358 49922
rect 27410 49870 27412 49922
rect 27356 49858 27412 49870
rect 27580 49924 27636 49934
rect 27580 49830 27636 49868
rect 27468 49810 27524 49822
rect 27468 49758 27470 49810
rect 27522 49758 27524 49810
rect 27188 49196 27300 49252
rect 27356 49588 27412 49598
rect 27356 49364 27412 49532
rect 26908 49026 26964 49038
rect 26908 48974 26910 49026
rect 26962 48974 26964 49026
rect 26908 48916 26964 48974
rect 27132 49026 27188 49196
rect 27132 48974 27134 49026
rect 27186 48974 27188 49026
rect 27132 48962 27188 48974
rect 26908 48692 26964 48860
rect 26796 48636 26964 48692
rect 27244 48804 27300 48814
rect 26572 48468 26628 48478
rect 26796 48468 26852 48636
rect 26572 48466 26852 48468
rect 26572 48414 26574 48466
rect 26626 48414 26852 48466
rect 26572 48412 26852 48414
rect 26572 48402 26628 48412
rect 27020 48356 27076 48366
rect 27020 48262 27076 48300
rect 27244 48130 27300 48748
rect 27356 48242 27412 49308
rect 27468 49028 27524 49758
rect 27468 48802 27524 48972
rect 27468 48750 27470 48802
rect 27522 48750 27524 48802
rect 27468 48356 27524 48750
rect 27692 48802 27748 50092
rect 27804 49588 27860 49598
rect 27804 49250 27860 49532
rect 27804 49198 27806 49250
rect 27858 49198 27860 49250
rect 27804 49186 27860 49198
rect 27916 48916 27972 51100
rect 28028 51090 28084 51100
rect 28140 50820 28196 50830
rect 28140 50428 28196 50764
rect 28252 50596 28308 50606
rect 28252 50502 28308 50540
rect 28140 50372 28308 50428
rect 28028 49924 28084 49934
rect 28028 49830 28084 49868
rect 28140 49812 28196 49822
rect 28028 48916 28084 48926
rect 27916 48914 28084 48916
rect 27916 48862 28030 48914
rect 28082 48862 28084 48914
rect 27916 48860 28084 48862
rect 27692 48750 27694 48802
rect 27746 48750 27748 48802
rect 27692 48468 27748 48750
rect 27692 48402 27748 48412
rect 27468 48290 27524 48300
rect 27356 48190 27358 48242
rect 27410 48190 27412 48242
rect 27356 48178 27412 48190
rect 28028 48244 28084 48860
rect 28140 48804 28196 49756
rect 28252 49810 28308 50372
rect 28252 49758 28254 49810
rect 28306 49758 28308 49810
rect 28252 49746 28308 49758
rect 28364 50372 28420 51324
rect 29036 51266 29092 52332
rect 29148 52164 29204 52174
rect 29372 52164 29428 52174
rect 29148 52070 29204 52108
rect 29260 52162 29428 52164
rect 29260 52110 29374 52162
rect 29426 52110 29428 52162
rect 29260 52108 29428 52110
rect 29036 51214 29038 51266
rect 29090 51214 29092 51266
rect 29036 51202 29092 51214
rect 29260 51044 29316 52108
rect 29372 52098 29428 52108
rect 28588 50988 29316 51044
rect 28588 50818 28644 50988
rect 28588 50766 28590 50818
rect 28642 50766 28644 50818
rect 28588 50754 28644 50766
rect 28476 50708 28532 50718
rect 28476 50614 28532 50652
rect 28364 49252 28420 50316
rect 28812 50596 28868 50606
rect 28812 50034 28868 50540
rect 28812 49982 28814 50034
rect 28866 49982 28868 50034
rect 28812 49970 28868 49982
rect 29148 50482 29204 50494
rect 29148 50430 29150 50482
rect 29202 50430 29204 50482
rect 28700 49810 28756 49822
rect 28700 49758 28702 49810
rect 28754 49758 28756 49810
rect 28700 49364 28756 49758
rect 28924 49812 28980 49822
rect 28924 49718 28980 49756
rect 28700 49298 28756 49308
rect 28812 49476 28868 49486
rect 28364 49186 28420 49196
rect 28588 49140 28644 49150
rect 28588 49046 28644 49084
rect 28252 49028 28308 49038
rect 28252 48934 28308 48972
rect 28812 48916 28868 49420
rect 28812 48850 28868 48860
rect 29036 49364 29092 49374
rect 28476 48804 28532 48814
rect 28140 48748 28308 48804
rect 28252 48580 28308 48748
rect 28252 48524 28420 48580
rect 28252 48356 28308 48366
rect 28252 48262 28308 48300
rect 28140 48244 28196 48254
rect 28028 48242 28196 48244
rect 28028 48190 28142 48242
rect 28194 48190 28196 48242
rect 28028 48188 28196 48190
rect 28140 48178 28196 48188
rect 27244 48078 27246 48130
rect 27298 48078 27300 48130
rect 27244 48066 27300 48078
rect 28252 47684 28308 47694
rect 28364 47684 28420 48524
rect 28252 47682 28420 47684
rect 28252 47630 28254 47682
rect 28306 47630 28420 47682
rect 28252 47628 28420 47630
rect 28252 47618 28308 47628
rect 28028 47460 28084 47470
rect 28476 47460 28532 48748
rect 28588 48356 28644 48366
rect 28588 47682 28644 48300
rect 29036 48130 29092 49308
rect 29148 49140 29204 50430
rect 29260 50372 29316 50382
rect 29260 50370 29428 50372
rect 29260 50318 29262 50370
rect 29314 50318 29428 50370
rect 29260 50316 29428 50318
rect 29260 50306 29316 50316
rect 29372 50036 29428 50316
rect 29372 49970 29428 49980
rect 29484 50034 29540 52332
rect 30044 52294 30100 52332
rect 30268 52274 30324 52780
rect 30940 52724 30996 52734
rect 31276 52724 31332 52734
rect 30380 52722 31108 52724
rect 30380 52670 30942 52722
rect 30994 52670 31108 52722
rect 30380 52668 31108 52670
rect 30380 52386 30436 52668
rect 30940 52658 30996 52668
rect 30380 52334 30382 52386
rect 30434 52334 30436 52386
rect 30380 52322 30436 52334
rect 30268 52222 30270 52274
rect 30322 52222 30324 52274
rect 30268 52210 30324 52222
rect 31052 52274 31108 52668
rect 31052 52222 31054 52274
rect 31106 52222 31108 52274
rect 31052 52210 31108 52222
rect 29596 52162 29652 52174
rect 29596 52110 29598 52162
rect 29650 52110 29652 52162
rect 29596 51268 29652 52110
rect 31276 52162 31332 52668
rect 31500 52164 31556 52174
rect 31276 52110 31278 52162
rect 31330 52110 31332 52162
rect 31276 52098 31332 52110
rect 31388 52162 31556 52164
rect 31388 52110 31502 52162
rect 31554 52110 31556 52162
rect 31388 52108 31556 52110
rect 29596 51202 29652 51212
rect 29708 51604 29764 51614
rect 29708 50594 29764 51548
rect 30604 51604 30660 51614
rect 30268 51268 30324 51278
rect 30324 51212 30436 51268
rect 30268 51202 30324 51212
rect 30268 50820 30324 50830
rect 29708 50542 29710 50594
rect 29762 50542 29764 50594
rect 29708 50530 29764 50542
rect 29932 50708 29988 50718
rect 29484 49982 29486 50034
rect 29538 49982 29540 50034
rect 29484 49970 29540 49982
rect 29820 50484 29876 50494
rect 29372 49812 29428 49822
rect 29372 49718 29428 49756
rect 29596 49810 29652 49822
rect 29596 49758 29598 49810
rect 29650 49758 29652 49810
rect 29596 49476 29652 49758
rect 29596 49410 29652 49420
rect 29260 49252 29316 49262
rect 29260 49158 29316 49196
rect 29148 49074 29204 49084
rect 29820 49138 29876 50428
rect 29932 50484 29988 50652
rect 30268 50594 30324 50764
rect 30380 50818 30436 51212
rect 30380 50766 30382 50818
rect 30434 50766 30436 50818
rect 30380 50754 30436 50766
rect 30268 50542 30270 50594
rect 30322 50542 30324 50594
rect 29932 50482 30212 50484
rect 29932 50430 29934 50482
rect 29986 50430 30212 50482
rect 29932 50428 30212 50430
rect 29932 50418 29988 50428
rect 29820 49086 29822 49138
rect 29874 49086 29876 49138
rect 29820 49074 29876 49086
rect 29932 50036 29988 50046
rect 29372 49028 29428 49038
rect 29372 48914 29428 48972
rect 29932 49026 29988 49980
rect 30044 49810 30100 49822
rect 30044 49758 30046 49810
rect 30098 49758 30100 49810
rect 30044 49700 30100 49758
rect 30044 49634 30100 49644
rect 29932 48974 29934 49026
rect 29986 48974 29988 49026
rect 29932 48962 29988 48974
rect 29372 48862 29374 48914
rect 29426 48862 29428 48914
rect 29260 48804 29316 48814
rect 29260 48710 29316 48748
rect 29036 48078 29038 48130
rect 29090 48078 29092 48130
rect 29036 48066 29092 48078
rect 28588 47630 28590 47682
rect 28642 47630 28644 47682
rect 28588 47618 28644 47630
rect 28028 47458 28532 47460
rect 28028 47406 28030 47458
rect 28082 47406 28532 47458
rect 28028 47404 28532 47406
rect 29260 47460 29316 47470
rect 29372 47460 29428 48862
rect 30156 48914 30212 50428
rect 30268 49252 30324 50542
rect 30492 50484 30548 50494
rect 30492 50390 30548 50428
rect 30380 49922 30436 49934
rect 30380 49870 30382 49922
rect 30434 49870 30436 49922
rect 30380 49812 30436 49870
rect 30380 49746 30436 49756
rect 30604 49810 30660 51548
rect 31276 50708 31332 50718
rect 31276 50594 31332 50652
rect 31276 50542 31278 50594
rect 31330 50542 31332 50594
rect 31276 50530 31332 50542
rect 30940 50482 30996 50494
rect 30940 50430 30942 50482
rect 30994 50430 30996 50482
rect 30604 49758 30606 49810
rect 30658 49758 30660 49810
rect 30604 49746 30660 49758
rect 30716 50370 30772 50382
rect 30716 50318 30718 50370
rect 30770 50318 30772 50370
rect 30716 49812 30772 50318
rect 30716 49746 30772 49756
rect 30940 49700 30996 50430
rect 31388 50428 31444 52108
rect 31500 52098 31556 52108
rect 32172 51602 32228 53564
rect 32620 53554 32676 53564
rect 33180 52948 33236 53676
rect 33180 52946 33572 52948
rect 33180 52894 33182 52946
rect 33234 52894 33572 52946
rect 33180 52892 33572 52894
rect 33180 52882 33236 52892
rect 33292 52276 33348 52286
rect 33292 52050 33348 52220
rect 33292 51998 33294 52050
rect 33346 51998 33348 52050
rect 33292 51986 33348 51998
rect 33404 52164 33460 52174
rect 32284 51940 32340 51950
rect 32284 51846 32340 51884
rect 33180 51940 33236 51950
rect 32172 51550 32174 51602
rect 32226 51550 32228 51602
rect 32172 51538 32228 51550
rect 33180 51604 33236 51884
rect 33180 51602 33348 51604
rect 33180 51550 33182 51602
rect 33234 51550 33348 51602
rect 33180 51548 33348 51550
rect 33180 51538 33236 51548
rect 31836 51492 31892 51502
rect 31836 51490 32116 51492
rect 31836 51438 31838 51490
rect 31890 51438 32116 51490
rect 31836 51436 32116 51438
rect 31836 51426 31892 51436
rect 31724 51380 31780 51390
rect 31612 51378 31780 51380
rect 31612 51326 31726 51378
rect 31778 51326 31780 51378
rect 31612 51324 31780 51326
rect 31276 50372 31444 50428
rect 31500 50484 31556 50494
rect 31612 50484 31668 51324
rect 31724 51314 31780 51324
rect 31836 51156 31892 51166
rect 31836 51154 32004 51156
rect 31836 51102 31838 51154
rect 31890 51102 32004 51154
rect 31836 51100 32004 51102
rect 31836 51090 31892 51100
rect 31948 50820 32004 51100
rect 31948 50754 32004 50764
rect 31836 50708 31892 50718
rect 31836 50614 31892 50652
rect 31500 50482 31668 50484
rect 31500 50430 31502 50482
rect 31554 50430 31668 50482
rect 31500 50428 31668 50430
rect 32060 50428 32116 51436
rect 32396 51490 32452 51502
rect 32396 51438 32398 51490
rect 32450 51438 32452 51490
rect 32172 50596 32228 50606
rect 32172 50502 32228 50540
rect 31164 49924 31220 49934
rect 31164 49810 31220 49868
rect 31164 49758 31166 49810
rect 31218 49758 31220 49810
rect 31164 49746 31220 49758
rect 31276 49922 31332 50372
rect 31276 49870 31278 49922
rect 31330 49870 31332 49922
rect 31052 49700 31108 49710
rect 30940 49644 31052 49700
rect 31052 49634 31108 49644
rect 31164 49588 31220 49598
rect 31052 49476 31108 49486
rect 30268 49186 30324 49196
rect 30940 49252 30996 49262
rect 30828 49140 30884 49150
rect 30828 49046 30884 49084
rect 30156 48862 30158 48914
rect 30210 48862 30212 48914
rect 29708 48804 29764 48814
rect 29708 48710 29764 48748
rect 30156 48692 30212 48862
rect 30940 48914 30996 49196
rect 30940 48862 30942 48914
rect 30994 48862 30996 48914
rect 30940 48850 30996 48862
rect 30604 48804 30660 48814
rect 30604 48710 30660 48748
rect 30828 48802 30884 48814
rect 30828 48750 30830 48802
rect 30882 48750 30884 48802
rect 30156 48626 30212 48636
rect 30828 48692 30884 48750
rect 31052 48692 31108 49420
rect 30828 48626 30884 48636
rect 30940 48636 31108 48692
rect 29260 47458 29428 47460
rect 29260 47406 29262 47458
rect 29314 47406 29428 47458
rect 29260 47404 29428 47406
rect 29820 48244 29876 48254
rect 29820 47458 29876 48188
rect 30828 47572 30884 47582
rect 30940 47572 30996 48636
rect 31052 48468 31108 48478
rect 31052 48242 31108 48412
rect 31052 48190 31054 48242
rect 31106 48190 31108 48242
rect 31052 48178 31108 48190
rect 30828 47570 30996 47572
rect 30828 47518 30830 47570
rect 30882 47518 30996 47570
rect 30828 47516 30996 47518
rect 31164 47570 31220 49532
rect 31276 49364 31332 49870
rect 31276 49298 31332 49308
rect 31388 50148 31444 50158
rect 31388 49026 31444 50092
rect 31388 48974 31390 49026
rect 31442 48974 31444 49026
rect 31388 48962 31444 48974
rect 31276 47684 31332 47694
rect 31500 47684 31556 50428
rect 31724 50372 31780 50382
rect 31612 50370 31780 50372
rect 31612 50318 31726 50370
rect 31778 50318 31780 50370
rect 31612 50316 31780 50318
rect 31612 49924 31668 50316
rect 31724 50306 31780 50316
rect 31836 50372 31892 50382
rect 31836 50036 31892 50316
rect 31612 49858 31668 49868
rect 31724 49980 31892 50036
rect 31948 50372 32116 50428
rect 31724 49476 31780 49980
rect 31724 49410 31780 49420
rect 31836 49812 31892 49822
rect 31612 49364 31668 49374
rect 31612 49252 31668 49308
rect 31612 49196 31780 49252
rect 31612 49028 31668 49038
rect 31612 48244 31668 48972
rect 31724 49026 31780 49196
rect 31724 48974 31726 49026
rect 31778 48974 31780 49026
rect 31724 48962 31780 48974
rect 31612 48150 31668 48188
rect 31836 48020 31892 49756
rect 31948 49028 32004 50372
rect 32284 50260 32340 50270
rect 32284 49924 32340 50204
rect 32396 50148 32452 51438
rect 32508 51378 32564 51390
rect 32508 51326 32510 51378
rect 32562 51326 32564 51378
rect 32508 50706 32564 51326
rect 32508 50654 32510 50706
rect 32562 50654 32564 50706
rect 32508 50642 32564 50654
rect 33068 51378 33124 51390
rect 33068 51326 33070 51378
rect 33122 51326 33124 51378
rect 33068 50708 33124 51326
rect 33292 51044 33348 51548
rect 33404 51602 33460 52108
rect 33516 51716 33572 52892
rect 33852 52834 33908 52846
rect 33852 52782 33854 52834
rect 33906 52782 33908 52834
rect 33852 52164 33908 52782
rect 34076 52276 34132 52286
rect 34076 52182 34132 52220
rect 33852 52098 33908 52108
rect 33628 51940 33684 51950
rect 33628 51938 33796 51940
rect 33628 51886 33630 51938
rect 33682 51886 33796 51938
rect 33628 51884 33796 51886
rect 33628 51874 33684 51884
rect 33516 51660 33684 51716
rect 33404 51550 33406 51602
rect 33458 51550 33460 51602
rect 33404 51538 33460 51550
rect 33292 50988 33572 51044
rect 33068 50642 33124 50652
rect 33404 50820 33460 50830
rect 33180 50482 33236 50494
rect 33180 50430 33182 50482
rect 33234 50430 33236 50482
rect 32508 50372 32564 50382
rect 32508 50278 32564 50316
rect 32732 50372 32788 50382
rect 33068 50372 33124 50382
rect 32732 50370 33124 50372
rect 32732 50318 32734 50370
rect 32786 50318 33070 50370
rect 33122 50318 33124 50370
rect 32732 50316 33124 50318
rect 32732 50306 32788 50316
rect 32452 50092 32676 50148
rect 32396 50054 32452 50092
rect 32620 50034 32676 50092
rect 32620 49982 32622 50034
rect 32674 49982 32676 50034
rect 32620 49970 32676 49982
rect 33068 50034 33124 50316
rect 33180 50372 33236 50430
rect 33180 50306 33236 50316
rect 33292 50484 33348 50494
rect 33292 50148 33348 50428
rect 33068 49982 33070 50034
rect 33122 49982 33124 50034
rect 33068 49970 33124 49982
rect 33180 50092 33348 50148
rect 33180 50034 33236 50092
rect 33180 49982 33182 50034
rect 33234 49982 33236 50034
rect 33180 49970 33236 49982
rect 32060 49810 32116 49822
rect 32060 49758 32062 49810
rect 32114 49758 32116 49810
rect 32060 49476 32116 49758
rect 32060 49410 32116 49420
rect 32172 49700 32228 49710
rect 32172 49138 32228 49644
rect 32172 49086 32174 49138
rect 32226 49086 32228 49138
rect 32172 49074 32228 49086
rect 31948 49026 32116 49028
rect 31948 48974 31950 49026
rect 32002 48974 32116 49026
rect 31948 48972 32116 48974
rect 31948 48962 32004 48972
rect 32060 48580 32116 48972
rect 32284 49026 32340 49868
rect 33292 49922 33348 49934
rect 33292 49870 33294 49922
rect 33346 49870 33348 49922
rect 32284 48974 32286 49026
rect 32338 48974 32340 49026
rect 32284 48962 32340 48974
rect 32732 49700 32788 49710
rect 32732 49028 32788 49644
rect 32732 48934 32788 48972
rect 32956 48804 33012 48814
rect 33292 48804 33348 49870
rect 33404 49922 33460 50764
rect 33516 50428 33572 50988
rect 33628 50594 33684 51660
rect 33740 51604 33796 51884
rect 33852 51604 33908 51614
rect 33740 51548 33852 51604
rect 33852 51510 33908 51548
rect 34188 51604 34244 53900
rect 34748 53842 34804 55246
rect 34860 55188 34916 56028
rect 35196 55692 35460 55702
rect 34972 55636 35028 55646
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 34972 55468 35028 55580
rect 34972 55412 35140 55468
rect 35084 55410 35140 55412
rect 35084 55358 35086 55410
rect 35138 55358 35140 55410
rect 35084 55346 35140 55358
rect 34860 55122 34916 55132
rect 35756 54516 35812 54526
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 34748 53790 34750 53842
rect 34802 53790 34804 53842
rect 34748 53778 34804 53790
rect 35756 53844 35812 54460
rect 35756 53778 35812 53788
rect 35980 53844 36036 53854
rect 35644 53618 35700 53630
rect 35644 53566 35646 53618
rect 35698 53566 35700 53618
rect 34300 52612 34356 52622
rect 34300 52162 34356 52556
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 34972 52276 35028 52286
rect 34972 52182 35028 52220
rect 35644 52276 35700 53566
rect 35980 53618 36036 53788
rect 35980 53566 35982 53618
rect 36034 53566 36036 53618
rect 35980 53554 36036 53566
rect 35980 52836 36036 52846
rect 36092 52836 36148 56030
rect 37100 55298 37156 55310
rect 37100 55246 37102 55298
rect 37154 55246 37156 55298
rect 36204 55188 36260 55198
rect 36204 55094 36260 55132
rect 37100 54516 37156 55246
rect 37156 54460 37268 54516
rect 37100 54450 37156 54460
rect 36428 54404 36484 54414
rect 36428 54402 36932 54404
rect 36428 54350 36430 54402
rect 36482 54350 36932 54402
rect 36428 54348 36932 54350
rect 36428 54338 36484 54348
rect 36876 53732 36932 54348
rect 37100 53844 37156 53854
rect 37100 53750 37156 53788
rect 36988 53732 37044 53742
rect 36876 53730 37044 53732
rect 36876 53678 36990 53730
rect 37042 53678 37044 53730
rect 36876 53676 37044 53678
rect 36988 53666 37044 53676
rect 35980 52834 36148 52836
rect 35980 52782 35982 52834
rect 36034 52782 36148 52834
rect 35980 52780 36148 52782
rect 36428 53060 36484 53070
rect 35980 52770 36036 52780
rect 35644 52210 35700 52220
rect 34300 52110 34302 52162
rect 34354 52110 34356 52162
rect 34300 52098 34356 52110
rect 34188 51602 34468 51604
rect 34188 51550 34190 51602
rect 34242 51550 34468 51602
rect 34188 51548 34468 51550
rect 34188 51538 34244 51548
rect 33628 50542 33630 50594
rect 33682 50542 33684 50594
rect 33628 50530 33684 50542
rect 34300 50484 34356 50494
rect 33516 50372 33684 50428
rect 34300 50390 34356 50428
rect 33404 49870 33406 49922
rect 33458 49870 33460 49922
rect 33404 49858 33460 49870
rect 33628 49922 33684 50372
rect 33628 49870 33630 49922
rect 33682 49870 33684 49922
rect 33628 49858 33684 49870
rect 34412 49810 34468 51548
rect 36204 51492 36260 51502
rect 36204 51490 36372 51492
rect 36204 51438 36206 51490
rect 36258 51438 36372 51490
rect 36204 51436 36372 51438
rect 36204 51426 36260 51436
rect 34412 49758 34414 49810
rect 34466 49758 34468 49810
rect 34412 49746 34468 49758
rect 35084 51380 35140 51390
rect 34188 49700 34244 49710
rect 34188 49606 34244 49644
rect 32956 48802 33348 48804
rect 32956 48750 32958 48802
rect 33010 48750 33348 48802
rect 32956 48748 33348 48750
rect 32956 48580 33012 48748
rect 32060 48524 33012 48580
rect 32060 48466 32116 48524
rect 32060 48414 32062 48466
rect 32114 48414 32116 48466
rect 32060 48402 32116 48414
rect 31948 48356 32004 48366
rect 31948 48262 32004 48300
rect 32956 48132 33012 48142
rect 32060 48020 32116 48030
rect 31836 48018 32116 48020
rect 31836 47966 32062 48018
rect 32114 47966 32116 48018
rect 31836 47964 32116 47966
rect 32060 47954 32116 47964
rect 31276 47682 31556 47684
rect 31276 47630 31278 47682
rect 31330 47630 31556 47682
rect 31276 47628 31556 47630
rect 31276 47618 31332 47628
rect 31164 47518 31166 47570
rect 31218 47518 31220 47570
rect 30828 47506 30884 47516
rect 31164 47506 31220 47518
rect 29820 47406 29822 47458
rect 29874 47406 29876 47458
rect 28028 47394 28084 47404
rect 29260 47394 29316 47404
rect 29820 47394 29876 47406
rect 32956 47236 33012 48076
rect 31724 46786 31780 46798
rect 31724 46734 31726 46786
rect 31778 46734 31780 46786
rect 28140 46674 28196 46686
rect 28140 46622 28142 46674
rect 28194 46622 28196 46674
rect 27356 46564 27412 46574
rect 28140 46564 28196 46622
rect 30156 46676 30212 46686
rect 28588 46564 28644 46574
rect 28140 46562 28644 46564
rect 28140 46510 28590 46562
rect 28642 46510 28644 46562
rect 28140 46508 28644 46510
rect 27356 46470 27412 46508
rect 27916 46004 27972 46014
rect 26684 45668 26740 45678
rect 26684 45574 26740 45612
rect 27132 44994 27188 45006
rect 27132 44942 27134 44994
rect 27186 44942 27188 44994
rect 27132 43540 27188 44942
rect 27580 44884 27636 44894
rect 27580 44434 27636 44828
rect 27580 44382 27582 44434
rect 27634 44382 27636 44434
rect 27580 44370 27636 44382
rect 27244 43652 27300 43662
rect 27244 43558 27300 43596
rect 27916 43650 27972 45948
rect 28364 44322 28420 44334
rect 28364 44270 28366 44322
rect 28418 44270 28420 44322
rect 28364 44100 28420 44270
rect 28588 44100 28644 46508
rect 29820 46004 29876 46014
rect 29820 45892 29876 45948
rect 29820 45890 30100 45892
rect 29820 45838 29822 45890
rect 29874 45838 30100 45890
rect 29820 45836 30100 45838
rect 29820 45826 29876 45836
rect 28924 45668 28980 45678
rect 28700 44100 28756 44110
rect 28364 44044 28700 44100
rect 28700 44034 28756 44044
rect 28924 43988 28980 45612
rect 29596 45106 29652 45118
rect 29596 45054 29598 45106
rect 29650 45054 29652 45106
rect 29260 44996 29316 45006
rect 29260 44902 29316 44940
rect 28812 43932 28980 43988
rect 29260 44100 29316 44110
rect 29596 44100 29652 45054
rect 29316 44044 29652 44100
rect 27916 43598 27918 43650
rect 27970 43598 27972 43650
rect 27916 43586 27972 43598
rect 28252 43650 28308 43662
rect 28252 43598 28254 43650
rect 28306 43598 28308 43650
rect 27132 43474 27188 43484
rect 27580 43540 27636 43550
rect 27580 43538 27748 43540
rect 27580 43486 27582 43538
rect 27634 43486 27748 43538
rect 27580 43484 27748 43486
rect 27580 43474 27636 43484
rect 26460 42814 26462 42866
rect 26514 42814 26516 42866
rect 26460 42308 26516 42814
rect 26460 42242 26516 42252
rect 27692 43316 27748 43484
rect 28252 43316 28308 43598
rect 28700 43652 28756 43662
rect 28700 43558 28756 43596
rect 28588 43540 28644 43550
rect 28588 43426 28644 43484
rect 28588 43374 28590 43426
rect 28642 43374 28644 43426
rect 28588 43362 28644 43374
rect 27692 43260 28308 43316
rect 27692 42532 27748 43260
rect 28812 43092 28868 43932
rect 28924 43316 28980 43326
rect 28924 43314 29092 43316
rect 28924 43262 28926 43314
rect 28978 43262 29092 43314
rect 28924 43260 29092 43262
rect 28924 43250 28980 43260
rect 28812 43036 28980 43092
rect 27804 42532 27860 42542
rect 27692 42530 27860 42532
rect 27692 42478 27806 42530
rect 27858 42478 27860 42530
rect 27692 42476 27860 42478
rect 25564 41972 25620 41982
rect 25900 41972 25956 41982
rect 25340 41970 25956 41972
rect 25340 41918 25566 41970
rect 25618 41918 25902 41970
rect 25954 41918 25956 41970
rect 25340 41916 25956 41918
rect 25340 41186 25396 41916
rect 25564 41906 25620 41916
rect 25900 41906 25956 41916
rect 26684 41860 26740 41870
rect 26460 41858 26740 41860
rect 26460 41806 26686 41858
rect 26738 41806 26740 41858
rect 26460 41804 26740 41806
rect 25340 41134 25342 41186
rect 25394 41134 25396 41186
rect 25340 41122 25396 41134
rect 25676 41298 25732 41310
rect 25676 41246 25678 41298
rect 25730 41246 25732 41298
rect 25676 40516 25732 41246
rect 26460 40626 26516 41804
rect 26684 41794 26740 41804
rect 26460 40574 26462 40626
rect 26514 40574 26516 40626
rect 26460 40562 26516 40574
rect 25676 40450 25732 40460
rect 27580 40514 27636 40526
rect 27580 40462 27582 40514
rect 27634 40462 27636 40514
rect 26348 40402 26404 40414
rect 26348 40350 26350 40402
rect 26402 40350 26404 40402
rect 26348 39956 26404 40350
rect 26348 39890 26404 39900
rect 26460 40404 26516 40414
rect 26348 39732 26404 39742
rect 26460 39732 26516 40348
rect 26572 40402 26628 40414
rect 26572 40350 26574 40402
rect 26626 40350 26628 40402
rect 26572 40292 26628 40350
rect 26908 40402 26964 40414
rect 26908 40350 26910 40402
rect 26962 40350 26964 40402
rect 26628 40236 26740 40292
rect 26572 40226 26628 40236
rect 26348 39730 26516 39732
rect 26348 39678 26350 39730
rect 26402 39678 26516 39730
rect 26348 39676 26516 39678
rect 26572 39956 26628 39966
rect 26348 39666 26404 39676
rect 26572 39618 26628 39900
rect 26572 39566 26574 39618
rect 26626 39566 26628 39618
rect 25228 39508 25284 39518
rect 25228 39172 25284 39452
rect 26236 39394 26292 39406
rect 26236 39342 26238 39394
rect 26290 39342 26292 39394
rect 26236 39284 26292 39342
rect 26236 39218 26292 39228
rect 26460 39394 26516 39406
rect 26460 39342 26462 39394
rect 26514 39342 26516 39394
rect 25228 38946 25284 39116
rect 26460 39060 26516 39342
rect 25228 38894 25230 38946
rect 25282 38894 25284 38946
rect 25228 38882 25284 38894
rect 25900 39004 26516 39060
rect 25340 38836 25396 38846
rect 25340 38742 25396 38780
rect 25004 38612 25172 38668
rect 25228 38724 25284 38734
rect 24892 38276 24948 38286
rect 24892 38050 24948 38220
rect 24892 37998 24894 38050
rect 24946 37998 24948 38050
rect 24892 37986 24948 37998
rect 24892 37826 24948 37838
rect 24892 37774 24894 37826
rect 24946 37774 24948 37826
rect 24892 35700 24948 37774
rect 24892 35634 24948 35644
rect 24892 35364 24948 35374
rect 24892 34804 24948 35308
rect 24892 34738 24948 34748
rect 24780 32722 24836 32732
rect 25004 32676 25060 38612
rect 25228 38050 25284 38668
rect 25228 37998 25230 38050
rect 25282 37998 25284 38050
rect 25228 37986 25284 37998
rect 25676 38050 25732 38062
rect 25676 37998 25678 38050
rect 25730 37998 25732 38050
rect 25676 37604 25732 37998
rect 25676 37538 25732 37548
rect 25900 37826 25956 39004
rect 26572 38948 26628 39566
rect 26684 39060 26740 40236
rect 26908 39956 26964 40350
rect 27580 40292 27636 40462
rect 27580 40226 27636 40236
rect 27692 40180 27748 42476
rect 27804 42466 27860 42476
rect 27916 41860 27972 41870
rect 27804 41074 27860 41086
rect 27804 41022 27806 41074
rect 27858 41022 27860 41074
rect 27804 40404 27860 41022
rect 27916 40628 27972 41804
rect 28812 41860 28868 41870
rect 28812 41766 28868 41804
rect 28588 41188 28644 41198
rect 28588 41094 28644 41132
rect 28924 40852 28980 43036
rect 29036 40964 29092 43260
rect 29148 41972 29204 41982
rect 29148 41858 29204 41916
rect 29148 41806 29150 41858
rect 29202 41806 29204 41858
rect 29148 41794 29204 41806
rect 29260 41188 29316 44044
rect 30044 43652 30100 45836
rect 30156 45778 30212 46620
rect 30156 45726 30158 45778
rect 30210 45726 30212 45778
rect 30156 45714 30212 45726
rect 30828 46676 30884 46686
rect 30380 44994 30436 45006
rect 30380 44942 30382 44994
rect 30434 44942 30436 44994
rect 30380 44436 30436 44942
rect 30380 44370 30436 44380
rect 30156 43652 30212 43662
rect 30044 43650 30212 43652
rect 30044 43598 30158 43650
rect 30210 43598 30212 43650
rect 30044 43596 30212 43598
rect 30156 43586 30212 43596
rect 30492 43652 30548 43662
rect 30492 43558 30548 43596
rect 30828 42868 30884 46620
rect 31388 46676 31444 46686
rect 31388 46582 31444 46620
rect 31052 46564 31108 46574
rect 31052 45668 31108 46508
rect 31724 46116 31780 46734
rect 32060 46674 32116 46686
rect 32060 46622 32062 46674
rect 32114 46622 32116 46674
rect 32060 46564 32116 46622
rect 32060 46498 32116 46508
rect 32284 46562 32340 46574
rect 32284 46510 32286 46562
rect 32338 46510 32340 46562
rect 32284 46116 32340 46510
rect 32396 46452 32452 46462
rect 32396 46358 32452 46396
rect 32284 46060 32676 46116
rect 31724 46050 31780 46060
rect 32620 46002 32676 46060
rect 32620 45950 32622 46002
rect 32674 45950 32676 46002
rect 32620 45938 32676 45950
rect 31948 45892 32004 45902
rect 31948 45798 32004 45836
rect 31052 45602 31108 45612
rect 31388 44996 31444 45006
rect 31052 44434 31108 44446
rect 31052 44382 31054 44434
rect 31106 44382 31108 44434
rect 31052 44212 31108 44382
rect 31388 44324 31444 44940
rect 32508 44994 32564 45006
rect 32508 44942 32510 44994
rect 32562 44942 32564 44994
rect 32508 44434 32564 44942
rect 32508 44382 32510 44434
rect 32562 44382 32564 44434
rect 31388 44230 31444 44268
rect 32172 44324 32228 44334
rect 32172 44230 32228 44268
rect 32508 44324 32564 44382
rect 32508 44258 32564 44268
rect 31052 44146 31108 44156
rect 32844 44210 32900 44222
rect 32844 44158 32846 44210
rect 32898 44158 32900 44210
rect 31948 43652 32004 43662
rect 30828 42812 30996 42868
rect 30716 42756 30772 42766
rect 30772 42700 30884 42756
rect 30716 42690 30772 42700
rect 30604 42642 30660 42654
rect 30604 42590 30606 42642
rect 30658 42590 30660 42642
rect 30604 41298 30660 42590
rect 30828 42642 30884 42700
rect 30828 42590 30830 42642
rect 30882 42590 30884 42642
rect 30828 41972 30884 42590
rect 30828 41906 30884 41916
rect 30604 41246 30606 41298
rect 30658 41246 30660 41298
rect 30604 41234 30660 41246
rect 29260 41094 29316 41132
rect 30828 41074 30884 41086
rect 30828 41022 30830 41074
rect 30882 41022 30884 41074
rect 29036 40908 30212 40964
rect 28924 40796 29428 40852
rect 27916 40626 28084 40628
rect 27916 40574 27918 40626
rect 27970 40574 28084 40626
rect 27916 40572 28084 40574
rect 27916 40562 27972 40572
rect 27804 40338 27860 40348
rect 27692 40124 27972 40180
rect 26796 39900 26964 39956
rect 26796 39508 26852 39900
rect 26908 39732 26964 39742
rect 27580 39732 27636 39742
rect 26908 39730 27636 39732
rect 26908 39678 26910 39730
rect 26962 39678 27582 39730
rect 27634 39678 27636 39730
rect 26908 39676 27636 39678
rect 26908 39666 26964 39676
rect 27580 39666 27636 39676
rect 27804 39618 27860 39630
rect 27804 39566 27806 39618
rect 27858 39566 27860 39618
rect 26796 39452 27076 39508
rect 26684 38994 26740 39004
rect 26796 39284 26852 39294
rect 26572 38882 26628 38892
rect 26348 38836 26404 38846
rect 26236 38724 26292 38734
rect 26236 38050 26292 38668
rect 26236 37998 26238 38050
rect 26290 37998 26292 38050
rect 26236 37986 26292 37998
rect 25900 37774 25902 37826
rect 25954 37774 25956 37826
rect 25788 37266 25844 37278
rect 25788 37214 25790 37266
rect 25842 37214 25844 37266
rect 25788 36484 25844 37214
rect 25900 36820 25956 37774
rect 26348 37828 26404 38780
rect 26684 38836 26740 38846
rect 26796 38836 26852 39228
rect 27020 39058 27076 39452
rect 27020 39006 27022 39058
rect 27074 39006 27076 39058
rect 27020 38994 27076 39006
rect 27692 39172 27748 39182
rect 26684 38834 26852 38836
rect 26684 38782 26686 38834
rect 26738 38782 26852 38834
rect 26684 38780 26852 38782
rect 27132 38948 27188 38958
rect 26684 38770 26740 38780
rect 26460 38722 26516 38734
rect 26460 38670 26462 38722
rect 26514 38670 26516 38722
rect 26460 38668 26516 38670
rect 26460 38612 26852 38668
rect 27132 38612 27188 38892
rect 27580 38946 27636 38958
rect 27580 38894 27582 38946
rect 27634 38894 27636 38946
rect 27468 38836 27524 38846
rect 27468 38742 27524 38780
rect 26796 38556 27188 38612
rect 27580 38612 27636 38894
rect 26572 37828 26628 37838
rect 26684 37828 26740 37838
rect 26348 37826 26516 37828
rect 26348 37774 26350 37826
rect 26402 37774 26516 37826
rect 26348 37772 26516 37774
rect 26348 37762 26404 37772
rect 26348 37604 26404 37614
rect 26348 37154 26404 37548
rect 26460 37266 26516 37772
rect 26572 37826 26684 37828
rect 26572 37774 26574 37826
rect 26626 37774 26684 37826
rect 26572 37772 26684 37774
rect 26572 37762 26628 37772
rect 26460 37214 26462 37266
rect 26514 37214 26516 37266
rect 26460 37202 26516 37214
rect 26348 37102 26350 37154
rect 26402 37102 26404 37154
rect 26348 37090 26404 37102
rect 26236 36820 26292 36830
rect 25900 36764 26236 36820
rect 26236 36754 26292 36764
rect 26236 36484 26292 36494
rect 25788 36482 26292 36484
rect 25788 36430 26238 36482
rect 26290 36430 26292 36482
rect 25788 36428 26292 36430
rect 25676 36372 25732 36382
rect 25452 36316 25676 36372
rect 25340 34692 25396 34702
rect 25340 34598 25396 34636
rect 25340 34356 25396 34366
rect 25452 34356 25508 36316
rect 25676 36306 25732 36316
rect 25676 35698 25732 35710
rect 25676 35646 25678 35698
rect 25730 35646 25732 35698
rect 25676 35140 25732 35646
rect 25900 35308 25956 36428
rect 26236 36418 26292 36428
rect 26460 36484 26516 36494
rect 26684 36484 26740 37772
rect 26796 37268 26852 38556
rect 27580 38546 27636 38556
rect 27692 37938 27748 39116
rect 27804 39058 27860 39566
rect 27804 39006 27806 39058
rect 27858 39006 27860 39058
rect 27804 38994 27860 39006
rect 27692 37886 27694 37938
rect 27746 37886 27748 37938
rect 27692 37874 27748 37886
rect 27804 37940 27860 37950
rect 27804 37846 27860 37884
rect 27468 37826 27524 37838
rect 27468 37774 27470 37826
rect 27522 37774 27524 37826
rect 27356 37268 27412 37278
rect 26796 37212 27076 37268
rect 26796 37042 26852 37054
rect 26796 36990 26798 37042
rect 26850 36990 26852 37042
rect 26796 36708 26852 36990
rect 26796 36642 26852 36652
rect 26908 36820 26964 36830
rect 26460 36260 26516 36428
rect 26124 36204 26516 36260
rect 26572 36428 26740 36484
rect 26908 36482 26964 36764
rect 26908 36430 26910 36482
rect 26962 36430 26964 36482
rect 26124 35308 26180 36204
rect 26572 36036 26628 36428
rect 26796 36372 26852 36382
rect 26796 36278 26852 36316
rect 26684 36258 26740 36270
rect 26684 36206 26686 36258
rect 26738 36206 26740 36258
rect 26684 36148 26740 36206
rect 26684 36082 26740 36092
rect 26348 35980 26628 36036
rect 25788 35252 25956 35308
rect 26012 35252 26180 35308
rect 26236 35924 26292 35934
rect 25788 35140 25844 35252
rect 25900 35140 25956 35150
rect 25788 35084 25900 35140
rect 25676 35074 25732 35084
rect 25900 35074 25956 35084
rect 25676 34916 25732 34926
rect 25676 34822 25732 34860
rect 26012 34916 26068 35252
rect 26012 34850 26068 34860
rect 25340 34354 25508 34356
rect 25340 34302 25342 34354
rect 25394 34302 25508 34354
rect 25340 34300 25508 34302
rect 26012 34692 26068 34702
rect 25340 34290 25396 34300
rect 25676 34244 25732 34254
rect 25564 34188 25676 34244
rect 25228 34130 25284 34142
rect 25228 34078 25230 34130
rect 25282 34078 25284 34130
rect 24556 32622 24558 32674
rect 24610 32622 24612 32674
rect 24556 32004 24612 32622
rect 24892 32620 25060 32676
rect 25116 33348 25172 33358
rect 25228 33348 25284 34078
rect 25564 34130 25620 34188
rect 25676 34178 25732 34188
rect 25564 34078 25566 34130
rect 25618 34078 25620 34130
rect 25564 34066 25620 34078
rect 26012 33908 26068 34636
rect 26236 34130 26292 35868
rect 26348 34802 26404 35980
rect 26796 35812 26852 35822
rect 26796 35718 26852 35756
rect 26684 35700 26740 35710
rect 26572 35698 26740 35700
rect 26572 35646 26686 35698
rect 26738 35646 26740 35698
rect 26572 35644 26740 35646
rect 26460 34916 26516 34926
rect 26460 34822 26516 34860
rect 26348 34750 26350 34802
rect 26402 34750 26404 34802
rect 26348 34738 26404 34750
rect 26236 34078 26238 34130
rect 26290 34078 26292 34130
rect 26236 34066 26292 34078
rect 25340 33348 25396 33358
rect 25228 33346 25396 33348
rect 25228 33294 25342 33346
rect 25394 33294 25396 33346
rect 25228 33292 25396 33294
rect 24556 31938 24612 31948
rect 24780 32564 24836 32574
rect 24332 31612 24500 31668
rect 24668 31890 24724 31902
rect 24668 31838 24670 31890
rect 24722 31838 24724 31890
rect 22540 29708 22932 29764
rect 22092 29650 22708 29652
rect 22092 29598 22094 29650
rect 22146 29598 22708 29650
rect 22092 29596 22708 29598
rect 22092 29586 22148 29596
rect 22540 29426 22596 29438
rect 22540 29374 22542 29426
rect 22594 29374 22596 29426
rect 22540 29316 22596 29374
rect 22540 29250 22596 29260
rect 22092 28644 22148 28654
rect 21868 28642 22148 28644
rect 21868 28590 22094 28642
rect 22146 28590 22148 28642
rect 21868 28588 22148 28590
rect 22092 28578 22148 28588
rect 22652 28642 22708 29596
rect 22876 29650 22932 29708
rect 22876 29598 22878 29650
rect 22930 29598 22932 29650
rect 22876 29586 22932 29598
rect 23548 29650 23604 30156
rect 23996 30996 24052 31006
rect 24332 30996 24388 31612
rect 24556 31444 24612 31454
rect 23996 30882 24052 30940
rect 23996 30830 23998 30882
rect 24050 30830 24052 30882
rect 23996 30210 24052 30830
rect 24220 30940 24388 30996
rect 24444 31332 24500 31342
rect 24220 30660 24276 30940
rect 24332 30772 24388 30782
rect 24332 30678 24388 30716
rect 24220 30594 24276 30604
rect 23996 30158 23998 30210
rect 24050 30158 24052 30210
rect 23996 30146 24052 30158
rect 24332 30212 24388 30222
rect 24444 30212 24500 31276
rect 24556 31106 24612 31388
rect 24556 31054 24558 31106
rect 24610 31054 24612 31106
rect 24556 31042 24612 31054
rect 24332 30210 24500 30212
rect 24332 30158 24334 30210
rect 24386 30158 24500 30210
rect 24332 30156 24500 30158
rect 24668 30436 24724 31838
rect 24780 31778 24836 32508
rect 24780 31726 24782 31778
rect 24834 31726 24836 31778
rect 24780 31714 24836 31726
rect 24892 31220 24948 32620
rect 25116 32564 25172 33292
rect 25340 33282 25396 33292
rect 25676 33234 25732 33246
rect 25676 33182 25678 33234
rect 25730 33182 25732 33234
rect 25452 33124 25508 33134
rect 25116 32498 25172 32508
rect 25228 32900 25284 32910
rect 25228 32786 25284 32844
rect 25228 32734 25230 32786
rect 25282 32734 25284 32786
rect 25004 32452 25060 32462
rect 25004 32002 25060 32396
rect 25004 31950 25006 32002
rect 25058 31950 25060 32002
rect 25004 31938 25060 31950
rect 24892 31154 24948 31164
rect 25004 31444 25060 31454
rect 24892 30772 24948 30782
rect 24780 30436 24836 30446
rect 24668 30434 24836 30436
rect 24668 30382 24782 30434
rect 24834 30382 24836 30434
rect 24668 30380 24836 30382
rect 24332 30146 24388 30156
rect 24108 29988 24164 29998
rect 24668 29988 24724 30380
rect 24780 30370 24836 30380
rect 24892 30324 24948 30716
rect 24892 30210 24948 30268
rect 24892 30158 24894 30210
rect 24946 30158 24948 30210
rect 24892 30146 24948 30158
rect 24108 29986 24724 29988
rect 24108 29934 24110 29986
rect 24162 29934 24724 29986
rect 24108 29932 24724 29934
rect 24780 29988 24836 29998
rect 25004 29988 25060 31388
rect 25228 30996 25284 32734
rect 25452 32676 25508 33068
rect 25564 33122 25620 33134
rect 25564 33070 25566 33122
rect 25618 33070 25620 33122
rect 25564 32788 25620 33070
rect 25676 33124 25732 33182
rect 26012 33234 26068 33852
rect 26012 33182 26014 33234
rect 26066 33182 26068 33234
rect 26012 33170 26068 33182
rect 26236 33346 26292 33358
rect 26236 33294 26238 33346
rect 26290 33294 26292 33346
rect 26236 33236 26292 33294
rect 26236 33170 26292 33180
rect 25676 33058 25732 33068
rect 26124 32788 26180 32798
rect 25564 32786 26404 32788
rect 25564 32734 26126 32786
rect 26178 32734 26404 32786
rect 25564 32732 26404 32734
rect 25452 32610 25508 32620
rect 25340 32562 25396 32574
rect 25788 32564 25844 32574
rect 25340 32510 25342 32562
rect 25394 32510 25396 32562
rect 25340 31780 25396 32510
rect 25340 31220 25396 31724
rect 25340 31154 25396 31164
rect 25564 32508 25788 32564
rect 25340 30996 25396 31006
rect 25228 30994 25396 30996
rect 25228 30942 25342 30994
rect 25394 30942 25396 30994
rect 25228 30940 25396 30942
rect 25340 30930 25396 30940
rect 25564 30324 25620 32508
rect 25788 32470 25844 32508
rect 25900 32004 25956 32014
rect 25900 31890 25956 31948
rect 25900 31838 25902 31890
rect 25954 31838 25956 31890
rect 25788 31778 25844 31790
rect 25788 31726 25790 31778
rect 25842 31726 25844 31778
rect 25788 31444 25844 31726
rect 25900 31780 25956 31838
rect 25900 31714 25956 31724
rect 25788 31378 25844 31388
rect 26012 31218 26068 32732
rect 26124 32722 26180 32732
rect 26348 32674 26404 32732
rect 26348 32622 26350 32674
rect 26402 32622 26404 32674
rect 26348 32610 26404 32622
rect 26012 31166 26014 31218
rect 26066 31166 26068 31218
rect 26012 31154 26068 31166
rect 26124 32564 26180 32574
rect 25340 30268 25620 30324
rect 25788 30994 25844 31006
rect 25788 30942 25790 30994
rect 25842 30942 25844 30994
rect 25228 30212 25284 30222
rect 25228 30118 25284 30156
rect 25340 30210 25396 30268
rect 25788 30212 25844 30942
rect 25900 30996 25956 31006
rect 26124 30996 26180 32508
rect 26572 31892 26628 35644
rect 26684 35634 26740 35644
rect 26908 35364 26964 36430
rect 27020 36148 27076 37212
rect 27020 36082 27076 36092
rect 27244 37266 27412 37268
rect 27244 37214 27358 37266
rect 27410 37214 27412 37266
rect 27244 37212 27412 37214
rect 27244 37156 27300 37212
rect 27356 37202 27412 37212
rect 26796 35308 26964 35364
rect 26796 34916 26852 35308
rect 26796 34850 26852 34860
rect 27132 34916 27188 34926
rect 27244 34916 27300 37100
rect 27468 36932 27524 37774
rect 27580 37380 27636 37418
rect 27580 37314 27636 37324
rect 27804 37380 27860 37390
rect 27692 37266 27748 37278
rect 27692 37214 27694 37266
rect 27746 37214 27748 37266
rect 27692 36932 27748 37214
rect 27468 36876 27748 36932
rect 27580 36484 27636 36876
rect 27804 36820 27860 37324
rect 27580 36418 27636 36428
rect 27692 36764 27860 36820
rect 27692 35698 27748 36764
rect 27804 36260 27860 36270
rect 27804 36166 27860 36204
rect 27804 36036 27860 36046
rect 27804 35810 27860 35980
rect 27804 35758 27806 35810
rect 27858 35758 27860 35810
rect 27804 35746 27860 35758
rect 27692 35646 27694 35698
rect 27746 35646 27748 35698
rect 27692 35634 27748 35646
rect 27468 35586 27524 35598
rect 27468 35534 27470 35586
rect 27522 35534 27524 35586
rect 27356 34916 27412 34926
rect 27244 34914 27412 34916
rect 27244 34862 27358 34914
rect 27410 34862 27412 34914
rect 27244 34860 27412 34862
rect 27132 34822 27188 34860
rect 27356 34850 27412 34860
rect 26796 34692 26852 34702
rect 26684 34690 26852 34692
rect 26684 34638 26798 34690
rect 26850 34638 26852 34690
rect 26684 34636 26852 34638
rect 26684 33346 26740 34636
rect 26796 34626 26852 34636
rect 26908 34692 26964 34702
rect 26908 34598 26964 34636
rect 26908 34244 26964 34254
rect 26908 34150 26964 34188
rect 26796 34130 26852 34142
rect 26796 34078 26798 34130
rect 26850 34078 26852 34130
rect 26796 33796 26852 34078
rect 26796 33730 26852 33740
rect 27020 33908 27076 33918
rect 26684 33294 26686 33346
rect 26738 33294 26740 33346
rect 26684 33282 26740 33294
rect 26908 33684 26964 33694
rect 26908 33346 26964 33628
rect 26908 33294 26910 33346
rect 26962 33294 26964 33346
rect 26908 33282 26964 33294
rect 27020 33124 27076 33852
rect 27468 33572 27524 35534
rect 27804 35588 27860 35598
rect 27804 34916 27860 35532
rect 27916 35140 27972 40124
rect 28028 39844 28084 40572
rect 28084 39788 28308 39844
rect 28028 39778 28084 39788
rect 28028 39620 28084 39630
rect 28084 39564 28196 39620
rect 28028 39526 28084 39564
rect 28028 39172 28084 39182
rect 28028 39058 28084 39116
rect 28028 39006 28030 39058
rect 28082 39006 28084 39058
rect 28028 38994 28084 39006
rect 28140 37492 28196 39564
rect 28252 38164 28308 39788
rect 28364 38946 28420 38958
rect 28364 38894 28366 38946
rect 28418 38894 28420 38946
rect 28364 38668 28420 38894
rect 28924 38948 28980 38958
rect 28924 38854 28980 38892
rect 29260 38834 29316 38846
rect 29260 38782 29262 38834
rect 29314 38782 29316 38834
rect 28364 38612 28644 38668
rect 28364 38546 28420 38556
rect 28476 38164 28532 38174
rect 28252 38162 28532 38164
rect 28252 38110 28478 38162
rect 28530 38110 28532 38162
rect 28252 38108 28532 38110
rect 28476 38098 28532 38108
rect 28588 38052 28644 38612
rect 28364 37940 28420 37950
rect 28364 37846 28420 37884
rect 28252 37492 28308 37502
rect 28140 37436 28252 37492
rect 28252 37398 28308 37436
rect 28476 37266 28532 37278
rect 28476 37214 28478 37266
rect 28530 37214 28532 37266
rect 28364 37154 28420 37166
rect 28364 37102 28366 37154
rect 28418 37102 28420 37154
rect 28364 36708 28420 37102
rect 28476 37156 28532 37214
rect 28588 37156 28644 37996
rect 29148 38050 29204 38062
rect 29148 37998 29150 38050
rect 29202 37998 29204 38050
rect 29148 37492 29204 37998
rect 29260 37940 29316 38782
rect 29260 37846 29316 37884
rect 29148 37426 29204 37436
rect 28924 37266 28980 37278
rect 28924 37214 28926 37266
rect 28978 37214 28980 37266
rect 28476 37100 28756 37156
rect 28140 36652 28420 36708
rect 28140 36370 28196 36652
rect 28588 36594 28644 36606
rect 28588 36542 28590 36594
rect 28642 36542 28644 36594
rect 28140 36318 28142 36370
rect 28194 36318 28196 36370
rect 28140 36306 28196 36318
rect 28476 36482 28532 36494
rect 28476 36430 28478 36482
rect 28530 36430 28532 36482
rect 28028 36258 28084 36270
rect 28028 36206 28030 36258
rect 28082 36206 28084 36258
rect 28028 35700 28084 36206
rect 28252 35700 28308 35710
rect 28028 35698 28308 35700
rect 28028 35646 28254 35698
rect 28306 35646 28308 35698
rect 28028 35644 28308 35646
rect 28252 35364 28308 35644
rect 28476 35476 28532 36430
rect 28588 36484 28644 36542
rect 28588 36418 28644 36428
rect 28588 35700 28644 35710
rect 28588 35606 28644 35644
rect 28476 35420 28644 35476
rect 28252 35298 28308 35308
rect 28588 35140 28644 35420
rect 27916 35084 28196 35140
rect 27916 34916 27972 34926
rect 27804 34914 27972 34916
rect 27804 34862 27918 34914
rect 27970 34862 27972 34914
rect 27804 34860 27972 34862
rect 27916 34850 27972 34860
rect 27580 34692 27636 34702
rect 27804 34692 27860 34702
rect 27580 34690 27748 34692
rect 27580 34638 27582 34690
rect 27634 34638 27748 34690
rect 27580 34636 27748 34638
rect 27580 34626 27636 34636
rect 27692 34356 27748 34636
rect 27804 34598 27860 34636
rect 27692 34300 27860 34356
rect 27580 34242 27636 34254
rect 27580 34190 27582 34242
rect 27634 34190 27636 34242
rect 27580 33908 27636 34190
rect 27580 33842 27636 33852
rect 27804 33572 27860 34300
rect 27468 33516 27636 33572
rect 27468 33348 27524 33358
rect 27468 33254 27524 33292
rect 27356 33236 27412 33246
rect 27356 33142 27412 33180
rect 26908 33068 27076 33124
rect 27132 33124 27188 33134
rect 27580 33124 27636 33516
rect 27804 33506 27860 33516
rect 27916 34130 27972 34142
rect 27916 34078 27918 34130
rect 27970 34078 27972 34130
rect 27692 33460 27748 33470
rect 27692 33236 27748 33404
rect 27692 33170 27748 33180
rect 27132 33122 27300 33124
rect 27132 33070 27134 33122
rect 27186 33070 27300 33122
rect 27132 33068 27300 33070
rect 26684 32676 26740 32686
rect 26684 32674 26852 32676
rect 26684 32622 26686 32674
rect 26738 32622 26852 32674
rect 26684 32620 26852 32622
rect 26684 32610 26740 32620
rect 26348 31836 26628 31892
rect 26796 32562 26852 32620
rect 26796 32510 26798 32562
rect 26850 32510 26852 32562
rect 26236 31668 26292 31678
rect 26236 31574 26292 31612
rect 25900 30994 26180 30996
rect 25900 30942 25902 30994
rect 25954 30942 26180 30994
rect 25900 30940 26180 30942
rect 25900 30930 25956 30940
rect 25340 30158 25342 30210
rect 25394 30158 25396 30210
rect 24780 29986 25060 29988
rect 24780 29934 24782 29986
rect 24834 29934 25060 29986
rect 24780 29932 25060 29934
rect 24108 29922 24164 29932
rect 24780 29922 24836 29932
rect 25340 29764 25396 30158
rect 23548 29598 23550 29650
rect 23602 29598 23604 29650
rect 23548 29586 23604 29598
rect 25228 29708 25396 29764
rect 25452 30210 25844 30212
rect 25452 30158 25790 30210
rect 25842 30158 25844 30210
rect 25452 30156 25844 30158
rect 23660 29540 23716 29550
rect 23436 28868 23492 28878
rect 22652 28590 22654 28642
rect 22706 28590 22708 28642
rect 22652 28578 22708 28590
rect 23100 28866 23492 28868
rect 23100 28814 23438 28866
rect 23490 28814 23492 28866
rect 23100 28812 23492 28814
rect 23100 28642 23156 28812
rect 23436 28802 23492 28812
rect 23660 28644 23716 29484
rect 25228 29316 25284 29708
rect 25228 29250 25284 29260
rect 25340 29540 25396 29550
rect 25452 29540 25508 30156
rect 25788 30146 25844 30156
rect 26348 30212 26404 31836
rect 26796 31778 26852 32510
rect 26796 31726 26798 31778
rect 26850 31726 26852 31778
rect 26796 31714 26852 31726
rect 26460 31666 26516 31678
rect 26460 31614 26462 31666
rect 26514 31614 26516 31666
rect 26460 31220 26516 31614
rect 26572 31556 26628 31566
rect 26572 31462 26628 31500
rect 26460 31154 26516 31164
rect 26348 30146 26404 30156
rect 26684 30994 26740 31006
rect 26684 30942 26686 30994
rect 26738 30942 26740 30994
rect 26684 30324 26740 30942
rect 26908 30772 26964 33068
rect 27132 33058 27188 33068
rect 27020 32788 27076 32798
rect 27244 32788 27300 33068
rect 27468 33068 27636 33124
rect 27804 33122 27860 33134
rect 27804 33070 27806 33122
rect 27858 33070 27860 33122
rect 27356 32788 27412 32798
rect 27244 32786 27412 32788
rect 27244 32734 27358 32786
rect 27410 32734 27412 32786
rect 27244 32732 27412 32734
rect 27020 32450 27076 32732
rect 27356 32722 27412 32732
rect 27020 32398 27022 32450
rect 27074 32398 27076 32450
rect 27020 32386 27076 32398
rect 27020 31780 27076 31790
rect 27020 30994 27076 31724
rect 27356 31780 27412 31790
rect 27356 31666 27412 31724
rect 27356 31614 27358 31666
rect 27410 31614 27412 31666
rect 27356 31602 27412 31614
rect 27468 31666 27524 33068
rect 27804 32900 27860 33070
rect 27580 32844 27860 32900
rect 27580 32730 27636 32844
rect 27580 32678 27582 32730
rect 27634 32678 27636 32730
rect 27804 32788 27860 32844
rect 27916 32788 27972 34078
rect 28028 34018 28084 34030
rect 28028 33966 28030 34018
rect 28082 33966 28084 34018
rect 28028 33460 28084 33966
rect 28028 33394 28084 33404
rect 27916 32732 28084 32788
rect 27580 32666 27636 32678
rect 27692 32676 27748 32686
rect 27692 32582 27748 32620
rect 27468 31614 27470 31666
rect 27522 31614 27524 31666
rect 27468 31602 27524 31614
rect 27132 31554 27188 31566
rect 27132 31502 27134 31554
rect 27186 31502 27188 31554
rect 27132 31332 27188 31502
rect 27132 31266 27188 31276
rect 27244 31554 27300 31566
rect 27244 31502 27246 31554
rect 27298 31502 27300 31554
rect 27020 30942 27022 30994
rect 27074 30942 27076 30994
rect 27020 30930 27076 30942
rect 27020 30772 27076 30782
rect 26908 30770 27076 30772
rect 26908 30718 27022 30770
rect 27074 30718 27076 30770
rect 26908 30716 27076 30718
rect 27020 30706 27076 30716
rect 26684 30098 26740 30268
rect 26684 30046 26686 30098
rect 26738 30046 26740 30098
rect 26684 30034 26740 30046
rect 25396 29484 25508 29540
rect 27020 29986 27076 29998
rect 27020 29934 27022 29986
rect 27074 29934 27076 29986
rect 23100 28590 23102 28642
rect 23154 28590 23156 28642
rect 23100 28578 23156 28590
rect 23436 28588 23716 28644
rect 24444 29204 24500 29214
rect 24444 28754 24500 29148
rect 24444 28702 24446 28754
rect 24498 28702 24500 28754
rect 21420 28466 21476 28476
rect 22428 28532 22484 28542
rect 22428 28438 22484 28476
rect 23324 28532 23380 28570
rect 23324 28466 23380 28476
rect 23436 28530 23492 28588
rect 23436 28478 23438 28530
rect 23490 28478 23492 28530
rect 23436 28466 23492 28478
rect 21868 28420 21924 28430
rect 21868 28326 21924 28364
rect 21980 28418 22036 28430
rect 21980 28366 21982 28418
rect 22034 28366 22036 28418
rect 21980 28084 22036 28366
rect 22540 28418 22596 28430
rect 22540 28366 22542 28418
rect 22594 28366 22596 28418
rect 22540 28308 22596 28366
rect 24108 28418 24164 28430
rect 24108 28366 24110 28418
rect 24162 28366 24164 28418
rect 22540 28242 22596 28252
rect 23324 28308 23380 28318
rect 21980 28028 22820 28084
rect 22764 27970 22820 28028
rect 22764 27918 22766 27970
rect 22818 27918 22820 27970
rect 22764 27906 22820 27918
rect 22876 27860 22932 27870
rect 20636 27748 20692 27758
rect 20524 27746 20692 27748
rect 20524 27694 20638 27746
rect 20690 27694 20692 27746
rect 20524 27692 20692 27694
rect 20300 27682 20356 27692
rect 20636 27682 20692 27692
rect 19292 27188 19348 27198
rect 18732 27186 19348 27188
rect 18732 27134 18734 27186
rect 18786 27134 19294 27186
rect 19346 27134 19348 27186
rect 18732 27132 19348 27134
rect 17948 27122 18004 27132
rect 18732 27122 18788 27132
rect 19292 27122 19348 27132
rect 22428 27188 22484 27198
rect 22876 27188 22932 27804
rect 22428 27186 22932 27188
rect 22428 27134 22430 27186
rect 22482 27134 22932 27186
rect 22428 27132 22932 27134
rect 17836 27010 17892 27020
rect 18060 26964 18116 26974
rect 17388 26852 17556 26908
rect 17724 26852 17892 26908
rect 16492 26516 16548 26526
rect 16380 26514 16548 26516
rect 16380 26462 16494 26514
rect 16546 26462 16548 26514
rect 16380 26460 16548 26462
rect 16492 26450 16548 26460
rect 17500 26402 17556 26852
rect 17500 26350 17502 26402
rect 17554 26350 17556 26402
rect 17500 26338 17556 26350
rect 15820 26290 15988 26292
rect 15820 26238 15822 26290
rect 15874 26238 15988 26290
rect 15820 26236 15988 26238
rect 16044 26290 16100 26302
rect 16044 26238 16046 26290
rect 16098 26238 16100 26290
rect 15820 26226 15876 26236
rect 15932 25508 15988 25518
rect 15708 25506 15988 25508
rect 15708 25454 15934 25506
rect 15986 25454 15988 25506
rect 15708 25452 15988 25454
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 15036 24658 15092 24670
rect 15148 25228 15428 25284
rect 14812 24612 14868 24622
rect 14700 24556 14812 24612
rect 14588 24164 14644 24174
rect 14700 24164 14756 24556
rect 14812 24546 14868 24556
rect 15148 24276 15204 25228
rect 15932 24948 15988 25452
rect 16044 25284 16100 26238
rect 16716 26292 16772 26302
rect 16716 26198 16772 26236
rect 17388 26292 17444 26302
rect 16604 26180 16660 26190
rect 16604 26086 16660 26124
rect 17388 26066 17444 26236
rect 17388 26014 17390 26066
rect 17442 26014 17444 26066
rect 17276 25618 17332 25630
rect 17276 25566 17278 25618
rect 17330 25566 17332 25618
rect 16044 25190 16100 25228
rect 16604 25506 16660 25518
rect 16604 25454 16606 25506
rect 16658 25454 16660 25506
rect 15932 24892 16212 24948
rect 16044 24724 16100 24734
rect 15484 24612 15540 24622
rect 15484 24610 15988 24612
rect 15484 24558 15486 24610
rect 15538 24558 15988 24610
rect 15484 24556 15988 24558
rect 15484 24546 15540 24556
rect 14588 24162 14756 24164
rect 14588 24110 14590 24162
rect 14642 24110 14756 24162
rect 14588 24108 14756 24110
rect 14812 24220 15204 24276
rect 14588 24098 14644 24108
rect 14028 24052 14084 24062
rect 14084 23996 14308 24052
rect 14028 23958 14084 23996
rect 13804 22390 13860 22428
rect 14140 23380 14196 23390
rect 14140 22594 14196 23324
rect 14252 23266 14308 23996
rect 14812 23938 14868 24220
rect 14812 23886 14814 23938
rect 14866 23886 14868 23938
rect 14476 23828 14532 23838
rect 14476 23734 14532 23772
rect 14252 23214 14254 23266
rect 14306 23214 14308 23266
rect 14252 23202 14308 23214
rect 14140 22542 14142 22594
rect 14194 22542 14196 22594
rect 11116 22318 11118 22370
rect 11170 22318 11172 22370
rect 11116 22306 11172 22318
rect 14140 22372 14196 22542
rect 14140 22306 14196 22316
rect 14252 22596 14308 22606
rect 14252 22482 14308 22540
rect 14252 22430 14254 22482
rect 14306 22430 14308 22482
rect 11676 22258 11732 22270
rect 11676 22206 11678 22258
rect 11730 22206 11732 22258
rect 11676 21924 11732 22206
rect 11676 21858 11732 21868
rect 14028 21924 14084 21934
rect 11340 21812 11396 21822
rect 11340 21698 11396 21756
rect 11340 21646 11342 21698
rect 11394 21646 11396 21698
rect 11340 21634 11396 21646
rect 12124 21812 12180 21822
rect 12124 21586 12180 21756
rect 12124 21534 12126 21586
rect 12178 21534 12180 21586
rect 12124 21522 12180 21534
rect 12012 21476 12068 21486
rect 11452 20692 11508 20702
rect 11788 20692 11844 20702
rect 11452 20690 11844 20692
rect 11452 20638 11454 20690
rect 11506 20638 11790 20690
rect 11842 20638 11844 20690
rect 11452 20636 11844 20638
rect 11452 20626 11508 20636
rect 11788 20626 11844 20636
rect 11228 20578 11284 20590
rect 11228 20526 11230 20578
rect 11282 20526 11284 20578
rect 11228 20468 11284 20526
rect 11340 20580 11396 20590
rect 11340 20486 11396 20524
rect 11228 20402 11284 20412
rect 12012 20468 12068 21420
rect 12572 21474 12628 21486
rect 12572 21422 12574 21474
rect 12626 21422 12628 21474
rect 12460 20916 12516 20926
rect 12460 20822 12516 20860
rect 12572 20804 12628 21422
rect 13020 21476 13076 21486
rect 13020 21382 13076 21420
rect 13468 21364 13524 21374
rect 13468 20916 13524 21308
rect 12572 20802 13412 20804
rect 12572 20750 12574 20802
rect 12626 20750 13412 20802
rect 12572 20748 13412 20750
rect 12572 20738 12628 20748
rect 10220 19294 10222 19346
rect 10274 19294 10276 19346
rect 10220 19282 10276 19294
rect 10668 20130 11060 20132
rect 10668 20078 11006 20130
rect 11058 20078 11060 20130
rect 10668 20076 11060 20078
rect 10668 19346 10724 20076
rect 11004 20066 11060 20076
rect 10668 19294 10670 19346
rect 10722 19294 10724 19346
rect 7420 19182 7422 19234
rect 7474 19182 7476 19234
rect 7420 18452 7476 19182
rect 7420 18386 7476 18396
rect 8428 18452 8484 18462
rect 7868 18228 7924 18238
rect 7868 17666 7924 18172
rect 7868 17614 7870 17666
rect 7922 17614 7924 17666
rect 7868 17602 7924 17614
rect 8428 17666 8484 18396
rect 9660 18452 9716 18462
rect 9660 18358 9716 18396
rect 10668 18452 10724 19294
rect 12012 19236 12068 20412
rect 13356 20242 13412 20748
rect 13356 20190 13358 20242
rect 13410 20190 13412 20242
rect 12124 20132 13188 20188
rect 12124 19906 12180 20132
rect 13132 20130 13188 20132
rect 13132 20078 13134 20130
rect 13186 20078 13188 20130
rect 13132 20066 13188 20078
rect 13356 20132 13412 20190
rect 13356 20066 13412 20076
rect 13468 20130 13524 20860
rect 13580 20914 13636 20926
rect 13580 20862 13582 20914
rect 13634 20862 13636 20914
rect 13580 20468 13636 20862
rect 14028 20804 14084 21868
rect 14252 21476 14308 22430
rect 14252 20804 14308 21420
rect 14588 22146 14644 22158
rect 14588 22094 14590 22146
rect 14642 22094 14644 22146
rect 14588 21364 14644 22094
rect 14812 21588 14868 23886
rect 15036 23940 15092 23950
rect 15820 23940 15876 23950
rect 15036 23938 15316 23940
rect 15036 23886 15038 23938
rect 15090 23886 15316 23938
rect 15036 23884 15316 23886
rect 15036 23874 15092 23884
rect 15260 23716 15316 23884
rect 15820 23846 15876 23884
rect 15932 23938 15988 24556
rect 15932 23886 15934 23938
rect 15986 23886 15988 23938
rect 15932 23828 15988 23886
rect 16044 24052 16100 24668
rect 16156 24388 16212 24892
rect 16380 24612 16436 24622
rect 16604 24612 16660 25454
rect 16380 24610 16660 24612
rect 16380 24558 16382 24610
rect 16434 24558 16660 24610
rect 16380 24556 16660 24558
rect 16380 24546 16436 24556
rect 16156 24322 16212 24332
rect 16492 24388 16548 24398
rect 16044 23938 16100 23996
rect 16044 23886 16046 23938
rect 16098 23886 16100 23938
rect 16044 23874 16100 23886
rect 16268 24164 16324 24174
rect 15932 23762 15988 23772
rect 15372 23716 15428 23726
rect 15260 23714 15428 23716
rect 15260 23662 15374 23714
rect 15426 23662 15428 23714
rect 15260 23660 15428 23662
rect 15148 23268 15204 23278
rect 15260 23268 15316 23660
rect 15372 23650 15428 23660
rect 14924 23266 15316 23268
rect 14924 23214 15150 23266
rect 15202 23214 15316 23266
rect 14924 23212 15316 23214
rect 15372 23266 15428 23278
rect 15372 23214 15374 23266
rect 15426 23214 15428 23266
rect 14924 22594 14980 23212
rect 15148 23174 15204 23212
rect 14924 22542 14926 22594
rect 14978 22542 14980 22594
rect 14924 22530 14980 22542
rect 15148 22596 15204 22606
rect 15148 22482 15204 22540
rect 15148 22430 15150 22482
rect 15202 22430 15204 22482
rect 15148 22418 15204 22430
rect 15372 21924 15428 23214
rect 15484 22930 15540 22942
rect 15484 22878 15486 22930
rect 15538 22878 15540 22930
rect 15484 22148 15540 22878
rect 15708 22372 15764 22382
rect 15708 22278 15764 22316
rect 15484 22082 15540 22092
rect 14812 21522 14868 21532
rect 15036 21868 15428 21924
rect 14588 21298 14644 21308
rect 14924 20916 14980 20926
rect 15036 20916 15092 21868
rect 16268 21700 16324 24108
rect 16492 23938 16548 24332
rect 16492 23886 16494 23938
rect 16546 23886 16548 23938
rect 16492 23874 16548 23886
rect 16268 21634 16324 21644
rect 16492 23266 16548 23278
rect 16492 23214 16494 23266
rect 16546 23214 16548 23266
rect 15820 21588 15876 21598
rect 15148 21474 15204 21486
rect 15148 21422 15150 21474
rect 15202 21422 15204 21474
rect 15148 21252 15204 21422
rect 15148 21186 15204 21196
rect 15596 20916 15652 20926
rect 14980 20860 15092 20916
rect 15148 20914 15652 20916
rect 15148 20862 15598 20914
rect 15650 20862 15652 20914
rect 15148 20860 15652 20862
rect 14924 20822 14980 20860
rect 14364 20804 14420 20814
rect 14252 20802 14420 20804
rect 14252 20750 14366 20802
rect 14418 20750 14420 20802
rect 14252 20748 14420 20750
rect 14028 20710 14084 20748
rect 14364 20738 14420 20748
rect 13580 20402 13636 20412
rect 15148 20188 15204 20860
rect 15596 20850 15652 20860
rect 15372 20690 15428 20702
rect 15372 20638 15374 20690
rect 15426 20638 15428 20690
rect 15372 20468 15428 20638
rect 15372 20402 15428 20412
rect 13468 20078 13470 20130
rect 13522 20078 13524 20130
rect 13468 20066 13524 20078
rect 14924 20132 15204 20188
rect 14924 20066 14980 20076
rect 12348 20020 12404 20030
rect 12348 19926 12404 19964
rect 15036 20018 15092 20132
rect 15820 20130 15876 21532
rect 15820 20078 15822 20130
rect 15874 20078 15876 20130
rect 15820 20066 15876 20078
rect 15932 21586 15988 21598
rect 15932 21534 15934 21586
rect 15986 21534 15988 21586
rect 15036 19966 15038 20018
rect 15090 19966 15092 20018
rect 15036 19954 15092 19966
rect 12908 19908 12964 19918
rect 12124 19854 12126 19906
rect 12178 19854 12180 19906
rect 12124 19842 12180 19854
rect 12460 19906 12964 19908
rect 12460 19854 12910 19906
rect 12962 19854 12964 19906
rect 12460 19852 12964 19854
rect 12124 19460 12180 19470
rect 12124 19366 12180 19404
rect 12460 19458 12516 19852
rect 12908 19842 12964 19852
rect 15148 19572 15204 19582
rect 12460 19406 12462 19458
rect 12514 19406 12516 19458
rect 12460 19394 12516 19406
rect 15036 19516 15148 19572
rect 12124 19236 12180 19246
rect 12012 19234 12180 19236
rect 12012 19182 12126 19234
rect 12178 19182 12180 19234
rect 12012 19180 12180 19182
rect 12124 19170 12180 19180
rect 14476 19234 14532 19246
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 12124 19012 12180 19022
rect 14140 19012 14196 19022
rect 10668 18386 10724 18396
rect 11788 18562 11844 18574
rect 11788 18510 11790 18562
rect 11842 18510 11844 18562
rect 8876 18338 8932 18350
rect 8876 18286 8878 18338
rect 8930 18286 8932 18338
rect 8876 18116 8932 18286
rect 10780 18228 10836 18238
rect 10780 18134 10836 18172
rect 11116 18226 11172 18238
rect 11116 18174 11118 18226
rect 11170 18174 11172 18226
rect 8876 18050 8932 18060
rect 11116 17892 11172 18174
rect 8428 17614 8430 17666
rect 8482 17614 8484 17666
rect 8428 17602 8484 17614
rect 10780 17836 11116 17892
rect 9212 17556 9268 17566
rect 9212 17554 9604 17556
rect 9212 17502 9214 17554
rect 9266 17502 9604 17554
rect 9212 17500 9604 17502
rect 9212 17490 9268 17500
rect 8092 17444 8148 17454
rect 8092 17442 8372 17444
rect 8092 17390 8094 17442
rect 8146 17390 8372 17442
rect 8092 17388 8372 17390
rect 8092 17378 8148 17388
rect 8316 16772 8372 17388
rect 9548 17106 9604 17500
rect 9548 17054 9550 17106
rect 9602 17054 9604 17106
rect 9548 17042 9604 17054
rect 9884 16882 9940 16894
rect 9884 16830 9886 16882
rect 9938 16830 9940 16882
rect 8316 16716 8708 16772
rect 8652 16210 8708 16716
rect 9884 16324 9940 16830
rect 9884 16258 9940 16268
rect 8652 16158 8654 16210
rect 8706 16158 8708 16210
rect 8652 16146 8708 16158
rect 10780 16210 10836 17836
rect 11116 17826 11172 17836
rect 11340 17778 11396 17790
rect 11340 17726 11342 17778
rect 11394 17726 11396 17778
rect 11340 17108 11396 17726
rect 11564 17108 11620 17118
rect 11340 17052 11564 17108
rect 11228 16324 11284 16334
rect 11228 16230 11284 16268
rect 11564 16322 11620 17052
rect 11564 16270 11566 16322
rect 11618 16270 11620 16322
rect 11564 16258 11620 16270
rect 11788 16324 11844 18510
rect 10780 16158 10782 16210
rect 10834 16158 10836 16210
rect 10780 16146 10836 16158
rect 6748 15426 6916 15428
rect 6748 15374 6750 15426
rect 6802 15374 6916 15426
rect 6748 15372 6916 15374
rect 7980 16098 8036 16110
rect 7980 16046 7982 16098
rect 8034 16046 8036 16098
rect 6748 15362 6804 15372
rect 7980 15204 8036 16046
rect 8876 15540 8932 15550
rect 7980 15138 8036 15148
rect 8540 15204 8596 15214
rect 8540 14532 8596 15148
rect 8876 15202 8932 15484
rect 11788 15428 11844 16268
rect 11900 18450 11956 18462
rect 11900 18398 11902 18450
rect 11954 18398 11956 18450
rect 11900 17220 11956 18398
rect 11900 15986 11956 17164
rect 12012 18452 12068 18462
rect 12012 17778 12068 18396
rect 12012 17726 12014 17778
rect 12066 17726 12068 17778
rect 12012 16770 12068 17726
rect 12012 16718 12014 16770
rect 12066 16718 12068 16770
rect 12012 16706 12068 16718
rect 11900 15934 11902 15986
rect 11954 15934 11956 15986
rect 11900 15922 11956 15934
rect 12124 15986 12180 18956
rect 13804 19010 14196 19012
rect 13804 18958 14142 19010
rect 14194 18958 14196 19010
rect 13804 18956 14196 18958
rect 12348 18452 12404 18462
rect 12348 17780 12404 18396
rect 13132 18340 13188 18350
rect 13132 18338 13524 18340
rect 13132 18286 13134 18338
rect 13186 18286 13524 18338
rect 13132 18284 13524 18286
rect 13132 18274 13188 18284
rect 12460 17780 12516 17790
rect 12348 17724 12460 17780
rect 12460 17686 12516 17724
rect 13468 17554 13524 18284
rect 13804 17666 13860 18956
rect 14140 18946 14196 18956
rect 14476 19012 14532 19182
rect 15036 19234 15092 19516
rect 15036 19182 15038 19234
rect 15090 19182 15092 19234
rect 15036 19170 15092 19182
rect 14476 18946 14532 18956
rect 14476 17892 14532 17902
rect 14476 17798 14532 17836
rect 13804 17614 13806 17666
rect 13858 17614 13860 17666
rect 13804 17602 13860 17614
rect 13468 17502 13470 17554
rect 13522 17502 13524 17554
rect 13468 17490 13524 17502
rect 14588 17444 14644 17454
rect 14588 17350 14644 17388
rect 14700 17444 14756 17454
rect 14700 17442 14868 17444
rect 14700 17390 14702 17442
rect 14754 17390 14868 17442
rect 14700 17388 14868 17390
rect 14700 17378 14756 17388
rect 13132 16884 13188 16894
rect 12908 16828 13132 16884
rect 12124 15934 12126 15986
rect 12178 15934 12180 15986
rect 11900 15428 11956 15438
rect 11788 15426 11956 15428
rect 11788 15374 11902 15426
rect 11954 15374 11956 15426
rect 11788 15372 11956 15374
rect 11900 15362 11956 15372
rect 10556 15316 10612 15326
rect 10444 15314 10612 15316
rect 10444 15262 10558 15314
rect 10610 15262 10612 15314
rect 10444 15260 10612 15262
rect 8876 15150 8878 15202
rect 8930 15150 8932 15202
rect 8876 15138 8932 15150
rect 9660 15204 9716 15242
rect 9660 15138 9716 15148
rect 10444 15204 10500 15260
rect 10556 15250 10612 15260
rect 12012 15314 12068 15326
rect 12012 15262 12014 15314
rect 12066 15262 12068 15314
rect 11340 15202 11396 15214
rect 11340 15150 11342 15202
rect 11394 15150 11396 15202
rect 11340 15148 11396 15150
rect 11900 15204 11956 15214
rect 10444 15138 10500 15148
rect 11004 15092 11060 15102
rect 6412 13806 6414 13858
rect 6466 13806 6468 13858
rect 6412 13794 6468 13806
rect 8428 14530 8596 14532
rect 8428 14478 8542 14530
rect 8594 14478 8596 14530
rect 8428 14476 8596 14478
rect 8428 13860 8484 14476
rect 8540 14466 8596 14476
rect 10556 15090 11060 15092
rect 10556 15038 11006 15090
rect 11058 15038 11060 15090
rect 10556 15036 11060 15038
rect 9212 14420 9268 14430
rect 9212 14418 9604 14420
rect 9212 14366 9214 14418
rect 9266 14366 9604 14418
rect 9212 14364 9604 14366
rect 9212 14354 9268 14364
rect 9548 13970 9604 14364
rect 9548 13918 9550 13970
rect 9602 13918 9604 13970
rect 9548 13906 9604 13918
rect 8988 13860 9044 13870
rect 8428 13858 9044 13860
rect 8428 13806 8990 13858
rect 9042 13806 9044 13858
rect 8428 13804 9044 13806
rect 5740 13746 6020 13748
rect 5740 13694 5742 13746
rect 5794 13694 6020 13746
rect 5740 13692 6020 13694
rect 5740 13682 5796 13692
rect 8428 13524 8484 13804
rect 8988 13794 9044 13804
rect 10220 13858 10276 13870
rect 10220 13806 10222 13858
rect 10274 13806 10276 13858
rect 9884 13748 9940 13758
rect 9884 13654 9940 13692
rect 8316 13468 8484 13524
rect 8540 13634 8596 13646
rect 8540 13582 8542 13634
rect 8594 13582 8596 13634
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 8316 12962 8372 13468
rect 8316 12910 8318 12962
rect 8370 12910 8372 12962
rect 8316 12898 8372 12910
rect 8540 12740 8596 13582
rect 8988 13524 9044 13534
rect 8988 13074 9044 13468
rect 10220 13524 10276 13806
rect 10556 13858 10612 15036
rect 11004 15026 11060 15036
rect 11228 15092 11396 15148
rect 11788 15092 11956 15148
rect 10556 13806 10558 13858
rect 10610 13806 10612 13858
rect 10556 13794 10612 13806
rect 11116 13748 11172 13758
rect 11116 13654 11172 13692
rect 10220 13458 10276 13468
rect 11228 13636 11284 15092
rect 11340 14642 11396 14654
rect 11788 14644 11844 15092
rect 12012 14756 12068 15262
rect 12124 15148 12180 15934
rect 12796 16772 12852 16782
rect 12796 15314 12852 16716
rect 12908 16210 12964 16828
rect 13132 16790 13188 16828
rect 14700 16324 14756 16334
rect 14700 16230 14756 16268
rect 12908 16158 12910 16210
rect 12962 16158 12964 16210
rect 12908 16146 12964 16158
rect 13804 15988 13860 15998
rect 13580 15876 13636 15886
rect 13468 15874 13636 15876
rect 13468 15822 13582 15874
rect 13634 15822 13636 15874
rect 13468 15820 13636 15822
rect 13468 15426 13524 15820
rect 13580 15810 13636 15820
rect 13468 15374 13470 15426
rect 13522 15374 13524 15426
rect 13468 15362 13524 15374
rect 12796 15262 12798 15314
rect 12850 15262 12852 15314
rect 12796 15204 12852 15262
rect 13804 15148 13860 15932
rect 13916 15988 13972 15998
rect 14364 15988 14420 15998
rect 13916 15986 14420 15988
rect 13916 15934 13918 15986
rect 13970 15934 14366 15986
rect 14418 15934 14420 15986
rect 13916 15932 14420 15934
rect 13916 15922 13972 15932
rect 14364 15922 14420 15932
rect 14812 15988 14868 17388
rect 15036 17332 15092 17342
rect 14924 16772 14980 16782
rect 14924 16678 14980 16716
rect 15036 16324 15092 17276
rect 15036 16258 15092 16268
rect 15148 16098 15204 19516
rect 15932 19348 15988 21534
rect 16380 21476 16436 21486
rect 16380 21382 16436 21420
rect 16268 21362 16324 21374
rect 16268 21310 16270 21362
rect 16322 21310 16324 21362
rect 16268 21252 16324 21310
rect 16268 21186 16324 21196
rect 16492 20804 16548 23214
rect 16604 23156 16660 24556
rect 16828 24836 16884 24846
rect 16828 23826 16884 24780
rect 17276 24052 17332 25566
rect 17388 25506 17444 26014
rect 17388 25454 17390 25506
rect 17442 25454 17444 25506
rect 17388 25442 17444 25454
rect 17836 25506 17892 26796
rect 17948 26068 18004 26078
rect 18060 26068 18116 26908
rect 22428 26964 22484 27132
rect 22876 27074 22932 27132
rect 22876 27022 22878 27074
rect 22930 27022 22932 27074
rect 22876 27010 22932 27022
rect 23324 27076 23380 28252
rect 23436 27860 23492 27870
rect 23436 27766 23492 27804
rect 24108 27860 24164 28366
rect 24444 28420 24500 28702
rect 25340 28530 25396 29484
rect 26460 29426 26516 29438
rect 26460 29374 26462 29426
rect 26514 29374 26516 29426
rect 25452 29316 25508 29326
rect 25452 29222 25508 29260
rect 25900 29316 25956 29326
rect 25900 29222 25956 29260
rect 26460 29316 26516 29374
rect 26908 29428 26964 29438
rect 26908 29334 26964 29372
rect 26460 29250 26516 29260
rect 27020 28868 27076 29934
rect 27244 29652 27300 31502
rect 27244 29586 27300 29596
rect 27468 31444 27524 31454
rect 27468 29650 27524 31388
rect 27692 31220 27748 31230
rect 27804 31220 27860 32732
rect 27916 31780 27972 31790
rect 27916 31686 27972 31724
rect 28028 31444 28084 32732
rect 28028 31378 28084 31388
rect 27692 31218 27860 31220
rect 27692 31166 27694 31218
rect 27746 31166 27860 31218
rect 27692 31164 27860 31166
rect 27692 31154 27748 31164
rect 28140 30772 28196 35084
rect 28588 34802 28644 35084
rect 28700 34916 28756 37100
rect 28924 36260 28980 37214
rect 29260 36708 29316 36718
rect 29260 36594 29316 36652
rect 29260 36542 29262 36594
rect 29314 36542 29316 36594
rect 29148 36260 29204 36270
rect 28924 36258 29204 36260
rect 28924 36206 29150 36258
rect 29202 36206 29204 36258
rect 28924 36204 29204 36206
rect 29148 36036 29204 36204
rect 29148 35970 29204 35980
rect 29260 35700 29316 36542
rect 29260 35634 29316 35644
rect 28924 35364 28980 35374
rect 28812 34916 28868 34926
rect 28700 34860 28812 34916
rect 28812 34850 28868 34860
rect 28588 34750 28590 34802
rect 28642 34750 28644 34802
rect 28588 34738 28644 34750
rect 28252 34690 28308 34702
rect 28252 34638 28254 34690
rect 28306 34638 28308 34690
rect 28252 33236 28308 34638
rect 28924 34354 28980 35308
rect 29372 35140 29428 40796
rect 30044 39060 30100 39070
rect 30044 38966 30100 39004
rect 29708 38948 29764 38958
rect 29708 38854 29764 38892
rect 30044 38052 30100 38090
rect 30044 37986 30100 37996
rect 30044 37828 30100 37838
rect 29932 37826 30100 37828
rect 29932 37774 30046 37826
rect 30098 37774 30100 37826
rect 29932 37772 30100 37774
rect 29596 36484 29652 36494
rect 29820 36484 29876 36494
rect 29596 36390 29652 36428
rect 29708 36482 29876 36484
rect 29708 36430 29822 36482
rect 29874 36430 29876 36482
rect 29708 36428 29876 36430
rect 28924 34302 28926 34354
rect 28978 34302 28980 34354
rect 28924 34290 28980 34302
rect 29036 35084 29428 35140
rect 29484 35698 29540 35710
rect 29484 35646 29486 35698
rect 29538 35646 29540 35698
rect 29484 35140 29540 35646
rect 29708 35476 29764 36428
rect 29820 36418 29876 36428
rect 29820 35700 29876 35710
rect 29820 35606 29876 35644
rect 29932 35698 29988 37772
rect 30044 37762 30100 37772
rect 30156 36594 30212 40908
rect 30492 40516 30548 40526
rect 30156 36542 30158 36594
rect 30210 36542 30212 36594
rect 30156 36530 30212 36542
rect 30268 39732 30324 39742
rect 30044 36484 30100 36494
rect 30268 36484 30324 39676
rect 30492 39732 30548 40460
rect 30492 39730 30772 39732
rect 30492 39678 30494 39730
rect 30546 39678 30772 39730
rect 30492 39676 30772 39678
rect 30492 39666 30548 39676
rect 30716 39620 30772 39676
rect 30716 39526 30772 39564
rect 30828 39396 30884 41022
rect 30828 39330 30884 39340
rect 30940 40402 30996 42812
rect 31276 42754 31332 42766
rect 31948 42756 32004 43596
rect 32844 43540 32900 44158
rect 32844 43474 32900 43484
rect 31276 42702 31278 42754
rect 31330 42702 31332 42754
rect 31052 42530 31108 42542
rect 31052 42478 31054 42530
rect 31106 42478 31108 42530
rect 31052 42196 31108 42478
rect 31276 42532 31332 42702
rect 31500 42754 32004 42756
rect 31500 42702 31950 42754
rect 32002 42702 32004 42754
rect 31500 42700 32004 42702
rect 31332 42476 31444 42532
rect 31276 42466 31332 42476
rect 31052 42140 31332 42196
rect 31276 42082 31332 42140
rect 31276 42030 31278 42082
rect 31330 42030 31332 42082
rect 31276 42018 31332 42030
rect 31164 41972 31220 41982
rect 30940 40350 30942 40402
rect 30994 40350 30996 40402
rect 30940 39060 30996 40350
rect 31052 41074 31108 41086
rect 31052 41022 31054 41074
rect 31106 41022 31108 41074
rect 31052 40404 31108 41022
rect 31164 41074 31220 41916
rect 31388 41186 31444 42476
rect 31388 41134 31390 41186
rect 31442 41134 31444 41186
rect 31388 41122 31444 41134
rect 31164 41022 31166 41074
rect 31218 41022 31220 41074
rect 31164 41010 31220 41022
rect 31052 40338 31108 40348
rect 31164 40514 31220 40526
rect 31164 40462 31166 40514
rect 31218 40462 31220 40514
rect 31164 40292 31220 40462
rect 31164 39732 31220 40236
rect 31164 39666 31220 39676
rect 31052 39396 31108 39406
rect 31052 39302 31108 39340
rect 30940 38966 30996 39004
rect 31388 38836 31444 38846
rect 31500 38836 31556 42700
rect 31948 42690 32004 42700
rect 32508 42754 32564 42766
rect 32508 42702 32510 42754
rect 32562 42702 32564 42754
rect 32508 42196 32564 42702
rect 32508 42130 32564 42140
rect 31948 41972 32004 41982
rect 32508 41972 32564 41982
rect 31948 41970 32564 41972
rect 31948 41918 31950 41970
rect 32002 41918 32510 41970
rect 32562 41918 32564 41970
rect 31948 41916 32564 41918
rect 31724 41188 31780 41198
rect 31948 41188 32004 41916
rect 32508 41906 32564 41916
rect 31780 41132 32004 41188
rect 31612 40290 31668 40302
rect 31612 40238 31614 40290
rect 31666 40238 31668 40290
rect 31612 39396 31668 40238
rect 31612 39330 31668 39340
rect 31276 38834 31556 38836
rect 31276 38782 31390 38834
rect 31442 38782 31556 38834
rect 31276 38780 31556 38782
rect 31612 39172 31668 39182
rect 30380 38722 30436 38734
rect 30380 38670 30382 38722
rect 30434 38670 30436 38722
rect 30380 38612 30436 38670
rect 30380 38546 30436 38556
rect 30940 38052 30996 38062
rect 30268 36428 30436 36484
rect 30044 36390 30100 36428
rect 30268 36260 30324 36270
rect 30268 36166 30324 36204
rect 30380 35700 30436 36428
rect 29932 35646 29934 35698
rect 29986 35646 29988 35698
rect 29932 35588 29988 35646
rect 29932 35522 29988 35532
rect 30268 35644 30436 35700
rect 30268 35476 30324 35644
rect 28476 34244 28532 34254
rect 28476 34242 28644 34244
rect 28476 34190 28478 34242
rect 28530 34190 28644 34242
rect 28476 34188 28644 34190
rect 28476 34178 28532 34188
rect 28364 34130 28420 34142
rect 28364 34078 28366 34130
rect 28418 34078 28420 34130
rect 28364 33908 28420 34078
rect 28588 34020 28644 34188
rect 28588 33954 28644 33964
rect 28364 33842 28420 33852
rect 28252 33170 28308 33180
rect 28476 33684 28532 33694
rect 28476 32674 28532 33628
rect 28476 32622 28478 32674
rect 28530 32622 28532 32674
rect 28476 32610 28532 32622
rect 28812 33572 28868 33582
rect 28588 32564 28644 32574
rect 28588 32470 28644 32508
rect 28812 32562 28868 33516
rect 28812 32510 28814 32562
rect 28866 32510 28868 32562
rect 28812 32498 28868 32510
rect 28252 32450 28308 32462
rect 28252 32398 28254 32450
rect 28306 32398 28308 32450
rect 28252 31780 28308 32398
rect 28252 31714 28308 31724
rect 29036 30884 29092 35084
rect 29484 35074 29540 35084
rect 29596 35420 29764 35476
rect 30156 35420 30324 35476
rect 30380 35474 30436 35486
rect 30380 35422 30382 35474
rect 30434 35422 30436 35474
rect 29148 34916 29204 34926
rect 29148 34822 29204 34860
rect 29372 34916 29428 34926
rect 29596 34916 29652 35420
rect 29372 34822 29428 34860
rect 29484 34860 29652 34916
rect 29708 35252 29764 35262
rect 29708 34914 29764 35196
rect 29708 34862 29710 34914
rect 29762 34862 29764 34914
rect 29372 34130 29428 34142
rect 29372 34078 29374 34130
rect 29426 34078 29428 34130
rect 29148 33236 29204 33246
rect 29148 33142 29204 33180
rect 29372 32788 29428 34078
rect 29484 33796 29540 34860
rect 29708 34850 29764 34862
rect 30156 34916 30212 35420
rect 30268 35252 30324 35262
rect 30268 35138 30324 35196
rect 30268 35086 30270 35138
rect 30322 35086 30324 35138
rect 30268 35074 30324 35086
rect 30156 34860 30324 34916
rect 29596 34690 29652 34702
rect 29596 34638 29598 34690
rect 29650 34638 29652 34690
rect 29596 34244 29652 34638
rect 30044 34468 30100 34478
rect 29932 34244 29988 34254
rect 29596 34242 29988 34244
rect 29596 34190 29934 34242
rect 29986 34190 29988 34242
rect 29596 34188 29988 34190
rect 29932 34178 29988 34188
rect 29484 33740 29876 33796
rect 29372 32722 29428 32732
rect 29484 33122 29540 33134
rect 29484 33070 29486 33122
rect 29538 33070 29540 33122
rect 29260 32564 29316 32574
rect 29260 32470 29316 32508
rect 29372 32564 29428 32574
rect 29484 32564 29540 33070
rect 29372 32562 29540 32564
rect 29372 32510 29374 32562
rect 29426 32510 29540 32562
rect 29372 32508 29540 32510
rect 29820 32786 29876 33740
rect 29820 32734 29822 32786
rect 29874 32734 29876 32786
rect 29260 31780 29316 31790
rect 29372 31780 29428 32508
rect 29820 32452 29876 32734
rect 30044 32786 30100 34412
rect 30044 32734 30046 32786
rect 30098 32734 30100 32786
rect 30044 32722 30100 32734
rect 30268 32786 30324 34860
rect 30268 32734 30270 32786
rect 30322 32734 30324 32786
rect 30268 32722 30324 32734
rect 29820 32386 29876 32396
rect 29932 32450 29988 32462
rect 29932 32398 29934 32450
rect 29986 32398 29988 32450
rect 29316 31724 29428 31780
rect 29820 32228 29876 32238
rect 29148 31668 29204 31678
rect 29148 31574 29204 31612
rect 29260 31666 29316 31724
rect 29260 31614 29262 31666
rect 29314 31614 29316 31666
rect 29260 31602 29316 31614
rect 29484 31556 29540 31566
rect 29484 31462 29540 31500
rect 29484 30996 29540 31006
rect 29484 30902 29540 30940
rect 29820 30884 29876 32172
rect 29932 32004 29988 32398
rect 29932 31948 30212 32004
rect 30044 31780 30100 31790
rect 30156 31780 30212 31948
rect 30268 31780 30324 31790
rect 30156 31778 30324 31780
rect 30156 31726 30270 31778
rect 30322 31726 30324 31778
rect 30156 31724 30324 31726
rect 30044 31686 30100 31724
rect 30268 31714 30324 31724
rect 30268 31554 30324 31566
rect 30268 31502 30270 31554
rect 30322 31502 30324 31554
rect 30156 31108 30212 31118
rect 30268 31108 30324 31502
rect 30156 31106 30324 31108
rect 30156 31054 30158 31106
rect 30210 31054 30324 31106
rect 30156 31052 30324 31054
rect 30156 31042 30212 31052
rect 29036 30828 29316 30884
rect 28140 30716 28420 30772
rect 27468 29598 27470 29650
rect 27522 29598 27524 29650
rect 27468 29586 27524 29598
rect 28364 29652 28420 30716
rect 28700 30212 28756 30222
rect 29148 30212 29204 30222
rect 28700 30210 29204 30212
rect 28700 30158 28702 30210
rect 28754 30158 29150 30210
rect 29202 30158 29204 30210
rect 28700 30156 29204 30158
rect 28700 29988 28756 30156
rect 29148 30146 29204 30156
rect 28700 29922 28756 29932
rect 28700 29652 28756 29662
rect 28364 29650 28756 29652
rect 28364 29598 28366 29650
rect 28418 29598 28702 29650
rect 28754 29598 28756 29650
rect 28364 29596 28756 29598
rect 27804 29428 27860 29438
rect 27132 29316 27188 29326
rect 27132 29314 27748 29316
rect 27132 29262 27134 29314
rect 27186 29262 27748 29314
rect 27132 29260 27748 29262
rect 27132 29250 27188 29260
rect 26908 28812 27076 28868
rect 25340 28478 25342 28530
rect 25394 28478 25396 28530
rect 25340 28466 25396 28478
rect 25676 28644 25732 28654
rect 26348 28644 26404 28654
rect 25676 28642 26404 28644
rect 25676 28590 25678 28642
rect 25730 28590 26350 28642
rect 26402 28590 26404 28642
rect 25676 28588 26404 28590
rect 24444 28354 24500 28364
rect 24780 28084 24836 28094
rect 24780 27990 24836 28028
rect 25452 28084 25508 28094
rect 25452 27990 25508 28028
rect 24108 27794 24164 27804
rect 24668 27860 24724 27870
rect 24332 27746 24388 27758
rect 24332 27694 24334 27746
rect 24386 27694 24388 27746
rect 24332 27412 24388 27694
rect 24332 27346 24388 27356
rect 23548 27076 23604 27086
rect 23324 27074 23604 27076
rect 23324 27022 23550 27074
rect 23602 27022 23604 27074
rect 23324 27020 23604 27022
rect 23548 27010 23604 27020
rect 22428 26898 22484 26908
rect 18620 26850 18676 26862
rect 18620 26798 18622 26850
rect 18674 26798 18676 26850
rect 18620 26402 18676 26798
rect 20524 26852 20580 26862
rect 20580 26796 21028 26852
rect 20524 26758 20580 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20972 26516 21028 26796
rect 22092 26516 22148 26526
rect 20972 26514 21364 26516
rect 20972 26462 20974 26514
rect 21026 26462 21364 26514
rect 20972 26460 21364 26462
rect 20972 26450 21028 26460
rect 18620 26350 18622 26402
rect 18674 26350 18676 26402
rect 18620 26338 18676 26350
rect 19180 26404 19236 26414
rect 18284 26292 18340 26302
rect 18284 26198 18340 26236
rect 18844 26292 18900 26302
rect 18732 26178 18788 26190
rect 18732 26126 18734 26178
rect 18786 26126 18788 26178
rect 17948 26066 18116 26068
rect 17948 26014 17950 26066
rect 18002 26014 18116 26066
rect 17948 26012 18116 26014
rect 17948 26002 18004 26012
rect 17836 25454 17838 25506
rect 17890 25454 17892 25506
rect 17836 25442 17892 25454
rect 17500 25396 17556 25406
rect 17500 25302 17556 25340
rect 17836 24834 17892 24846
rect 17836 24782 17838 24834
rect 17890 24782 17892 24834
rect 17612 24724 17668 24734
rect 17612 24630 17668 24668
rect 17836 24500 17892 24782
rect 17836 24434 17892 24444
rect 18060 24722 18116 26012
rect 18284 26068 18340 26078
rect 18284 25974 18340 26012
rect 18620 25620 18676 25630
rect 18732 25620 18788 26126
rect 18620 25618 18788 25620
rect 18620 25566 18622 25618
rect 18674 25566 18788 25618
rect 18620 25564 18788 25566
rect 18620 25554 18676 25564
rect 18844 25060 18900 26236
rect 19180 26290 19236 26348
rect 19852 26404 19908 26414
rect 19852 26310 19908 26348
rect 19180 26238 19182 26290
rect 19234 26238 19236 26290
rect 19180 26226 19236 26238
rect 20300 26178 20356 26190
rect 20300 26126 20302 26178
rect 20354 26126 20356 26178
rect 19068 26068 19124 26078
rect 19068 25974 19124 26012
rect 20300 25396 20356 26126
rect 20300 25330 20356 25340
rect 20748 25618 20804 25630
rect 20748 25566 20750 25618
rect 20802 25566 20804 25618
rect 18620 25004 18900 25060
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20748 25060 20804 25566
rect 21308 25506 21364 26460
rect 22092 25618 22148 26460
rect 24668 26178 24724 27804
rect 25228 27634 25284 27646
rect 25228 27582 25230 27634
rect 25282 27582 25284 27634
rect 25228 27412 25284 27582
rect 25228 27346 25284 27356
rect 25564 27634 25620 27646
rect 25564 27582 25566 27634
rect 25618 27582 25620 27634
rect 25564 26908 25620 27582
rect 25676 27186 25732 28588
rect 26348 28578 26404 28588
rect 26908 28642 26964 28812
rect 27468 28756 27524 28766
rect 27468 28662 27524 28700
rect 26908 28590 26910 28642
rect 26962 28590 26964 28642
rect 25676 27134 25678 27186
rect 25730 27134 25732 27186
rect 25676 27122 25732 27134
rect 26908 26908 26964 28590
rect 27020 28644 27076 28654
rect 27356 28644 27412 28654
rect 27020 28642 27412 28644
rect 27020 28590 27022 28642
rect 27074 28590 27358 28642
rect 27410 28590 27412 28642
rect 27020 28588 27412 28590
rect 27020 28578 27076 28588
rect 27356 28578 27412 28588
rect 27692 28642 27748 29260
rect 27692 28590 27694 28642
rect 27746 28590 27748 28642
rect 27692 28578 27748 28590
rect 27804 26908 27860 29372
rect 28364 29092 28420 29596
rect 28700 29540 28756 29596
rect 28700 29474 28756 29484
rect 29260 29428 29316 30828
rect 29820 30818 29876 30828
rect 30380 30212 30436 35422
rect 30604 35028 30660 35038
rect 30604 35026 30772 35028
rect 30604 34974 30606 35026
rect 30658 34974 30772 35026
rect 30604 34972 30772 34974
rect 30604 34962 30660 34972
rect 30492 34690 30548 34702
rect 30492 34638 30494 34690
rect 30546 34638 30548 34690
rect 30492 34132 30548 34638
rect 30604 34132 30660 34142
rect 30492 34130 30660 34132
rect 30492 34078 30606 34130
rect 30658 34078 30660 34130
rect 30492 34076 30660 34078
rect 30604 34020 30660 34076
rect 30604 33954 30660 33964
rect 30716 33796 30772 34972
rect 30828 34916 30884 34926
rect 30828 34822 30884 34860
rect 30940 34692 30996 37996
rect 31276 38050 31332 38780
rect 31388 38770 31444 38780
rect 31276 37998 31278 38050
rect 31330 37998 31332 38050
rect 31276 37492 31332 37998
rect 31612 38052 31668 39116
rect 31724 38668 31780 41132
rect 32508 41076 32564 41086
rect 32508 40982 32564 41020
rect 32060 40404 32116 40414
rect 32060 40310 32116 40348
rect 32508 40402 32564 40414
rect 32508 40350 32510 40402
rect 32562 40350 32564 40402
rect 32508 40292 32564 40350
rect 32508 40226 32564 40236
rect 31836 39172 31892 39182
rect 31836 38834 31892 39116
rect 31836 38782 31838 38834
rect 31890 38782 31892 38834
rect 31836 38770 31892 38782
rect 32284 38948 32340 38958
rect 31724 38612 32004 38668
rect 31612 37986 31668 37996
rect 31948 38050 32004 38612
rect 31948 37998 31950 38050
rect 32002 37998 32004 38050
rect 31276 37426 31332 37436
rect 31500 37938 31556 37950
rect 31500 37886 31502 37938
rect 31554 37886 31556 37938
rect 31500 37380 31556 37886
rect 31836 37492 31892 37502
rect 31500 37324 31668 37380
rect 31500 37154 31556 37166
rect 31500 37102 31502 37154
rect 31554 37102 31556 37154
rect 31388 36260 31444 36270
rect 31052 36148 31108 36158
rect 31052 35476 31108 36092
rect 31388 35922 31444 36204
rect 31388 35870 31390 35922
rect 31442 35870 31444 35922
rect 31388 35858 31444 35870
rect 31500 35924 31556 37102
rect 31500 35858 31556 35868
rect 31164 35700 31220 35710
rect 31164 35698 31332 35700
rect 31164 35646 31166 35698
rect 31218 35646 31332 35698
rect 31164 35644 31332 35646
rect 31164 35634 31220 35644
rect 31052 35420 31220 35476
rect 31164 34804 31220 35420
rect 31276 35140 31332 35644
rect 31276 34916 31332 35084
rect 31500 34916 31556 34926
rect 31276 34914 31556 34916
rect 31276 34862 31502 34914
rect 31554 34862 31556 34914
rect 31276 34860 31556 34862
rect 31500 34850 31556 34860
rect 31164 34802 31332 34804
rect 31164 34750 31166 34802
rect 31218 34750 31332 34802
rect 31164 34748 31332 34750
rect 31164 34738 31220 34748
rect 30716 33730 30772 33740
rect 30828 34636 30996 34692
rect 31052 34692 31108 34702
rect 30604 33348 30660 33358
rect 30604 33254 30660 33292
rect 30716 33122 30772 33134
rect 30716 33070 30718 33122
rect 30770 33070 30772 33122
rect 30492 32786 30548 32798
rect 30492 32734 30494 32786
rect 30546 32734 30548 32786
rect 30492 32676 30548 32734
rect 30604 32676 30660 32686
rect 30492 32674 30660 32676
rect 30492 32622 30606 32674
rect 30658 32622 30660 32674
rect 30492 32620 30660 32622
rect 30492 31780 30548 32620
rect 30604 32610 30660 32620
rect 30716 32228 30772 33070
rect 30828 32788 30884 34636
rect 31052 34598 31108 34636
rect 30940 34242 30996 34254
rect 30940 34190 30942 34242
rect 30994 34190 30996 34242
rect 30940 34132 30996 34190
rect 31276 34242 31332 34748
rect 31612 34580 31668 37324
rect 31836 37266 31892 37436
rect 31836 37214 31838 37266
rect 31890 37214 31892 37266
rect 31836 37202 31892 37214
rect 31948 37268 32004 37998
rect 31948 37044 32004 37212
rect 31724 36988 32004 37044
rect 31724 36482 31780 36988
rect 31724 36430 31726 36482
rect 31778 36430 31780 36482
rect 31724 36418 31780 36430
rect 32172 35698 32228 35710
rect 32172 35646 32174 35698
rect 32226 35646 32228 35698
rect 32172 35364 32228 35646
rect 32172 35298 32228 35308
rect 32284 35028 32340 38892
rect 32620 37938 32676 37950
rect 32620 37886 32622 37938
rect 32674 37886 32676 37938
rect 32396 36370 32452 36382
rect 32396 36318 32398 36370
rect 32450 36318 32452 36370
rect 32396 35922 32452 36318
rect 32396 35870 32398 35922
rect 32450 35870 32452 35922
rect 32396 35858 32452 35870
rect 32620 35700 32676 37886
rect 32284 34962 32340 34972
rect 32396 35644 32676 35700
rect 32732 35700 32788 35710
rect 32396 35026 32452 35644
rect 32508 35476 32564 35486
rect 32508 35382 32564 35420
rect 32396 34974 32398 35026
rect 32450 34974 32452 35026
rect 32396 34962 32452 34974
rect 32172 34914 32228 34926
rect 32172 34862 32174 34914
rect 32226 34862 32228 34914
rect 31836 34804 31892 34814
rect 31836 34710 31892 34748
rect 31276 34190 31278 34242
rect 31330 34190 31332 34242
rect 31276 34178 31332 34190
rect 31388 34524 31668 34580
rect 30940 34066 30996 34076
rect 30940 33908 30996 33918
rect 30940 33346 30996 33852
rect 30940 33294 30942 33346
rect 30994 33294 30996 33346
rect 30940 33282 30996 33294
rect 30828 32732 30996 32788
rect 30828 32564 30884 32574
rect 30828 32470 30884 32508
rect 30716 32162 30772 32172
rect 30492 31714 30548 31724
rect 30604 32004 30660 32014
rect 30940 32004 30996 32732
rect 31164 32562 31220 32574
rect 31164 32510 31166 32562
rect 31218 32510 31220 32562
rect 31164 32228 31220 32510
rect 31388 32340 31444 34524
rect 31724 34244 31780 34254
rect 31724 34150 31780 34188
rect 31500 34130 31556 34142
rect 31500 34078 31502 34130
rect 31554 34078 31556 34130
rect 31500 33796 31556 34078
rect 31948 34132 32004 34142
rect 32004 34076 32116 34132
rect 31948 34038 32004 34076
rect 31500 33730 31556 33740
rect 31612 34018 31668 34030
rect 31612 33966 31614 34018
rect 31666 33966 31668 34018
rect 31612 33572 31668 33966
rect 31948 33572 32004 33582
rect 31612 33570 32004 33572
rect 31612 33518 31950 33570
rect 32002 33518 32004 33570
rect 31612 33516 32004 33518
rect 31948 33506 32004 33516
rect 32060 33348 32116 34076
rect 32172 33908 32228 34862
rect 32620 34804 32676 34814
rect 32620 34710 32676 34748
rect 32172 33842 32228 33852
rect 32732 33684 32788 35644
rect 32844 35588 32900 35598
rect 32844 34914 32900 35532
rect 32844 34862 32846 34914
rect 32898 34862 32900 34914
rect 32844 34850 32900 34862
rect 31948 33292 32116 33348
rect 32172 33628 32788 33684
rect 31836 32564 31892 32574
rect 31836 32470 31892 32508
rect 31612 32452 31668 32462
rect 31612 32358 31668 32396
rect 31724 32450 31780 32462
rect 31724 32398 31726 32450
rect 31778 32398 31780 32450
rect 31388 32246 31444 32284
rect 31164 32162 31220 32172
rect 30604 31778 30660 31948
rect 30604 31726 30606 31778
rect 30658 31726 30660 31778
rect 30604 31714 30660 31726
rect 30828 31948 30996 32004
rect 30380 30146 30436 30156
rect 29596 29540 29652 29550
rect 29596 29446 29652 29484
rect 29932 29538 29988 29550
rect 29932 29486 29934 29538
rect 29986 29486 29988 29538
rect 29260 29426 29540 29428
rect 29260 29374 29262 29426
rect 29314 29374 29540 29426
rect 29260 29372 29540 29374
rect 29260 29362 29316 29372
rect 28364 28754 28420 29036
rect 28364 28702 28366 28754
rect 28418 28702 28420 28754
rect 28364 28690 28420 28702
rect 29260 28642 29316 28654
rect 29260 28590 29262 28642
rect 29314 28590 29316 28642
rect 29260 27076 29316 28590
rect 29484 28084 29540 29372
rect 29932 28756 29988 29486
rect 30828 29204 30884 31948
rect 31612 31892 31668 31902
rect 31724 31892 31780 32398
rect 31948 32452 32004 33292
rect 32060 33122 32116 33134
rect 32060 33070 32062 33122
rect 32114 33070 32116 33122
rect 32060 32788 32116 33070
rect 32172 32788 32228 33628
rect 32508 33460 32564 33470
rect 32956 33460 33012 47180
rect 33516 47458 33572 47470
rect 33516 47406 33518 47458
rect 33570 47406 33572 47458
rect 33516 46900 33572 47406
rect 34188 47346 34244 47358
rect 34188 47294 34190 47346
rect 34242 47294 34244 47346
rect 34188 47012 34244 47294
rect 34188 46946 34244 46956
rect 33180 46844 33516 46900
rect 33180 45892 33236 46844
rect 33516 46834 33572 46844
rect 34748 46004 34804 46014
rect 34748 45910 34804 45948
rect 33180 45330 33236 45836
rect 34636 45332 34692 45342
rect 33180 45278 33182 45330
rect 33234 45278 33236 45330
rect 33180 45266 33236 45278
rect 34300 45330 34692 45332
rect 34300 45278 34638 45330
rect 34690 45278 34692 45330
rect 34300 45276 34692 45278
rect 33292 44324 33348 44334
rect 33292 44230 33348 44268
rect 33964 44324 34020 44334
rect 34300 44324 34356 45276
rect 34636 45266 34692 45276
rect 34860 45220 34916 45230
rect 34748 45218 34916 45220
rect 34748 45166 34862 45218
rect 34914 45166 34916 45218
rect 34748 45164 34916 45166
rect 34412 45106 34468 45118
rect 34412 45054 34414 45106
rect 34466 45054 34468 45106
rect 34412 44772 34468 45054
rect 34524 45108 34580 45118
rect 34524 45014 34580 45052
rect 34412 44716 34692 44772
rect 33516 44100 33572 44110
rect 33516 44006 33572 44044
rect 33964 43650 34020 44268
rect 33964 43598 33966 43650
rect 34018 43598 34020 43650
rect 33964 43586 34020 43598
rect 34188 44322 34356 44324
rect 34188 44270 34302 44322
rect 34354 44270 34356 44322
rect 34188 44268 34356 44270
rect 34188 44212 34244 44268
rect 34300 44258 34356 44268
rect 33628 43540 33684 43550
rect 33628 43446 33684 43484
rect 33404 43426 33460 43438
rect 33404 43374 33406 43426
rect 33458 43374 33460 43426
rect 33404 42868 33460 43374
rect 33740 42868 33796 42878
rect 33404 42812 33740 42868
rect 33740 42774 33796 42812
rect 33740 41748 33796 41758
rect 33516 41076 33572 41086
rect 33404 40964 33460 40974
rect 33068 40402 33124 40414
rect 33068 40350 33070 40402
rect 33122 40350 33124 40402
rect 33068 40292 33124 40350
rect 33404 40402 33460 40908
rect 33516 40626 33572 41020
rect 33516 40574 33518 40626
rect 33570 40574 33572 40626
rect 33516 40562 33572 40574
rect 33404 40350 33406 40402
rect 33458 40350 33460 40402
rect 33404 40338 33460 40350
rect 33516 40404 33572 40414
rect 33068 40226 33124 40236
rect 33516 37380 33572 40348
rect 33740 40402 33796 41692
rect 33740 40350 33742 40402
rect 33794 40350 33796 40402
rect 33740 40338 33796 40350
rect 33516 37314 33572 37324
rect 33964 39620 34020 39630
rect 33628 36260 33684 36270
rect 33628 35922 33684 36204
rect 33628 35870 33630 35922
rect 33682 35870 33684 35922
rect 33628 35858 33684 35870
rect 33852 35812 33908 35822
rect 33852 35718 33908 35756
rect 33740 35588 33796 35598
rect 33740 35494 33796 35532
rect 33964 35028 34020 39564
rect 34076 36596 34132 36606
rect 34076 35922 34132 36540
rect 34188 36484 34244 44156
rect 34636 44210 34692 44716
rect 34636 44158 34638 44210
rect 34690 44158 34692 44210
rect 34636 44100 34692 44158
rect 34636 44034 34692 44044
rect 34748 43652 34804 45164
rect 34860 45154 34916 45164
rect 35084 44884 35140 51324
rect 35868 51380 35924 51390
rect 35868 51286 35924 51324
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 36316 50484 36372 51436
rect 36428 50706 36484 53004
rect 37100 51716 37156 51726
rect 37100 51490 37156 51660
rect 37100 51438 37102 51490
rect 37154 51438 37156 51490
rect 37100 51426 37156 51438
rect 36428 50654 36430 50706
rect 36482 50654 36484 50706
rect 36428 50642 36484 50654
rect 36540 51378 36596 51390
rect 36540 51326 36542 51378
rect 36594 51326 36596 51378
rect 36540 51156 36596 51326
rect 36540 50484 36596 51100
rect 36316 49588 36372 50428
rect 36428 50428 36596 50484
rect 36428 49700 36484 50428
rect 36540 49924 36596 49934
rect 36540 49922 36932 49924
rect 36540 49870 36542 49922
rect 36594 49870 36932 49922
rect 36540 49868 36932 49870
rect 36540 49858 36596 49868
rect 36652 49700 36708 49710
rect 36428 49644 36596 49700
rect 36316 49494 36372 49532
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 36540 49026 36596 49644
rect 36652 49606 36708 49644
rect 36540 48974 36542 49026
rect 36594 48974 36596 49026
rect 36540 48962 36596 48974
rect 36764 49588 36820 49598
rect 36204 48916 36260 48926
rect 35980 48914 36260 48916
rect 35980 48862 36206 48914
rect 36258 48862 36260 48914
rect 35980 48860 36260 48862
rect 35868 48802 35924 48814
rect 35868 48750 35870 48802
rect 35922 48750 35924 48802
rect 35644 48132 35700 48142
rect 35868 48132 35924 48750
rect 35700 48076 35924 48132
rect 35644 48038 35700 48076
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35532 46900 35588 46910
rect 35532 46562 35588 46844
rect 35532 46510 35534 46562
rect 35586 46510 35588 46562
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 46060 35364 46116
rect 35196 46002 35252 46060
rect 35196 45950 35198 46002
rect 35250 45950 35252 46002
rect 35196 45938 35252 45950
rect 35308 46004 35364 46060
rect 35532 46004 35588 46510
rect 35868 46676 35924 46686
rect 35980 46676 36036 48860
rect 36204 48850 36260 48860
rect 36316 48916 36372 48926
rect 36204 48130 36260 48142
rect 36204 48078 36206 48130
rect 36258 48078 36260 48130
rect 36204 46900 36260 48078
rect 36316 47572 36372 48860
rect 36316 47570 36484 47572
rect 36316 47518 36318 47570
rect 36370 47518 36484 47570
rect 36316 47516 36484 47518
rect 36316 47506 36372 47516
rect 36204 46834 36260 46844
rect 36428 46900 36484 47516
rect 36764 47460 36820 49532
rect 36764 47394 36820 47404
rect 36428 46834 36484 46844
rect 36764 46786 36820 46798
rect 36764 46734 36766 46786
rect 36818 46734 36820 46786
rect 36204 46676 36260 46686
rect 35868 46674 36036 46676
rect 35868 46622 35870 46674
rect 35922 46622 36036 46674
rect 35868 46620 36036 46622
rect 36092 46620 36204 46676
rect 35868 46004 35924 46620
rect 35980 46452 36036 46462
rect 36092 46452 36148 46620
rect 36204 46610 36260 46620
rect 36316 46676 36372 46686
rect 36764 46676 36820 46734
rect 36316 46674 36820 46676
rect 36316 46622 36318 46674
rect 36370 46622 36820 46674
rect 36316 46620 36820 46622
rect 36316 46610 36372 46620
rect 35980 46450 36148 46452
rect 35980 46398 35982 46450
rect 36034 46398 36148 46450
rect 35980 46396 36148 46398
rect 36428 46450 36484 46462
rect 36428 46398 36430 46450
rect 36482 46398 36484 46450
rect 35980 46386 36036 46396
rect 36428 46340 36484 46398
rect 36428 46274 36484 46284
rect 36764 46228 36820 46620
rect 36876 46676 36932 49868
rect 37212 49138 37268 54460
rect 37436 53956 37492 56140
rect 37436 53890 37492 53900
rect 37548 56082 37604 56094
rect 37548 56030 37550 56082
rect 37602 56030 37604 56082
rect 37548 53060 37604 56030
rect 37660 54740 37716 59200
rect 37996 57092 38052 57102
rect 37996 55970 38052 57036
rect 38108 56980 38164 59200
rect 38108 56914 38164 56924
rect 37996 55918 37998 55970
rect 38050 55918 38052 55970
rect 37996 55906 38052 55918
rect 38556 56084 38612 56094
rect 37660 54674 37716 54684
rect 37772 55186 37828 55198
rect 37772 55134 37774 55186
rect 37826 55134 37828 55186
rect 37772 53844 37828 55134
rect 38556 54402 38612 56028
rect 38892 54740 38948 54750
rect 39004 54740 39060 59200
rect 39116 56308 39172 56318
rect 39116 56214 39172 56252
rect 39452 55412 39508 59200
rect 39900 56308 39956 59200
rect 39900 56242 39956 56252
rect 39788 56084 39844 56094
rect 39788 55990 39844 56028
rect 40348 55972 40404 59200
rect 40572 56980 40628 56990
rect 40572 56306 40628 56924
rect 40572 56254 40574 56306
rect 40626 56254 40628 56306
rect 40572 56242 40628 56254
rect 40796 56084 40852 59200
rect 41132 56308 41188 56318
rect 41132 56214 41188 56252
rect 41244 56084 41300 59200
rect 41692 56420 41748 59200
rect 42140 57092 42196 59200
rect 42140 57036 42644 57092
rect 41692 56364 42308 56420
rect 41580 56308 41636 56318
rect 41636 56252 41748 56308
rect 41580 56242 41636 56252
rect 41356 56196 41412 56206
rect 41356 56102 41412 56140
rect 41692 56194 41748 56252
rect 41692 56142 41694 56194
rect 41746 56142 41748 56194
rect 41692 56130 41748 56142
rect 40796 56028 41188 56084
rect 40348 55906 40404 55916
rect 39452 55346 39508 55356
rect 39900 55412 39956 55422
rect 40684 55412 40740 55422
rect 39900 55410 40292 55412
rect 39900 55358 39902 55410
rect 39954 55358 40292 55410
rect 39900 55356 40292 55358
rect 39900 55346 39956 55356
rect 40236 55298 40292 55356
rect 40684 55318 40740 55356
rect 40236 55246 40238 55298
rect 40290 55246 40292 55298
rect 40236 55234 40292 55246
rect 41132 55300 41188 56028
rect 41244 56018 41300 56028
rect 41580 56084 41636 56094
rect 41580 55410 41636 56028
rect 42028 56084 42084 56094
rect 42028 55990 42084 56028
rect 42252 55522 42308 56364
rect 42252 55470 42254 55522
rect 42306 55470 42308 55522
rect 42252 55458 42308 55470
rect 42364 56194 42420 56206
rect 42364 56142 42366 56194
rect 42418 56142 42420 56194
rect 41580 55358 41582 55410
rect 41634 55358 41636 55410
rect 41580 55346 41636 55358
rect 41132 55244 41524 55300
rect 41468 55188 41524 55244
rect 41804 55188 41860 55198
rect 41468 55186 41860 55188
rect 41468 55134 41806 55186
rect 41858 55134 41860 55186
rect 41468 55132 41860 55134
rect 41804 55122 41860 55132
rect 39340 54740 39396 54750
rect 39004 54738 39396 54740
rect 39004 54686 39342 54738
rect 39394 54686 39396 54738
rect 39004 54684 39396 54686
rect 38892 54646 38948 54684
rect 39340 54674 39396 54684
rect 38556 54350 38558 54402
rect 38610 54350 38612 54402
rect 38556 54338 38612 54350
rect 38780 54516 38836 54526
rect 37772 53778 37828 53788
rect 38780 53730 38836 54460
rect 40908 54516 40964 54526
rect 40908 54422 40964 54460
rect 41692 54404 41748 54414
rect 38780 53678 38782 53730
rect 38834 53678 38836 53730
rect 38780 53666 38836 53678
rect 41468 54402 41748 54404
rect 41468 54350 41694 54402
rect 41746 54350 41748 54402
rect 41468 54348 41748 54350
rect 39564 53620 39620 53630
rect 39564 53618 39956 53620
rect 39564 53566 39566 53618
rect 39618 53566 39956 53618
rect 39564 53564 39956 53566
rect 39564 53554 39620 53564
rect 37548 52994 37604 53004
rect 39004 52946 39060 52958
rect 39004 52894 39006 52946
rect 39058 52894 39060 52946
rect 38892 52276 38948 52286
rect 37884 52164 37940 52174
rect 37436 51380 37492 51390
rect 37436 51286 37492 51324
rect 37884 51378 37940 52108
rect 38892 52162 38948 52220
rect 38892 52110 38894 52162
rect 38946 52110 38948 52162
rect 38892 52098 38948 52110
rect 39004 52274 39060 52894
rect 39452 52836 39508 52846
rect 39452 52742 39508 52780
rect 39004 52222 39006 52274
rect 39058 52222 39060 52274
rect 38108 51828 38164 51838
rect 37884 51326 37886 51378
rect 37938 51326 37940 51378
rect 37884 51314 37940 51326
rect 37996 51772 38108 51828
rect 37660 51156 37716 51166
rect 37660 51062 37716 51100
rect 37996 50706 38052 51772
rect 38108 51762 38164 51772
rect 38668 51716 38724 51726
rect 38108 51492 38164 51502
rect 38108 51378 38164 51436
rect 38108 51326 38110 51378
rect 38162 51326 38164 51378
rect 38108 51314 38164 51326
rect 38556 51156 38612 51166
rect 38556 51062 38612 51100
rect 38668 50818 38724 51660
rect 38668 50766 38670 50818
rect 38722 50766 38724 50818
rect 38668 50754 38724 50766
rect 39004 50818 39060 52222
rect 39452 52052 39508 52062
rect 39676 52052 39732 52062
rect 39452 52050 39676 52052
rect 39452 51998 39454 52050
rect 39506 51998 39676 52050
rect 39452 51996 39676 51998
rect 39452 51986 39508 51996
rect 39676 51986 39732 51996
rect 39788 51938 39844 51950
rect 39788 51886 39790 51938
rect 39842 51886 39844 51938
rect 39004 50766 39006 50818
rect 39058 50766 39060 50818
rect 39004 50754 39060 50766
rect 39116 51828 39172 51838
rect 37996 50654 37998 50706
rect 38050 50654 38052 50706
rect 37996 50642 38052 50654
rect 37548 50484 37604 50494
rect 37548 50390 37604 50428
rect 38444 50484 38500 50494
rect 38444 50390 38500 50428
rect 37884 50260 37940 50270
rect 37212 49086 37214 49138
rect 37266 49086 37268 49138
rect 37212 49074 37268 49086
rect 37324 49922 37380 49934
rect 37324 49870 37326 49922
rect 37378 49870 37380 49922
rect 37324 48916 37380 49870
rect 37884 49810 37940 50204
rect 39116 49924 39172 51772
rect 39676 51492 39732 51502
rect 39788 51492 39844 51886
rect 39900 51602 39956 53564
rect 41468 53170 41524 54348
rect 41692 54338 41748 54348
rect 42364 54068 42420 56142
rect 42588 55188 42644 57036
rect 43036 56642 43092 59200
rect 43484 56980 43540 59200
rect 43484 56924 44100 56980
rect 43036 56590 43038 56642
rect 43090 56590 43092 56642
rect 43036 56578 43092 56590
rect 43596 56642 43652 56654
rect 43596 56590 43598 56642
rect 43650 56590 43652 56642
rect 42700 55972 42756 55982
rect 42700 55878 42756 55916
rect 43596 55970 43652 56590
rect 44044 56306 44100 56924
rect 44044 56254 44046 56306
rect 44098 56254 44100 56306
rect 44044 56242 44100 56254
rect 43596 55918 43598 55970
rect 43650 55918 43652 55970
rect 43596 55906 43652 55918
rect 44380 55972 44436 59200
rect 44828 56308 44884 59200
rect 45052 56308 45108 56318
rect 44828 56306 45108 56308
rect 44828 56254 45054 56306
rect 45106 56254 45108 56306
rect 44828 56252 45108 56254
rect 45052 56242 45108 56252
rect 44604 55972 44660 55982
rect 44380 55970 44660 55972
rect 44380 55918 44606 55970
rect 44658 55918 44660 55970
rect 44380 55916 44660 55918
rect 45724 55972 45780 59200
rect 46172 56308 46228 59200
rect 46396 56308 46452 56318
rect 46172 56306 46452 56308
rect 46172 56254 46398 56306
rect 46450 56254 46452 56306
rect 46172 56252 46452 56254
rect 46396 56242 46452 56252
rect 45948 55972 46004 55982
rect 45724 55970 46004 55972
rect 45724 55918 45950 55970
rect 46002 55918 46004 55970
rect 45724 55916 46004 55918
rect 47068 55972 47124 59200
rect 47516 57764 47572 59200
rect 47516 57708 47908 57764
rect 47852 56306 47908 57708
rect 47852 56254 47854 56306
rect 47906 56254 47908 56306
rect 47852 56242 47908 56254
rect 47404 55972 47460 55982
rect 47068 55970 47460 55972
rect 47068 55918 47406 55970
rect 47458 55918 47460 55970
rect 47068 55916 47460 55918
rect 48412 55972 48468 59200
rect 48860 56308 48916 59200
rect 49084 56308 49140 56318
rect 48860 56306 49140 56308
rect 48860 56254 49086 56306
rect 49138 56254 49140 56306
rect 48860 56252 49140 56254
rect 49084 56242 49140 56252
rect 48636 55972 48692 55982
rect 48412 55970 48692 55972
rect 48412 55918 48638 55970
rect 48690 55918 48692 55970
rect 48412 55916 48692 55918
rect 49756 55972 49812 59200
rect 50204 56308 50260 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 50428 56308 50484 56318
rect 50204 56306 50484 56308
rect 50204 56254 50430 56306
rect 50482 56254 50484 56306
rect 50204 56252 50484 56254
rect 50428 56242 50484 56252
rect 49980 55972 50036 55982
rect 49756 55970 50036 55972
rect 49756 55918 49982 55970
rect 50034 55918 50036 55970
rect 49756 55916 50036 55918
rect 51100 55972 51156 59200
rect 51548 56308 51604 59200
rect 51772 56308 51828 56318
rect 51548 56306 51828 56308
rect 51548 56254 51774 56306
rect 51826 56254 51828 56306
rect 51548 56252 51828 56254
rect 51772 56242 51828 56252
rect 51324 55972 51380 55982
rect 51100 55970 51380 55972
rect 51100 55918 51326 55970
rect 51378 55918 51380 55970
rect 51100 55916 51380 55918
rect 52444 55972 52500 59200
rect 52892 56308 52948 59200
rect 53116 56308 53172 56318
rect 52892 56306 53172 56308
rect 52892 56254 53118 56306
rect 53170 56254 53172 56306
rect 52892 56252 53172 56254
rect 53116 56242 53172 56252
rect 52668 55972 52724 55982
rect 52444 55970 52724 55972
rect 52444 55918 52670 55970
rect 52722 55918 52724 55970
rect 52444 55916 52724 55918
rect 53788 55972 53844 59200
rect 54236 56866 54292 59200
rect 54236 56814 54238 56866
rect 54290 56814 54292 56866
rect 54236 56802 54292 56814
rect 55020 56866 55076 56878
rect 55020 56814 55022 56866
rect 55074 56814 55076 56866
rect 55020 56306 55076 56814
rect 55020 56254 55022 56306
rect 55074 56254 55076 56306
rect 55020 56242 55076 56254
rect 54012 55972 54068 55982
rect 53788 55970 54068 55972
rect 53788 55918 54014 55970
rect 54066 55918 54068 55970
rect 53788 55916 54068 55918
rect 55132 55972 55188 59200
rect 55580 57764 55636 59200
rect 55580 57708 55972 57764
rect 55916 56306 55972 57708
rect 55916 56254 55918 56306
rect 55970 56254 55972 56306
rect 55916 56242 55972 56254
rect 55468 55972 55524 55982
rect 55132 55970 55524 55972
rect 55132 55918 55470 55970
rect 55522 55918 55524 55970
rect 55132 55916 55524 55918
rect 44604 55906 44660 55916
rect 45948 55906 46004 55916
rect 47404 55906 47460 55916
rect 48636 55906 48692 55916
rect 49980 55906 50036 55916
rect 51324 55906 51380 55916
rect 52668 55906 52724 55916
rect 54012 55906 54068 55916
rect 55468 55906 55524 55916
rect 42700 55188 42756 55198
rect 42588 55186 42756 55188
rect 42588 55134 42702 55186
rect 42754 55134 42756 55186
rect 42588 55132 42756 55134
rect 42700 55122 42756 55132
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 47068 54514 47124 54526
rect 47068 54462 47070 54514
rect 47122 54462 47124 54514
rect 43820 54402 43876 54414
rect 43820 54350 43822 54402
rect 43874 54350 43876 54402
rect 42364 54012 42756 54068
rect 41468 53118 41470 53170
rect 41522 53118 41524 53170
rect 41468 53106 41524 53118
rect 41580 53844 41636 53854
rect 41356 53058 41412 53070
rect 41356 53006 41358 53058
rect 41410 53006 41412 53058
rect 40796 52948 40852 52958
rect 40460 52834 40516 52846
rect 40460 52782 40462 52834
rect 40514 52782 40516 52834
rect 40460 52276 40516 52782
rect 40236 52220 40516 52276
rect 40796 52276 40852 52892
rect 41356 52388 41412 53006
rect 41580 53058 41636 53788
rect 41580 53006 41582 53058
rect 41634 53006 41636 53058
rect 41580 52994 41636 53006
rect 41692 53842 41748 53854
rect 41692 53790 41694 53842
rect 41746 53790 41748 53842
rect 41692 52948 41748 53790
rect 42476 53844 42532 53854
rect 42476 53750 42532 53788
rect 42364 53732 42420 53742
rect 42364 53638 42420 53676
rect 42588 53508 42644 53518
rect 42588 53172 42644 53452
rect 42700 53284 42756 54012
rect 43036 53730 43092 53742
rect 43036 53678 43038 53730
rect 43090 53678 43092 53730
rect 43036 53620 43092 53678
rect 43036 53554 43092 53564
rect 43484 53732 43540 53742
rect 42700 53228 42868 53284
rect 42028 53116 42644 53172
rect 42028 53060 42084 53116
rect 41692 52882 41748 52892
rect 41916 53058 42084 53060
rect 41916 53006 42030 53058
rect 42082 53006 42084 53058
rect 41916 53004 42084 53006
rect 41356 52332 41524 52388
rect 39900 51550 39902 51602
rect 39954 51550 39956 51602
rect 39900 51538 39956 51550
rect 40124 52162 40180 52174
rect 40124 52110 40126 52162
rect 40178 52110 40180 52162
rect 40124 51604 40180 52110
rect 40124 51538 40180 51548
rect 39676 51490 39844 51492
rect 39676 51438 39678 51490
rect 39730 51438 39844 51490
rect 39676 51436 39844 51438
rect 39676 51426 39732 51436
rect 39452 51378 39508 51390
rect 40124 51380 40180 51390
rect 40236 51380 40292 52220
rect 40796 52182 40852 52220
rect 40908 52164 40964 52174
rect 41356 52164 41412 52174
rect 40908 52162 41412 52164
rect 40908 52110 40910 52162
rect 40962 52110 41358 52162
rect 41410 52110 41412 52162
rect 40908 52108 41412 52110
rect 40348 52052 40404 52062
rect 40348 51958 40404 51996
rect 40908 51828 40964 52108
rect 41356 52098 41412 52108
rect 40348 51772 40964 51828
rect 41020 51940 41076 51950
rect 40348 51490 40404 51772
rect 40348 51438 40350 51490
rect 40402 51438 40404 51490
rect 40348 51426 40404 51438
rect 40908 51604 40964 51614
rect 40908 51490 40964 51548
rect 40908 51438 40910 51490
rect 40962 51438 40964 51490
rect 39452 51326 39454 51378
rect 39506 51326 39508 51378
rect 39228 51268 39284 51278
rect 39452 51268 39508 51326
rect 39788 51324 40068 51380
rect 39788 51268 39844 51324
rect 39228 51266 39396 51268
rect 39228 51214 39230 51266
rect 39282 51214 39396 51266
rect 39228 51212 39396 51214
rect 39452 51212 39844 51268
rect 39228 51202 39284 51212
rect 39340 51156 39396 51212
rect 39900 51156 39956 51166
rect 39340 51154 39956 51156
rect 39340 51102 39902 51154
rect 39954 51102 39956 51154
rect 39340 51100 39956 51102
rect 39116 49868 39396 49924
rect 37884 49758 37886 49810
rect 37938 49758 37940 49810
rect 37884 49746 37940 49758
rect 38668 49812 38724 49822
rect 38668 49718 38724 49756
rect 39228 49698 39284 49710
rect 39228 49646 39230 49698
rect 39282 49646 39284 49698
rect 39004 49028 39060 49038
rect 37324 48850 37380 48860
rect 38892 49026 39060 49028
rect 38892 48974 39006 49026
rect 39058 48974 39060 49026
rect 38892 48972 39060 48974
rect 37996 48242 38052 48254
rect 37996 48190 37998 48242
rect 38050 48190 38052 48242
rect 37996 48132 38052 48190
rect 37996 48066 38052 48076
rect 38556 48244 38612 48254
rect 38556 47572 38612 48188
rect 38892 48020 38948 48972
rect 39004 48962 39060 48972
rect 39228 48354 39284 49646
rect 39228 48302 39230 48354
rect 39282 48302 39284 48354
rect 38892 47954 38948 47964
rect 39004 48242 39060 48254
rect 39004 48190 39006 48242
rect 39058 48190 39060 48242
rect 39004 47684 39060 48190
rect 39116 48244 39172 48254
rect 39116 48150 39172 48188
rect 38444 47570 38612 47572
rect 38444 47518 38558 47570
rect 38610 47518 38612 47570
rect 38444 47516 38612 47518
rect 37100 47460 37156 47470
rect 37100 47366 37156 47404
rect 37436 47458 37492 47470
rect 37436 47406 37438 47458
rect 37490 47406 37492 47458
rect 37100 46900 37156 46910
rect 37100 46806 37156 46844
rect 36876 46610 36932 46620
rect 36764 46162 36820 46172
rect 37212 46452 37268 46462
rect 35308 45948 35812 46004
rect 35308 45108 35364 45118
rect 35308 45014 35364 45052
rect 34972 44828 35140 44884
rect 35420 44884 35476 44894
rect 35420 44882 35700 44884
rect 35420 44830 35422 44882
rect 35474 44830 35700 44882
rect 35420 44828 35700 44830
rect 34860 44324 34916 44334
rect 34972 44324 35028 44828
rect 35420 44818 35476 44828
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34860 44322 35028 44324
rect 34860 44270 34862 44322
rect 34914 44270 35028 44322
rect 34860 44268 35028 44270
rect 35196 44322 35252 44334
rect 35196 44270 35198 44322
rect 35250 44270 35252 44322
rect 34860 44258 34916 44268
rect 35196 43988 35252 44270
rect 35308 44212 35364 44222
rect 35308 44118 35364 44156
rect 35644 44212 35700 44828
rect 35644 44146 35700 44156
rect 35196 43932 35364 43988
rect 35308 43652 35364 43932
rect 35644 43652 35700 43662
rect 35308 43596 35476 43652
rect 34412 43540 34468 43550
rect 34412 43446 34468 43484
rect 34636 42980 34692 42990
rect 34636 42868 34692 42924
rect 34524 42866 34692 42868
rect 34524 42814 34638 42866
rect 34690 42814 34692 42866
rect 34524 42812 34692 42814
rect 34300 42754 34356 42766
rect 34300 42702 34302 42754
rect 34354 42702 34356 42754
rect 34300 41858 34356 42702
rect 34300 41806 34302 41858
rect 34354 41806 34356 41858
rect 34300 41076 34356 41806
rect 34524 41970 34580 42812
rect 34636 42802 34692 42812
rect 34524 41918 34526 41970
rect 34578 41918 34580 41970
rect 34524 41300 34580 41918
rect 34748 41972 34804 43596
rect 34860 43540 34916 43550
rect 34860 43446 34916 43484
rect 35308 43428 35364 43438
rect 35308 43334 35364 43372
rect 35420 43316 35476 43596
rect 35644 43558 35700 43596
rect 35420 43250 35476 43260
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34860 41972 34916 41982
rect 34748 41970 34916 41972
rect 34748 41918 34862 41970
rect 34914 41918 34916 41970
rect 34748 41916 34916 41918
rect 34860 41906 34916 41916
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 34636 41300 34692 41310
rect 34524 41298 35140 41300
rect 34524 41246 34638 41298
rect 34690 41246 35140 41298
rect 34524 41244 35140 41246
rect 34636 41234 34692 41244
rect 34300 41020 34580 41076
rect 34412 40290 34468 40302
rect 34412 40238 34414 40290
rect 34466 40238 34468 40290
rect 34300 40068 34356 40078
rect 34300 39732 34356 40012
rect 34300 39060 34356 39676
rect 34412 39620 34468 40238
rect 34412 39554 34468 39564
rect 34300 38966 34356 39004
rect 34188 36418 34244 36428
rect 34412 37828 34468 37838
rect 34188 36260 34244 36270
rect 34244 36204 34356 36260
rect 34188 36194 34244 36204
rect 34076 35870 34078 35922
rect 34130 35870 34132 35922
rect 34076 35588 34132 35870
rect 34076 35522 34132 35532
rect 33964 34962 34020 34972
rect 32284 33348 32340 33358
rect 32284 33346 32452 33348
rect 32284 33294 32286 33346
rect 32338 33294 32452 33346
rect 32284 33292 32452 33294
rect 32284 33282 32340 33292
rect 32284 32788 32340 32798
rect 32172 32786 32340 32788
rect 32172 32734 32286 32786
rect 32338 32734 32340 32786
rect 32172 32732 32340 32734
rect 32396 32788 32452 33292
rect 32508 33346 32564 33404
rect 32508 33294 32510 33346
rect 32562 33294 32564 33346
rect 32508 33282 32564 33294
rect 32844 33404 33012 33460
rect 33068 34804 33124 34814
rect 32732 33236 32788 33246
rect 32732 33142 32788 33180
rect 32396 32732 32676 32788
rect 32060 32722 32116 32732
rect 31948 32386 32004 32396
rect 32060 32562 32116 32574
rect 32060 32510 32062 32562
rect 32114 32510 32116 32562
rect 32060 32004 32116 32510
rect 32060 31938 32116 31948
rect 31612 31890 31780 31892
rect 31612 31838 31614 31890
rect 31666 31838 31780 31890
rect 31612 31836 31780 31838
rect 31612 31826 31668 31836
rect 30940 31778 30996 31790
rect 30940 31726 30942 31778
rect 30994 31726 30996 31778
rect 30940 30996 30996 31726
rect 30940 30324 30996 30940
rect 32284 30882 32340 32732
rect 32396 32562 32452 32574
rect 32396 32510 32398 32562
rect 32450 32510 32452 32562
rect 32396 32452 32452 32510
rect 32396 31108 32452 32396
rect 32396 31042 32452 31052
rect 32284 30830 32286 30882
rect 32338 30830 32340 30882
rect 32284 30818 32340 30830
rect 30940 30258 30996 30268
rect 32620 29876 32676 32732
rect 32844 30100 32900 33404
rect 31948 29652 32004 29662
rect 31948 29426 32004 29596
rect 32284 29540 32340 29550
rect 32284 29446 32340 29484
rect 31948 29374 31950 29426
rect 32002 29374 32004 29426
rect 31948 29362 32004 29374
rect 32508 29428 32564 29438
rect 32508 29334 32564 29372
rect 30828 29138 30884 29148
rect 32396 29314 32452 29326
rect 32396 29262 32398 29314
rect 32450 29262 32452 29314
rect 32396 28866 32452 29262
rect 32396 28814 32398 28866
rect 32450 28814 32452 28866
rect 32396 28802 32452 28814
rect 29932 28690 29988 28700
rect 32060 28754 32116 28766
rect 32060 28702 32062 28754
rect 32114 28702 32116 28754
rect 30604 28644 30660 28654
rect 29932 28532 29988 28542
rect 29932 28530 30100 28532
rect 29932 28478 29934 28530
rect 29986 28478 30100 28530
rect 29932 28476 30100 28478
rect 29932 28466 29988 28476
rect 29596 28084 29652 28094
rect 29484 28082 29876 28084
rect 29484 28030 29598 28082
rect 29650 28030 29876 28082
rect 29484 28028 29876 28030
rect 29596 28018 29652 28028
rect 29820 27858 29876 28028
rect 30044 28082 30100 28476
rect 30044 28030 30046 28082
rect 30098 28030 30100 28082
rect 30044 28018 30100 28030
rect 30604 28082 30660 28588
rect 30604 28030 30606 28082
rect 30658 28030 30660 28082
rect 30604 28018 30660 28030
rect 30156 27972 30212 27982
rect 30156 27878 30212 27916
rect 30716 27972 30772 27982
rect 29820 27806 29822 27858
rect 29874 27806 29876 27858
rect 29820 27794 29876 27806
rect 30492 27636 30548 27646
rect 30268 27634 30548 27636
rect 30268 27582 30494 27634
rect 30546 27582 30548 27634
rect 30268 27580 30548 27582
rect 30268 27300 30324 27580
rect 30492 27570 30548 27580
rect 29932 27244 30324 27300
rect 29932 27186 29988 27244
rect 29932 27134 29934 27186
rect 29986 27134 29988 27186
rect 29932 27122 29988 27134
rect 29260 26982 29316 27020
rect 30716 26908 30772 27916
rect 32060 27972 32116 28702
rect 32620 28644 32676 29820
rect 32620 28530 32676 28588
rect 32620 28478 32622 28530
rect 32674 28478 32676 28530
rect 32620 28466 32676 28478
rect 32732 30098 32900 30100
rect 32732 30046 32846 30098
rect 32898 30046 32900 30098
rect 32732 30044 32900 30046
rect 32508 28420 32564 28430
rect 32508 28326 32564 28364
rect 32060 27906 32116 27916
rect 32284 27860 32340 27870
rect 32284 27766 32340 27804
rect 25564 26852 26068 26908
rect 26908 26852 27076 26908
rect 27804 26852 28308 26908
rect 26012 26402 26068 26852
rect 26012 26350 26014 26402
rect 26066 26350 26068 26402
rect 26012 26338 26068 26350
rect 24668 26126 24670 26178
rect 24722 26126 24724 26178
rect 22092 25566 22094 25618
rect 22146 25566 22148 25618
rect 22092 25554 22148 25566
rect 24220 25620 24276 25630
rect 24220 25618 24612 25620
rect 24220 25566 24222 25618
rect 24274 25566 24612 25618
rect 24220 25564 24612 25566
rect 24220 25554 24276 25564
rect 21308 25454 21310 25506
rect 21362 25454 21364 25506
rect 21308 25442 21364 25454
rect 20748 25004 21028 25060
rect 18060 24670 18062 24722
rect 18114 24670 18116 24722
rect 17276 23996 17780 24052
rect 17388 23828 17444 23838
rect 16828 23774 16830 23826
rect 16882 23774 16884 23826
rect 16828 23762 16884 23774
rect 17276 23826 17444 23828
rect 17276 23774 17390 23826
rect 17442 23774 17444 23826
rect 17276 23772 17444 23774
rect 16716 23156 16772 23166
rect 16604 23154 16884 23156
rect 16604 23102 16718 23154
rect 16770 23102 16884 23154
rect 16604 23100 16884 23102
rect 16716 23090 16772 23100
rect 16828 23044 16884 23100
rect 17276 23044 17332 23772
rect 17388 23762 17444 23772
rect 16828 22988 17332 23044
rect 17388 23154 17444 23166
rect 17388 23102 17390 23154
rect 17442 23102 17444 23154
rect 16716 22930 16772 22942
rect 16716 22878 16718 22930
rect 16770 22878 16772 22930
rect 16604 22148 16660 22158
rect 16604 21586 16660 22092
rect 16604 21534 16606 21586
rect 16658 21534 16660 21586
rect 16604 21522 16660 21534
rect 16716 21588 16772 22878
rect 16828 22260 16884 22270
rect 16828 22166 16884 22204
rect 16716 21522 16772 21532
rect 16716 21364 16772 21374
rect 16716 21270 16772 21308
rect 16492 20738 16548 20748
rect 16604 21140 16660 21150
rect 16604 20802 16660 21084
rect 16604 20750 16606 20802
rect 16658 20750 16660 20802
rect 16604 20020 16660 20750
rect 16940 20802 16996 22988
rect 17388 22596 17444 23102
rect 17388 22530 17444 22540
rect 16940 20750 16942 20802
rect 16994 20750 16996 20802
rect 16940 20738 16996 20750
rect 17388 22370 17444 22382
rect 17388 22318 17390 22370
rect 17442 22318 17444 22370
rect 17388 22260 17444 22318
rect 17388 21586 17444 22204
rect 17500 21700 17556 21710
rect 17500 21606 17556 21644
rect 17388 21534 17390 21586
rect 17442 21534 17444 21586
rect 17388 20804 17444 21534
rect 17500 20804 17556 20814
rect 17388 20802 17556 20804
rect 17388 20750 17502 20802
rect 17554 20750 17556 20802
rect 17388 20748 17556 20750
rect 16716 20692 16772 20702
rect 16716 20598 16772 20636
rect 16828 20580 16884 20590
rect 16828 20468 16884 20524
rect 16716 20412 16884 20468
rect 16716 20242 16772 20412
rect 16716 20190 16718 20242
rect 16770 20190 16772 20242
rect 16716 20188 16772 20190
rect 16716 20132 16884 20188
rect 16716 20020 16772 20030
rect 16604 19964 16716 20020
rect 16716 19926 16772 19964
rect 16828 19796 16884 20132
rect 17388 20020 17444 20030
rect 17388 19926 17444 19964
rect 16604 19740 16884 19796
rect 16156 19348 16212 19358
rect 15932 19292 16156 19348
rect 16156 19254 16212 19292
rect 15260 19122 15316 19134
rect 15260 19070 15262 19122
rect 15314 19070 15316 19122
rect 15260 18338 15316 19070
rect 15708 18340 15764 18350
rect 15260 18286 15262 18338
rect 15314 18286 15316 18338
rect 15260 17332 15316 18286
rect 15484 18338 15764 18340
rect 15484 18286 15710 18338
rect 15762 18286 15764 18338
rect 15484 18284 15764 18286
rect 15484 17668 15540 18284
rect 15708 18274 15764 18284
rect 15484 17574 15540 17612
rect 16156 17556 16212 17566
rect 16156 17554 16548 17556
rect 16156 17502 16158 17554
rect 16210 17502 16548 17554
rect 16156 17500 16548 17502
rect 16156 17490 16212 17500
rect 15260 17276 16212 17332
rect 16044 16884 16100 16894
rect 16044 16790 16100 16828
rect 15148 16046 15150 16098
rect 15202 16046 15204 16098
rect 15148 16034 15204 16046
rect 15820 16772 15876 16782
rect 14812 15922 14868 15932
rect 15484 15986 15540 15998
rect 15484 15934 15486 15986
rect 15538 15934 15540 15986
rect 15484 15204 15540 15934
rect 15820 15652 15876 16716
rect 15932 15988 15988 15998
rect 15932 15894 15988 15932
rect 16156 15986 16212 17276
rect 16492 17106 16548 17500
rect 16492 17054 16494 17106
rect 16546 17054 16548 17106
rect 16492 17042 16548 17054
rect 16268 16324 16324 16334
rect 16268 16230 16324 16268
rect 16156 15934 16158 15986
rect 16210 15934 16212 15986
rect 16156 15922 16212 15934
rect 15820 15596 16100 15652
rect 16044 15538 16100 15596
rect 16044 15486 16046 15538
rect 16098 15486 16100 15538
rect 16044 15474 16100 15486
rect 15596 15204 15652 15242
rect 15484 15148 15596 15204
rect 12124 15092 12292 15148
rect 12796 15138 12852 15148
rect 11340 14590 11342 14642
rect 11394 14590 11396 14642
rect 11340 13860 11396 14590
rect 11564 14642 11844 14644
rect 11564 14590 11790 14642
rect 11842 14590 11844 14642
rect 11564 14588 11844 14590
rect 11452 13860 11508 13870
rect 11340 13804 11452 13860
rect 11452 13746 11508 13804
rect 11452 13694 11454 13746
rect 11506 13694 11508 13746
rect 11452 13682 11508 13694
rect 11340 13636 11396 13646
rect 11228 13580 11340 13636
rect 8988 13022 8990 13074
rect 9042 13022 9044 13074
rect 8988 13010 9044 13022
rect 11004 13076 11060 13086
rect 8540 12674 8596 12684
rect 11004 12180 11060 13020
rect 11116 13076 11172 13086
rect 11228 13076 11284 13580
rect 11340 13570 11396 13580
rect 11116 13074 11284 13076
rect 11116 13022 11118 13074
rect 11170 13022 11284 13074
rect 11116 13020 11284 13022
rect 11564 13076 11620 14588
rect 11788 14578 11844 14588
rect 11900 14700 12068 14756
rect 11900 14420 11956 14700
rect 12236 14644 12292 15092
rect 11900 14354 11956 14364
rect 12012 14588 12292 14644
rect 13580 15092 13860 15148
rect 15596 15138 15652 15148
rect 12012 13858 12068 14588
rect 12012 13806 12014 13858
rect 12066 13806 12068 13858
rect 12012 13794 12068 13806
rect 12236 14420 12292 14430
rect 12236 13746 12292 14364
rect 13580 13748 13636 15092
rect 16604 14530 16660 19740
rect 17500 19236 17556 20748
rect 17724 19572 17780 23996
rect 18060 23940 18116 24670
rect 18508 24724 18564 24734
rect 18620 24724 18676 25004
rect 20076 24834 20132 24846
rect 20076 24782 20078 24834
rect 20130 24782 20132 24834
rect 18508 24722 18676 24724
rect 18508 24670 18510 24722
rect 18562 24670 18676 24722
rect 18508 24668 18676 24670
rect 18732 24722 18788 24734
rect 18732 24670 18734 24722
rect 18786 24670 18788 24722
rect 18284 24612 18340 24622
rect 18284 24518 18340 24556
rect 18508 24276 18564 24668
rect 18508 24210 18564 24220
rect 18732 24500 18788 24670
rect 19068 24724 19124 24734
rect 19068 24630 19124 24668
rect 19292 24724 19348 24734
rect 19292 24630 19348 24668
rect 19628 24724 19684 24734
rect 19684 24668 19796 24724
rect 19628 24658 19684 24668
rect 18396 24050 18452 24062
rect 18396 23998 18398 24050
rect 18450 23998 18452 24050
rect 18060 23874 18116 23884
rect 18172 23938 18228 23950
rect 18172 23886 18174 23938
rect 18226 23886 18228 23938
rect 18172 21924 18228 23886
rect 18396 23266 18452 23998
rect 18732 23940 18788 24444
rect 19628 24498 19684 24510
rect 19628 24446 19630 24498
rect 19682 24446 19684 24498
rect 19628 24164 19684 24446
rect 18732 23874 18788 23884
rect 18956 24108 19684 24164
rect 18396 23214 18398 23266
rect 18450 23214 18452 23266
rect 18172 21700 18228 21868
rect 18172 21634 18228 21644
rect 18284 22260 18340 22270
rect 18396 22260 18452 23214
rect 18956 23826 19012 24108
rect 19740 23938 19796 24668
rect 20076 24276 20132 24782
rect 20860 24834 20916 24846
rect 20860 24782 20862 24834
rect 20914 24782 20916 24834
rect 20412 24722 20468 24734
rect 20412 24670 20414 24722
rect 20466 24670 20468 24722
rect 20412 24500 20468 24670
rect 20748 24724 20804 24734
rect 20748 24630 20804 24668
rect 20860 24500 20916 24782
rect 20412 24444 20916 24500
rect 20076 24210 20132 24220
rect 19740 23886 19742 23938
rect 19794 23886 19796 23938
rect 19740 23874 19796 23886
rect 20412 23940 20468 23950
rect 18956 23774 18958 23826
rect 19010 23774 19012 23826
rect 18956 22596 19012 23774
rect 20188 23828 20244 23838
rect 19068 23714 19124 23726
rect 19068 23662 19070 23714
rect 19122 23662 19124 23714
rect 19068 22932 19124 23662
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19068 22866 19124 22876
rect 19180 23042 19236 23054
rect 19180 22990 19182 23042
rect 19234 22990 19236 23042
rect 18956 22530 19012 22540
rect 18284 22258 18452 22260
rect 18284 22206 18286 22258
rect 18338 22206 18452 22258
rect 18284 22204 18452 22206
rect 19068 22372 19124 22382
rect 19180 22372 19236 22990
rect 19740 23044 19796 23054
rect 19740 22950 19796 22988
rect 20188 22482 20244 23772
rect 20188 22430 20190 22482
rect 20242 22430 20244 22482
rect 20188 22418 20244 22430
rect 20300 23826 20356 23838
rect 20300 23774 20302 23826
rect 20354 23774 20356 23826
rect 19068 22370 19236 22372
rect 19068 22318 19070 22370
rect 19122 22318 19236 22370
rect 19068 22316 19236 22318
rect 17724 19506 17780 19516
rect 18284 20132 18340 22204
rect 18396 21588 18452 21598
rect 18396 20690 18452 21532
rect 19068 20916 19124 22316
rect 19628 22146 19684 22158
rect 19628 22094 19630 22146
rect 19682 22094 19684 22146
rect 19068 20850 19124 20860
rect 19180 21700 19236 21710
rect 19180 21588 19236 21644
rect 19404 21588 19460 21598
rect 19180 21586 19460 21588
rect 19180 21534 19406 21586
rect 19458 21534 19460 21586
rect 19180 21532 19460 21534
rect 19180 20914 19236 21532
rect 19404 21522 19460 21532
rect 19628 21588 19684 22094
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21522 19684 21532
rect 19180 20862 19182 20914
rect 19234 20862 19236 20914
rect 19180 20850 19236 20862
rect 18396 20638 18398 20690
rect 18450 20638 18452 20690
rect 18396 20626 18452 20638
rect 18508 20692 18564 20702
rect 18396 20132 18452 20142
rect 18284 20130 18452 20132
rect 18284 20078 18398 20130
rect 18450 20078 18452 20130
rect 18284 20076 18452 20078
rect 17724 19236 17780 19246
rect 17500 19234 17780 19236
rect 17500 19182 17726 19234
rect 17778 19182 17780 19234
rect 17500 19180 17780 19182
rect 17724 19170 17780 19180
rect 18284 19122 18340 20076
rect 18396 20066 18452 20076
rect 18284 19070 18286 19122
rect 18338 19070 18340 19122
rect 18284 19058 18340 19070
rect 18508 18788 18564 20636
rect 18956 20578 19012 20590
rect 18956 20526 18958 20578
rect 19010 20526 19012 20578
rect 18396 18732 18564 18788
rect 18844 19348 18900 19358
rect 17500 18562 17556 18574
rect 17500 18510 17502 18562
rect 17554 18510 17556 18562
rect 17500 17332 17556 18510
rect 17836 18450 17892 18462
rect 17836 18398 17838 18450
rect 17890 18398 17892 18450
rect 17836 17780 17892 18398
rect 18284 18450 18340 18462
rect 18284 18398 18286 18450
rect 18338 18398 18340 18450
rect 18284 18004 18340 18398
rect 18396 18116 18452 18732
rect 18508 18562 18564 18574
rect 18508 18510 18510 18562
rect 18562 18510 18564 18562
rect 18508 18340 18564 18510
rect 18844 18450 18900 19292
rect 18844 18398 18846 18450
rect 18898 18398 18900 18450
rect 18844 18386 18900 18398
rect 18508 18274 18564 18284
rect 18956 18228 19012 20526
rect 18396 18060 18564 18116
rect 18284 17938 18340 17948
rect 18396 17892 18452 17902
rect 18284 17780 18340 17790
rect 18396 17780 18452 17836
rect 17836 17714 17892 17724
rect 17948 17778 18452 17780
rect 17948 17726 18286 17778
rect 18338 17726 18452 17778
rect 17948 17724 18452 17726
rect 17500 17266 17556 17276
rect 16828 16996 16884 17006
rect 16828 16902 16884 16940
rect 17500 16996 17556 17006
rect 17500 16902 17556 16940
rect 16716 16884 16772 16894
rect 16716 16210 16772 16828
rect 17836 16884 17892 16894
rect 17948 16884 18004 17724
rect 18284 17714 18340 17724
rect 17836 16882 18004 16884
rect 17836 16830 17838 16882
rect 17890 16830 18004 16882
rect 17836 16828 18004 16830
rect 18284 17444 18340 17454
rect 17836 16818 17892 16828
rect 18284 16772 18340 17388
rect 18396 17332 18452 17342
rect 18396 16994 18452 17276
rect 18396 16942 18398 16994
rect 18450 16942 18452 16994
rect 18396 16930 18452 16942
rect 18284 16706 18340 16716
rect 16716 16158 16718 16210
rect 16770 16158 16772 16210
rect 16716 16146 16772 16158
rect 16604 14478 16606 14530
rect 16658 14478 16660 14530
rect 16380 14420 16436 14430
rect 16380 14326 16436 14364
rect 13692 13860 13748 13870
rect 15484 13860 15540 13870
rect 13692 13766 13748 13804
rect 15148 13858 15540 13860
rect 15148 13806 15486 13858
rect 15538 13806 15540 13858
rect 15148 13804 15540 13806
rect 12236 13694 12238 13746
rect 12290 13694 12292 13746
rect 12236 13682 12292 13694
rect 13468 13746 13636 13748
rect 13468 13694 13582 13746
rect 13634 13694 13636 13746
rect 13468 13692 13636 13694
rect 11116 13010 11172 13020
rect 11564 12982 11620 13020
rect 10444 12178 11060 12180
rect 10444 12126 11006 12178
rect 11058 12126 11060 12178
rect 10444 12124 11060 12126
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 10444 10610 10500 12124
rect 11004 12114 11060 12124
rect 11676 12066 11732 12078
rect 11676 12014 11678 12066
rect 11730 12014 11732 12066
rect 11676 11284 11732 12014
rect 12460 11956 12516 11966
rect 12460 11394 12516 11900
rect 12460 11342 12462 11394
rect 12514 11342 12516 11394
rect 12460 11330 12516 11342
rect 12124 11284 12180 11294
rect 11676 11282 12180 11284
rect 11676 11230 12126 11282
rect 12178 11230 12180 11282
rect 11676 11228 12180 11230
rect 12124 11218 12180 11228
rect 13468 10724 13524 13692
rect 13580 13682 13636 13692
rect 14364 13524 14420 13534
rect 14700 13524 14756 13534
rect 13804 13522 14644 13524
rect 13804 13470 14366 13522
rect 14418 13470 14644 13522
rect 13804 13468 14644 13470
rect 13804 12066 13860 13468
rect 14364 13458 14420 13468
rect 13804 12014 13806 12066
rect 13858 12014 13860 12066
rect 13804 12002 13860 12014
rect 14028 13076 14084 13086
rect 14028 11508 14084 13020
rect 14364 13076 14420 13086
rect 14364 12962 14420 13020
rect 14364 12910 14366 12962
rect 14418 12910 14420 12962
rect 14364 12898 14420 12910
rect 14588 12178 14644 13468
rect 14700 13430 14756 13468
rect 15148 13074 15204 13804
rect 15484 13794 15540 13804
rect 16492 13858 16548 13870
rect 16492 13806 16494 13858
rect 16546 13806 16548 13858
rect 15820 13746 15876 13758
rect 15820 13694 15822 13746
rect 15874 13694 15876 13746
rect 15148 13022 15150 13074
rect 15202 13022 15204 13074
rect 15148 13010 15204 13022
rect 15372 13188 15428 13198
rect 14588 12126 14590 12178
rect 14642 12126 14644 12178
rect 14588 12114 14644 12126
rect 15260 12290 15316 12302
rect 15260 12238 15262 12290
rect 15314 12238 15316 12290
rect 14252 11956 14308 11966
rect 14252 11862 14308 11900
rect 13468 10658 13524 10668
rect 13580 11506 14084 11508
rect 13580 11454 14030 11506
rect 14082 11454 14084 11506
rect 13580 11452 14084 11454
rect 10444 10558 10446 10610
rect 10498 10558 10500 10610
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 10444 9044 10500 10558
rect 11116 10500 11172 10510
rect 13244 10500 13300 10510
rect 11116 10498 11396 10500
rect 11116 10446 11118 10498
rect 11170 10446 11396 10498
rect 11116 10444 11396 10446
rect 11116 10434 11172 10444
rect 11340 9714 11396 10444
rect 13244 10406 13300 10444
rect 13580 9940 13636 11452
rect 14028 11442 14084 11452
rect 15148 11844 15204 11854
rect 15036 10836 15092 10846
rect 15148 10836 15204 11788
rect 15036 10834 15204 10836
rect 15036 10782 15038 10834
rect 15090 10782 15204 10834
rect 15036 10780 15204 10782
rect 15036 10770 15092 10780
rect 14140 10724 14196 10734
rect 14476 10724 14532 10734
rect 14140 10722 14308 10724
rect 14140 10670 14142 10722
rect 14194 10670 14308 10722
rect 14140 10668 14308 10670
rect 14140 10658 14196 10668
rect 13468 9938 13636 9940
rect 13468 9886 13582 9938
rect 13634 9886 13636 9938
rect 13468 9884 13636 9886
rect 11340 9662 11342 9714
rect 11394 9662 11396 9714
rect 11340 9650 11396 9662
rect 11676 9716 11732 9726
rect 11676 9622 11732 9660
rect 13468 9156 13524 9884
rect 13580 9874 13636 9884
rect 14028 9716 14084 9726
rect 14028 9622 14084 9660
rect 13356 9100 13524 9156
rect 10556 9044 10612 9054
rect 10444 9042 10612 9044
rect 10444 8990 10558 9042
rect 10610 8990 10612 9042
rect 10444 8988 10612 8990
rect 10556 8978 10612 8988
rect 11340 8930 11396 8942
rect 11340 8878 11342 8930
rect 11394 8878 11396 8930
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 11340 8428 11396 8878
rect 11900 8820 11956 8830
rect 11340 8372 11620 8428
rect 11564 8146 11620 8372
rect 11900 8258 11956 8764
rect 13356 8708 13412 9100
rect 14252 9044 14308 10668
rect 14476 10630 14532 10668
rect 14364 10500 14420 10510
rect 14364 10050 14420 10444
rect 14700 10500 14756 10510
rect 14700 10406 14756 10444
rect 14364 9998 14366 10050
rect 14418 9998 14420 10050
rect 14364 9986 14420 9998
rect 15260 10052 15316 12238
rect 15372 12178 15428 13132
rect 15820 12964 15876 13694
rect 16492 13636 16548 13806
rect 16604 13746 16660 14478
rect 16604 13694 16606 13746
rect 16658 13694 16660 13746
rect 16604 13682 16660 13694
rect 16940 15428 16996 15438
rect 16940 14418 16996 15372
rect 17612 15426 17668 15438
rect 17612 15374 17614 15426
rect 17666 15374 17668 15426
rect 17388 15204 17444 15242
rect 17388 15138 17444 15148
rect 17388 14756 17444 14766
rect 17388 14532 17444 14700
rect 16940 14366 16942 14418
rect 16994 14366 16996 14418
rect 16492 13570 16548 13580
rect 16716 13522 16772 13534
rect 16716 13470 16718 13522
rect 16770 13470 16772 13522
rect 16716 13188 16772 13470
rect 16716 13122 16772 13132
rect 15820 12898 15876 12908
rect 15372 12126 15374 12178
rect 15426 12126 15428 12178
rect 15372 12114 15428 12126
rect 16044 11732 16100 11742
rect 15708 11394 15764 11406
rect 15708 11342 15710 11394
rect 15762 11342 15764 11394
rect 15708 10724 15764 11342
rect 15708 10658 15764 10668
rect 15260 9986 15316 9996
rect 14812 9826 14868 9838
rect 14812 9774 14814 9826
rect 14866 9774 14868 9826
rect 14812 9716 14868 9774
rect 14812 9650 14868 9660
rect 14924 9714 14980 9726
rect 14924 9662 14926 9714
rect 14978 9662 14980 9714
rect 14924 9156 14980 9662
rect 15932 9604 15988 9614
rect 15596 9156 15652 9166
rect 14924 9062 14980 9100
rect 15372 9154 15652 9156
rect 15372 9102 15598 9154
rect 15650 9102 15652 9154
rect 15372 9100 15652 9102
rect 13804 9042 14308 9044
rect 13804 8990 14254 9042
rect 14306 8990 14308 9042
rect 13804 8988 14308 8990
rect 13468 8930 13524 8942
rect 13468 8878 13470 8930
rect 13522 8878 13524 8930
rect 13468 8820 13524 8878
rect 13804 8820 13860 8988
rect 14252 8978 14308 8988
rect 15036 9044 15092 9054
rect 15036 8950 15092 8988
rect 13468 8764 13860 8820
rect 13916 8820 13972 8830
rect 13916 8726 13972 8764
rect 13356 8652 13636 8708
rect 11900 8206 11902 8258
rect 11954 8206 11956 8258
rect 11900 8194 11956 8206
rect 11564 8094 11566 8146
rect 11618 8094 11620 8146
rect 11564 8082 11620 8094
rect 13580 8036 13636 8652
rect 15148 8372 15204 8382
rect 15036 8316 15148 8372
rect 13692 8036 13748 8046
rect 14812 8036 14868 8046
rect 13580 8034 13748 8036
rect 13580 7982 13694 8034
rect 13746 7982 13748 8034
rect 13580 7980 13748 7982
rect 12236 7476 12292 7486
rect 12236 7382 12292 7420
rect 13580 7476 13636 7980
rect 13692 7970 13748 7980
rect 13804 8034 14868 8036
rect 13804 7982 14814 8034
rect 14866 7982 14868 8034
rect 13804 7980 14868 7982
rect 12908 7364 12964 7374
rect 12908 7362 13524 7364
rect 12908 7310 12910 7362
rect 12962 7310 13524 7362
rect 12908 7308 13524 7310
rect 12908 7298 12964 7308
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 13468 6578 13524 7308
rect 13468 6526 13470 6578
rect 13522 6526 13524 6578
rect 13468 6514 13524 6526
rect 13356 5908 13412 5918
rect 13580 5908 13636 7420
rect 13804 6690 13860 7980
rect 14812 7970 14868 7980
rect 15036 7362 15092 8316
rect 15148 8278 15204 8316
rect 15036 7310 15038 7362
rect 15090 7310 15092 7362
rect 15036 7298 15092 7310
rect 15372 6916 15428 9100
rect 15596 9090 15652 9100
rect 15932 8258 15988 9548
rect 16044 9154 16100 11676
rect 16716 11284 16772 11294
rect 16268 11172 16324 11182
rect 16268 11078 16324 11116
rect 16716 9266 16772 11228
rect 16940 9716 16996 14366
rect 17164 14530 17444 14532
rect 17164 14478 17390 14530
rect 17442 14478 17444 14530
rect 17164 14476 17444 14478
rect 17164 12180 17220 14476
rect 17388 14466 17444 14476
rect 17612 14084 17668 15374
rect 18396 15426 18452 15438
rect 18396 15374 18398 15426
rect 18450 15374 18452 15426
rect 18396 15148 18452 15374
rect 17724 15092 17780 15102
rect 17724 14998 17780 15036
rect 18172 15092 18452 15148
rect 18172 14642 18228 15092
rect 18172 14590 18174 14642
rect 18226 14590 18228 14642
rect 18172 14578 18228 14590
rect 17612 14028 17780 14084
rect 17612 13860 17668 13870
rect 17612 13766 17668 13804
rect 17724 13746 17780 14028
rect 17724 13694 17726 13746
rect 17778 13694 17780 13746
rect 17724 13524 17780 13694
rect 18284 13524 18340 13534
rect 17612 13468 17780 13524
rect 18060 13522 18340 13524
rect 18060 13470 18286 13522
rect 18338 13470 18340 13522
rect 18060 13468 18340 13470
rect 17276 13300 17332 13310
rect 17276 13074 17332 13244
rect 17276 13022 17278 13074
rect 17330 13022 17332 13074
rect 17276 13010 17332 13022
rect 17500 13076 17556 13086
rect 17500 12402 17556 13020
rect 17500 12350 17502 12402
rect 17554 12350 17556 12402
rect 17500 12338 17556 12350
rect 17164 11396 17220 12124
rect 17500 11732 17556 11742
rect 17612 11732 17668 13468
rect 18060 13300 18116 13468
rect 18284 13458 18340 13468
rect 18508 13412 18564 18060
rect 18844 17780 18900 17790
rect 18844 17686 18900 17724
rect 18620 17556 18676 17566
rect 18620 16884 18676 17500
rect 18956 16996 19012 18172
rect 19068 20580 19124 20590
rect 19068 17668 19124 20524
rect 19180 20468 19236 20478
rect 19180 19906 19236 20412
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19740 20244 19796 20254
rect 19740 20150 19796 20188
rect 19180 19854 19182 19906
rect 19234 19854 19236 19906
rect 19180 19348 19236 19854
rect 19516 19348 19572 19358
rect 19180 19346 19572 19348
rect 19180 19294 19518 19346
rect 19570 19294 19572 19346
rect 19180 19292 19572 19294
rect 19516 19282 19572 19292
rect 19628 19010 19684 19022
rect 19628 18958 19630 19010
rect 19682 18958 19684 19010
rect 19628 18676 19684 18958
rect 20188 19012 20244 19022
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18610 19684 18620
rect 19628 18340 19684 18350
rect 19628 18246 19684 18284
rect 19292 18004 19348 18014
rect 19292 17890 19348 17948
rect 19292 17838 19294 17890
rect 19346 17838 19348 17890
rect 19292 17826 19348 17838
rect 19628 17668 19684 17678
rect 19068 17612 19348 17668
rect 19180 17220 19236 17230
rect 18956 16940 19124 16996
rect 18620 16882 19012 16884
rect 18620 16830 18622 16882
rect 18674 16830 19012 16882
rect 18620 16828 19012 16830
rect 18620 16818 18676 16828
rect 18956 16098 19012 16828
rect 18956 16046 18958 16098
rect 19010 16046 19012 16098
rect 18956 16034 19012 16046
rect 19068 16660 19124 16940
rect 19180 16994 19236 17164
rect 19180 16942 19182 16994
rect 19234 16942 19236 16994
rect 19180 16930 19236 16942
rect 19292 16882 19348 17612
rect 19628 17574 19684 17612
rect 19852 17556 19908 17566
rect 19852 17462 19908 17500
rect 20188 17554 20244 18956
rect 20188 17502 20190 17554
rect 20242 17502 20244 17554
rect 20188 17490 20244 17502
rect 19628 17444 19684 17454
rect 19628 16994 19684 17388
rect 20300 17444 20356 23774
rect 20412 23604 20468 23884
rect 20412 23538 20468 23548
rect 20636 23938 20692 24444
rect 20636 23886 20638 23938
rect 20690 23886 20692 23938
rect 20636 23380 20692 23886
rect 20860 24276 20916 24286
rect 20636 23314 20692 23324
rect 20748 23604 20804 23614
rect 20748 23266 20804 23548
rect 20748 23214 20750 23266
rect 20802 23214 20804 23266
rect 20748 23202 20804 23214
rect 20860 23266 20916 24220
rect 20972 23828 21028 25004
rect 21084 24724 21140 24734
rect 21084 24722 21252 24724
rect 21084 24670 21086 24722
rect 21138 24670 21252 24722
rect 21084 24668 21252 24670
rect 21084 24658 21140 24668
rect 20972 23762 21028 23772
rect 20860 23214 20862 23266
rect 20914 23214 20916 23266
rect 20860 23202 20916 23214
rect 20972 23156 21028 23166
rect 20412 22596 20468 22606
rect 20412 22502 20468 22540
rect 20748 22148 20804 22158
rect 20748 22146 20916 22148
rect 20748 22094 20750 22146
rect 20802 22094 20916 22146
rect 20748 22092 20916 22094
rect 20748 22082 20804 22092
rect 20524 21700 20580 21710
rect 20412 21698 20580 21700
rect 20412 21646 20526 21698
rect 20578 21646 20580 21698
rect 20412 21644 20580 21646
rect 20412 20804 20468 21644
rect 20524 21634 20580 21644
rect 20524 20916 20580 20926
rect 20524 20822 20580 20860
rect 20412 20710 20468 20748
rect 20412 20468 20468 20478
rect 20412 20018 20468 20412
rect 20412 19966 20414 20018
rect 20466 19966 20468 20018
rect 20412 19348 20468 19966
rect 20748 19348 20804 19358
rect 20468 19346 20804 19348
rect 20468 19294 20750 19346
rect 20802 19294 20804 19346
rect 20468 19292 20804 19294
rect 20412 19282 20468 19292
rect 20748 19282 20804 19292
rect 20524 18788 20580 18798
rect 20524 17780 20580 18732
rect 20860 18676 20916 22092
rect 20972 21812 21028 23100
rect 21196 22596 21252 24668
rect 23996 23938 24052 23950
rect 23996 23886 23998 23938
rect 24050 23886 24052 23938
rect 21308 23828 21364 23838
rect 21308 23734 21364 23772
rect 21756 23828 21812 23838
rect 21644 23714 21700 23726
rect 21644 23662 21646 23714
rect 21698 23662 21700 23714
rect 21532 23604 21588 23614
rect 21420 23492 21476 23502
rect 21420 23378 21476 23436
rect 21420 23326 21422 23378
rect 21474 23326 21476 23378
rect 21420 23314 21476 23326
rect 21308 22596 21364 22606
rect 21196 22594 21364 22596
rect 21196 22542 21310 22594
rect 21362 22542 21364 22594
rect 21196 22540 21364 22542
rect 21308 22530 21364 22540
rect 21532 22258 21588 23548
rect 21644 23380 21700 23662
rect 21644 22372 21700 23324
rect 21756 23042 21812 23772
rect 23548 23828 23604 23838
rect 23548 23734 23604 23772
rect 22204 23714 22260 23726
rect 22204 23662 22206 23714
rect 22258 23662 22260 23714
rect 22204 23156 22260 23662
rect 23212 23716 23268 23726
rect 23212 23622 23268 23660
rect 23660 23714 23716 23726
rect 23660 23662 23662 23714
rect 23714 23662 23716 23714
rect 23660 23268 23716 23662
rect 23996 23716 24052 23886
rect 23996 23650 24052 23660
rect 23660 23212 24052 23268
rect 22204 23090 22260 23100
rect 21756 22990 21758 23042
rect 21810 22990 21812 23042
rect 21756 22978 21812 22990
rect 22764 23044 22820 23054
rect 21980 22932 22036 22942
rect 21980 22594 22036 22876
rect 21980 22542 21982 22594
rect 22034 22542 22036 22594
rect 21980 22530 22036 22542
rect 21644 22316 22260 22372
rect 21532 22206 21534 22258
rect 21586 22206 21588 22258
rect 21532 22194 21588 22206
rect 21644 22204 22148 22260
rect 21420 22148 21476 22158
rect 21420 22054 21476 22092
rect 21084 21812 21140 21822
rect 20972 21810 21140 21812
rect 20972 21758 21086 21810
rect 21138 21758 21140 21810
rect 20972 21756 21140 21758
rect 21084 20804 21140 21756
rect 21644 20804 21700 22204
rect 22092 22146 22148 22204
rect 22204 22258 22260 22316
rect 22204 22206 22206 22258
rect 22258 22206 22260 22258
rect 22204 22194 22260 22206
rect 22092 22094 22094 22146
rect 22146 22094 22148 22146
rect 22092 22082 22148 22094
rect 22652 22148 22708 22158
rect 21980 22036 22036 22046
rect 21980 21810 22036 21980
rect 21980 21758 21982 21810
rect 22034 21758 22036 21810
rect 21980 21746 22036 21758
rect 21868 21698 21924 21710
rect 21868 21646 21870 21698
rect 21922 21646 21924 21698
rect 21868 21028 21924 21646
rect 21980 21588 22036 21598
rect 21980 21494 22036 21532
rect 22652 21586 22708 22092
rect 22652 21534 22654 21586
rect 22706 21534 22708 21586
rect 22652 21476 22708 21534
rect 22652 21410 22708 21420
rect 21868 20972 22036 21028
rect 21084 20738 21140 20748
rect 21420 20748 21700 20804
rect 21084 19908 21140 19918
rect 21084 19814 21140 19852
rect 21308 19012 21364 19022
rect 21308 18918 21364 18956
rect 20524 17714 20580 17724
rect 20636 18620 20916 18676
rect 20300 17378 20356 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16942 19630 16994
rect 19682 16942 19684 16994
rect 19628 16930 19684 16942
rect 20188 16996 20244 17006
rect 19292 16830 19294 16882
rect 19346 16830 19348 16882
rect 19292 16818 19348 16830
rect 19068 16604 19348 16660
rect 18732 15876 18788 15886
rect 19068 15876 19124 16604
rect 19292 16098 19348 16604
rect 20188 16324 20244 16940
rect 20188 16258 20244 16268
rect 20300 16548 20356 16558
rect 19292 16046 19294 16098
rect 19346 16046 19348 16098
rect 19292 16034 19348 16046
rect 20076 16212 20132 16222
rect 18732 15874 19124 15876
rect 18732 15822 18734 15874
rect 18786 15822 19124 15874
rect 18732 15820 19124 15822
rect 19180 15874 19236 15886
rect 19180 15822 19182 15874
rect 19234 15822 19236 15874
rect 18732 15810 18788 15820
rect 19180 15428 19236 15822
rect 20076 15876 20132 16156
rect 20076 15820 20244 15876
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19292 15428 19348 15438
rect 19180 15372 19292 15428
rect 19292 15334 19348 15372
rect 18732 15314 18788 15326
rect 18732 15262 18734 15314
rect 18786 15262 18788 15314
rect 18732 15148 18788 15262
rect 19628 15316 19684 15354
rect 19628 15250 19684 15260
rect 20076 15316 20132 15326
rect 20188 15316 20244 15820
rect 20076 15314 20244 15316
rect 20076 15262 20078 15314
rect 20130 15262 20244 15314
rect 20076 15260 20244 15262
rect 18732 15092 19684 15148
rect 19180 14532 19236 14542
rect 18620 13748 18676 13758
rect 18620 13654 18676 13692
rect 19180 13636 19236 14476
rect 19628 13972 19684 15092
rect 20076 14756 20132 15260
rect 20076 14690 20132 14700
rect 20300 14644 20356 16492
rect 20188 14642 20356 14644
rect 20188 14590 20302 14642
rect 20354 14590 20356 14642
rect 20188 14588 20356 14590
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19740 13972 19796 13982
rect 19628 13970 19796 13972
rect 19628 13918 19742 13970
rect 19794 13918 19796 13970
rect 19628 13916 19796 13918
rect 19740 13906 19796 13916
rect 20076 13748 20132 13758
rect 20188 13748 20244 14588
rect 20300 14578 20356 14588
rect 20636 14532 20692 18620
rect 20972 18228 21028 18238
rect 20972 17220 21028 18172
rect 20972 17106 21028 17164
rect 20972 17054 20974 17106
rect 21026 17054 21028 17106
rect 20972 17042 21028 17054
rect 21308 16994 21364 17006
rect 21308 16942 21310 16994
rect 21362 16942 21364 16994
rect 21308 16100 21364 16942
rect 20748 16044 21364 16100
rect 20748 15426 20804 16044
rect 21420 15988 21476 20748
rect 21868 20690 21924 20702
rect 21868 20638 21870 20690
rect 21922 20638 21924 20690
rect 21532 20578 21588 20590
rect 21532 20526 21534 20578
rect 21586 20526 21588 20578
rect 21532 20468 21588 20526
rect 21756 20580 21812 20590
rect 21868 20580 21924 20638
rect 21980 20692 22036 20972
rect 21980 20598 22036 20636
rect 22428 20802 22484 20814
rect 22428 20750 22430 20802
rect 22482 20750 22484 20802
rect 21812 20524 21924 20580
rect 22204 20580 22260 20590
rect 21756 20514 21812 20524
rect 21532 17778 21588 20412
rect 22204 20356 22260 20524
rect 21980 20300 22260 20356
rect 22428 20468 22484 20750
rect 21644 19236 21700 19246
rect 21644 19142 21700 19180
rect 21980 19234 22036 20300
rect 22092 19908 22148 19918
rect 22092 19346 22148 19852
rect 22092 19294 22094 19346
rect 22146 19294 22148 19346
rect 22092 19282 22148 19294
rect 22316 19796 22372 19806
rect 21980 19182 21982 19234
rect 22034 19182 22036 19234
rect 21980 19170 22036 19182
rect 22316 19234 22372 19740
rect 22428 19348 22484 20412
rect 22428 19282 22484 19292
rect 22540 20244 22596 20254
rect 22316 19182 22318 19234
rect 22370 19182 22372 19234
rect 22316 18452 22372 19182
rect 22540 19234 22596 20188
rect 22764 19460 22820 22988
rect 23884 23042 23940 23054
rect 23884 22990 23886 23042
rect 23938 22990 23940 23042
rect 23660 22596 23716 22606
rect 23436 22372 23492 22382
rect 23660 22372 23716 22540
rect 23436 22370 23716 22372
rect 23436 22318 23438 22370
rect 23490 22318 23662 22370
rect 23714 22318 23716 22370
rect 23436 22316 23716 22318
rect 23436 22306 23492 22316
rect 23660 22306 23716 22316
rect 23100 22258 23156 22270
rect 23100 22206 23102 22258
rect 23154 22206 23156 22258
rect 22876 22148 22932 22158
rect 23100 22148 23156 22206
rect 22876 22146 23156 22148
rect 22876 22094 22878 22146
rect 22930 22094 23156 22146
rect 22876 22092 23156 22094
rect 23212 22146 23268 22158
rect 23212 22094 23214 22146
rect 23266 22094 23268 22146
rect 22876 20916 22932 22092
rect 22876 20850 22932 20860
rect 22988 21476 23044 21486
rect 23212 21476 23268 22094
rect 23884 22146 23940 22990
rect 23884 22094 23886 22146
rect 23938 22094 23940 22146
rect 23884 22082 23940 22094
rect 23996 22258 24052 23212
rect 24220 23044 24276 23054
rect 23996 22206 23998 22258
rect 24050 22206 24052 22258
rect 23996 21812 24052 22206
rect 23884 21756 24052 21812
rect 24108 22372 24164 22382
rect 22988 21474 23268 21476
rect 22988 21422 22990 21474
rect 23042 21422 23268 21474
rect 22988 21420 23268 21422
rect 23772 21474 23828 21486
rect 23772 21422 23774 21474
rect 23826 21422 23828 21474
rect 22988 20692 23044 21420
rect 23660 21362 23716 21374
rect 23660 21310 23662 21362
rect 23714 21310 23716 21362
rect 23212 20692 23268 20702
rect 22764 19404 22932 19460
rect 22876 19236 22932 19404
rect 22540 19182 22542 19234
rect 22594 19182 22596 19234
rect 22540 19170 22596 19182
rect 22652 19234 22932 19236
rect 22652 19182 22878 19234
rect 22930 19182 22932 19234
rect 22652 19180 22932 19182
rect 22540 18676 22596 18686
rect 22652 18676 22708 19180
rect 22876 19170 22932 19180
rect 22988 19122 23044 20636
rect 23100 20690 23268 20692
rect 23100 20638 23214 20690
rect 23266 20638 23268 20690
rect 23100 20636 23268 20638
rect 23100 20132 23156 20636
rect 23212 20626 23268 20636
rect 23660 20580 23716 21310
rect 23660 20514 23716 20524
rect 23772 20244 23828 21422
rect 23772 20178 23828 20188
rect 23100 20066 23156 20076
rect 23660 20020 23716 20030
rect 23212 20018 23716 20020
rect 23212 19966 23662 20018
rect 23714 19966 23716 20018
rect 23212 19964 23716 19966
rect 22988 19070 22990 19122
rect 23042 19070 23044 19122
rect 22988 19058 23044 19070
rect 23100 19908 23156 19918
rect 23100 18676 23156 19852
rect 23212 19906 23268 19964
rect 23660 19954 23716 19964
rect 23212 19854 23214 19906
rect 23266 19854 23268 19906
rect 23212 19842 23268 19854
rect 23548 19796 23604 19806
rect 23884 19796 23940 21756
rect 23996 21588 24052 21598
rect 24108 21588 24164 22316
rect 24220 22370 24276 22988
rect 24220 22318 24222 22370
rect 24274 22318 24276 22370
rect 24220 22306 24276 22318
rect 23996 21586 24164 21588
rect 23996 21534 23998 21586
rect 24050 21534 24164 21586
rect 23996 21532 24164 21534
rect 23996 21522 24052 21532
rect 24332 21362 24388 21374
rect 24332 21310 24334 21362
rect 24386 21310 24388 21362
rect 23996 20580 24052 20590
rect 24332 20580 24388 21310
rect 24052 20524 24388 20580
rect 23996 20018 24052 20524
rect 24220 20132 24276 20142
rect 24220 20038 24276 20076
rect 23996 19966 23998 20018
rect 24050 19966 24052 20018
rect 23996 19954 24052 19966
rect 24444 20020 24500 20030
rect 24444 19926 24500 19964
rect 23884 19740 24164 19796
rect 23548 19702 23604 19740
rect 23996 19348 24052 19358
rect 23996 19254 24052 19292
rect 23884 19124 23940 19134
rect 23436 19012 23492 19022
rect 23436 18918 23492 18956
rect 22540 18674 22708 18676
rect 22540 18622 22542 18674
rect 22594 18622 22708 18674
rect 22540 18620 22708 18622
rect 22540 18610 22596 18620
rect 22316 18396 22596 18452
rect 21532 17726 21534 17778
rect 21586 17726 21588 17778
rect 21532 17714 21588 17726
rect 21756 18338 21812 18350
rect 21756 18286 21758 18338
rect 21810 18286 21812 18338
rect 21756 17668 21812 18286
rect 21756 17602 21812 17612
rect 22428 18004 22484 18014
rect 22092 17444 22148 17454
rect 22092 17108 22148 17388
rect 21980 17106 22148 17108
rect 21980 17054 22094 17106
rect 22146 17054 22148 17106
rect 21980 17052 22148 17054
rect 20748 15374 20750 15426
rect 20802 15374 20804 15426
rect 20748 15362 20804 15374
rect 21308 15932 21476 15988
rect 21532 16882 21588 16894
rect 21532 16830 21534 16882
rect 21586 16830 21588 16882
rect 21308 15316 21364 15932
rect 20748 14756 20804 14766
rect 20748 14642 20804 14700
rect 20748 14590 20750 14642
rect 20802 14590 20804 14642
rect 20748 14578 20804 14590
rect 20636 14466 20692 14476
rect 20860 14420 20916 14430
rect 20636 13860 20692 13870
rect 20076 13746 20244 13748
rect 20076 13694 20078 13746
rect 20130 13694 20244 13746
rect 20076 13692 20244 13694
rect 20524 13858 20692 13860
rect 20524 13806 20638 13858
rect 20690 13806 20692 13858
rect 20524 13804 20692 13806
rect 20076 13682 20132 13692
rect 18508 13356 19124 13412
rect 18060 13186 18116 13244
rect 18060 13134 18062 13186
rect 18114 13134 18116 13186
rect 18060 13122 18116 13134
rect 18508 13188 18564 13198
rect 17724 12964 17780 12974
rect 17724 12870 17780 12908
rect 18508 12962 18564 13132
rect 18508 12910 18510 12962
rect 18562 12910 18564 12962
rect 18508 12898 18564 12910
rect 18732 12850 18788 12862
rect 18732 12798 18734 12850
rect 18786 12798 18788 12850
rect 18732 11788 18788 12798
rect 18732 11732 18900 11788
rect 17556 11676 17668 11732
rect 17500 11666 17556 11676
rect 17276 11396 17332 11406
rect 17164 11394 17332 11396
rect 17164 11342 17278 11394
rect 17330 11342 17332 11394
rect 17164 11340 17332 11342
rect 17276 11330 17332 11340
rect 17612 10836 17668 11676
rect 18060 11284 18116 11294
rect 18060 11282 18676 11284
rect 18060 11230 18062 11282
rect 18114 11230 18676 11282
rect 18060 11228 18676 11230
rect 18060 11218 18116 11228
rect 17612 10770 17668 10780
rect 18508 11060 18564 11070
rect 17836 10612 17892 10622
rect 18508 10612 18564 11004
rect 18620 10834 18676 11228
rect 18620 10782 18622 10834
rect 18674 10782 18676 10834
rect 18620 10770 18676 10782
rect 18620 10612 18676 10622
rect 18508 10556 18620 10612
rect 17836 10518 17892 10556
rect 17388 10500 17444 10510
rect 17052 9940 17108 9950
rect 17388 9940 17444 10444
rect 18284 10500 18340 10510
rect 18284 10406 18340 10444
rect 17052 9938 17444 9940
rect 17052 9886 17054 9938
rect 17106 9886 17444 9938
rect 17052 9884 17444 9886
rect 17052 9874 17108 9884
rect 16940 9650 16996 9660
rect 17388 9714 17444 9884
rect 17500 9940 17556 9950
rect 17500 9826 17556 9884
rect 17500 9774 17502 9826
rect 17554 9774 17556 9826
rect 17500 9762 17556 9774
rect 18060 9940 18116 9950
rect 18060 9826 18116 9884
rect 18060 9774 18062 9826
rect 18114 9774 18116 9826
rect 18060 9762 18116 9774
rect 17388 9662 17390 9714
rect 17442 9662 17444 9714
rect 17388 9650 17444 9662
rect 17948 9716 18004 9726
rect 17948 9622 18004 9660
rect 17164 9604 17220 9614
rect 17164 9510 17220 9548
rect 17724 9602 17780 9614
rect 17724 9550 17726 9602
rect 17778 9550 17780 9602
rect 16716 9214 16718 9266
rect 16770 9214 16772 9266
rect 16716 9202 16772 9214
rect 17612 9156 17668 9166
rect 16044 9102 16046 9154
rect 16098 9102 16100 9154
rect 16044 9090 16100 9102
rect 17388 9154 17668 9156
rect 17388 9102 17614 9154
rect 17666 9102 17668 9154
rect 17388 9100 17668 9102
rect 16156 9044 16212 9054
rect 16212 8988 16324 9044
rect 16156 8978 16212 8988
rect 15932 8206 15934 8258
rect 15986 8206 15988 8258
rect 15932 8194 15988 8206
rect 15820 8146 15876 8158
rect 15820 8094 15822 8146
rect 15874 8094 15876 8146
rect 15484 7364 15540 7374
rect 15484 7362 15652 7364
rect 15484 7310 15486 7362
rect 15538 7310 15652 7362
rect 15484 7308 15652 7310
rect 15484 7298 15540 7308
rect 15484 6916 15540 6926
rect 15372 6860 15484 6916
rect 15484 6822 15540 6860
rect 13804 6638 13806 6690
rect 13858 6638 13860 6690
rect 13804 6626 13860 6638
rect 13356 5906 13636 5908
rect 13356 5854 13358 5906
rect 13410 5854 13636 5906
rect 13356 5852 13636 5854
rect 15148 6466 15204 6478
rect 15148 6414 15150 6466
rect 15202 6414 15204 6466
rect 13356 5842 13412 5852
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 13468 5012 13524 5852
rect 14028 5796 14084 5806
rect 14028 5794 14308 5796
rect 14028 5742 14030 5794
rect 14082 5742 14308 5794
rect 14028 5740 14308 5742
rect 14028 5730 14084 5740
rect 13468 4946 13524 4956
rect 14028 5012 14084 5022
rect 14028 4338 14084 4956
rect 14252 5010 14308 5740
rect 14476 5124 14532 5134
rect 14476 5030 14532 5068
rect 15148 5124 15204 6414
rect 15148 5058 15204 5068
rect 15484 5124 15540 5134
rect 15596 5124 15652 7308
rect 15820 6580 15876 8094
rect 15932 6916 15988 6926
rect 15988 6860 16212 6916
rect 15932 6850 15988 6860
rect 16044 6580 16100 6590
rect 15820 6578 16100 6580
rect 15820 6526 16046 6578
rect 16098 6526 16100 6578
rect 15820 6524 16100 6526
rect 16044 6020 16100 6524
rect 16044 5954 16100 5964
rect 16156 5794 16212 6860
rect 16268 6690 16324 8988
rect 16380 8818 16436 8830
rect 16380 8766 16382 8818
rect 16434 8766 16436 8818
rect 16380 8372 16436 8766
rect 16380 8306 16436 8316
rect 16716 8372 16772 8382
rect 16716 8258 16772 8316
rect 17388 8370 17444 9100
rect 17612 9090 17668 9100
rect 17724 9044 17780 9550
rect 18396 9604 18452 9614
rect 18396 9602 18564 9604
rect 18396 9550 18398 9602
rect 18450 9550 18564 9602
rect 18396 9548 18564 9550
rect 18396 9538 18452 9548
rect 17724 8978 17780 8988
rect 17948 9042 18004 9054
rect 17948 8990 17950 9042
rect 18002 8990 18004 9042
rect 17836 8372 17892 8382
rect 17388 8318 17390 8370
rect 17442 8318 17444 8370
rect 17388 8306 17444 8318
rect 17724 8316 17836 8372
rect 16716 8206 16718 8258
rect 16770 8206 16772 8258
rect 16716 8194 16772 8206
rect 16268 6638 16270 6690
rect 16322 6638 16324 6690
rect 16268 6626 16324 6638
rect 16156 5742 16158 5794
rect 16210 5742 16212 5794
rect 16156 5730 16212 5742
rect 16604 5796 16660 5806
rect 16940 5796 16996 5806
rect 16604 5794 16772 5796
rect 16604 5742 16606 5794
rect 16658 5742 16772 5794
rect 16604 5740 16772 5742
rect 16604 5730 16660 5740
rect 15540 5068 15652 5124
rect 15484 5058 15540 5068
rect 14252 4958 14254 5010
rect 14306 4958 14308 5010
rect 14252 4946 14308 4958
rect 16716 5012 16772 5740
rect 16828 5012 16884 5022
rect 16716 4956 16828 5012
rect 16828 4946 16884 4956
rect 16940 4788 16996 5740
rect 17500 5684 17556 5694
rect 17500 5682 17668 5684
rect 17500 5630 17502 5682
rect 17554 5630 17668 5682
rect 17500 5628 17668 5630
rect 17500 5618 17556 5628
rect 16828 4732 16996 4788
rect 17164 5012 17220 5022
rect 14700 4452 14756 4462
rect 14700 4358 14756 4396
rect 14028 4286 14030 4338
rect 14082 4286 14084 4338
rect 14028 4274 14084 4286
rect 16828 4226 16884 4732
rect 16828 4174 16830 4226
rect 16882 4174 16884 4226
rect 16828 4162 16884 4174
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17164 3666 17220 4956
rect 17388 4452 17444 4462
rect 17388 4358 17444 4396
rect 17612 4338 17668 5628
rect 17724 5122 17780 8316
rect 17836 8306 17892 8316
rect 17836 7700 17892 7710
rect 17948 7700 18004 8990
rect 17836 7698 18004 7700
rect 17836 7646 17838 7698
rect 17890 7646 18004 7698
rect 17836 7644 18004 7646
rect 18172 8260 18228 8270
rect 17836 7634 17892 7644
rect 18172 7474 18228 8204
rect 18172 7422 18174 7474
rect 18226 7422 18228 7474
rect 18172 7410 18228 7422
rect 18508 6580 18564 9548
rect 18620 9602 18676 10556
rect 18620 9550 18622 9602
rect 18674 9550 18676 9602
rect 18620 9492 18676 9550
rect 18620 9266 18676 9436
rect 18620 9214 18622 9266
rect 18674 9214 18676 9266
rect 18620 9202 18676 9214
rect 18732 9828 18788 9838
rect 18732 8818 18788 9772
rect 18732 8766 18734 8818
rect 18786 8766 18788 8818
rect 18732 8754 18788 8766
rect 18844 7588 18900 11732
rect 19068 10724 19124 13356
rect 19180 11060 19236 13580
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19852 12180 19908 12190
rect 19852 11732 19908 12124
rect 19852 11666 19908 11676
rect 20188 11508 20244 11518
rect 19180 10994 19236 11004
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 10836 20244 11452
rect 19964 10780 20244 10836
rect 19068 10668 19348 10724
rect 18956 10612 19012 10622
rect 18956 10518 19012 10556
rect 19292 9826 19348 10668
rect 19628 10612 19684 10622
rect 19628 10518 19684 10556
rect 19964 10610 20020 10780
rect 19964 10558 19966 10610
rect 20018 10558 20020 10610
rect 19964 10546 20020 10558
rect 20524 10722 20580 13804
rect 20636 13794 20692 13804
rect 20860 13746 20916 14364
rect 21308 13970 21364 15260
rect 21420 14756 21476 14766
rect 21532 14756 21588 16830
rect 21420 14754 21588 14756
rect 21420 14702 21422 14754
rect 21474 14702 21588 14754
rect 21420 14700 21588 14702
rect 21756 15204 21812 15214
rect 21756 14754 21812 15148
rect 21756 14702 21758 14754
rect 21810 14702 21812 14754
rect 21420 14690 21476 14700
rect 21756 14690 21812 14702
rect 21980 14644 22036 17052
rect 22092 17042 22148 17052
rect 22428 17220 22484 17948
rect 22204 16884 22260 16894
rect 22428 16884 22484 17164
rect 22540 16994 22596 18396
rect 22540 16942 22542 16994
rect 22594 16942 22596 16994
rect 22540 16930 22596 16942
rect 22204 16882 22484 16884
rect 22204 16830 22206 16882
rect 22258 16830 22484 16882
rect 22204 16828 22484 16830
rect 22204 16818 22260 16828
rect 22652 16772 22708 18620
rect 22988 18620 23156 18676
rect 22988 18004 23044 18620
rect 23324 18562 23380 18574
rect 23324 18510 23326 18562
rect 23378 18510 23380 18562
rect 22988 17938 23044 17948
rect 23100 18450 23156 18462
rect 23100 18398 23102 18450
rect 23154 18398 23156 18450
rect 23100 17332 23156 18398
rect 23324 17556 23380 18510
rect 23324 17490 23380 17500
rect 23660 18562 23716 18574
rect 23660 18510 23662 18562
rect 23714 18510 23716 18562
rect 23660 17332 23716 18510
rect 23884 17666 23940 19068
rect 23996 18450 24052 18462
rect 23996 18398 23998 18450
rect 24050 18398 24052 18450
rect 23996 18116 24052 18398
rect 23996 18050 24052 18060
rect 23884 17614 23886 17666
rect 23938 17614 23940 17666
rect 23100 17276 23716 17332
rect 23772 17556 23828 17566
rect 22428 16716 22708 16772
rect 22764 17106 22820 17118
rect 22764 17054 22766 17106
rect 22818 17054 22820 17106
rect 22092 16658 22148 16670
rect 22092 16606 22094 16658
rect 22146 16606 22148 16658
rect 22092 15148 22148 16606
rect 22092 15092 22260 15148
rect 21980 14588 22148 14644
rect 21980 14420 22036 14430
rect 21980 14326 22036 14364
rect 21308 13918 21310 13970
rect 21362 13918 21364 13970
rect 21308 13906 21364 13918
rect 21756 13860 21812 13870
rect 20860 13694 20862 13746
rect 20914 13694 20916 13746
rect 20860 13682 20916 13694
rect 21644 13804 21756 13860
rect 21532 12964 21588 12974
rect 21420 12962 21588 12964
rect 21420 12910 21534 12962
rect 21586 12910 21588 12962
rect 21420 12908 21588 12910
rect 21308 12740 21364 12750
rect 20636 12738 21364 12740
rect 20636 12686 21310 12738
rect 21362 12686 21364 12738
rect 20636 12684 21364 12686
rect 20636 12290 20692 12684
rect 21308 12674 21364 12684
rect 20636 12238 20638 12290
rect 20690 12238 20692 12290
rect 20636 12226 20692 12238
rect 20524 10670 20526 10722
rect 20578 10670 20580 10722
rect 19292 9774 19294 9826
rect 19346 9774 19348 9826
rect 19180 9716 19236 9726
rect 19180 9622 19236 9660
rect 18956 9602 19012 9614
rect 18956 9550 18958 9602
rect 19010 9550 19012 9602
rect 18956 9156 19012 9550
rect 19292 9604 19348 9774
rect 19628 10052 19684 10062
rect 19292 9538 19348 9548
rect 19516 9716 19572 9726
rect 19516 9492 19572 9660
rect 19516 9426 19572 9436
rect 18956 9100 19236 9156
rect 19180 9044 19236 9100
rect 19628 9154 19684 9996
rect 20524 10052 20580 10670
rect 20524 9986 20580 9996
rect 20636 11732 20692 11742
rect 20636 11506 20692 11676
rect 21420 11618 21476 12908
rect 21532 12898 21588 12908
rect 21420 11566 21422 11618
rect 21474 11566 21476 11618
rect 21420 11554 21476 11566
rect 20636 11454 20638 11506
rect 20690 11454 20692 11506
rect 19740 9716 19796 9726
rect 19740 9622 19796 9660
rect 20188 9604 20244 9614
rect 20188 9510 20244 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19628 9102 19630 9154
rect 19682 9102 19684 9154
rect 19628 9090 19684 9102
rect 19404 9044 19460 9054
rect 19180 9042 19460 9044
rect 19180 8990 19406 9042
rect 19458 8990 19460 9042
rect 19180 8988 19460 8990
rect 19068 8930 19124 8942
rect 19068 8878 19070 8930
rect 19122 8878 19124 8930
rect 19068 8818 19124 8878
rect 19068 8766 19070 8818
rect 19122 8766 19124 8818
rect 19068 8754 19124 8766
rect 18844 7494 18900 7532
rect 18956 7476 19012 7486
rect 19292 7476 19348 8988
rect 19404 8978 19460 8988
rect 19964 8820 20020 8830
rect 18956 7474 19348 7476
rect 18956 7422 18958 7474
rect 19010 7422 19348 7474
rect 18956 7420 19348 7422
rect 19404 8372 19460 8382
rect 19404 7474 19460 8316
rect 19516 8370 19572 8382
rect 19516 8318 19518 8370
rect 19570 8318 19572 8370
rect 19516 8260 19572 8318
rect 19516 8194 19572 8204
rect 19964 8258 20020 8764
rect 20188 8818 20244 8830
rect 20188 8766 20190 8818
rect 20242 8766 20244 8818
rect 20188 8596 20244 8766
rect 20524 8820 20580 8830
rect 20524 8726 20580 8764
rect 20188 8540 20468 8596
rect 19964 8206 19966 8258
rect 20018 8206 20020 8258
rect 19964 8194 20020 8206
rect 20188 8034 20244 8046
rect 20188 7982 20190 8034
rect 20242 7982 20244 8034
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20188 7586 20244 7982
rect 20188 7534 20190 7586
rect 20242 7534 20244 7586
rect 20188 7522 20244 7534
rect 19404 7422 19406 7474
rect 19458 7422 19460 7474
rect 18956 7410 19012 7420
rect 19404 7410 19460 7422
rect 20412 7364 20468 8540
rect 20636 8372 20692 11454
rect 21644 11508 21700 13804
rect 21756 13794 21812 13804
rect 21756 13636 21812 13646
rect 21756 13634 21924 13636
rect 21756 13582 21758 13634
rect 21810 13582 21924 13634
rect 21756 13580 21924 13582
rect 21756 13570 21812 13580
rect 21756 12068 21812 12078
rect 21756 11618 21812 12012
rect 21756 11566 21758 11618
rect 21810 11566 21812 11618
rect 21756 11554 21812 11566
rect 21644 11442 21700 11452
rect 20748 10612 20804 10622
rect 20748 10518 20804 10556
rect 21196 10052 21252 10062
rect 21196 9266 21252 9996
rect 21868 9716 21924 13580
rect 21980 11396 22036 11406
rect 21980 11282 22036 11340
rect 21980 11230 21982 11282
rect 22034 11230 22036 11282
rect 21980 10612 22036 11230
rect 21980 10546 22036 10556
rect 22092 10724 22148 14588
rect 22204 14420 22260 15092
rect 22204 14354 22260 14364
rect 22316 14418 22372 14430
rect 22316 14366 22318 14418
rect 22370 14366 22372 14418
rect 22316 11284 22372 14366
rect 22092 10610 22148 10668
rect 22092 10558 22094 10610
rect 22146 10558 22148 10610
rect 22092 10546 22148 10558
rect 22204 11282 22372 11284
rect 22204 11230 22318 11282
rect 22370 11230 22372 11282
rect 22204 11228 22372 11230
rect 22204 10500 22260 11228
rect 22316 11218 22372 11228
rect 22316 10724 22372 10734
rect 22316 10630 22372 10668
rect 22204 10444 22372 10500
rect 22092 9828 22148 9838
rect 22092 9734 22148 9772
rect 21868 9660 22036 9716
rect 21196 9214 21198 9266
rect 21250 9214 21252 9266
rect 21196 9202 21252 9214
rect 21644 9602 21700 9614
rect 21644 9550 21646 9602
rect 21698 9550 21700 9602
rect 21532 9044 21588 9054
rect 21644 9044 21700 9550
rect 21532 9042 21700 9044
rect 21532 8990 21534 9042
rect 21586 8990 21700 9042
rect 21532 8988 21700 8990
rect 21868 9156 21924 9166
rect 21532 8932 21588 8988
rect 21532 8866 21588 8876
rect 20636 8278 20692 8316
rect 20412 7298 20468 7308
rect 18284 6524 18564 6580
rect 21756 6692 21812 6702
rect 18284 5906 18340 6524
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 18396 6020 18452 6030
rect 19068 6020 19124 6030
rect 18396 5926 18452 5964
rect 18508 6018 19124 6020
rect 18508 5966 19070 6018
rect 19122 5966 19124 6018
rect 18508 5964 19124 5966
rect 18284 5854 18286 5906
rect 18338 5854 18340 5906
rect 17836 5796 17892 5806
rect 17836 5702 17892 5740
rect 17724 5070 17726 5122
rect 17778 5070 17780 5122
rect 17724 5058 17780 5070
rect 18284 5124 18340 5854
rect 18508 5234 18564 5964
rect 19068 5954 19124 5964
rect 20636 6020 20692 6030
rect 21756 6020 21812 6636
rect 20636 6018 21252 6020
rect 20636 5966 20638 6018
rect 20690 5966 21252 6018
rect 20636 5964 21252 5966
rect 20636 5954 20692 5964
rect 19404 5908 19460 5918
rect 19404 5906 19684 5908
rect 19404 5854 19406 5906
rect 19458 5854 19684 5906
rect 19404 5852 19684 5854
rect 19404 5842 19460 5852
rect 18508 5182 18510 5234
rect 18562 5182 18564 5234
rect 18508 5170 18564 5182
rect 19292 5348 19348 5358
rect 18284 5068 18452 5124
rect 18396 5012 18452 5068
rect 18396 4956 18564 5012
rect 17612 4286 17614 4338
rect 17666 4286 17668 4338
rect 17612 4274 17668 4286
rect 18508 4338 18564 4956
rect 18732 4452 18788 4462
rect 18732 4358 18788 4396
rect 18508 4286 18510 4338
rect 18562 4286 18564 4338
rect 18508 4274 18564 4286
rect 19292 4338 19348 5292
rect 19628 4562 19684 5852
rect 20412 5906 20468 5918
rect 20412 5854 20414 5906
rect 20466 5854 20468 5906
rect 20412 5796 20468 5854
rect 21084 5796 21140 5806
rect 20412 5794 21140 5796
rect 20412 5742 21086 5794
rect 21138 5742 21140 5794
rect 20412 5740 21140 5742
rect 21084 5730 21140 5740
rect 20636 5348 20692 5358
rect 20636 5234 20692 5292
rect 20636 5182 20638 5234
rect 20690 5182 20692 5234
rect 20636 5170 20692 5182
rect 20412 5012 20468 5022
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4510 19630 4562
rect 19682 4510 19684 4562
rect 19628 4498 19684 4510
rect 19292 4286 19294 4338
rect 19346 4286 19348 4338
rect 19292 4274 19348 4286
rect 20412 4338 20468 4956
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20412 4274 20468 4286
rect 20972 5012 21028 5022
rect 17164 3614 17166 3666
rect 17218 3614 17220 3666
rect 17164 3602 17220 3614
rect 20972 3666 21028 4956
rect 21084 4452 21140 4462
rect 21196 4452 21252 5964
rect 21420 5684 21476 5694
rect 21420 5590 21476 5628
rect 21756 5010 21812 5964
rect 21756 4958 21758 5010
rect 21810 4958 21812 5010
rect 21756 4946 21812 4958
rect 21868 6020 21924 9100
rect 21980 8148 22036 9660
rect 22204 9042 22260 9054
rect 22204 8990 22206 9042
rect 22258 8990 22260 9042
rect 22204 8932 22260 8990
rect 22204 8866 22260 8876
rect 21980 8054 22036 8092
rect 22316 8034 22372 10444
rect 22428 10388 22484 16716
rect 22764 16436 22820 17054
rect 22652 16380 22820 16436
rect 22876 16882 22932 16894
rect 22876 16830 22878 16882
rect 22930 16830 22932 16882
rect 22876 16436 22932 16830
rect 23324 16882 23380 16894
rect 23324 16830 23326 16882
rect 23378 16830 23380 16882
rect 22988 16772 23044 16782
rect 22988 16678 23044 16716
rect 23324 16660 23380 16830
rect 23324 16594 23380 16604
rect 22652 15988 22708 16380
rect 22876 16370 22932 16380
rect 22764 16212 22820 16222
rect 22764 16118 22820 16156
rect 23324 16212 23380 16222
rect 22652 15932 23044 15988
rect 22876 15204 22932 15242
rect 22876 15138 22932 15148
rect 22988 14308 23044 15932
rect 23324 15538 23380 16156
rect 23324 15486 23326 15538
rect 23378 15486 23380 15538
rect 23324 15474 23380 15486
rect 22876 14252 23044 14308
rect 22540 13748 22596 13758
rect 22540 13654 22596 13692
rect 22764 13746 22820 13758
rect 22764 13694 22766 13746
rect 22818 13694 22820 13746
rect 22540 12738 22596 12750
rect 22540 12686 22542 12738
rect 22594 12686 22596 12738
rect 22540 11732 22596 12686
rect 22764 12404 22820 13694
rect 22876 13748 22932 14252
rect 23324 13972 23380 13982
rect 23324 13878 23380 13916
rect 22988 13748 23044 13758
rect 22876 13746 23044 13748
rect 22876 13694 22990 13746
rect 23042 13694 23044 13746
rect 22876 13692 23044 13694
rect 22988 13682 23044 13692
rect 23324 13748 23380 13758
rect 23324 12850 23380 13692
rect 23324 12798 23326 12850
rect 23378 12798 23380 12850
rect 23324 12786 23380 12798
rect 22988 12740 23044 12750
rect 22988 12646 23044 12684
rect 22764 12338 22820 12348
rect 22988 12516 23044 12526
rect 22764 12068 22820 12078
rect 22764 11974 22820 12012
rect 22540 11666 22596 11676
rect 22988 11396 23044 12460
rect 23212 12404 23268 12414
rect 23212 12310 23268 12348
rect 23436 12178 23492 17276
rect 23660 16996 23716 17006
rect 23660 16882 23716 16940
rect 23660 16830 23662 16882
rect 23714 16830 23716 16882
rect 23660 16818 23716 16830
rect 23772 15148 23828 17500
rect 23884 16884 23940 17614
rect 23884 16100 23940 16828
rect 24108 16882 24164 19740
rect 24444 19124 24500 19134
rect 24444 19030 24500 19068
rect 24332 18450 24388 18462
rect 24332 18398 24334 18450
rect 24386 18398 24388 18450
rect 24332 18116 24388 18398
rect 24332 18050 24388 18060
rect 24444 17554 24500 17566
rect 24444 17502 24446 17554
rect 24498 17502 24500 17554
rect 24444 17108 24500 17502
rect 24556 17332 24612 25564
rect 24668 25284 24724 26126
rect 24668 23716 24724 25228
rect 25340 26290 25396 26302
rect 25340 26238 25342 26290
rect 25394 26238 25396 26290
rect 25340 25284 25396 26238
rect 25340 25190 25396 25228
rect 25788 25506 25844 25518
rect 25788 25454 25790 25506
rect 25842 25454 25844 25506
rect 25788 25284 25844 25454
rect 25788 25218 25844 25228
rect 26460 25394 26516 25406
rect 26460 25342 26462 25394
rect 26514 25342 26516 25394
rect 26460 24052 26516 25342
rect 26908 24610 26964 24622
rect 26908 24558 26910 24610
rect 26962 24558 26964 24610
rect 26460 23986 26516 23996
rect 26796 24498 26852 24510
rect 26796 24446 26798 24498
rect 26850 24446 26852 24498
rect 24668 23154 24724 23660
rect 24780 23826 24836 23838
rect 24780 23774 24782 23826
rect 24834 23774 24836 23826
rect 24780 23380 24836 23774
rect 24780 23314 24836 23324
rect 25564 23380 25620 23390
rect 25564 23286 25620 23324
rect 25228 23156 25284 23166
rect 24668 23102 24670 23154
rect 24722 23102 24724 23154
rect 24668 22148 24724 23102
rect 25116 23154 25284 23156
rect 25116 23102 25230 23154
rect 25282 23102 25284 23154
rect 25116 23100 25284 23102
rect 24780 22596 24836 22606
rect 24780 22502 24836 22540
rect 25116 22594 25172 23100
rect 25228 23090 25284 23100
rect 25564 23154 25620 23166
rect 25564 23102 25566 23154
rect 25618 23102 25620 23154
rect 25116 22542 25118 22594
rect 25170 22542 25172 22594
rect 25116 22530 25172 22542
rect 25452 22484 25508 22494
rect 25116 22372 25172 22382
rect 25116 22278 25172 22316
rect 25452 22148 25508 22428
rect 25564 22372 25620 23102
rect 25900 23156 25956 23166
rect 26124 23156 26180 23166
rect 25900 23154 26180 23156
rect 25900 23102 25902 23154
rect 25954 23102 26126 23154
rect 26178 23102 26180 23154
rect 25900 23100 26180 23102
rect 25900 22596 25956 23100
rect 26124 23090 26180 23100
rect 26460 23156 26516 23194
rect 26460 23090 26516 23100
rect 26236 23044 26292 23054
rect 26236 22950 26292 22988
rect 25900 22530 25956 22540
rect 26796 22372 26852 24446
rect 26908 24050 26964 24558
rect 26908 23998 26910 24050
rect 26962 23998 26964 24050
rect 26908 23986 26964 23998
rect 27020 23828 27076 26852
rect 28140 26178 28196 26190
rect 28140 26126 28142 26178
rect 28194 26126 28196 26178
rect 27804 24052 27860 24062
rect 25564 22316 26852 22372
rect 25564 22148 25620 22158
rect 25452 22092 25564 22148
rect 24668 22082 24724 22092
rect 24668 21924 24724 21934
rect 24668 21586 24724 21868
rect 24668 21534 24670 21586
rect 24722 21534 24724 21586
rect 24668 21522 24724 21534
rect 25340 21476 25396 21486
rect 25564 21476 25620 22092
rect 25228 21474 25732 21476
rect 25228 21422 25342 21474
rect 25394 21422 25732 21474
rect 25228 21420 25732 21422
rect 24668 21362 24724 21374
rect 24668 21310 24670 21362
rect 24722 21310 24724 21362
rect 24668 20130 24724 21310
rect 24668 20078 24670 20130
rect 24722 20078 24724 20130
rect 24668 20066 24724 20078
rect 25116 19348 25172 19358
rect 25228 19348 25284 21420
rect 25340 21410 25396 21420
rect 25340 20916 25396 20926
rect 25340 20914 25620 20916
rect 25340 20862 25342 20914
rect 25394 20862 25620 20914
rect 25340 20860 25620 20862
rect 25340 20850 25396 20860
rect 25564 20130 25620 20860
rect 25676 20802 25732 21420
rect 25676 20750 25678 20802
rect 25730 20750 25732 20802
rect 25676 20738 25732 20750
rect 25564 20078 25566 20130
rect 25618 20078 25620 20130
rect 25564 20066 25620 20078
rect 26460 20690 26516 20702
rect 26460 20638 26462 20690
rect 26514 20638 26516 20690
rect 26460 20132 26516 20638
rect 26460 20066 26516 20076
rect 25452 20020 25508 20030
rect 25172 19292 25284 19348
rect 25340 19964 25452 20020
rect 25116 19282 25172 19292
rect 24668 18564 24724 18574
rect 24668 18470 24724 18508
rect 25228 18564 25284 18574
rect 25340 18564 25396 19964
rect 25452 19926 25508 19964
rect 26348 19908 26404 19918
rect 26348 19814 26404 19852
rect 26684 19906 26740 19918
rect 26684 19854 26686 19906
rect 26738 19854 26740 19906
rect 26124 19012 26180 19022
rect 26124 18918 26180 18956
rect 26684 19012 26740 19854
rect 26684 18946 26740 18956
rect 26348 18676 26404 18686
rect 26348 18674 26740 18676
rect 26348 18622 26350 18674
rect 26402 18622 26740 18674
rect 26348 18620 26740 18622
rect 26348 18610 26404 18620
rect 25228 18562 25396 18564
rect 25228 18510 25230 18562
rect 25282 18510 25396 18562
rect 25228 18508 25396 18510
rect 25228 18498 25284 18508
rect 25564 18450 25620 18462
rect 25564 18398 25566 18450
rect 25618 18398 25620 18450
rect 25340 18338 25396 18350
rect 25340 18286 25342 18338
rect 25394 18286 25396 18338
rect 24780 18228 24836 18238
rect 24780 17890 24836 18172
rect 24780 17838 24782 17890
rect 24834 17838 24836 17890
rect 24780 17826 24836 17838
rect 24780 17668 24836 17678
rect 24780 17666 24948 17668
rect 24780 17614 24782 17666
rect 24834 17614 24948 17666
rect 24780 17612 24948 17614
rect 24780 17602 24836 17612
rect 24556 17266 24612 17276
rect 24892 17444 24948 17612
rect 25228 17444 25284 17454
rect 24892 17442 25284 17444
rect 24892 17390 25230 17442
rect 25282 17390 25284 17442
rect 24892 17388 25284 17390
rect 24444 17042 24500 17052
rect 24108 16830 24110 16882
rect 24162 16830 24164 16882
rect 24108 16818 24164 16830
rect 24332 16882 24388 16894
rect 24332 16830 24334 16882
rect 24386 16830 24388 16882
rect 23996 16660 24052 16670
rect 24052 16604 24276 16660
rect 23996 16566 24052 16604
rect 24220 16100 24276 16604
rect 23884 16098 24164 16100
rect 23884 16046 23886 16098
rect 23938 16046 24164 16098
rect 23884 16044 24164 16046
rect 23884 16034 23940 16044
rect 24108 15540 24164 16044
rect 24220 16034 24276 16044
rect 24220 15540 24276 15550
rect 24108 15538 24276 15540
rect 24108 15486 24222 15538
rect 24274 15486 24276 15538
rect 24108 15484 24276 15486
rect 24220 15474 24276 15484
rect 24220 15316 24276 15326
rect 23772 15092 24164 15148
rect 23772 13860 23828 15092
rect 24108 14530 24164 15092
rect 24108 14478 24110 14530
rect 24162 14478 24164 14530
rect 24108 14466 24164 14478
rect 23884 14420 23940 14430
rect 23884 14326 23940 14364
rect 23996 14306 24052 14318
rect 23996 14254 23998 14306
rect 24050 14254 24052 14306
rect 23884 13860 23940 13870
rect 23772 13858 23940 13860
rect 23772 13806 23886 13858
rect 23938 13806 23940 13858
rect 23772 13804 23940 13806
rect 23884 13794 23940 13804
rect 23660 13748 23716 13758
rect 23660 13746 23828 13748
rect 23660 13694 23662 13746
rect 23714 13694 23828 13746
rect 23660 13692 23828 13694
rect 23660 13682 23716 13692
rect 23548 12962 23604 12974
rect 23548 12910 23550 12962
rect 23602 12910 23604 12962
rect 23548 12740 23604 12910
rect 23548 12674 23604 12684
rect 23436 12126 23438 12178
rect 23490 12126 23492 12178
rect 23436 11956 23492 12126
rect 23436 11890 23492 11900
rect 22652 11394 23044 11396
rect 22652 11342 22990 11394
rect 23042 11342 23044 11394
rect 22652 11340 23044 11342
rect 22428 10332 22596 10388
rect 22428 10164 22484 10174
rect 22428 9938 22484 10108
rect 22428 9886 22430 9938
rect 22482 9886 22484 9938
rect 22428 9874 22484 9886
rect 22540 9828 22596 10332
rect 22652 10052 22708 11340
rect 22988 11330 23044 11340
rect 23100 11618 23156 11630
rect 23100 11566 23102 11618
rect 23154 11566 23156 11618
rect 23100 11396 23156 11566
rect 23100 11330 23156 11340
rect 23100 11170 23156 11182
rect 23100 11118 23102 11170
rect 23154 11118 23156 11170
rect 22764 10724 22820 10734
rect 22764 10500 22820 10668
rect 23100 10500 23156 11118
rect 23212 11172 23268 11182
rect 23548 11172 23604 11182
rect 23268 11170 23604 11172
rect 23268 11118 23550 11170
rect 23602 11118 23604 11170
rect 23268 11116 23604 11118
rect 23212 10612 23268 11116
rect 23548 11106 23604 11116
rect 23212 10518 23268 10556
rect 23548 10836 23604 10846
rect 22764 10498 23156 10500
rect 22764 10446 22766 10498
rect 22818 10446 23156 10498
rect 22764 10444 23156 10446
rect 23548 10498 23604 10780
rect 23548 10446 23550 10498
rect 23602 10446 23604 10498
rect 22764 10434 22820 10444
rect 22652 9986 22708 9996
rect 22652 9828 22708 9838
rect 22596 9826 22820 9828
rect 22596 9774 22654 9826
rect 22706 9774 22820 9826
rect 22596 9772 22820 9774
rect 22540 9734 22596 9772
rect 22652 9762 22708 9772
rect 22764 9268 22820 9772
rect 22652 9154 22708 9166
rect 22652 9102 22654 9154
rect 22706 9102 22708 9154
rect 22316 7982 22318 8034
rect 22370 7982 22372 8034
rect 22316 7588 22372 7982
rect 22316 7522 22372 7532
rect 22428 9042 22484 9054
rect 22428 8990 22430 9042
rect 22482 8990 22484 9042
rect 22316 7364 22372 7374
rect 22316 7270 22372 7308
rect 21980 6020 22036 6030
rect 21868 6018 22036 6020
rect 21868 5966 21982 6018
rect 22034 5966 22036 6018
rect 21868 5964 22036 5966
rect 21084 4450 21252 4452
rect 21084 4398 21086 4450
rect 21138 4398 21252 4450
rect 21084 4396 21252 4398
rect 21868 4452 21924 5964
rect 21980 5954 22036 5964
rect 22204 5908 22260 5918
rect 22428 5908 22484 8990
rect 22652 8708 22708 9102
rect 22764 9154 22820 9212
rect 22764 9102 22766 9154
rect 22818 9102 22820 9154
rect 22764 9090 22820 9102
rect 22876 9156 22932 10444
rect 23548 10434 23604 10446
rect 22988 9716 23044 9726
rect 22988 9622 23044 9660
rect 23660 9268 23716 9278
rect 23660 9174 23716 9212
rect 22988 9156 23044 9166
rect 22876 9100 22988 9156
rect 22988 9090 23044 9100
rect 23212 8932 23268 8942
rect 23212 8838 23268 8876
rect 22652 8652 23268 8708
rect 22540 8372 22596 8382
rect 22540 6690 22596 8316
rect 23212 8148 23268 8652
rect 23772 8596 23828 13692
rect 23884 13636 23940 13646
rect 23996 13636 24052 14254
rect 24108 13972 24164 13982
rect 24220 13972 24276 15260
rect 24332 14754 24388 16830
rect 24444 16882 24500 16894
rect 24444 16830 24446 16882
rect 24498 16830 24500 16882
rect 24444 16324 24500 16830
rect 24668 16436 24724 16446
rect 24724 16380 24836 16436
rect 24668 16370 24724 16380
rect 24444 16258 24500 16268
rect 24780 16212 24836 16380
rect 24444 16100 24500 16110
rect 24444 16006 24500 16044
rect 24556 16100 24612 16110
rect 24556 16098 24724 16100
rect 24556 16046 24558 16098
rect 24610 16046 24724 16098
rect 24556 16044 24724 16046
rect 24556 16034 24612 16044
rect 24332 14702 24334 14754
rect 24386 14702 24388 14754
rect 24332 14690 24388 14702
rect 24556 15874 24612 15886
rect 24556 15822 24558 15874
rect 24610 15822 24612 15874
rect 24444 14530 24500 14542
rect 24444 14478 24446 14530
rect 24498 14478 24500 14530
rect 24108 13970 24276 13972
rect 24108 13918 24110 13970
rect 24162 13918 24276 13970
rect 24108 13916 24276 13918
rect 24332 14420 24388 14430
rect 24108 13906 24164 13916
rect 23996 13580 24164 13636
rect 23884 12404 23940 13580
rect 23996 13412 24052 13422
rect 23996 12962 24052 13356
rect 24108 13300 24164 13580
rect 24220 13524 24276 13534
rect 24220 13430 24276 13468
rect 24108 13234 24164 13244
rect 23996 12910 23998 12962
rect 24050 12910 24052 12962
rect 23996 12898 24052 12910
rect 24220 12850 24276 12862
rect 24220 12798 24222 12850
rect 24274 12798 24276 12850
rect 23996 12404 24052 12414
rect 23884 12402 24052 12404
rect 23884 12350 23998 12402
rect 24050 12350 24052 12402
rect 23884 12348 24052 12350
rect 23996 12338 24052 12348
rect 24220 12404 24276 12798
rect 24332 12404 24388 14364
rect 24444 13748 24500 14478
rect 24444 12964 24500 13692
rect 24556 13524 24612 15822
rect 24556 13458 24612 13468
rect 24556 13188 24612 13198
rect 24556 13094 24612 13132
rect 24556 12964 24612 12974
rect 24444 12962 24612 12964
rect 24444 12910 24558 12962
rect 24610 12910 24612 12962
rect 24444 12908 24612 12910
rect 24556 12898 24612 12908
rect 24332 12348 24612 12404
rect 24220 12292 24276 12348
rect 24220 12290 24388 12292
rect 24220 12238 24222 12290
rect 24274 12238 24388 12290
rect 24220 12236 24388 12238
rect 24220 12226 24276 12236
rect 23884 12178 23940 12190
rect 23884 12126 23886 12178
rect 23938 12126 23940 12178
rect 23884 11844 23940 12126
rect 24332 11956 24388 12236
rect 24444 12180 24500 12190
rect 24444 12086 24500 12124
rect 24332 11900 24500 11956
rect 23884 11778 23940 11788
rect 23884 11508 23940 11518
rect 23884 11396 23940 11452
rect 24332 11396 24388 11406
rect 23884 11394 24164 11396
rect 23884 11342 23886 11394
rect 23938 11342 24164 11394
rect 23884 11340 24164 11342
rect 23884 11330 23940 11340
rect 24108 10836 24164 11340
rect 24332 11302 24388 11340
rect 24444 11394 24500 11900
rect 24444 11342 24446 11394
rect 24498 11342 24500 11394
rect 24444 11330 24500 11342
rect 24220 11284 24276 11294
rect 24220 11190 24276 11228
rect 24220 10836 24276 10846
rect 24108 10834 24276 10836
rect 24108 10782 24222 10834
rect 24274 10782 24276 10834
rect 24108 10780 24276 10782
rect 24220 10770 24276 10780
rect 24332 10612 24388 10622
rect 23660 8540 23828 8596
rect 23996 9938 24052 9950
rect 23996 9886 23998 9938
rect 24050 9886 24052 9938
rect 23548 8372 23604 8382
rect 23548 8278 23604 8316
rect 23212 8082 23268 8092
rect 22652 8036 22708 8046
rect 23100 8036 23156 8046
rect 22652 8034 23156 8036
rect 22652 7982 22654 8034
rect 22706 7982 23102 8034
rect 23154 7982 23156 8034
rect 22652 7980 23156 7982
rect 22652 7970 22708 7980
rect 22540 6638 22542 6690
rect 22594 6638 22596 6690
rect 22540 6356 22596 6638
rect 22652 7586 22708 7598
rect 22652 7534 22654 7586
rect 22706 7534 22708 7586
rect 22652 6692 22708 7534
rect 22652 6626 22708 6636
rect 22988 7476 23044 7486
rect 23100 7476 23156 7980
rect 23548 7586 23604 7598
rect 23548 7534 23550 7586
rect 23602 7534 23604 7586
rect 23436 7476 23492 7486
rect 22988 7474 23156 7476
rect 22988 7422 22990 7474
rect 23042 7422 23156 7474
rect 22988 7420 23156 7422
rect 23324 7420 23436 7476
rect 22988 6580 23044 7420
rect 23212 6580 23268 6590
rect 22988 6524 23212 6580
rect 23212 6486 23268 6524
rect 22540 6290 22596 6300
rect 23212 6356 23268 6366
rect 22092 5906 22484 5908
rect 22092 5854 22206 5906
rect 22258 5854 22484 5906
rect 22092 5852 22484 5854
rect 22988 6018 23044 6030
rect 22988 5966 22990 6018
rect 23042 5966 23044 6018
rect 22092 5010 22148 5852
rect 22204 5842 22260 5852
rect 22988 5684 23044 5966
rect 22316 5236 22372 5246
rect 22316 5142 22372 5180
rect 22092 4958 22094 5010
rect 22146 4958 22148 5010
rect 22092 4946 22148 4958
rect 22876 5012 22932 5022
rect 22652 4900 22708 4910
rect 22652 4806 22708 4844
rect 21084 4386 21140 4396
rect 21868 4386 21924 4396
rect 20972 3614 20974 3666
rect 21026 3614 21028 3666
rect 20972 3602 21028 3614
rect 22876 3666 22932 4956
rect 22988 4228 23044 5628
rect 23212 5122 23268 6300
rect 23324 6018 23380 7420
rect 23436 7382 23492 7420
rect 23548 7364 23604 7534
rect 23548 7298 23604 7308
rect 23660 6692 23716 8540
rect 23772 8372 23828 8382
rect 23772 8260 23828 8316
rect 23884 8260 23940 8270
rect 23772 8258 23940 8260
rect 23772 8206 23886 8258
rect 23938 8206 23940 8258
rect 23772 8204 23940 8206
rect 23884 6804 23940 8204
rect 23996 7476 24052 9886
rect 24332 9826 24388 10556
rect 24332 9774 24334 9826
rect 24386 9774 24388 9826
rect 24332 9762 24388 9774
rect 24556 7698 24612 12348
rect 24668 10500 24724 16044
rect 24780 16098 24836 16156
rect 24780 16046 24782 16098
rect 24834 16046 24836 16098
rect 24780 16034 24836 16046
rect 24892 15148 24948 17388
rect 25228 17378 25284 17388
rect 25340 17108 25396 18286
rect 25564 18004 25620 18398
rect 26012 18450 26068 18462
rect 26012 18398 26014 18450
rect 26066 18398 26068 18450
rect 25676 18228 25732 18238
rect 25676 18134 25732 18172
rect 26012 18116 26068 18398
rect 26572 18450 26628 18462
rect 26572 18398 26574 18450
rect 26626 18398 26628 18450
rect 26460 18338 26516 18350
rect 26460 18286 26462 18338
rect 26514 18286 26516 18338
rect 26348 18228 26404 18238
rect 26012 18050 26068 18060
rect 26236 18172 26348 18228
rect 25564 17938 25620 17948
rect 25900 17668 25956 17678
rect 25900 17574 25956 17612
rect 26236 17554 26292 18172
rect 26348 18162 26404 18172
rect 26236 17502 26238 17554
rect 26290 17502 26292 17554
rect 26236 17490 26292 17502
rect 26348 17556 26404 17566
rect 26348 17462 26404 17500
rect 25564 17442 25620 17454
rect 25564 17390 25566 17442
rect 25618 17390 25620 17442
rect 25564 17332 25620 17390
rect 25564 17266 25620 17276
rect 25788 17444 25844 17454
rect 25340 17052 25732 17108
rect 25228 16884 25284 16894
rect 25116 16882 25284 16884
rect 25116 16830 25230 16882
rect 25282 16830 25284 16882
rect 25116 16828 25284 16830
rect 25004 16772 25060 16782
rect 25004 16098 25060 16716
rect 25004 16046 25006 16098
rect 25058 16046 25060 16098
rect 25004 16034 25060 16046
rect 24892 15092 25060 15148
rect 24780 12852 24836 12862
rect 24780 12738 24836 12796
rect 24780 12686 24782 12738
rect 24834 12686 24836 12738
rect 24780 12674 24836 12686
rect 25004 12740 25060 15092
rect 25116 13860 25172 16828
rect 25228 16818 25284 16828
rect 25452 16884 25508 16894
rect 25452 16790 25508 16828
rect 25340 16770 25396 16782
rect 25340 16718 25342 16770
rect 25394 16718 25396 16770
rect 25340 15428 25396 16718
rect 25340 15372 25508 15428
rect 25116 13794 25172 13804
rect 25228 15314 25284 15326
rect 25228 15262 25230 15314
rect 25282 15262 25284 15314
rect 25228 13636 25284 15262
rect 25452 15314 25508 15372
rect 25452 15262 25454 15314
rect 25506 15262 25508 15314
rect 25452 15250 25508 15262
rect 25340 15202 25396 15214
rect 25340 15150 25342 15202
rect 25394 15150 25396 15202
rect 25340 15148 25396 15150
rect 25676 15148 25732 17052
rect 25788 16882 25844 17388
rect 25788 16830 25790 16882
rect 25842 16830 25844 16882
rect 25788 16818 25844 16830
rect 26012 17442 26068 17454
rect 26012 17390 26014 17442
rect 26066 17390 26068 17442
rect 26012 16882 26068 17390
rect 26012 16830 26014 16882
rect 26066 16830 26068 16882
rect 26012 16818 26068 16830
rect 26124 17442 26180 17454
rect 26124 17390 26126 17442
rect 26178 17390 26180 17442
rect 26124 17332 26180 17390
rect 26124 16884 26180 17276
rect 26348 17108 26404 17118
rect 26460 17108 26516 18286
rect 26572 17332 26628 18398
rect 26572 17266 26628 17276
rect 26348 17106 26516 17108
rect 26348 17054 26350 17106
rect 26402 17054 26516 17106
rect 26348 17052 26516 17054
rect 26348 17042 26404 17052
rect 26572 16996 26628 17006
rect 26572 16902 26628 16940
rect 26124 16818 26180 16828
rect 26236 16660 26292 16670
rect 26012 16658 26292 16660
rect 26012 16606 26238 16658
rect 26290 16606 26292 16658
rect 26012 16604 26292 16606
rect 25900 15874 25956 15886
rect 25900 15822 25902 15874
rect 25954 15822 25956 15874
rect 25900 15428 25956 15822
rect 25900 15362 25956 15372
rect 25788 15316 25844 15354
rect 25788 15250 25844 15260
rect 26012 15148 26068 16604
rect 26236 16594 26292 16604
rect 26684 16548 26740 18620
rect 26684 16482 26740 16492
rect 26684 15540 26740 15550
rect 25340 15092 25508 15148
rect 25452 14530 25508 15092
rect 25452 14478 25454 14530
rect 25506 14478 25508 14530
rect 25452 14466 25508 14478
rect 25564 15092 25732 15148
rect 25900 15092 26068 15148
rect 26124 15428 26180 15438
rect 25564 14084 25620 15092
rect 25900 14530 25956 15092
rect 26124 14644 26180 15372
rect 26460 15426 26516 15438
rect 26460 15374 26462 15426
rect 26514 15374 26516 15426
rect 26460 15148 26516 15374
rect 26460 15092 26628 15148
rect 25900 14478 25902 14530
rect 25954 14478 25956 14530
rect 25900 14466 25956 14478
rect 26012 14588 26180 14644
rect 25452 14028 25620 14084
rect 25676 14420 25732 14430
rect 25676 14306 25732 14364
rect 25676 14254 25678 14306
rect 25730 14254 25732 14306
rect 25340 13972 25396 13982
rect 25340 13858 25396 13916
rect 25340 13806 25342 13858
rect 25394 13806 25396 13858
rect 25340 13794 25396 13806
rect 25228 13570 25284 13580
rect 25340 13412 25396 13422
rect 25340 13074 25396 13356
rect 25452 13188 25508 14028
rect 25452 13122 25508 13132
rect 25564 13858 25620 13870
rect 25564 13806 25566 13858
rect 25618 13806 25620 13858
rect 25340 13022 25342 13074
rect 25394 13022 25396 13074
rect 25340 13010 25396 13022
rect 25564 13076 25620 13806
rect 25676 13748 25732 14254
rect 25788 14308 25844 14318
rect 25788 14214 25844 14252
rect 25676 13682 25732 13692
rect 25788 14084 25844 14094
rect 25676 13524 25732 13534
rect 25676 13430 25732 13468
rect 25564 13010 25620 13020
rect 25788 13074 25844 14028
rect 26012 13970 26068 14588
rect 26124 14418 26180 14430
rect 26124 14366 26126 14418
rect 26178 14366 26180 14418
rect 26124 14084 26180 14366
rect 26124 14018 26180 14028
rect 26460 14418 26516 14430
rect 26460 14366 26462 14418
rect 26514 14366 26516 14418
rect 26012 13918 26014 13970
rect 26066 13918 26068 13970
rect 26012 13412 26068 13918
rect 26460 13524 26516 14366
rect 26572 14308 26628 15092
rect 26684 14530 26740 15484
rect 26796 15428 26852 22316
rect 26908 23772 27076 23828
rect 27132 23828 27188 23838
rect 27468 23828 27524 23838
rect 26908 21028 26964 23772
rect 27020 22932 27076 22942
rect 27020 22036 27076 22876
rect 27020 21970 27076 21980
rect 26908 20972 27076 21028
rect 26908 19908 26964 19918
rect 26908 19814 26964 19852
rect 27020 19684 27076 20972
rect 26908 19628 27076 19684
rect 27132 19684 27188 23772
rect 27356 23826 27524 23828
rect 27356 23774 27470 23826
rect 27522 23774 27524 23826
rect 27356 23772 27524 23774
rect 27244 23266 27300 23278
rect 27244 23214 27246 23266
rect 27298 23214 27300 23266
rect 27244 23156 27300 23214
rect 27244 21700 27300 23100
rect 27356 23042 27412 23772
rect 27468 23762 27524 23772
rect 27692 23828 27748 23838
rect 27692 23734 27748 23772
rect 27804 23714 27860 23996
rect 27804 23662 27806 23714
rect 27858 23662 27860 23714
rect 27804 23650 27860 23662
rect 28028 23826 28084 23838
rect 28028 23774 28030 23826
rect 28082 23774 28084 23826
rect 27692 23156 27748 23166
rect 27356 22990 27358 23042
rect 27410 22990 27412 23042
rect 27356 22978 27412 22990
rect 27468 23154 27748 23156
rect 27468 23102 27694 23154
rect 27746 23102 27748 23154
rect 27468 23100 27748 23102
rect 27356 22484 27412 22494
rect 27468 22484 27524 23100
rect 27692 23090 27748 23100
rect 28028 22932 28084 23774
rect 28028 22866 28084 22876
rect 27412 22428 27524 22484
rect 27356 22390 27412 22428
rect 28028 21812 28084 21822
rect 28028 21718 28084 21756
rect 27244 21634 27300 21644
rect 27916 21586 27972 21598
rect 27916 21534 27918 21586
rect 27970 21534 27972 21586
rect 27916 20356 27972 21534
rect 27580 20300 27972 20356
rect 27244 20244 27300 20254
rect 27580 20244 27636 20300
rect 27244 20242 27636 20244
rect 27244 20190 27246 20242
rect 27298 20190 27582 20242
rect 27634 20190 27636 20242
rect 27244 20188 27636 20190
rect 27244 20178 27300 20188
rect 27580 20178 27636 20188
rect 27692 20132 27748 20142
rect 27692 20038 27748 20076
rect 27916 20132 27972 20300
rect 28028 21362 28084 21374
rect 28028 21310 28030 21362
rect 28082 21310 28084 21362
rect 28028 20242 28084 21310
rect 28028 20190 28030 20242
rect 28082 20190 28084 20242
rect 28028 20178 28084 20190
rect 27916 20066 27972 20076
rect 26908 17332 26964 19628
rect 27132 19618 27188 19628
rect 27804 20018 27860 20030
rect 27804 19966 27806 20018
rect 27858 19966 27860 20018
rect 27804 19796 27860 19966
rect 28140 19908 28196 26126
rect 27020 19460 27076 19470
rect 27020 18788 27076 19404
rect 27580 19236 27636 19246
rect 27020 18722 27076 18732
rect 27244 19234 27636 19236
rect 27244 19182 27582 19234
rect 27634 19182 27636 19234
rect 27244 19180 27636 19182
rect 27244 18564 27300 19180
rect 27580 19170 27636 19180
rect 27356 19012 27412 19050
rect 27804 19012 27860 19740
rect 27356 18946 27412 18956
rect 27468 18956 27860 19012
rect 27916 19852 28196 19908
rect 27244 18498 27300 18508
rect 27356 18562 27412 18574
rect 27356 18510 27358 18562
rect 27410 18510 27412 18562
rect 27020 18450 27076 18462
rect 27020 18398 27022 18450
rect 27074 18398 27076 18450
rect 27020 18340 27076 18398
rect 27356 18452 27412 18510
rect 27468 18562 27524 18956
rect 27916 18900 27972 19852
rect 27692 18844 27972 18900
rect 28028 19684 28084 19694
rect 27468 18510 27470 18562
rect 27522 18510 27524 18562
rect 27468 18498 27524 18510
rect 27580 18788 27636 18798
rect 27356 18386 27412 18396
rect 27020 18274 27076 18284
rect 27356 18228 27412 18238
rect 27580 18228 27636 18732
rect 27356 18134 27412 18172
rect 27468 18172 27636 18228
rect 27468 18004 27524 18172
rect 27356 17948 27524 18004
rect 27020 17668 27076 17678
rect 27020 17574 27076 17612
rect 27356 17554 27412 17948
rect 27580 17668 27636 17678
rect 27356 17502 27358 17554
rect 27410 17502 27412 17554
rect 27356 17490 27412 17502
rect 27468 17556 27524 17566
rect 27468 17462 27524 17500
rect 27244 17442 27300 17454
rect 27244 17390 27246 17442
rect 27298 17390 27300 17442
rect 27132 17332 27188 17342
rect 26908 17276 27132 17332
rect 27132 17266 27188 17276
rect 27132 17108 27188 17118
rect 27020 17052 27132 17108
rect 27020 16994 27076 17052
rect 27132 17042 27188 17052
rect 27020 16942 27022 16994
rect 27074 16942 27076 16994
rect 27020 16930 27076 16942
rect 26796 15362 26852 15372
rect 26908 16882 26964 16894
rect 26908 16830 26910 16882
rect 26962 16830 26964 16882
rect 26908 15204 26964 16830
rect 27132 16884 27188 16894
rect 27132 16790 27188 16828
rect 26908 15138 26964 15148
rect 27244 14756 27300 17390
rect 27468 17332 27524 17342
rect 27468 14980 27524 17276
rect 27580 16882 27636 17612
rect 27580 16830 27582 16882
rect 27634 16830 27636 16882
rect 27580 16818 27636 16830
rect 27692 15148 27748 18844
rect 28028 18788 28084 19628
rect 27916 18732 28084 18788
rect 28140 19012 28196 19022
rect 28140 18788 28196 18956
rect 27804 18564 27860 18574
rect 27916 18564 27972 18732
rect 28140 18722 28196 18732
rect 27804 18562 27972 18564
rect 27804 18510 27806 18562
rect 27858 18510 27972 18562
rect 27804 18508 27972 18510
rect 27804 18498 27860 18508
rect 28028 18452 28084 18462
rect 27916 18338 27972 18350
rect 27916 18286 27918 18338
rect 27970 18286 27972 18338
rect 27804 17778 27860 17790
rect 27804 17726 27806 17778
rect 27858 17726 27860 17778
rect 27804 16994 27860 17726
rect 27916 17444 27972 18286
rect 28028 18228 28084 18396
rect 28252 18228 28308 26852
rect 30604 26852 30772 26908
rect 30828 27634 30884 27646
rect 30828 27582 30830 27634
rect 30882 27582 30884 27634
rect 30828 26908 30884 27582
rect 32732 27524 32788 30044
rect 32844 30034 32900 30044
rect 32956 33236 33012 33246
rect 33068 33236 33124 34748
rect 34188 34356 34244 34366
rect 34300 34356 34356 36204
rect 34412 35812 34468 37772
rect 34524 37380 34580 41020
rect 35084 41074 35140 41244
rect 35084 41022 35086 41074
rect 35138 41022 35140 41074
rect 35084 41010 35140 41022
rect 35196 41074 35252 41086
rect 35196 41022 35198 41074
rect 35250 41022 35252 41074
rect 34860 40964 34916 40974
rect 34860 40870 34916 40908
rect 35196 40964 35252 41022
rect 35196 40898 35252 40908
rect 35644 40964 35700 40974
rect 35756 40964 35812 45948
rect 35868 45938 35924 45948
rect 36540 46116 36596 46126
rect 36540 46002 36596 46060
rect 36540 45950 36542 46002
rect 36594 45950 36596 46002
rect 36540 45938 36596 45950
rect 37212 46002 37268 46396
rect 37212 45950 37214 46002
rect 37266 45950 37268 46002
rect 37212 45938 37268 45950
rect 37324 46004 37380 46014
rect 37436 46004 37492 47406
rect 37548 47012 37604 47022
rect 37548 46898 37604 46956
rect 37548 46846 37550 46898
rect 37602 46846 37604 46898
rect 37548 46834 37604 46846
rect 37996 47012 38052 47022
rect 37548 46674 37604 46686
rect 37548 46622 37550 46674
rect 37602 46622 37604 46674
rect 37548 46452 37604 46622
rect 37996 46674 38052 46956
rect 38332 46900 38388 46910
rect 38332 46786 38388 46844
rect 38332 46734 38334 46786
rect 38386 46734 38388 46786
rect 38332 46722 38388 46734
rect 37996 46622 37998 46674
rect 38050 46622 38052 46674
rect 37884 46564 37940 46574
rect 37884 46470 37940 46508
rect 37548 46116 37604 46396
rect 37996 46340 38052 46622
rect 37996 46274 38052 46284
rect 38444 46116 38500 47516
rect 38556 47506 38612 47516
rect 38668 47628 39060 47684
rect 38668 47012 38724 47628
rect 39228 47572 39284 48302
rect 39004 47516 39284 47572
rect 39340 47572 39396 49868
rect 39452 48244 39508 51100
rect 39900 51090 39956 51100
rect 40012 50932 40068 51324
rect 40124 51378 40236 51380
rect 40124 51326 40126 51378
rect 40178 51326 40236 51378
rect 40124 51324 40236 51326
rect 40124 51314 40180 51324
rect 40236 51286 40292 51324
rect 40012 50876 40292 50932
rect 40012 50708 40068 50718
rect 40012 50594 40068 50652
rect 40236 50706 40292 50876
rect 40236 50654 40238 50706
rect 40290 50654 40292 50706
rect 40236 50642 40292 50654
rect 40012 50542 40014 50594
rect 40066 50542 40068 50594
rect 40012 50530 40068 50542
rect 40124 50596 40180 50606
rect 39564 50484 39620 50494
rect 39788 50484 39844 50494
rect 39564 50482 39844 50484
rect 39564 50430 39566 50482
rect 39618 50430 39790 50482
rect 39842 50430 39844 50482
rect 39564 50428 39844 50430
rect 40124 50428 40180 50540
rect 40684 50594 40740 50606
rect 40684 50542 40686 50594
rect 40738 50542 40740 50594
rect 40348 50484 40404 50522
rect 40684 50428 40740 50542
rect 39564 50418 39620 50428
rect 39788 50372 39956 50428
rect 40124 50372 40292 50428
rect 40348 50418 40404 50428
rect 39676 49028 39732 49038
rect 39676 48466 39732 48972
rect 39676 48414 39678 48466
rect 39730 48414 39732 48466
rect 39676 48402 39732 48414
rect 39900 48356 39956 50372
rect 40012 50260 40068 50270
rect 40012 49588 40068 50204
rect 40236 50034 40292 50372
rect 40460 50372 40740 50428
rect 40796 50484 40852 50494
rect 40908 50428 40964 51438
rect 41020 51490 41076 51884
rect 41020 51438 41022 51490
rect 41074 51438 41076 51490
rect 41020 50820 41076 51438
rect 41020 50754 41076 50764
rect 41244 51378 41300 51390
rect 41244 51326 41246 51378
rect 41298 51326 41300 51378
rect 41244 50596 41300 51326
rect 41244 50530 41300 50540
rect 40796 50372 40964 50428
rect 41356 50484 41412 50494
rect 40460 50148 40516 50372
rect 40236 49982 40238 50034
rect 40290 49982 40292 50034
rect 40236 49970 40292 49982
rect 40348 50092 40516 50148
rect 40124 49922 40180 49934
rect 40124 49870 40126 49922
rect 40178 49870 40180 49922
rect 40124 49812 40180 49870
rect 40348 49812 40404 50092
rect 40796 50034 40852 50372
rect 40796 49982 40798 50034
rect 40850 49982 40852 50034
rect 40796 49970 40852 49982
rect 40124 49746 40180 49756
rect 40236 49756 40404 49812
rect 40012 49532 40180 49588
rect 40012 49028 40068 49038
rect 40012 48934 40068 48972
rect 39900 48300 40068 48356
rect 39452 48188 39956 48244
rect 39564 47572 39620 47582
rect 39340 47570 39620 47572
rect 39340 47518 39566 47570
rect 39618 47518 39620 47570
rect 39340 47516 39620 47518
rect 37548 46050 37604 46060
rect 38220 46114 38500 46116
rect 38220 46062 38446 46114
rect 38498 46062 38500 46114
rect 38220 46060 38500 46062
rect 37380 45948 37492 46004
rect 37324 45890 37380 45948
rect 37324 45838 37326 45890
rect 37378 45838 37380 45890
rect 37324 45826 37380 45838
rect 37548 45890 37604 45902
rect 37548 45838 37550 45890
rect 37602 45838 37604 45890
rect 37548 45780 37604 45838
rect 37548 45714 37604 45724
rect 37772 45890 37828 45902
rect 37772 45838 37774 45890
rect 37826 45838 37828 45890
rect 37100 45668 37156 45678
rect 37100 45574 37156 45612
rect 37660 45668 37716 45678
rect 36876 44994 36932 45006
rect 36876 44942 36878 44994
rect 36930 44942 36932 44994
rect 36876 44660 36932 44942
rect 37660 44660 37716 45612
rect 37772 45332 37828 45838
rect 38108 45780 38164 45790
rect 38108 45686 38164 45724
rect 37884 45332 37940 45342
rect 37772 45330 37940 45332
rect 37772 45278 37886 45330
rect 37938 45278 37940 45330
rect 37772 45276 37940 45278
rect 37884 45266 37940 45276
rect 37996 45332 38052 45342
rect 37996 45238 38052 45276
rect 37772 45108 37828 45118
rect 38220 45108 38276 46060
rect 38444 46050 38500 46060
rect 38556 46956 38724 47012
rect 38892 47458 38948 47470
rect 38892 47406 38894 47458
rect 38946 47406 38948 47458
rect 38892 47012 38948 47406
rect 38556 45668 38612 46956
rect 38892 46946 38948 46956
rect 38668 46788 38724 46798
rect 38668 46786 38948 46788
rect 38668 46734 38670 46786
rect 38722 46734 38948 46786
rect 38668 46732 38948 46734
rect 38668 46722 38724 46732
rect 38780 46564 38836 46574
rect 38780 46470 38836 46508
rect 38892 46452 38948 46732
rect 39004 46786 39060 47516
rect 39228 47460 39284 47516
rect 39564 47506 39620 47516
rect 39228 47404 39508 47460
rect 39452 47236 39508 47404
rect 39452 47180 39844 47236
rect 39676 46900 39732 46910
rect 39004 46734 39006 46786
rect 39058 46734 39060 46786
rect 39004 46722 39060 46734
rect 39228 46898 39732 46900
rect 39228 46846 39678 46898
rect 39730 46846 39732 46898
rect 39228 46844 39732 46846
rect 39228 46786 39284 46844
rect 39676 46834 39732 46844
rect 39788 46898 39844 47180
rect 39788 46846 39790 46898
rect 39842 46846 39844 46898
rect 39788 46834 39844 46846
rect 39228 46734 39230 46786
rect 39282 46734 39284 46786
rect 39228 46722 39284 46734
rect 39564 46674 39620 46686
rect 39900 46676 39956 48188
rect 40012 47684 40068 48300
rect 40124 48242 40180 49532
rect 40236 49138 40292 49756
rect 40348 49588 40404 49598
rect 41356 49588 41412 50428
rect 41468 50428 41524 52332
rect 41580 52162 41636 52174
rect 41580 52110 41582 52162
rect 41634 52110 41636 52162
rect 41580 51828 41636 52110
rect 41804 52162 41860 52174
rect 41804 52110 41806 52162
rect 41858 52110 41860 52162
rect 41580 51762 41636 51772
rect 41692 51938 41748 51950
rect 41692 51886 41694 51938
rect 41746 51886 41748 51938
rect 41692 51602 41748 51886
rect 41692 51550 41694 51602
rect 41746 51550 41748 51602
rect 41692 51538 41748 51550
rect 41804 51604 41860 52110
rect 41804 51538 41860 51548
rect 41916 51378 41972 53004
rect 42028 52994 42084 53004
rect 42140 52948 42196 52958
rect 42140 52854 42196 52892
rect 42364 52836 42420 52846
rect 42028 52722 42084 52734
rect 42028 52670 42030 52722
rect 42082 52670 42084 52722
rect 42028 52164 42084 52670
rect 42140 52164 42196 52174
rect 42028 52108 42140 52164
rect 42140 52070 42196 52108
rect 42364 52164 42420 52780
rect 42140 51940 42196 51950
rect 41916 51326 41918 51378
rect 41970 51326 41972 51378
rect 41804 51268 41860 51278
rect 41804 51174 41860 51212
rect 41916 51044 41972 51326
rect 41916 50978 41972 50988
rect 42028 51884 42140 51940
rect 41692 50708 41748 50718
rect 41692 50594 41748 50652
rect 41692 50542 41694 50594
rect 41746 50542 41748 50594
rect 41692 50530 41748 50542
rect 41916 50484 41972 50494
rect 42028 50484 42084 51884
rect 42140 51874 42196 51884
rect 42140 51380 42196 51390
rect 42140 51286 42196 51324
rect 42364 51378 42420 52108
rect 42364 51326 42366 51378
rect 42418 51326 42420 51378
rect 41916 50482 42084 50484
rect 41916 50430 41918 50482
rect 41970 50430 42084 50482
rect 41916 50428 42084 50430
rect 41468 50372 41860 50428
rect 41916 50418 41972 50428
rect 41804 50370 41860 50372
rect 41804 50318 41806 50370
rect 41858 50318 41860 50370
rect 41804 50306 41860 50318
rect 41692 50148 41748 50158
rect 41580 50092 41692 50148
rect 40348 49586 41412 49588
rect 40348 49534 40350 49586
rect 40402 49534 41412 49586
rect 40348 49532 41412 49534
rect 40348 49522 40404 49532
rect 40236 49086 40238 49138
rect 40290 49086 40292 49138
rect 40236 49074 40292 49086
rect 40348 49026 40404 49038
rect 40348 48974 40350 49026
rect 40402 48974 40404 49026
rect 40348 48580 40404 48974
rect 41244 48916 41300 48926
rect 41356 48916 41412 49532
rect 41244 48914 41412 48916
rect 41244 48862 41246 48914
rect 41298 48862 41412 48914
rect 41244 48860 41412 48862
rect 41468 49810 41524 49822
rect 41468 49758 41470 49810
rect 41522 49758 41524 49810
rect 41244 48850 41300 48860
rect 40348 48524 40628 48580
rect 40348 48356 40404 48366
rect 40348 48354 40516 48356
rect 40348 48302 40350 48354
rect 40402 48302 40516 48354
rect 40348 48300 40516 48302
rect 40348 48290 40404 48300
rect 40124 48190 40126 48242
rect 40178 48190 40180 48242
rect 40124 48178 40180 48190
rect 40012 47628 40180 47684
rect 40012 47458 40068 47470
rect 40012 47406 40014 47458
rect 40066 47406 40068 47458
rect 40012 46900 40068 47406
rect 40012 46834 40068 46844
rect 39564 46622 39566 46674
rect 39618 46622 39620 46674
rect 39564 46452 39620 46622
rect 38892 46396 39620 46452
rect 39564 46114 39620 46396
rect 39564 46062 39566 46114
rect 39618 46062 39620 46114
rect 39564 46050 39620 46062
rect 39676 46620 39956 46676
rect 38668 45892 38724 45902
rect 38668 45890 38836 45892
rect 38668 45838 38670 45890
rect 38722 45838 38836 45890
rect 38668 45836 38836 45838
rect 38668 45826 38724 45836
rect 38556 45612 38724 45668
rect 38668 45218 38724 45612
rect 38780 45332 38836 45836
rect 39228 45890 39284 45902
rect 39228 45838 39230 45890
rect 39282 45838 39284 45890
rect 39004 45780 39060 45790
rect 39004 45686 39060 45724
rect 39228 45444 39284 45838
rect 39228 45378 39284 45388
rect 38780 45238 38836 45276
rect 38668 45166 38670 45218
rect 38722 45166 38724 45218
rect 37772 45106 38276 45108
rect 37772 45054 37774 45106
rect 37826 45054 38276 45106
rect 37772 45052 38276 45054
rect 38444 45108 38500 45118
rect 37772 45042 37828 45052
rect 38444 45014 38500 45052
rect 37660 44604 37828 44660
rect 35980 44324 36036 44334
rect 35980 44230 36036 44268
rect 36876 44212 36932 44604
rect 37100 44322 37156 44334
rect 37100 44270 37102 44322
rect 37154 44270 37156 44322
rect 37100 44212 37156 44270
rect 37660 44324 37716 44334
rect 37660 44230 37716 44268
rect 37772 44324 37828 44604
rect 38668 44548 38724 45166
rect 39004 45106 39060 45118
rect 39004 45054 39006 45106
rect 39058 45054 39060 45106
rect 39004 44884 39060 45054
rect 39452 44996 39508 45006
rect 39452 44902 39508 44940
rect 39004 44818 39060 44828
rect 38668 44492 38836 44548
rect 38220 44436 38276 44446
rect 38220 44342 38276 44380
rect 38668 44324 38724 44334
rect 37772 44322 38052 44324
rect 37772 44270 37774 44322
rect 37826 44270 38052 44322
rect 37772 44268 38052 44270
rect 37772 44258 37828 44268
rect 36764 44156 37156 44212
rect 36652 44100 36708 44110
rect 36652 43650 36708 44044
rect 36652 43598 36654 43650
rect 36706 43598 36708 43650
rect 36652 43586 36708 43598
rect 35868 43538 35924 43550
rect 35868 43486 35870 43538
rect 35922 43486 35924 43538
rect 35868 42868 35924 43486
rect 36092 43540 36148 43550
rect 36092 43446 36148 43484
rect 36204 43538 36260 43550
rect 36204 43486 36206 43538
rect 36258 43486 36260 43538
rect 35868 42754 35924 42812
rect 35868 42702 35870 42754
rect 35922 42702 35924 42754
rect 35868 42690 35924 42702
rect 36204 43316 36260 43486
rect 36204 42756 36260 43260
rect 36540 43538 36596 43550
rect 36540 43486 36542 43538
rect 36594 43486 36596 43538
rect 36540 42980 36596 43486
rect 36540 42914 36596 42924
rect 36316 42868 36372 42878
rect 36316 42774 36372 42812
rect 36204 42662 36260 42700
rect 35644 40962 35812 40964
rect 35644 40910 35646 40962
rect 35698 40910 35812 40962
rect 35644 40908 35812 40910
rect 36092 40964 36148 40974
rect 35644 40516 35700 40908
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34636 39060 34692 39070
rect 34636 38966 34692 39004
rect 35196 38836 35252 38846
rect 35196 38742 35252 38780
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34748 38162 34804 38174
rect 34748 38110 34750 38162
rect 34802 38110 34804 38162
rect 34748 38052 34804 38110
rect 34748 37986 34804 37996
rect 35420 38052 35476 38062
rect 35420 37958 35476 37996
rect 35084 37828 35140 37838
rect 35644 37828 35700 40460
rect 36092 40404 36148 40908
rect 36540 40964 36596 40974
rect 36540 40514 36596 40908
rect 36540 40462 36542 40514
rect 36594 40462 36596 40514
rect 36540 40450 36596 40462
rect 36092 40338 36148 40348
rect 36092 39620 36148 39630
rect 35980 39284 36036 39294
rect 35756 38834 35812 38846
rect 35756 38782 35758 38834
rect 35810 38782 35812 38834
rect 35756 38052 35812 38782
rect 35756 37986 35812 37996
rect 35980 38836 36036 39228
rect 35868 37828 35924 37838
rect 35084 37734 35140 37772
rect 35532 37826 35924 37828
rect 35532 37774 35870 37826
rect 35922 37774 35924 37826
rect 35532 37772 35924 37774
rect 34748 37380 34804 37390
rect 34524 37378 34804 37380
rect 34524 37326 34750 37378
rect 34802 37326 34804 37378
rect 34524 37324 34804 37326
rect 34524 36708 34580 36718
rect 34524 36594 34580 36652
rect 34524 36542 34526 36594
rect 34578 36542 34580 36594
rect 34524 36530 34580 36542
rect 34412 35746 34468 35756
rect 34636 35588 34692 35598
rect 34636 35494 34692 35532
rect 34412 35028 34468 35038
rect 34748 35028 34804 37324
rect 34972 37378 35028 37390
rect 34972 37326 34974 37378
rect 35026 37326 35028 37378
rect 34860 36484 34916 36494
rect 34972 36484 35028 37326
rect 35532 37268 35588 37772
rect 35868 37762 35924 37772
rect 35980 37492 36036 38780
rect 36092 38722 36148 39564
rect 36652 39620 36708 39630
rect 36428 39394 36484 39406
rect 36428 39342 36430 39394
rect 36482 39342 36484 39394
rect 36428 38948 36484 39342
rect 36540 38948 36596 38958
rect 36428 38892 36540 38948
rect 36092 38670 36094 38722
rect 36146 38670 36148 38722
rect 36092 38668 36148 38670
rect 36316 38836 36372 38846
rect 36092 38612 36260 38668
rect 36204 38050 36260 38612
rect 36316 38274 36372 38780
rect 36316 38222 36318 38274
rect 36370 38222 36372 38274
rect 36316 38210 36372 38222
rect 36204 37998 36206 38050
rect 36258 37998 36260 38050
rect 36204 37986 36260 37998
rect 36540 38052 36596 38892
rect 36652 38946 36708 39564
rect 36652 38894 36654 38946
rect 36706 38894 36708 38946
rect 36652 38500 36708 38894
rect 36652 38434 36708 38444
rect 36540 37996 36708 38052
rect 36316 37828 36372 37838
rect 36372 37772 36484 37828
rect 36316 37734 36372 37772
rect 35532 37174 35588 37212
rect 35644 37490 36036 37492
rect 35644 37438 35982 37490
rect 36034 37438 36036 37490
rect 35644 37436 36036 37438
rect 34916 36428 35028 36484
rect 35084 37042 35140 37054
rect 35084 36990 35086 37042
rect 35138 36990 35140 37042
rect 35084 36484 35140 36990
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 34860 36418 34916 36428
rect 35084 36418 35140 36428
rect 35308 36708 35364 36718
rect 34860 36260 34916 36270
rect 34860 36166 34916 36204
rect 34972 36258 35028 36270
rect 34972 36206 34974 36258
rect 35026 36206 35028 36258
rect 34972 35476 35028 36206
rect 35084 36260 35140 36270
rect 35308 36260 35364 36652
rect 35084 36258 35364 36260
rect 35084 36206 35086 36258
rect 35138 36206 35364 36258
rect 35084 36204 35364 36206
rect 35420 36484 35476 36494
rect 35084 36194 35140 36204
rect 34972 35410 35028 35420
rect 35084 36036 35140 36046
rect 35084 35588 35140 35980
rect 35196 35698 35252 36204
rect 35308 35812 35364 35822
rect 35308 35718 35364 35756
rect 35196 35646 35198 35698
rect 35250 35646 35252 35698
rect 35196 35634 35252 35646
rect 35420 35700 35476 36428
rect 35532 36484 35588 36494
rect 35644 36484 35700 37436
rect 35980 37426 36036 37436
rect 36316 37492 36372 37502
rect 36316 36706 36372 37436
rect 36428 37378 36484 37772
rect 36428 37326 36430 37378
rect 36482 37326 36484 37378
rect 36428 37314 36484 37326
rect 36652 37266 36708 37996
rect 36652 37214 36654 37266
rect 36706 37214 36708 37266
rect 36652 37202 36708 37214
rect 36316 36654 36318 36706
rect 36370 36654 36372 36706
rect 36316 36642 36372 36654
rect 35532 36482 35700 36484
rect 35532 36430 35534 36482
rect 35586 36430 35700 36482
rect 35532 36428 35700 36430
rect 35980 36484 36036 36494
rect 35532 36418 35588 36428
rect 35980 36390 36036 36428
rect 35756 36370 35812 36382
rect 35756 36318 35758 36370
rect 35810 36318 35812 36370
rect 35756 35924 35812 36318
rect 36204 36260 36260 36270
rect 36092 36258 36260 36260
rect 36092 36206 36206 36258
rect 36258 36206 36260 36258
rect 36092 36204 36260 36206
rect 35756 35922 36036 35924
rect 35756 35870 35758 35922
rect 35810 35870 36036 35922
rect 35756 35868 36036 35870
rect 35756 35858 35812 35868
rect 35420 35644 35924 35700
rect 34412 34934 34468 34972
rect 34636 34972 34804 35028
rect 34860 35028 34916 35038
rect 34188 34354 34356 34356
rect 34188 34302 34190 34354
rect 34242 34302 34356 34354
rect 34188 34300 34356 34302
rect 34188 34290 34244 34300
rect 34412 34130 34468 34142
rect 34412 34078 34414 34130
rect 34466 34078 34468 34130
rect 33180 34020 33236 34030
rect 33180 33346 33236 33964
rect 34300 34020 34356 34030
rect 34300 33926 34356 33964
rect 33180 33294 33182 33346
rect 33234 33294 33236 33346
rect 33180 33282 33236 33294
rect 33628 33346 33684 33358
rect 33628 33294 33630 33346
rect 33682 33294 33684 33346
rect 32956 33234 33124 33236
rect 32956 33182 32958 33234
rect 33010 33182 33124 33234
rect 32956 33180 33124 33182
rect 32956 29876 33012 33180
rect 33628 33124 33684 33294
rect 34300 33236 34356 33246
rect 34300 33142 34356 33180
rect 33628 33058 33684 33068
rect 33180 33012 33236 33022
rect 33180 32674 33236 32956
rect 33180 32622 33182 32674
rect 33234 32622 33236 32674
rect 33180 32610 33236 32622
rect 33740 33012 33796 33022
rect 33068 32564 33124 32574
rect 33068 32470 33124 32508
rect 33628 32450 33684 32462
rect 33628 32398 33630 32450
rect 33682 32398 33684 32450
rect 33628 32340 33684 32398
rect 33628 32274 33684 32284
rect 33740 31890 33796 32956
rect 33740 31838 33742 31890
rect 33794 31838 33796 31890
rect 33740 31826 33796 31838
rect 33068 31780 33124 31790
rect 33068 31106 33124 31724
rect 34188 31780 34244 31790
rect 34188 31686 34244 31724
rect 34412 31668 34468 34078
rect 34524 33124 34580 33134
rect 34524 32564 34580 33068
rect 34636 33012 34692 34972
rect 34860 34914 34916 34972
rect 34860 34862 34862 34914
rect 34914 34862 34916 34914
rect 34860 34850 34916 34862
rect 35084 35028 35140 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 35028 35252 35038
rect 35644 35028 35700 35038
rect 35084 35026 35364 35028
rect 35084 34974 35198 35026
rect 35250 34974 35364 35026
rect 35084 34972 35364 34974
rect 34860 34132 34916 34142
rect 35084 34132 35140 34972
rect 35196 34962 35252 34972
rect 35308 34354 35364 34972
rect 35308 34302 35310 34354
rect 35362 34302 35364 34354
rect 35308 34290 35364 34302
rect 34860 34130 35140 34132
rect 34860 34078 34862 34130
rect 34914 34078 35140 34130
rect 34860 34076 35140 34078
rect 34860 34066 34916 34076
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34636 32946 34692 32956
rect 35196 32788 35252 32798
rect 35196 32674 35252 32732
rect 35196 32622 35198 32674
rect 35250 32622 35252 32674
rect 35196 32610 35252 32622
rect 34524 32562 34692 32564
rect 34524 32510 34526 32562
rect 34578 32510 34692 32562
rect 34524 32508 34692 32510
rect 34524 32498 34580 32508
rect 33068 31054 33070 31106
rect 33122 31054 33124 31106
rect 33068 31042 33124 31054
rect 33292 31556 33348 31566
rect 33292 31106 33348 31500
rect 33292 31054 33294 31106
rect 33346 31054 33348 31106
rect 33292 31042 33348 31054
rect 33964 31108 34020 31118
rect 33964 31014 34020 31052
rect 34076 31108 34132 31118
rect 34076 31106 34244 31108
rect 34076 31054 34078 31106
rect 34130 31054 34244 31106
rect 34076 31052 34244 31054
rect 34076 31042 34132 31052
rect 33740 30994 33796 31006
rect 33740 30942 33742 30994
rect 33794 30942 33796 30994
rect 33516 30882 33572 30894
rect 33516 30830 33518 30882
rect 33570 30830 33572 30882
rect 33404 30436 33460 30446
rect 33180 30324 33236 30334
rect 32844 29820 33012 29876
rect 33068 30212 33124 30222
rect 32844 29428 32900 29820
rect 32844 29362 32900 29372
rect 33068 29426 33124 30156
rect 33068 29374 33070 29426
rect 33122 29374 33124 29426
rect 33068 29362 33124 29374
rect 33180 28642 33236 30268
rect 33180 28590 33182 28642
rect 33234 28590 33236 28642
rect 32284 27468 32788 27524
rect 32844 27860 32900 27870
rect 33180 27860 33236 28590
rect 32900 27858 33236 27860
rect 32900 27806 33182 27858
rect 33234 27806 33236 27858
rect 32900 27804 33236 27806
rect 32060 27186 32116 27198
rect 32060 27134 32062 27186
rect 32114 27134 32116 27186
rect 32060 26908 32116 27134
rect 30828 26852 31108 26908
rect 30604 26292 30660 26852
rect 31052 26402 31108 26852
rect 31052 26350 31054 26402
rect 31106 26350 31108 26402
rect 31052 26338 31108 26350
rect 31388 26852 32116 26908
rect 30492 26290 30660 26292
rect 30492 26238 30606 26290
rect 30658 26238 30660 26290
rect 30492 26236 30660 26238
rect 28588 25620 28644 25630
rect 28588 25618 28980 25620
rect 28588 25566 28590 25618
rect 28642 25566 28980 25618
rect 28588 25564 28980 25566
rect 28588 25554 28644 25564
rect 28924 24834 28980 25564
rect 30492 25618 30548 26236
rect 30604 26226 30660 26236
rect 30716 26180 30772 26190
rect 30716 25730 30772 26124
rect 30828 26180 30884 26190
rect 31388 26180 31444 26852
rect 30828 26178 31444 26180
rect 30828 26126 30830 26178
rect 30882 26126 31390 26178
rect 31442 26126 31444 26178
rect 30828 26124 31444 26126
rect 30828 26114 30884 26124
rect 31388 26114 31444 26124
rect 31612 26180 31668 26190
rect 31612 26086 31668 26124
rect 30716 25678 30718 25730
rect 30770 25678 30772 25730
rect 30716 25666 30772 25678
rect 31948 26066 32004 26078
rect 31948 26014 31950 26066
rect 32002 26014 32004 26066
rect 30492 25566 30494 25618
rect 30546 25566 30548 25618
rect 30492 25554 30548 25566
rect 31052 25284 31108 25294
rect 31052 25282 31332 25284
rect 31052 25230 31054 25282
rect 31106 25230 31332 25282
rect 31052 25228 31332 25230
rect 31052 25218 31108 25228
rect 28924 24782 28926 24834
rect 28978 24782 28980 24834
rect 28924 24770 28980 24782
rect 28812 24498 28868 24510
rect 28812 24446 28814 24498
rect 28866 24446 28868 24498
rect 28812 23828 28868 24446
rect 29484 24052 29540 24062
rect 29484 24050 29652 24052
rect 29484 23998 29486 24050
rect 29538 23998 29652 24050
rect 29484 23996 29652 23998
rect 29484 23986 29540 23996
rect 28812 23762 28868 23772
rect 29148 23826 29204 23838
rect 29148 23774 29150 23826
rect 29202 23774 29204 23826
rect 28476 23044 28532 23054
rect 28476 22950 28532 22988
rect 29036 22932 29092 22942
rect 29148 22932 29204 23774
rect 29372 23716 29428 23726
rect 29372 23714 29540 23716
rect 29372 23662 29374 23714
rect 29426 23662 29540 23714
rect 29372 23660 29540 23662
rect 29372 23650 29428 23660
rect 29092 22876 29204 22932
rect 29260 23044 29316 23054
rect 29036 22370 29092 22876
rect 29260 22482 29316 22988
rect 29260 22430 29262 22482
rect 29314 22430 29316 22482
rect 29260 22418 29316 22430
rect 29484 22484 29540 23660
rect 29036 22318 29038 22370
rect 29090 22318 29092 22370
rect 29036 22306 29092 22318
rect 29372 22372 29428 22382
rect 28588 21812 28644 21822
rect 29372 21812 29428 22316
rect 29484 22036 29540 22428
rect 29596 22370 29652 23996
rect 31052 23156 31108 23166
rect 30604 23154 31108 23156
rect 30604 23102 31054 23154
rect 31106 23102 31108 23154
rect 30604 23100 31108 23102
rect 30604 23042 30660 23100
rect 31052 23090 31108 23100
rect 30604 22990 30606 23042
rect 30658 22990 30660 23042
rect 30604 22978 30660 22990
rect 29596 22318 29598 22370
rect 29650 22318 29652 22370
rect 29596 22306 29652 22318
rect 30940 22930 30996 22942
rect 30940 22878 30942 22930
rect 30994 22878 30996 22930
rect 30940 22372 30996 22878
rect 30940 22306 30996 22316
rect 31052 22370 31108 22382
rect 31052 22318 31054 22370
rect 31106 22318 31108 22370
rect 29484 21970 29540 21980
rect 30268 22148 30324 22158
rect 28588 21718 28644 21756
rect 29148 21756 29428 21812
rect 28588 20914 28644 20926
rect 28588 20862 28590 20914
rect 28642 20862 28644 20914
rect 28588 20130 28644 20862
rect 28588 20078 28590 20130
rect 28642 20078 28644 20130
rect 28588 20066 28644 20078
rect 28476 19906 28532 19918
rect 28476 19854 28478 19906
rect 28530 19854 28532 19906
rect 28364 19796 28420 19806
rect 28476 19796 28532 19854
rect 28420 19740 28532 19796
rect 28364 19730 28420 19740
rect 29036 18676 29092 18686
rect 28364 18452 28420 18462
rect 28364 18358 28420 18396
rect 28812 18452 28868 18462
rect 28812 18358 28868 18396
rect 29036 18450 29092 18620
rect 29148 18564 29204 21756
rect 29484 21698 29540 21710
rect 29484 21646 29486 21698
rect 29538 21646 29540 21698
rect 29260 21588 29316 21598
rect 29260 20802 29316 21532
rect 29260 20750 29262 20802
rect 29314 20750 29316 20802
rect 29260 20738 29316 20750
rect 29372 21586 29428 21598
rect 29372 21534 29374 21586
rect 29426 21534 29428 21586
rect 29372 20242 29428 21534
rect 29484 21140 29540 21646
rect 29708 21588 29764 21598
rect 29708 21586 29988 21588
rect 29708 21534 29710 21586
rect 29762 21534 29988 21586
rect 29708 21532 29988 21534
rect 29708 21522 29764 21532
rect 29484 21074 29540 21084
rect 29932 20916 29988 21532
rect 30044 21474 30100 21486
rect 30044 21422 30046 21474
rect 30098 21422 30100 21474
rect 30044 21140 30100 21422
rect 30044 21074 30100 21084
rect 29932 20860 30100 20916
rect 29932 20692 29988 20702
rect 29372 20190 29374 20242
rect 29426 20190 29428 20242
rect 29372 20132 29428 20190
rect 29484 20690 29988 20692
rect 29484 20638 29934 20690
rect 29986 20638 29988 20690
rect 29484 20636 29988 20638
rect 29484 20242 29540 20636
rect 29932 20626 29988 20636
rect 29484 20190 29486 20242
rect 29538 20190 29540 20242
rect 29484 20178 29540 20190
rect 29372 20066 29428 20076
rect 29596 20020 29652 20030
rect 29596 19926 29652 19964
rect 29932 20020 29988 20030
rect 29932 19234 29988 19964
rect 30044 20018 30100 20860
rect 30044 19966 30046 20018
rect 30098 19966 30100 20018
rect 30044 19954 30100 19966
rect 29932 19182 29934 19234
rect 29986 19182 29988 19234
rect 29932 19170 29988 19182
rect 29596 19012 29652 19022
rect 29596 18918 29652 18956
rect 29820 19010 29876 19022
rect 29820 18958 29822 19010
rect 29874 18958 29876 19010
rect 29820 18676 29876 18958
rect 29820 18610 29876 18620
rect 30156 18900 30212 18910
rect 29260 18564 29316 18574
rect 29148 18562 29316 18564
rect 29148 18510 29262 18562
rect 29314 18510 29316 18562
rect 29148 18508 29316 18510
rect 29260 18498 29316 18508
rect 29484 18564 29540 18574
rect 29036 18398 29038 18450
rect 29090 18398 29092 18450
rect 29036 18386 29092 18398
rect 28028 18162 28084 18172
rect 28140 18172 28308 18228
rect 29148 18338 29204 18350
rect 29148 18286 29150 18338
rect 29202 18286 29204 18338
rect 27916 17378 27972 17388
rect 28028 17108 28084 17118
rect 28028 17014 28084 17052
rect 27804 16942 27806 16994
rect 27858 16942 27860 16994
rect 27804 16930 27860 16942
rect 27916 16658 27972 16670
rect 27916 16606 27918 16658
rect 27970 16606 27972 16658
rect 27916 15540 27972 16606
rect 27916 15474 27972 15484
rect 28028 15428 28084 15438
rect 28028 15334 28084 15372
rect 27692 15092 27972 15148
rect 27468 14924 27860 14980
rect 27692 14756 27748 14766
rect 27244 14700 27636 14756
rect 27020 14642 27076 14654
rect 27020 14590 27022 14642
rect 27074 14590 27076 14642
rect 26684 14478 26686 14530
rect 26738 14478 26740 14530
rect 26684 14466 26740 14478
rect 26796 14532 26852 14542
rect 27020 14532 27076 14590
rect 27468 14532 27524 14542
rect 27020 14530 27524 14532
rect 27020 14478 27470 14530
rect 27522 14478 27524 14530
rect 27020 14476 27524 14478
rect 26572 14252 26740 14308
rect 26572 13748 26628 13758
rect 26572 13654 26628 13692
rect 26460 13458 26516 13468
rect 26684 13412 26740 14252
rect 26012 13346 26068 13356
rect 26572 13356 26740 13412
rect 26348 13300 26404 13310
rect 26348 13186 26404 13244
rect 26348 13134 26350 13186
rect 26402 13134 26404 13186
rect 26348 13122 26404 13134
rect 25788 13022 25790 13074
rect 25842 13022 25844 13074
rect 25788 13010 25844 13022
rect 25900 12964 25956 12974
rect 25900 12870 25956 12908
rect 26572 12964 26628 13356
rect 26684 13188 26740 13198
rect 26796 13188 26852 14476
rect 27468 14466 27524 14476
rect 26908 14420 26964 14430
rect 26908 14326 26964 14364
rect 27020 14308 27076 14318
rect 27468 14308 27524 14318
rect 27020 14306 27188 14308
rect 27020 14254 27022 14306
rect 27074 14254 27188 14306
rect 27020 14252 27188 14254
rect 27020 14242 27076 14252
rect 26684 13186 26852 13188
rect 26684 13134 26686 13186
rect 26738 13134 26852 13186
rect 26684 13132 26852 13134
rect 26684 13122 26740 13132
rect 25564 12852 25620 12862
rect 25564 12758 25620 12796
rect 26572 12850 26628 12908
rect 26572 12798 26574 12850
rect 26626 12798 26628 12850
rect 26572 12786 26628 12798
rect 25228 12740 25284 12750
rect 25004 12684 25172 12740
rect 24780 12180 24836 12190
rect 24780 11394 24836 12124
rect 25116 12068 25172 12684
rect 25228 12290 25284 12684
rect 25900 12740 25956 12750
rect 25900 12404 25956 12684
rect 25900 12310 25956 12348
rect 25228 12238 25230 12290
rect 25282 12238 25284 12290
rect 25228 12226 25284 12238
rect 25340 12180 25396 12190
rect 25340 12086 25396 12124
rect 25116 12012 25284 12068
rect 24780 11342 24782 11394
rect 24834 11342 24836 11394
rect 24780 11330 24836 11342
rect 25228 11956 25284 12012
rect 25116 11282 25172 11294
rect 25116 11230 25118 11282
rect 25170 11230 25172 11282
rect 25116 10724 25172 11230
rect 25228 11284 25284 11900
rect 25452 11284 25508 11294
rect 25228 11282 25508 11284
rect 25228 11230 25454 11282
rect 25506 11230 25508 11282
rect 25228 11228 25508 11230
rect 27132 11284 27188 14252
rect 27468 13746 27524 14252
rect 27468 13694 27470 13746
rect 27522 13694 27524 13746
rect 27468 13682 27524 13694
rect 27244 13634 27300 13646
rect 27244 13582 27246 13634
rect 27298 13582 27300 13634
rect 27244 12738 27300 13582
rect 27580 13524 27636 14700
rect 27244 12686 27246 12738
rect 27298 12686 27300 12738
rect 27244 12404 27300 12686
rect 27244 12338 27300 12348
rect 27468 13468 27636 13524
rect 27468 12516 27524 13468
rect 27468 12402 27524 12460
rect 27468 12350 27470 12402
rect 27522 12350 27524 12402
rect 27468 12338 27524 12350
rect 27580 12852 27636 12862
rect 27580 12404 27636 12796
rect 27580 12338 27636 12348
rect 27692 12402 27748 14700
rect 27804 13634 27860 14924
rect 27916 14418 27972 15092
rect 28140 14642 28196 18172
rect 28252 16996 28308 17006
rect 28308 16940 28532 16996
rect 28252 16902 28308 16940
rect 28364 16212 28420 16222
rect 28364 15314 28420 16156
rect 28476 15764 28532 16940
rect 28476 15708 28756 15764
rect 28364 15262 28366 15314
rect 28418 15262 28420 15314
rect 28364 15250 28420 15262
rect 28476 15538 28532 15550
rect 28476 15486 28478 15538
rect 28530 15486 28532 15538
rect 28140 14590 28142 14642
rect 28194 14590 28196 14642
rect 28140 14578 28196 14590
rect 28364 14532 28420 14542
rect 27916 14366 27918 14418
rect 27970 14366 27972 14418
rect 27916 13860 27972 14366
rect 28252 14530 28420 14532
rect 28252 14478 28366 14530
rect 28418 14478 28420 14530
rect 28252 14476 28420 14478
rect 28252 13972 28308 14476
rect 28364 14466 28420 14476
rect 28252 13906 28308 13916
rect 28364 14308 28420 14318
rect 27916 13766 27972 13804
rect 28364 13746 28420 14252
rect 28364 13694 28366 13746
rect 28418 13694 28420 13746
rect 28364 13682 28420 13694
rect 27804 13582 27806 13634
rect 27858 13582 27860 13634
rect 27804 13570 27860 13582
rect 28252 12852 28308 12862
rect 28252 12758 28308 12796
rect 27692 12350 27694 12402
rect 27746 12350 27748 12402
rect 27692 12338 27748 12350
rect 27916 12738 27972 12750
rect 27916 12686 27918 12738
rect 27970 12686 27972 12738
rect 27916 12404 27972 12686
rect 28364 12404 28420 12414
rect 27916 12348 28364 12404
rect 27244 12180 27300 12190
rect 27244 12086 27300 12124
rect 28364 12178 28420 12348
rect 28364 12126 28366 12178
rect 28418 12126 28420 12178
rect 28364 12114 28420 12126
rect 28476 12178 28532 15486
rect 28588 15092 28644 15102
rect 28588 14998 28644 15036
rect 28700 14196 28756 15708
rect 28812 15316 28868 15326
rect 28812 15222 28868 15260
rect 29148 14756 29204 18286
rect 29484 17668 29540 18508
rect 29708 18452 29764 18462
rect 29484 17666 29652 17668
rect 29484 17614 29486 17666
rect 29538 17614 29652 17666
rect 29484 17612 29652 17614
rect 29484 17602 29540 17612
rect 29596 17108 29652 17612
rect 29708 17556 29764 18396
rect 29820 18450 29876 18462
rect 29820 18398 29822 18450
rect 29874 18398 29876 18450
rect 29820 18228 29876 18398
rect 30044 18340 30100 18350
rect 30044 18246 30100 18284
rect 29820 18162 29876 18172
rect 30156 18116 30212 18844
rect 30268 18450 30324 22092
rect 31052 21588 31108 22318
rect 31052 21522 31108 21532
rect 31164 21924 31220 21934
rect 30940 20916 30996 20926
rect 30940 20130 30996 20860
rect 30940 20078 30942 20130
rect 30994 20078 30996 20130
rect 30940 20066 30996 20078
rect 30828 20020 30884 20030
rect 30828 19926 30884 19964
rect 30268 18398 30270 18450
rect 30322 18398 30324 18450
rect 30268 18386 30324 18398
rect 30492 18452 30548 18462
rect 30492 18358 30548 18396
rect 30716 18450 30772 18462
rect 30716 18398 30718 18450
rect 30770 18398 30772 18450
rect 30156 18050 30212 18060
rect 30380 18228 30436 18238
rect 29820 17556 29876 17566
rect 29708 17554 29876 17556
rect 29708 17502 29822 17554
rect 29874 17502 29876 17554
rect 29708 17500 29876 17502
rect 29820 17490 29876 17500
rect 29708 17108 29764 17118
rect 29596 17106 29764 17108
rect 29596 17054 29710 17106
rect 29762 17054 29764 17106
rect 29596 17052 29764 17054
rect 29484 16324 29540 16334
rect 29484 15428 29540 16268
rect 29596 16098 29652 17052
rect 29708 17042 29764 17052
rect 30380 17106 30436 18172
rect 30716 18228 30772 18398
rect 31164 18450 31220 21868
rect 31164 18398 31166 18450
rect 31218 18398 31220 18450
rect 31164 18386 31220 18398
rect 31276 20130 31332 25228
rect 31724 23266 31780 23278
rect 31724 23214 31726 23266
rect 31778 23214 31780 23266
rect 31724 22482 31780 23214
rect 31724 22430 31726 22482
rect 31778 22430 31780 22482
rect 31724 22418 31780 22430
rect 31276 20078 31278 20130
rect 31330 20078 31332 20130
rect 30716 18162 30772 18172
rect 30940 18338 30996 18350
rect 30940 18286 30942 18338
rect 30994 18286 30996 18338
rect 30940 17668 30996 18286
rect 30940 17602 30996 17612
rect 31052 18004 31108 18014
rect 31052 17556 31108 17948
rect 31052 17462 31108 17500
rect 30940 17220 30996 17230
rect 30380 17054 30382 17106
rect 30434 17054 30436 17106
rect 30380 17042 30436 17054
rect 30828 17164 30940 17220
rect 30996 17164 31108 17220
rect 29596 16046 29598 16098
rect 29650 16046 29652 16098
rect 29596 16034 29652 16046
rect 30044 16994 30100 17006
rect 30044 16942 30046 16994
rect 30098 16942 30100 16994
rect 30044 16100 30100 16942
rect 30716 16882 30772 16894
rect 30716 16830 30718 16882
rect 30770 16830 30772 16882
rect 30716 16436 30772 16830
rect 30716 16370 30772 16380
rect 30716 16212 30772 16222
rect 30828 16212 30884 17164
rect 30940 17154 30996 17164
rect 31052 16994 31108 17164
rect 31052 16942 31054 16994
rect 31106 16942 31108 16994
rect 31052 16930 31108 16942
rect 30044 16034 30100 16044
rect 30492 16210 30884 16212
rect 30492 16158 30718 16210
rect 30770 16158 30884 16210
rect 30492 16156 30884 16158
rect 29932 15876 29988 15886
rect 29484 15362 29540 15372
rect 29820 15874 29988 15876
rect 29820 15822 29934 15874
rect 29986 15822 29988 15874
rect 29820 15820 29988 15822
rect 29596 15316 29652 15326
rect 29820 15316 29876 15820
rect 29932 15810 29988 15820
rect 30156 15876 30212 15886
rect 29932 15428 29988 15438
rect 29932 15334 29988 15372
rect 30156 15426 30212 15820
rect 30156 15374 30158 15426
rect 30210 15374 30212 15426
rect 30156 15362 30212 15374
rect 29652 15260 29876 15316
rect 29596 15222 29652 15260
rect 30044 15202 30100 15214
rect 30044 15150 30046 15202
rect 30098 15150 30100 15202
rect 29148 14690 29204 14700
rect 29596 15090 29652 15102
rect 29596 15038 29598 15090
rect 29650 15038 29652 15090
rect 29148 14532 29204 14542
rect 29148 14438 29204 14476
rect 29036 14308 29092 14318
rect 29036 14214 29092 14252
rect 28588 12852 28644 12862
rect 28700 12852 28756 14140
rect 28812 13972 28868 13982
rect 28812 13878 28868 13916
rect 29260 13746 29316 13758
rect 29260 13694 29262 13746
rect 29314 13694 29316 13746
rect 29260 13074 29316 13694
rect 29260 13022 29262 13074
rect 29314 13022 29316 13074
rect 29260 13010 29316 13022
rect 29484 12964 29540 12974
rect 29484 12870 29540 12908
rect 29148 12852 29204 12862
rect 28588 12850 28756 12852
rect 28588 12798 28590 12850
rect 28642 12798 28756 12850
rect 28588 12796 28756 12798
rect 28812 12850 29204 12852
rect 28812 12798 29150 12850
rect 29202 12798 29204 12850
rect 28812 12796 29204 12798
rect 28588 12786 28644 12796
rect 28812 12402 28868 12796
rect 29148 12786 29204 12796
rect 28812 12350 28814 12402
rect 28866 12350 28868 12402
rect 28812 12338 28868 12350
rect 28476 12126 28478 12178
rect 28530 12126 28532 12178
rect 28476 12114 28532 12126
rect 28700 12180 28756 12190
rect 28700 12086 28756 12124
rect 28924 12178 28980 12190
rect 29260 12180 29316 12190
rect 28924 12126 28926 12178
rect 28978 12126 28980 12178
rect 27356 12066 27412 12078
rect 27356 12014 27358 12066
rect 27410 12014 27412 12066
rect 27356 11620 27412 12014
rect 27916 12068 27972 12078
rect 27916 11844 27972 12012
rect 27916 11778 27972 11788
rect 28140 11844 28196 11854
rect 27356 11564 27860 11620
rect 27468 11396 27524 11406
rect 27468 11302 27524 11340
rect 27804 11394 27860 11564
rect 27804 11342 27806 11394
rect 27858 11342 27860 11394
rect 27804 11330 27860 11342
rect 28140 11394 28196 11788
rect 28140 11342 28142 11394
rect 28194 11342 28196 11394
rect 28140 11330 28196 11342
rect 27132 11228 27412 11284
rect 25452 11218 25508 11228
rect 25900 11172 25956 11182
rect 27020 11172 27076 11182
rect 25788 11170 26516 11172
rect 25788 11118 25902 11170
rect 25954 11118 26516 11170
rect 25788 11116 26516 11118
rect 25228 10836 25284 10846
rect 25284 10780 25396 10836
rect 25228 10770 25284 10780
rect 25116 10658 25172 10668
rect 25340 10722 25396 10780
rect 25340 10670 25342 10722
rect 25394 10670 25396 10722
rect 25340 10658 25396 10670
rect 25228 10500 25284 10510
rect 24668 10498 25284 10500
rect 24668 10446 25230 10498
rect 25282 10446 25284 10498
rect 24668 10444 25284 10446
rect 25228 10434 25284 10444
rect 25564 10388 25620 10398
rect 25564 10294 25620 10332
rect 25116 9716 25172 9726
rect 25564 9716 25620 9726
rect 25116 9714 25620 9716
rect 25116 9662 25118 9714
rect 25170 9662 25566 9714
rect 25618 9662 25620 9714
rect 25116 9660 25620 9662
rect 25116 9650 25172 9660
rect 25564 9650 25620 9660
rect 24780 9604 24836 9614
rect 24668 9602 24836 9604
rect 24668 9550 24782 9602
rect 24834 9550 24836 9602
rect 24668 9548 24836 9550
rect 24668 8370 24724 9548
rect 24780 9538 24836 9548
rect 25676 9604 25732 9614
rect 25788 9604 25844 11116
rect 25900 11106 25956 11116
rect 26124 10836 26180 10846
rect 26124 10500 26180 10780
rect 26460 10610 26516 11116
rect 26908 11170 27076 11172
rect 26908 11118 27022 11170
rect 27074 11118 27076 11170
rect 26908 11116 27076 11118
rect 27356 11172 27412 11228
rect 27692 11172 27748 11182
rect 27356 11170 27748 11172
rect 27356 11118 27694 11170
rect 27746 11118 27748 11170
rect 27356 11116 27748 11118
rect 26572 10836 26628 10846
rect 26572 10722 26628 10780
rect 26572 10670 26574 10722
rect 26626 10670 26628 10722
rect 26572 10658 26628 10670
rect 26908 10836 26964 11116
rect 27020 11106 27076 11116
rect 27692 11106 27748 11116
rect 26460 10558 26462 10610
rect 26514 10558 26516 10610
rect 26460 10546 26516 10558
rect 26124 10434 26180 10444
rect 26236 10388 26292 10398
rect 26292 10332 26516 10388
rect 26236 10322 26292 10332
rect 25900 10164 25956 10174
rect 25900 10050 25956 10108
rect 25900 9998 25902 10050
rect 25954 9998 25956 10050
rect 25900 9986 25956 9998
rect 26124 9716 26180 9726
rect 26124 9622 26180 9660
rect 26460 9716 26516 10332
rect 26908 10164 26964 10780
rect 27580 10724 27636 10734
rect 27132 10722 27636 10724
rect 27132 10670 27582 10722
rect 27634 10670 27636 10722
rect 27132 10668 27636 10670
rect 26908 10098 26964 10108
rect 27020 10498 27076 10510
rect 27020 10446 27022 10498
rect 27074 10446 27076 10498
rect 26460 9714 26852 9716
rect 26460 9662 26462 9714
rect 26514 9662 26852 9714
rect 26460 9660 26852 9662
rect 26460 9650 26516 9660
rect 25732 9548 25844 9604
rect 25676 9538 25732 9548
rect 26348 9042 26404 9054
rect 26348 8990 26350 9042
rect 26402 8990 26404 9042
rect 26012 8932 26068 8942
rect 26348 8932 26404 8990
rect 26012 8930 26404 8932
rect 26012 8878 26014 8930
rect 26066 8878 26404 8930
rect 26012 8876 26404 8878
rect 25676 8484 25732 8494
rect 26012 8484 26068 8876
rect 25732 8428 26068 8484
rect 25676 8418 25732 8428
rect 24668 8318 24670 8370
rect 24722 8318 24724 8370
rect 24668 8306 24724 8318
rect 26796 8370 26852 9660
rect 26796 8318 26798 8370
rect 26850 8318 26852 8370
rect 26796 8306 26852 8318
rect 24556 7646 24558 7698
rect 24610 7646 24612 7698
rect 24556 7634 24612 7646
rect 23996 7410 24052 7420
rect 24220 7252 24276 7262
rect 24220 7158 24276 7196
rect 26796 7252 26852 7262
rect 23996 6804 24052 6814
rect 23884 6802 24388 6804
rect 23884 6750 23998 6802
rect 24050 6750 24388 6802
rect 23884 6748 24388 6750
rect 23996 6738 24052 6748
rect 23660 6636 23940 6692
rect 23884 6130 23940 6636
rect 23884 6078 23886 6130
rect 23938 6078 23940 6130
rect 23884 6066 23940 6078
rect 24332 6690 24388 6748
rect 24332 6638 24334 6690
rect 24386 6638 24388 6690
rect 23324 5966 23326 6018
rect 23378 5966 23380 6018
rect 23324 5954 23380 5966
rect 23548 5682 23604 5694
rect 23548 5630 23550 5682
rect 23602 5630 23604 5682
rect 23548 5348 23604 5630
rect 23548 5282 23604 5292
rect 23212 5070 23214 5122
rect 23266 5070 23268 5122
rect 23212 5012 23268 5070
rect 23212 4946 23268 4956
rect 23884 5010 23940 5022
rect 23884 4958 23886 5010
rect 23938 4958 23940 5010
rect 23548 4900 23604 4910
rect 23548 4450 23604 4844
rect 23884 4562 23940 4958
rect 23884 4510 23886 4562
rect 23938 4510 23940 4562
rect 23884 4498 23940 4510
rect 24332 4564 24388 6638
rect 25116 6580 25172 6590
rect 25116 6578 25620 6580
rect 25116 6526 25118 6578
rect 25170 6526 25620 6578
rect 25116 6524 25620 6526
rect 25116 6514 25172 6524
rect 25564 6130 25620 6524
rect 25564 6078 25566 6130
rect 25618 6078 25620 6130
rect 25564 6066 25620 6078
rect 25900 5908 25956 5918
rect 26460 5908 26516 5918
rect 25900 5906 26516 5908
rect 25900 5854 25902 5906
rect 25954 5854 26462 5906
rect 26514 5854 26516 5906
rect 25900 5852 26516 5854
rect 25900 5842 25956 5852
rect 26460 5842 26516 5852
rect 26796 5906 26852 7196
rect 27020 6020 27076 10446
rect 27132 9154 27188 10668
rect 27580 10658 27636 10668
rect 28812 10724 28868 10734
rect 27804 10612 27860 10622
rect 27692 10610 27860 10612
rect 27692 10558 27806 10610
rect 27858 10558 27860 10610
rect 27692 10556 27860 10558
rect 27692 10164 27748 10556
rect 27804 10546 27860 10556
rect 27356 10108 27748 10164
rect 27356 10050 27412 10108
rect 27356 9998 27358 10050
rect 27410 9998 27412 10050
rect 27356 9986 27412 9998
rect 27692 9940 27748 9950
rect 27692 9846 27748 9884
rect 28812 9940 28868 10668
rect 28812 9874 28868 9884
rect 27916 9716 27972 9726
rect 27916 9622 27972 9660
rect 28476 9716 28532 9726
rect 28476 9622 28532 9660
rect 27132 9102 27134 9154
rect 27186 9102 27188 9154
rect 27132 9090 27188 9102
rect 27804 8260 27860 8270
rect 27804 7586 27860 8204
rect 28812 7700 28868 7710
rect 28924 7700 28980 12126
rect 28812 7698 28980 7700
rect 28812 7646 28814 7698
rect 28866 7646 28980 7698
rect 28812 7644 28980 7646
rect 29036 12178 29316 12180
rect 29036 12126 29262 12178
rect 29314 12126 29316 12178
rect 29036 12124 29316 12126
rect 28812 7634 28868 7644
rect 27804 7534 27806 7586
rect 27858 7534 27860 7586
rect 27804 7522 27860 7534
rect 28252 7588 28308 7598
rect 28252 7494 28308 7532
rect 27244 7252 27300 7262
rect 27244 6802 27300 7196
rect 27244 6750 27246 6802
rect 27298 6750 27300 6802
rect 27244 6738 27300 6750
rect 28476 7250 28532 7262
rect 28476 7198 28478 7250
rect 28530 7198 28532 7250
rect 28364 6468 28420 6478
rect 27580 6020 27636 6030
rect 27020 6018 27300 6020
rect 27020 5966 27022 6018
rect 27074 5966 27300 6018
rect 27020 5964 27300 5966
rect 27020 5954 27076 5964
rect 26796 5854 26798 5906
rect 26850 5854 26852 5906
rect 26796 5842 26852 5854
rect 27244 5796 27300 5964
rect 27580 5926 27636 5964
rect 28252 6018 28308 6030
rect 28252 5966 28254 6018
rect 28306 5966 28308 6018
rect 27244 5740 27972 5796
rect 26012 5236 26068 5246
rect 26012 5142 26068 5180
rect 27692 5122 27748 5134
rect 27692 5070 27694 5122
rect 27746 5070 27748 5122
rect 27692 5012 27748 5070
rect 27692 4946 27748 4956
rect 27916 5010 27972 5740
rect 28252 5236 28308 5966
rect 28252 5170 28308 5180
rect 27916 4958 27918 5010
rect 27970 4958 27972 5010
rect 27916 4946 27972 4958
rect 28364 5010 28420 6412
rect 28364 4958 28366 5010
rect 28418 4958 28420 5010
rect 28364 4946 28420 4958
rect 28476 5012 28532 7198
rect 28700 6132 28756 6142
rect 29036 6132 29092 12124
rect 29260 12114 29316 12124
rect 29484 12180 29540 12190
rect 29484 12086 29540 12124
rect 29372 12066 29428 12078
rect 29372 12014 29374 12066
rect 29426 12014 29428 12066
rect 29372 11844 29428 12014
rect 29372 11778 29428 11788
rect 29484 10052 29540 10062
rect 29596 10052 29652 15038
rect 29932 14308 29988 14318
rect 29932 13746 29988 14252
rect 30044 14084 30100 15150
rect 30156 14644 30212 14654
rect 30156 14530 30212 14588
rect 30156 14478 30158 14530
rect 30210 14478 30212 14530
rect 30156 14466 30212 14478
rect 30268 14418 30324 14430
rect 30268 14366 30270 14418
rect 30322 14366 30324 14418
rect 30044 14028 30212 14084
rect 29932 13694 29934 13746
rect 29986 13694 29988 13746
rect 29932 13682 29988 13694
rect 30044 13412 30100 13422
rect 30044 12404 30100 13356
rect 30044 12178 30100 12348
rect 30044 12126 30046 12178
rect 30098 12126 30100 12178
rect 30044 12114 30100 12126
rect 29820 11956 29876 11966
rect 30156 11956 30212 14028
rect 30268 13860 30324 14366
rect 30268 13766 30324 13804
rect 30492 12740 30548 16156
rect 30716 16146 30772 16156
rect 31052 14530 31108 14542
rect 31052 14478 31054 14530
rect 31106 14478 31108 14530
rect 31052 14420 31108 14478
rect 30828 13858 30884 13870
rect 30828 13806 30830 13858
rect 30882 13806 30884 13858
rect 30828 13076 30884 13806
rect 31052 13746 31108 14364
rect 31052 13694 31054 13746
rect 31106 13694 31108 13746
rect 31052 13682 31108 13694
rect 31164 14418 31220 14430
rect 31164 14366 31166 14418
rect 31218 14366 31220 14418
rect 30828 13010 30884 13020
rect 31052 13300 31108 13310
rect 30604 12908 30772 12964
rect 30604 12740 30660 12908
rect 30716 12852 30772 12908
rect 30940 12852 30996 12862
rect 30716 12850 30996 12852
rect 30716 12798 30942 12850
rect 30994 12798 30996 12850
rect 30716 12796 30996 12798
rect 30940 12786 30996 12796
rect 30492 12738 30660 12740
rect 30492 12686 30606 12738
rect 30658 12686 30660 12738
rect 30492 12684 30660 12686
rect 30380 12290 30436 12302
rect 30380 12238 30382 12290
rect 30434 12238 30436 12290
rect 30380 12180 30436 12238
rect 30380 12114 30436 12124
rect 29820 11954 30212 11956
rect 29820 11902 29822 11954
rect 29874 11902 30212 11954
rect 29820 11900 30212 11902
rect 29820 11890 29876 11900
rect 30268 11508 30324 11518
rect 30492 11508 30548 12684
rect 30604 12674 30660 12684
rect 30716 12628 30772 12638
rect 30604 12180 30660 12190
rect 30716 12180 30772 12572
rect 31052 12516 31108 13244
rect 31164 12628 31220 14366
rect 31164 12562 31220 12572
rect 31052 12402 31108 12460
rect 31052 12350 31054 12402
rect 31106 12350 31108 12402
rect 31052 12338 31108 12350
rect 30604 12178 30772 12180
rect 30604 12126 30606 12178
rect 30658 12126 30772 12178
rect 30604 12124 30772 12126
rect 30604 12068 30660 12124
rect 30604 12002 30660 12012
rect 30324 11452 30548 11508
rect 30716 11508 30772 11518
rect 30268 11414 30324 11452
rect 30716 11394 30772 11452
rect 30716 11342 30718 11394
rect 30770 11342 30772 11394
rect 30716 11330 30772 11342
rect 31052 11506 31108 11518
rect 31052 11454 31054 11506
rect 31106 11454 31108 11506
rect 29484 10050 29652 10052
rect 29484 9998 29486 10050
rect 29538 9998 29652 10050
rect 29484 9996 29652 9998
rect 31052 10612 31108 11454
rect 29484 9986 29540 9996
rect 29148 9716 29204 9726
rect 29148 8932 29204 9660
rect 29372 9602 29428 9614
rect 29372 9550 29374 9602
rect 29426 9550 29428 9602
rect 29260 8932 29316 8942
rect 29148 8930 29316 8932
rect 29148 8878 29262 8930
rect 29314 8878 29316 8930
rect 29148 8876 29316 8878
rect 29260 8866 29316 8876
rect 29372 7588 29428 9550
rect 29372 7522 29428 7532
rect 29708 9042 29764 9054
rect 29708 8990 29710 9042
rect 29762 8990 29764 9042
rect 29708 8820 29764 8990
rect 30380 8932 30436 8942
rect 30380 8930 30996 8932
rect 30380 8878 30382 8930
rect 30434 8878 30996 8930
rect 30380 8876 30996 8878
rect 30380 8866 30436 8876
rect 29708 7474 29764 8764
rect 30940 8146 30996 8876
rect 30940 8094 30942 8146
rect 30994 8094 30996 8146
rect 30940 8082 30996 8094
rect 29708 7422 29710 7474
rect 29762 7422 29764 7474
rect 29708 7410 29764 7422
rect 30380 7364 30436 7374
rect 30380 7362 30996 7364
rect 30380 7310 30382 7362
rect 30434 7310 30996 7362
rect 30380 7308 30996 7310
rect 30380 7298 30436 7308
rect 29372 6690 29428 6702
rect 29372 6638 29374 6690
rect 29426 6638 29428 6690
rect 29372 6580 29428 6638
rect 29372 6514 29428 6524
rect 29932 6580 29988 6590
rect 29932 6486 29988 6524
rect 30940 6578 30996 7308
rect 30940 6526 30942 6578
rect 30994 6526 30996 6578
rect 30940 6514 30996 6526
rect 29148 6468 29204 6478
rect 29148 6374 29204 6412
rect 29260 6132 29316 6142
rect 29036 6130 29316 6132
rect 29036 6078 29262 6130
rect 29314 6078 29316 6130
rect 29036 6076 29316 6078
rect 28700 6018 28756 6076
rect 29260 6066 29316 6076
rect 31052 6132 31108 10556
rect 31164 10612 31220 10622
rect 31276 10612 31332 20078
rect 31612 20130 31668 20142
rect 31612 20078 31614 20130
rect 31666 20078 31668 20130
rect 31612 20020 31668 20078
rect 31612 19236 31668 19964
rect 31612 19170 31668 19180
rect 31948 20130 32004 26014
rect 32172 24722 32228 24734
rect 32172 24670 32174 24722
rect 32226 24670 32228 24722
rect 32060 24164 32116 24174
rect 32172 24164 32228 24670
rect 32060 24162 32228 24164
rect 32060 24110 32062 24162
rect 32114 24110 32228 24162
rect 32060 24108 32228 24110
rect 32060 24098 32116 24108
rect 32060 23268 32116 23278
rect 32060 23174 32116 23212
rect 32284 23044 32340 27468
rect 32396 27076 32452 27086
rect 32732 27076 32788 27086
rect 32844 27076 32900 27804
rect 33180 27794 33236 27804
rect 33292 29988 33348 29998
rect 33292 27188 33348 29932
rect 33404 29652 33460 30380
rect 33516 29876 33572 30830
rect 33740 30772 33796 30942
rect 34076 30772 34132 30782
rect 33740 30770 34132 30772
rect 33740 30718 34078 30770
rect 34130 30718 34132 30770
rect 33740 30716 34132 30718
rect 34076 30706 34132 30716
rect 34188 30100 34244 31052
rect 34300 30100 34356 30110
rect 34188 30044 34300 30100
rect 34300 30034 34356 30044
rect 33516 29820 33908 29876
rect 33404 29596 33572 29652
rect 33404 29426 33460 29438
rect 33404 29374 33406 29426
rect 33458 29374 33460 29426
rect 33404 29316 33460 29374
rect 33516 29426 33572 29596
rect 33516 29374 33518 29426
rect 33570 29374 33572 29426
rect 33516 29362 33572 29374
rect 33628 29428 33684 29438
rect 33628 29334 33684 29372
rect 33404 29250 33460 29260
rect 33852 28754 33908 29820
rect 34300 29540 34356 29550
rect 34412 29540 34468 31612
rect 34636 31890 34692 32508
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34636 31838 34638 31890
rect 34690 31838 34692 31890
rect 34636 31218 34692 31838
rect 34636 31166 34638 31218
rect 34690 31166 34692 31218
rect 34636 30324 34692 31166
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34748 30436 34804 30446
rect 34748 30342 34804 30380
rect 34636 30258 34692 30268
rect 35420 30212 35476 30222
rect 35476 30156 35588 30212
rect 35420 30146 35476 30156
rect 34860 29988 34916 29998
rect 34860 29894 34916 29932
rect 34972 29986 35028 29998
rect 34972 29934 34974 29986
rect 35026 29934 35028 29986
rect 34972 29876 35028 29934
rect 34972 29810 35028 29820
rect 35084 29988 35140 29998
rect 34300 29538 34468 29540
rect 34300 29486 34302 29538
rect 34354 29486 34468 29538
rect 34300 29484 34468 29486
rect 34300 29474 34356 29484
rect 33852 28702 33854 28754
rect 33906 28702 33908 28754
rect 33852 28690 33908 28702
rect 33852 28420 33908 28430
rect 33852 27970 33908 28364
rect 35084 28084 35140 29932
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35532 28532 35588 30156
rect 35532 28466 35588 28476
rect 35084 28018 35140 28028
rect 33852 27918 33854 27970
rect 33906 27918 33908 27970
rect 33852 27906 33908 27918
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 33404 27188 33460 27198
rect 33292 27186 33460 27188
rect 33292 27134 33406 27186
rect 33458 27134 33460 27186
rect 33292 27132 33460 27134
rect 33404 27122 33460 27132
rect 35532 27188 35588 27198
rect 35532 27094 35588 27132
rect 32452 27074 32900 27076
rect 32452 27022 32734 27074
rect 32786 27022 32900 27074
rect 32452 27020 32900 27022
rect 35644 27076 35700 34972
rect 35868 34914 35924 35644
rect 35868 34862 35870 34914
rect 35922 34862 35924 34914
rect 35868 34850 35924 34862
rect 35980 34914 36036 35868
rect 35980 34862 35982 34914
rect 36034 34862 36036 34914
rect 35980 34850 36036 34862
rect 35756 34802 35812 34814
rect 35756 34750 35758 34802
rect 35810 34750 35812 34802
rect 35756 34580 35812 34750
rect 36092 34580 36148 36204
rect 36204 36194 36260 36204
rect 35756 34524 36148 34580
rect 36204 35698 36260 35710
rect 36204 35646 36206 35698
rect 36258 35646 36260 35698
rect 35756 29650 35812 34524
rect 36204 34244 36260 35646
rect 36428 35028 36484 35038
rect 36428 34934 36484 34972
rect 36204 34178 36260 34188
rect 36764 34580 36820 44156
rect 37548 44100 37604 44110
rect 37548 44006 37604 44044
rect 37996 43762 38052 44268
rect 38668 44230 38724 44268
rect 37996 43710 37998 43762
rect 38050 43710 38052 43762
rect 37996 43698 38052 43710
rect 38108 44210 38164 44222
rect 38108 44158 38110 44210
rect 38162 44158 38164 44210
rect 36876 43540 36932 43550
rect 36876 43446 36932 43484
rect 37548 42980 37604 42990
rect 38108 42980 38164 44158
rect 38444 44212 38500 44222
rect 38444 44118 38500 44156
rect 38780 43988 38836 44492
rect 39116 44100 39172 44110
rect 39116 44006 39172 44044
rect 38668 43932 38836 43988
rect 38556 43314 38612 43326
rect 38556 43262 38558 43314
rect 38610 43262 38612 43314
rect 37548 42978 37940 42980
rect 37548 42926 37550 42978
rect 37602 42926 37940 42978
rect 37548 42924 37940 42926
rect 38108 42924 38276 42980
rect 37548 42914 37604 42924
rect 36988 42756 37044 42766
rect 36988 41972 37044 42700
rect 37660 42756 37716 42766
rect 37660 42662 37716 42700
rect 37548 42530 37604 42542
rect 37548 42478 37550 42530
rect 37602 42478 37604 42530
rect 37548 42308 37604 42478
rect 37548 42242 37604 42252
rect 37884 42082 37940 42924
rect 38108 42754 38164 42766
rect 38108 42702 38110 42754
rect 38162 42702 38164 42754
rect 37996 42196 38052 42206
rect 37996 42102 38052 42140
rect 37884 42030 37886 42082
rect 37938 42030 37940 42082
rect 37884 42018 37940 42030
rect 36988 41906 37044 41916
rect 38108 41860 38164 42702
rect 38220 41970 38276 42924
rect 38556 42868 38612 43262
rect 38556 42802 38612 42812
rect 38668 42866 38724 43932
rect 39228 43876 39284 43886
rect 39004 43652 39060 43662
rect 38780 43596 39004 43652
rect 38780 43538 38836 43596
rect 38780 43486 38782 43538
rect 38834 43486 38836 43538
rect 38780 43474 38836 43486
rect 38668 42814 38670 42866
rect 38722 42814 38724 42866
rect 38668 42756 38724 42814
rect 38780 42868 38836 42878
rect 38780 42774 38836 42812
rect 38668 42690 38724 42700
rect 38220 41918 38222 41970
rect 38274 41918 38276 41970
rect 38220 41906 38276 41918
rect 38444 42642 38500 42654
rect 38444 42590 38446 42642
rect 38498 42590 38500 42642
rect 38108 41794 38164 41804
rect 38444 41858 38500 42590
rect 38780 41972 38836 41982
rect 38892 41972 38948 43596
rect 39004 43586 39060 43596
rect 39228 43538 39284 43820
rect 39228 43486 39230 43538
rect 39282 43486 39284 43538
rect 39228 43474 39284 43486
rect 39004 43426 39060 43438
rect 39004 43374 39006 43426
rect 39058 43374 39060 43426
rect 39004 42196 39060 43374
rect 39340 43428 39396 43438
rect 39228 42756 39284 42766
rect 39340 42756 39396 43372
rect 39228 42754 39396 42756
rect 39228 42702 39230 42754
rect 39282 42702 39396 42754
rect 39228 42700 39396 42702
rect 39228 42690 39284 42700
rect 39004 42130 39060 42140
rect 39452 42084 39508 42094
rect 39116 42082 39508 42084
rect 39116 42030 39454 42082
rect 39506 42030 39508 42082
rect 39116 42028 39508 42030
rect 39004 41972 39060 41982
rect 39116 41972 39172 42028
rect 39452 42018 39508 42028
rect 39564 42084 39620 42094
rect 39564 41990 39620 42028
rect 38892 41970 39172 41972
rect 38892 41918 39006 41970
rect 39058 41918 39172 41970
rect 38892 41916 39172 41918
rect 39676 41972 39732 46620
rect 40012 46340 40068 46350
rect 40012 46002 40068 46284
rect 40012 45950 40014 46002
rect 40066 45950 40068 46002
rect 40012 45668 40068 45950
rect 40012 45602 40068 45612
rect 40012 44324 40068 44334
rect 39900 44100 39956 44110
rect 39788 43652 39844 43662
rect 39788 43558 39844 43596
rect 39900 43428 39956 44044
rect 40012 43762 40068 44268
rect 40124 43876 40180 47628
rect 40348 47348 40404 47358
rect 40348 47254 40404 47292
rect 40236 46674 40292 46686
rect 40236 46622 40238 46674
rect 40290 46622 40292 46674
rect 40236 45668 40292 46622
rect 40460 46676 40516 48300
rect 40460 46610 40516 46620
rect 40460 45668 40516 45678
rect 40236 45666 40516 45668
rect 40236 45614 40462 45666
rect 40514 45614 40516 45666
rect 40236 45612 40516 45614
rect 40460 44996 40516 45612
rect 40124 43820 40292 43876
rect 40012 43710 40014 43762
rect 40066 43710 40068 43762
rect 40012 43698 40068 43710
rect 39900 43372 40068 43428
rect 38444 41806 38446 41858
rect 38498 41806 38500 41858
rect 38444 41076 38500 41806
rect 38444 41010 38500 41020
rect 38556 41860 38612 41870
rect 38556 41748 38612 41804
rect 38668 41748 38724 41758
rect 38556 41746 38724 41748
rect 38556 41694 38670 41746
rect 38722 41694 38724 41746
rect 38556 41692 38724 41694
rect 37548 40962 37604 40974
rect 37548 40910 37550 40962
rect 37602 40910 37604 40962
rect 37212 40516 37268 40526
rect 37548 40516 37604 40910
rect 37268 40460 37604 40516
rect 37212 40402 37268 40460
rect 37884 40404 37940 40414
rect 37212 40350 37214 40402
rect 37266 40350 37268 40402
rect 37212 40338 37268 40350
rect 37772 40402 37940 40404
rect 37772 40350 37886 40402
rect 37938 40350 37940 40402
rect 37772 40348 37940 40350
rect 37772 39620 37828 40348
rect 37884 40338 37940 40348
rect 37772 39526 37828 39564
rect 38108 40290 38164 40302
rect 38108 40238 38110 40290
rect 38162 40238 38164 40290
rect 38108 39618 38164 40238
rect 38220 39732 38276 39742
rect 38556 39732 38612 41692
rect 38668 41682 38724 41692
rect 38780 41524 38836 41916
rect 39004 41906 39060 41916
rect 39676 41906 39732 41916
rect 39788 41970 39844 41982
rect 39788 41918 39790 41970
rect 39842 41918 39844 41970
rect 38220 39730 38612 39732
rect 38220 39678 38222 39730
rect 38274 39678 38612 39730
rect 38220 39676 38612 39678
rect 38668 41468 38836 41524
rect 39228 41860 39284 41870
rect 38220 39666 38276 39676
rect 38108 39566 38110 39618
rect 38162 39566 38164 39618
rect 36988 39060 37044 39070
rect 36988 38966 37044 39004
rect 37212 39060 37268 39070
rect 37772 39060 37828 39070
rect 37212 39058 37604 39060
rect 37212 39006 37214 39058
rect 37266 39006 37604 39058
rect 37212 39004 37604 39006
rect 37212 38994 37268 39004
rect 37324 38836 37380 38846
rect 36988 38834 37380 38836
rect 36988 38782 37326 38834
rect 37378 38782 37380 38834
rect 36988 38780 37380 38782
rect 36988 38276 37044 38780
rect 37324 38770 37380 38780
rect 37548 38612 37604 39004
rect 37828 39004 37940 39060
rect 37772 38966 37828 39004
rect 37660 38836 37716 38846
rect 37660 38742 37716 38780
rect 37548 38556 37828 38612
rect 37100 38500 37156 38510
rect 37100 38276 37156 38444
rect 37324 38276 37380 38286
rect 37100 38274 37380 38276
rect 37100 38222 37326 38274
rect 37378 38222 37380 38274
rect 37100 38220 37380 38222
rect 36988 37268 37044 38220
rect 37324 38210 37380 38220
rect 37660 38276 37716 38286
rect 37660 38182 37716 38220
rect 37660 38050 37716 38062
rect 37660 37998 37662 38050
rect 37714 37998 37716 38050
rect 37660 37940 37716 37998
rect 37660 37874 37716 37884
rect 37436 37268 37492 37278
rect 36988 37266 37492 37268
rect 36988 37214 37438 37266
rect 37490 37214 37492 37266
rect 36988 37212 37492 37214
rect 37436 37202 37492 37212
rect 37772 37266 37828 38556
rect 37884 38050 37940 39004
rect 37884 37998 37886 38050
rect 37938 37998 37940 38050
rect 37884 37986 37940 37998
rect 37996 38834 38052 38846
rect 37996 38782 37998 38834
rect 38050 38782 38052 38834
rect 37772 37214 37774 37266
rect 37826 37214 37828 37266
rect 36988 37042 37044 37054
rect 36988 36990 36990 37042
rect 37042 36990 37044 37042
rect 36988 36260 37044 36990
rect 37772 36708 37828 37214
rect 37772 36642 37828 36652
rect 37996 36482 38052 38782
rect 38108 38274 38164 39566
rect 38556 38834 38612 38846
rect 38556 38782 38558 38834
rect 38610 38782 38612 38834
rect 38556 38500 38612 38782
rect 38668 38668 38724 41468
rect 39228 41188 39284 41804
rect 39228 41094 39284 41132
rect 39788 41186 39844 41918
rect 39788 41134 39790 41186
rect 39842 41134 39844 41186
rect 39788 41122 39844 41134
rect 39900 41188 39956 41198
rect 39900 41094 39956 41132
rect 39452 41076 39508 41086
rect 39452 41074 39732 41076
rect 39452 41022 39454 41074
rect 39506 41022 39732 41074
rect 39452 41020 39732 41022
rect 39452 41010 39508 41020
rect 39676 40626 39732 41020
rect 39788 40964 39844 40974
rect 39788 40870 39844 40908
rect 39676 40574 39678 40626
rect 39730 40574 39732 40626
rect 39676 40562 39732 40574
rect 39900 40516 39956 40526
rect 39900 40422 39956 40460
rect 38780 40404 38836 40414
rect 39452 40404 39508 40414
rect 38780 40402 39508 40404
rect 38780 40350 38782 40402
rect 38834 40350 39454 40402
rect 39506 40350 39508 40402
rect 38780 40348 39508 40350
rect 38780 40338 38836 40348
rect 39452 40338 39508 40348
rect 40012 40180 40068 43372
rect 40124 43314 40180 43326
rect 40124 43262 40126 43314
rect 40178 43262 40180 43314
rect 40124 42754 40180 43262
rect 40236 43204 40292 43820
rect 40460 43764 40516 44940
rect 40572 44100 40628 48524
rect 41468 48356 41524 49758
rect 41468 48290 41524 48300
rect 40908 48244 40964 48254
rect 40908 48150 40964 48188
rect 41580 48132 41636 50092
rect 41692 50082 41748 50092
rect 41804 49812 41860 49822
rect 41804 49718 41860 49756
rect 41916 49698 41972 49710
rect 41916 49646 41918 49698
rect 41970 49646 41972 49698
rect 41916 49028 41972 49646
rect 42028 49252 42084 50428
rect 42364 50148 42420 51326
rect 42700 52050 42756 52062
rect 42700 51998 42702 52050
rect 42754 51998 42756 52050
rect 42700 51380 42756 51998
rect 42700 51314 42756 51324
rect 42588 51268 42644 51278
rect 42588 50708 42644 51212
rect 42476 50596 42532 50606
rect 42476 50502 42532 50540
rect 42364 50082 42420 50092
rect 42588 49922 42644 50652
rect 42700 50482 42756 50494
rect 42700 50430 42702 50482
rect 42754 50430 42756 50482
rect 42700 50034 42756 50430
rect 42812 50260 42868 53228
rect 43484 53172 43540 53676
rect 43708 53620 43764 53630
rect 43484 53106 43540 53116
rect 43596 53564 43708 53620
rect 43484 52948 43540 52958
rect 42924 52164 42980 52174
rect 42924 51378 42980 52108
rect 43148 52164 43204 52174
rect 43148 51602 43204 52108
rect 43260 51940 43316 51950
rect 43260 51846 43316 51884
rect 43148 51550 43150 51602
rect 43202 51550 43204 51602
rect 43148 51538 43204 51550
rect 42924 51326 42926 51378
rect 42978 51326 42980 51378
rect 42924 51314 42980 51326
rect 43260 51380 43316 51390
rect 43260 51286 43316 51324
rect 43260 50482 43316 50494
rect 43260 50430 43262 50482
rect 43314 50430 43316 50482
rect 43260 50428 43316 50430
rect 42812 50194 42868 50204
rect 43036 50372 43316 50428
rect 42700 49982 42702 50034
rect 42754 49982 42756 50034
rect 42700 49970 42756 49982
rect 42588 49870 42590 49922
rect 42642 49870 42644 49922
rect 42588 49858 42644 49870
rect 42476 49812 42532 49822
rect 42028 49196 42308 49252
rect 42140 49028 42196 49038
rect 41972 49026 42196 49028
rect 41972 48974 42142 49026
rect 42194 48974 42196 49026
rect 41972 48972 42196 48974
rect 41916 48934 41972 48972
rect 42140 48962 42196 48972
rect 41244 48076 41636 48132
rect 41692 48356 41748 48366
rect 41020 47458 41076 47470
rect 41020 47406 41022 47458
rect 41074 47406 41076 47458
rect 41020 47348 41076 47406
rect 40908 47292 41020 47348
rect 40908 46674 40964 47292
rect 41020 47282 41076 47292
rect 41244 47346 41300 48076
rect 41244 47294 41246 47346
rect 41298 47294 41300 47346
rect 41244 46786 41300 47294
rect 41244 46734 41246 46786
rect 41298 46734 41300 46786
rect 41244 46722 41300 46734
rect 40908 46622 40910 46674
rect 40962 46622 40964 46674
rect 40908 46610 40964 46622
rect 41468 45780 41524 45790
rect 41356 45724 41468 45780
rect 41244 45668 41300 45678
rect 41132 45666 41300 45668
rect 41132 45614 41246 45666
rect 41298 45614 41300 45666
rect 41132 45612 41300 45614
rect 41020 45108 41076 45118
rect 41132 45108 41188 45612
rect 41244 45602 41300 45612
rect 41020 45106 41188 45108
rect 41020 45054 41022 45106
rect 41074 45054 41188 45106
rect 41020 45052 41188 45054
rect 41244 45332 41300 45342
rect 41356 45332 41412 45724
rect 41468 45714 41524 45724
rect 41580 45780 41636 45790
rect 41692 45780 41748 48300
rect 41916 48244 41972 48254
rect 41804 47348 41860 47358
rect 41804 47254 41860 47292
rect 41916 46898 41972 48188
rect 42140 48242 42196 48254
rect 42140 48190 42142 48242
rect 42194 48190 42196 48242
rect 42140 47570 42196 48190
rect 42140 47518 42142 47570
rect 42194 47518 42196 47570
rect 42140 47506 42196 47518
rect 41916 46846 41918 46898
rect 41970 46846 41972 46898
rect 41916 46834 41972 46846
rect 42028 47348 42084 47358
rect 41804 46676 41860 46686
rect 41804 45892 41860 46620
rect 41804 45798 41860 45836
rect 41580 45778 41748 45780
rect 41580 45726 41582 45778
rect 41634 45726 41748 45778
rect 41580 45724 41748 45726
rect 41580 45714 41636 45724
rect 41692 45556 41748 45724
rect 41692 45490 41748 45500
rect 41244 45330 41412 45332
rect 41244 45278 41246 45330
rect 41298 45278 41412 45330
rect 41244 45276 41412 45278
rect 42028 45332 42084 47292
rect 42140 46228 42196 46238
rect 42140 45892 42196 46172
rect 42252 46116 42308 49196
rect 42476 49026 42532 49756
rect 42588 49140 42644 49150
rect 42588 49046 42644 49084
rect 42476 48974 42478 49026
rect 42530 48974 42532 49026
rect 42476 48354 42532 48974
rect 42476 48302 42478 48354
rect 42530 48302 42532 48354
rect 42476 48290 42532 48302
rect 42700 48244 42756 48254
rect 42700 48150 42756 48188
rect 42924 47572 42980 47582
rect 42924 47458 42980 47516
rect 42924 47406 42926 47458
rect 42978 47406 42980 47458
rect 42924 47394 42980 47406
rect 43036 47570 43092 50372
rect 43148 49924 43204 49934
rect 43148 49922 43428 49924
rect 43148 49870 43150 49922
rect 43202 49870 43428 49922
rect 43148 49868 43428 49870
rect 43148 49858 43204 49868
rect 43036 47518 43038 47570
rect 43090 47518 43092 47570
rect 43036 47068 43092 47518
rect 43372 47570 43428 49868
rect 43484 49812 43540 52892
rect 43596 50596 43652 53564
rect 43708 53554 43764 53564
rect 43820 53508 43876 54350
rect 44156 54404 44212 54414
rect 45500 54404 45556 54414
rect 44156 54402 44548 54404
rect 44156 54350 44158 54402
rect 44210 54350 44548 54402
rect 44156 54348 44548 54350
rect 44156 54338 44212 54348
rect 43820 53442 43876 53452
rect 43932 53508 43988 53518
rect 44156 53508 44212 53518
rect 43932 53506 44156 53508
rect 43932 53454 43934 53506
rect 43986 53454 44156 53506
rect 43932 53452 44156 53454
rect 43932 53442 43988 53452
rect 44156 53442 44212 53452
rect 44380 53284 44436 53294
rect 44156 53172 44212 53182
rect 44044 53170 44212 53172
rect 44044 53118 44158 53170
rect 44210 53118 44212 53170
rect 44044 53116 44212 53118
rect 44044 52836 44100 53116
rect 44156 53106 44212 53116
rect 44380 53058 44436 53228
rect 44380 53006 44382 53058
rect 44434 53006 44436 53058
rect 44380 52948 44436 53006
rect 44492 53060 44548 54348
rect 44828 53842 44884 53854
rect 44828 53790 44830 53842
rect 44882 53790 44884 53842
rect 44828 53284 44884 53790
rect 44828 53218 44884 53228
rect 44828 53060 44884 53070
rect 44492 53058 44884 53060
rect 44492 53006 44494 53058
rect 44546 53006 44830 53058
rect 44882 53006 44884 53058
rect 44492 53004 44884 53006
rect 44492 52994 44548 53004
rect 44828 52994 44884 53004
rect 43932 52780 44100 52836
rect 44156 52892 44436 52948
rect 43708 51492 43764 51502
rect 43932 51492 43988 52780
rect 44044 52162 44100 52174
rect 44044 52110 44046 52162
rect 44098 52110 44100 52162
rect 44044 51716 44100 52110
rect 44156 51716 44212 52892
rect 44940 52722 44996 52734
rect 44940 52670 44942 52722
rect 44994 52670 44996 52722
rect 44940 52388 44996 52670
rect 44940 52332 45332 52388
rect 44940 52164 44996 52174
rect 44940 52070 44996 52108
rect 45164 52162 45220 52174
rect 45164 52110 45166 52162
rect 45218 52110 45220 52162
rect 44268 51940 44324 51950
rect 45164 51940 45220 52110
rect 44268 51938 45220 51940
rect 44268 51886 44270 51938
rect 44322 51886 45220 51938
rect 44268 51884 45220 51886
rect 44268 51874 44324 51884
rect 44156 51660 44324 51716
rect 44044 51650 44100 51660
rect 43764 51436 43988 51492
rect 43708 51398 43764 51436
rect 43932 51044 43988 51054
rect 43596 50540 43764 50596
rect 43596 50370 43652 50382
rect 43596 50318 43598 50370
rect 43650 50318 43652 50370
rect 43596 50260 43652 50318
rect 43596 50194 43652 50204
rect 43596 49812 43652 49822
rect 43484 49810 43652 49812
rect 43484 49758 43598 49810
rect 43650 49758 43652 49810
rect 43484 49756 43652 49758
rect 43596 49746 43652 49756
rect 43708 49588 43764 50540
rect 43820 50484 43876 50522
rect 43820 50418 43876 50428
rect 43932 50148 43988 50988
rect 44044 50820 44100 50830
rect 44044 50482 44100 50764
rect 44156 50708 44212 50718
rect 44156 50594 44212 50652
rect 44156 50542 44158 50594
rect 44210 50542 44212 50594
rect 44156 50530 44212 50542
rect 44044 50430 44046 50482
rect 44098 50430 44100 50482
rect 44044 50418 44100 50430
rect 43932 50092 44100 50148
rect 44044 49810 44100 50092
rect 44044 49758 44046 49810
rect 44098 49758 44100 49810
rect 44044 49746 44100 49758
rect 43372 47518 43374 47570
rect 43426 47518 43428 47570
rect 43372 47506 43428 47518
rect 43596 49532 43764 49588
rect 44156 49698 44212 49710
rect 44156 49646 44158 49698
rect 44210 49646 44212 49698
rect 42924 47012 43092 47068
rect 42476 46900 42532 46910
rect 42476 46806 42532 46844
rect 42700 46676 42756 46686
rect 42252 46050 42308 46060
rect 42364 46674 42756 46676
rect 42364 46622 42702 46674
rect 42754 46622 42756 46674
rect 42364 46620 42756 46622
rect 42364 45892 42420 46620
rect 42700 46610 42756 46620
rect 42924 46676 42980 47012
rect 42924 46582 42980 46620
rect 43260 46674 43316 46686
rect 43260 46622 43262 46674
rect 43314 46622 43316 46674
rect 42812 46562 42868 46574
rect 42812 46510 42814 46562
rect 42866 46510 42868 46562
rect 42140 45890 42420 45892
rect 42140 45838 42142 45890
rect 42194 45838 42420 45890
rect 42140 45836 42420 45838
rect 42140 45826 42196 45836
rect 42140 45668 42196 45678
rect 42140 45574 42196 45612
rect 42140 45332 42196 45342
rect 42028 45330 42196 45332
rect 42028 45278 42142 45330
rect 42194 45278 42196 45330
rect 42028 45276 42196 45278
rect 41020 44884 41076 45052
rect 41020 44818 41076 44828
rect 41244 44660 41300 45276
rect 42140 45266 42196 45276
rect 42364 45330 42420 45836
rect 42476 45892 42532 45902
rect 42812 45892 42868 46510
rect 42476 45890 42868 45892
rect 42476 45838 42478 45890
rect 42530 45838 42868 45890
rect 42476 45836 42868 45838
rect 42924 46004 42980 46014
rect 42476 45826 42532 45836
rect 42812 45668 42868 45678
rect 42924 45668 42980 45948
rect 43036 45892 43092 45902
rect 43260 45892 43316 46622
rect 43092 45836 43316 45892
rect 43036 45798 43092 45836
rect 42364 45278 42366 45330
rect 42418 45278 42420 45330
rect 42364 45266 42420 45278
rect 42476 45666 42980 45668
rect 42476 45614 42814 45666
rect 42866 45614 42980 45666
rect 42476 45612 42980 45614
rect 43260 45668 43316 45678
rect 43316 45612 43540 45668
rect 42252 45108 42308 45118
rect 42252 45014 42308 45052
rect 40796 44604 41300 44660
rect 40796 44324 40852 44604
rect 42252 44548 42308 44558
rect 40796 44230 40852 44268
rect 42028 44492 42252 44548
rect 40572 44034 40628 44044
rect 41020 44100 41076 44110
rect 41020 44098 41300 44100
rect 41020 44046 41022 44098
rect 41074 44046 41300 44098
rect 41020 44044 41300 44046
rect 41020 44034 41076 44044
rect 41244 43876 41300 44044
rect 40460 43698 40516 43708
rect 41132 43764 41188 43774
rect 40236 43138 40292 43148
rect 40460 42980 40516 42990
rect 40124 42702 40126 42754
rect 40178 42702 40180 42754
rect 40124 42690 40180 42702
rect 40236 42978 40516 42980
rect 40236 42926 40462 42978
rect 40514 42926 40516 42978
rect 40236 42924 40516 42926
rect 40124 42532 40180 42542
rect 40124 42194 40180 42476
rect 40124 42142 40126 42194
rect 40178 42142 40180 42194
rect 40124 42130 40180 42142
rect 40236 42082 40292 42924
rect 40460 42914 40516 42924
rect 40572 42868 40628 42878
rect 40572 42774 40628 42812
rect 40236 42030 40238 42082
rect 40290 42030 40292 42082
rect 40236 42018 40292 42030
rect 41020 41972 41076 41982
rect 41020 41878 41076 41916
rect 40236 41860 40292 41870
rect 40124 41748 40180 41758
rect 40124 41654 40180 41692
rect 40124 41412 40180 41422
rect 40124 41298 40180 41356
rect 40124 41246 40126 41298
rect 40178 41246 40180 41298
rect 40124 41234 40180 41246
rect 40124 40964 40180 40974
rect 40124 40514 40180 40908
rect 40124 40462 40126 40514
rect 40178 40462 40180 40514
rect 40124 40450 40180 40462
rect 39340 40124 40068 40180
rect 39228 38834 39284 38846
rect 39228 38782 39230 38834
rect 39282 38782 39284 38834
rect 38668 38612 38948 38668
rect 38556 38444 38724 38500
rect 38108 38222 38110 38274
rect 38162 38222 38164 38274
rect 38108 38210 38164 38222
rect 38220 38276 38276 38286
rect 38276 38220 38500 38276
rect 38220 38210 38276 38220
rect 37996 36430 37998 36482
rect 38050 36430 38052 36482
rect 37996 36418 38052 36430
rect 38444 36482 38500 38220
rect 38668 38052 38724 38444
rect 38780 38052 38836 38062
rect 38668 38050 38836 38052
rect 38668 37998 38782 38050
rect 38834 37998 38836 38050
rect 38668 37996 38836 37998
rect 38780 37940 38836 37996
rect 38780 37268 38836 37884
rect 38780 37174 38836 37212
rect 38892 37044 38948 38612
rect 39228 37154 39284 38782
rect 39228 37102 39230 37154
rect 39282 37102 39284 37154
rect 39228 37044 39284 37102
rect 38444 36430 38446 36482
rect 38498 36430 38500 36482
rect 38108 36260 38164 36270
rect 36988 36258 38164 36260
rect 36988 36206 38110 36258
rect 38162 36206 38164 36258
rect 36988 36204 38164 36206
rect 38108 36194 38164 36204
rect 38220 36258 38276 36270
rect 38220 36206 38222 36258
rect 38274 36206 38276 36258
rect 36988 35924 37044 35934
rect 37996 35924 38052 35934
rect 36876 35810 36932 35822
rect 36876 35758 36878 35810
rect 36930 35758 36932 35810
rect 36876 35588 36932 35758
rect 36876 35522 36932 35532
rect 36428 33458 36484 33470
rect 36428 33406 36430 33458
rect 36482 33406 36484 33458
rect 36428 32676 36484 33406
rect 36428 32610 36484 32620
rect 35756 29598 35758 29650
rect 35810 29598 35812 29650
rect 35756 29586 35812 29598
rect 35868 30210 35924 30222
rect 35868 30158 35870 30210
rect 35922 30158 35924 30210
rect 35868 30100 35924 30158
rect 36428 30100 36484 30110
rect 35868 29428 35924 30044
rect 35868 29334 35924 29372
rect 35980 30044 36428 30100
rect 35980 28754 36036 30044
rect 36428 30006 36484 30044
rect 36316 29540 36372 29550
rect 36316 29426 36372 29484
rect 36316 29374 36318 29426
rect 36370 29374 36372 29426
rect 36316 29362 36372 29374
rect 35980 28702 35982 28754
rect 36034 28702 36036 28754
rect 35980 28690 36036 28702
rect 36428 28532 36484 28542
rect 36428 28084 36484 28476
rect 36428 28082 36596 28084
rect 36428 28030 36430 28082
rect 36482 28030 36596 28082
rect 36428 28028 36596 28030
rect 36428 28018 36484 28028
rect 35980 27748 36036 27758
rect 35980 27654 36036 27692
rect 36428 27412 36484 27422
rect 36428 27186 36484 27356
rect 36428 27134 36430 27186
rect 36482 27134 36484 27186
rect 36428 27122 36484 27134
rect 35868 27076 35924 27086
rect 35644 27074 35924 27076
rect 35644 27022 35870 27074
rect 35922 27022 35924 27074
rect 35644 27020 35924 27022
rect 32396 26178 32452 27020
rect 32732 27010 32788 27020
rect 35532 26516 35588 26526
rect 35644 26516 35700 27020
rect 35868 27010 35924 27020
rect 36540 27076 36596 28028
rect 36764 27412 36820 34524
rect 36988 32900 37044 35868
rect 37772 35922 38052 35924
rect 37772 35870 37998 35922
rect 38050 35870 38052 35922
rect 37772 35868 38052 35870
rect 37100 34916 37156 34926
rect 37100 34244 37156 34860
rect 37772 34580 37828 35868
rect 37996 35858 38052 35868
rect 37884 35698 37940 35710
rect 37884 35646 37886 35698
rect 37938 35646 37940 35698
rect 37884 35252 37940 35646
rect 38108 35700 38164 35710
rect 38220 35700 38276 36206
rect 38332 36260 38388 36270
rect 38332 36166 38388 36204
rect 38332 35700 38388 35710
rect 38220 35698 38388 35700
rect 38220 35646 38334 35698
rect 38386 35646 38388 35698
rect 38220 35644 38388 35646
rect 37996 35476 38052 35486
rect 38108 35476 38164 35644
rect 38332 35634 38388 35644
rect 37996 35474 38164 35476
rect 37996 35422 37998 35474
rect 38050 35422 38164 35474
rect 37996 35420 38164 35422
rect 37996 35410 38052 35420
rect 38444 35364 38500 36430
rect 38668 36988 38948 37044
rect 39004 36988 39284 37044
rect 38556 35476 38612 35486
rect 38668 35476 38724 36988
rect 38892 36372 38948 36382
rect 39004 36372 39060 36988
rect 39228 36932 39284 36988
rect 39340 37044 39396 40124
rect 40236 40068 40292 41804
rect 40908 41748 40964 41758
rect 40348 41746 40964 41748
rect 40348 41694 40910 41746
rect 40962 41694 40964 41746
rect 40348 41692 40964 41694
rect 40348 41186 40404 41692
rect 40908 41682 40964 41692
rect 41132 41524 41188 43708
rect 41244 41748 41300 43820
rect 41244 41682 41300 41692
rect 41356 42644 41412 42654
rect 41132 41468 41300 41524
rect 41132 41300 41188 41310
rect 40348 41134 40350 41186
rect 40402 41134 40404 41186
rect 40348 41122 40404 41134
rect 40684 41244 41132 41300
rect 40572 40962 40628 40974
rect 40572 40910 40574 40962
rect 40626 40910 40628 40962
rect 40572 40516 40628 40910
rect 40572 40450 40628 40460
rect 39900 40012 40292 40068
rect 39900 39284 39956 40012
rect 40348 39844 40404 39854
rect 39900 39218 39956 39228
rect 40012 39618 40068 39630
rect 40012 39566 40014 39618
rect 40066 39566 40068 39618
rect 39564 38948 39620 38958
rect 40012 38948 40068 39566
rect 40124 39508 40180 39518
rect 40124 39506 40292 39508
rect 40124 39454 40126 39506
rect 40178 39454 40292 39506
rect 40124 39452 40292 39454
rect 40124 39442 40180 39452
rect 40236 39058 40292 39452
rect 40236 39006 40238 39058
rect 40290 39006 40292 39058
rect 40124 38948 40180 38958
rect 39564 38946 40180 38948
rect 39564 38894 39566 38946
rect 39618 38894 40126 38946
rect 40178 38894 40180 38946
rect 39564 38892 40180 38894
rect 39564 38882 39620 38892
rect 40124 38882 40180 38892
rect 39452 38834 39508 38846
rect 39452 38782 39454 38834
rect 39506 38782 39508 38834
rect 39452 38276 39508 38782
rect 39564 38276 39620 38286
rect 39452 38274 39620 38276
rect 39452 38222 39566 38274
rect 39618 38222 39620 38274
rect 39452 38220 39620 38222
rect 39452 37268 39508 37278
rect 39452 37174 39508 37212
rect 39564 37044 39620 38220
rect 39788 37938 39844 37950
rect 39788 37886 39790 37938
rect 39842 37886 39844 37938
rect 39676 37044 39732 37054
rect 39564 37042 39732 37044
rect 39564 36990 39678 37042
rect 39730 36990 39732 37042
rect 39564 36988 39732 36990
rect 39340 36978 39396 36988
rect 39228 36866 39284 36876
rect 39564 36482 39620 36494
rect 39564 36430 39566 36482
rect 39618 36430 39620 36482
rect 38556 35474 38724 35476
rect 38556 35422 38558 35474
rect 38610 35422 38724 35474
rect 38556 35420 38724 35422
rect 38780 36370 39060 36372
rect 38780 36318 38894 36370
rect 38946 36318 39060 36370
rect 38780 36316 39060 36318
rect 39116 36372 39172 36382
rect 38556 35410 38612 35420
rect 38108 35308 38500 35364
rect 38108 35252 38164 35308
rect 37884 35196 38164 35252
rect 38780 35026 38836 36316
rect 38892 36306 38948 36316
rect 38892 35700 38948 35710
rect 38892 35606 38948 35644
rect 38780 34974 38782 35026
rect 38834 34974 38836 35026
rect 38780 34962 38836 34974
rect 38220 34916 38276 34926
rect 38220 34822 38276 34860
rect 38668 34914 38724 34926
rect 38668 34862 38670 34914
rect 38722 34862 38724 34914
rect 37772 34524 38052 34580
rect 37100 34130 37156 34188
rect 37996 34244 38052 34524
rect 37996 34150 38052 34188
rect 37100 34078 37102 34130
rect 37154 34078 37156 34130
rect 37100 34066 37156 34078
rect 37660 34130 37716 34142
rect 37660 34078 37662 34130
rect 37714 34078 37716 34130
rect 37660 33796 37716 34078
rect 38444 34130 38500 34142
rect 38444 34078 38446 34130
rect 38498 34078 38500 34130
rect 38444 33796 38500 34078
rect 38668 34132 38724 34862
rect 38668 34020 38724 34076
rect 38780 34020 38836 34030
rect 38668 34018 38836 34020
rect 38668 33966 38782 34018
rect 38834 33966 38836 34018
rect 38668 33964 38836 33966
rect 38780 33954 38836 33964
rect 37660 33740 38500 33796
rect 37100 33124 37156 33134
rect 37548 33124 37604 33134
rect 37156 33122 37604 33124
rect 37156 33070 37550 33122
rect 37602 33070 37604 33122
rect 37156 33068 37604 33070
rect 37100 33030 37156 33068
rect 37548 33058 37604 33068
rect 37660 32900 37716 33740
rect 39116 33236 39172 36316
rect 39228 36260 39284 36270
rect 39228 36166 39284 36204
rect 39228 35700 39284 35710
rect 39228 35698 39508 35700
rect 39228 35646 39230 35698
rect 39282 35646 39508 35698
rect 39228 35644 39508 35646
rect 39228 35634 39284 35644
rect 39340 34914 39396 34926
rect 39340 34862 39342 34914
rect 39394 34862 39396 34914
rect 39340 33570 39396 34862
rect 39452 34130 39508 35644
rect 39452 34078 39454 34130
rect 39506 34078 39508 34130
rect 39452 33908 39508 34078
rect 39452 33842 39508 33852
rect 39564 35140 39620 36430
rect 39340 33518 39342 33570
rect 39394 33518 39396 33570
rect 39340 33506 39396 33518
rect 39452 33348 39508 33358
rect 39564 33348 39620 35084
rect 39676 35026 39732 36988
rect 39788 36932 39844 37886
rect 40124 37492 40180 37502
rect 40236 37492 40292 39006
rect 40124 37490 40292 37492
rect 40124 37438 40126 37490
rect 40178 37438 40292 37490
rect 40124 37436 40292 37438
rect 40124 37426 40180 37436
rect 39788 36866 39844 36876
rect 40124 35812 40180 35822
rect 39676 34974 39678 35026
rect 39730 34974 39732 35026
rect 39676 34962 39732 34974
rect 40012 35756 40124 35812
rect 39788 34802 39844 34814
rect 39788 34750 39790 34802
rect 39842 34750 39844 34802
rect 39788 34132 39844 34750
rect 39788 34130 39956 34132
rect 39788 34078 39790 34130
rect 39842 34078 39956 34130
rect 39788 34076 39956 34078
rect 39788 34066 39844 34076
rect 39900 33570 39956 34076
rect 39900 33518 39902 33570
rect 39954 33518 39956 33570
rect 39900 33506 39956 33518
rect 39452 33346 39620 33348
rect 39452 33294 39454 33346
rect 39506 33294 39620 33346
rect 39452 33292 39620 33294
rect 39788 33348 39844 33358
rect 40012 33348 40068 35756
rect 40124 35718 40180 35756
rect 39788 33346 40068 33348
rect 39788 33294 39790 33346
rect 39842 33294 40068 33346
rect 39788 33292 40068 33294
rect 40124 34914 40180 34926
rect 40124 34862 40126 34914
rect 40178 34862 40180 34914
rect 39452 33282 39508 33292
rect 39788 33282 39844 33292
rect 39340 33236 39396 33246
rect 39116 33234 39396 33236
rect 39116 33182 39342 33234
rect 39394 33182 39396 33234
rect 39116 33180 39396 33182
rect 39340 33170 39396 33180
rect 36988 32844 37156 32900
rect 36988 31780 37044 31790
rect 36988 31686 37044 31724
rect 37100 31444 37156 32844
rect 37548 32844 37716 32900
rect 37212 32676 37268 32686
rect 37212 31666 37268 32620
rect 37324 32452 37380 32462
rect 37548 32452 37604 32844
rect 39788 32788 39844 32798
rect 39564 32786 39844 32788
rect 39564 32734 39790 32786
rect 39842 32734 39844 32786
rect 39564 32732 39844 32734
rect 37660 32676 37716 32686
rect 37660 32582 37716 32620
rect 39116 32676 39172 32686
rect 39564 32676 39620 32732
rect 39788 32722 39844 32732
rect 39116 32674 39620 32676
rect 39116 32622 39118 32674
rect 39170 32622 39620 32674
rect 39116 32620 39620 32622
rect 39116 32610 39172 32620
rect 38780 32562 38836 32574
rect 38780 32510 38782 32562
rect 38834 32510 38836 32562
rect 37324 32450 37604 32452
rect 37324 32398 37326 32450
rect 37378 32398 37604 32450
rect 37324 32396 37604 32398
rect 38108 32450 38164 32462
rect 38108 32398 38110 32450
rect 38162 32398 38164 32450
rect 37324 32386 37380 32396
rect 37884 31778 37940 31790
rect 37884 31726 37886 31778
rect 37938 31726 37940 31778
rect 37212 31614 37214 31666
rect 37266 31614 37268 31666
rect 37212 31602 37268 31614
rect 37324 31666 37380 31678
rect 37324 31614 37326 31666
rect 37378 31614 37380 31666
rect 37324 31556 37380 31614
rect 37660 31668 37716 31678
rect 37660 31574 37716 31612
rect 37324 31490 37380 31500
rect 37884 31556 37940 31726
rect 38108 31780 38164 32398
rect 38108 31724 38388 31780
rect 38108 31668 38164 31724
rect 38108 31602 38164 31612
rect 37100 31388 37268 31444
rect 37100 29540 37156 29550
rect 36988 29316 37044 29326
rect 36988 28754 37044 29260
rect 36988 28702 36990 28754
rect 37042 28702 37044 28754
rect 36988 28084 37044 28702
rect 36988 28018 37044 28028
rect 37100 27970 37156 29484
rect 37212 29092 37268 31388
rect 37548 31220 37604 31230
rect 37548 31126 37604 31164
rect 37324 31108 37380 31118
rect 37772 31108 37828 31118
rect 37324 31014 37380 31052
rect 37660 31106 37828 31108
rect 37660 31054 37774 31106
rect 37826 31054 37828 31106
rect 37660 31052 37828 31054
rect 37884 31108 37940 31500
rect 38220 31554 38276 31566
rect 38220 31502 38222 31554
rect 38274 31502 38276 31554
rect 38108 31108 38164 31118
rect 37884 31106 38164 31108
rect 37884 31054 38110 31106
rect 38162 31054 38164 31106
rect 37884 31052 38164 31054
rect 37324 30100 37380 30110
rect 37660 30100 37716 31052
rect 37772 31042 37828 31052
rect 38108 31042 38164 31052
rect 38220 31108 38276 31502
rect 38220 31042 38276 31052
rect 38332 30994 38388 31724
rect 38332 30942 38334 30994
rect 38386 30942 38388 30994
rect 38332 30930 38388 30942
rect 38556 31778 38612 31790
rect 38556 31726 38558 31778
rect 38610 31726 38612 31778
rect 37884 30770 37940 30782
rect 37884 30718 37886 30770
rect 37938 30718 37940 30770
rect 37324 30098 37716 30100
rect 37324 30046 37326 30098
rect 37378 30046 37716 30098
rect 37324 30044 37716 30046
rect 37772 30210 37828 30222
rect 37772 30158 37774 30210
rect 37826 30158 37828 30210
rect 37772 30100 37828 30158
rect 37884 30212 37940 30718
rect 38220 30324 38276 30334
rect 38220 30230 38276 30268
rect 37884 30146 37940 30156
rect 37324 29652 37380 30044
rect 37772 30034 37828 30044
rect 37324 29586 37380 29596
rect 38556 29652 38612 31726
rect 38780 31780 38836 32510
rect 38780 31686 38836 31724
rect 38892 31668 38948 31678
rect 38892 31108 38948 31612
rect 39228 31220 39284 32620
rect 39676 32562 39732 32574
rect 39676 32510 39678 32562
rect 39730 32510 39732 32562
rect 39340 31780 39396 31790
rect 39340 31686 39396 31724
rect 39676 31668 39732 32510
rect 39676 31602 39732 31612
rect 39788 32338 39844 32350
rect 39788 32286 39790 32338
rect 39842 32286 39844 32338
rect 39788 31444 39844 32286
rect 39788 31378 39844 31388
rect 39900 31778 39956 31790
rect 39900 31726 39902 31778
rect 39954 31726 39956 31778
rect 39900 31220 39956 31726
rect 40012 31220 40068 31230
rect 39900 31218 40068 31220
rect 39900 31166 40014 31218
rect 40066 31166 40068 31218
rect 39900 31164 40068 31166
rect 39228 31154 39284 31164
rect 40012 31154 40068 31164
rect 38892 31042 38948 31052
rect 39116 30996 39172 31006
rect 39116 30994 39284 30996
rect 39116 30942 39118 30994
rect 39170 30942 39284 30994
rect 39116 30940 39284 30942
rect 39116 30930 39172 30940
rect 39228 30324 39284 30940
rect 38780 30212 38836 30222
rect 38780 30118 38836 30156
rect 39116 30210 39172 30222
rect 39116 30158 39118 30210
rect 39170 30158 39172 30210
rect 38556 29586 38612 29596
rect 37436 29538 37492 29550
rect 37436 29486 37438 29538
rect 37490 29486 37492 29538
rect 37324 29316 37380 29326
rect 37436 29316 37492 29486
rect 38780 29540 38836 29550
rect 38836 29484 38948 29540
rect 38780 29474 38836 29484
rect 37380 29260 37492 29316
rect 38892 29316 38948 29484
rect 38892 29314 39060 29316
rect 38892 29262 38894 29314
rect 38946 29262 39060 29314
rect 38892 29260 39060 29262
rect 37324 29250 37380 29260
rect 38892 29250 38948 29260
rect 38332 29204 38388 29214
rect 38668 29204 38724 29214
rect 38332 29202 38612 29204
rect 38332 29150 38334 29202
rect 38386 29150 38612 29202
rect 38332 29148 38612 29150
rect 38332 29138 38388 29148
rect 37212 29036 37604 29092
rect 37436 28642 37492 28654
rect 37436 28590 37438 28642
rect 37490 28590 37492 28642
rect 37100 27918 37102 27970
rect 37154 27918 37156 27970
rect 37100 27906 37156 27918
rect 37324 28532 37380 28542
rect 37324 27858 37380 28476
rect 37324 27806 37326 27858
rect 37378 27806 37380 27858
rect 37324 27794 37380 27806
rect 37436 28420 37492 28590
rect 36764 27346 36820 27356
rect 37212 27636 37268 27646
rect 36988 27076 37044 27086
rect 36540 27074 37044 27076
rect 36540 27022 36990 27074
rect 37042 27022 37044 27074
rect 36540 27020 37044 27022
rect 35532 26514 35700 26516
rect 35532 26462 35534 26514
rect 35586 26462 35700 26514
rect 35532 26460 35700 26462
rect 35980 26516 36036 26526
rect 36428 26516 36484 26526
rect 36540 26516 36596 27020
rect 36988 27010 37044 27020
rect 37100 26964 37156 26974
rect 35980 26514 36596 26516
rect 35980 26462 35982 26514
rect 36034 26462 36430 26514
rect 36482 26462 36596 26514
rect 35980 26460 36596 26462
rect 36764 26852 37156 26908
rect 35532 26450 35588 26460
rect 35980 26450 36036 26460
rect 32396 26126 32398 26178
rect 32450 26126 32452 26178
rect 32396 25060 32452 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 33628 25284 33684 25294
rect 33628 25282 33796 25284
rect 33628 25230 33630 25282
rect 33682 25230 33796 25282
rect 33628 25228 33796 25230
rect 33628 25218 33684 25228
rect 32396 25004 32676 25060
rect 32508 24836 32564 24846
rect 32508 24742 32564 24780
rect 32620 24724 32676 25004
rect 33180 24724 33236 24734
rect 32620 24722 33348 24724
rect 32620 24670 33182 24722
rect 33234 24670 33348 24722
rect 32620 24668 33348 24670
rect 33180 24658 33236 24668
rect 32396 23940 32452 23950
rect 32396 23846 32452 23884
rect 32620 23826 32676 23838
rect 32620 23774 32622 23826
rect 32674 23774 32676 23826
rect 32620 23492 32676 23774
rect 33180 23828 33236 23838
rect 33180 23734 33236 23772
rect 32620 23426 32676 23436
rect 33180 23268 33236 23278
rect 33180 23174 33236 23212
rect 32508 23044 32564 23054
rect 32284 23042 32564 23044
rect 32284 22990 32510 23042
rect 32562 22990 32564 23042
rect 32284 22988 32564 22990
rect 32508 22260 32564 22988
rect 33292 22484 33348 24668
rect 33628 23938 33684 23950
rect 33628 23886 33630 23938
rect 33682 23886 33684 23938
rect 33516 22932 33572 22942
rect 33292 22418 33348 22428
rect 33404 22876 33516 22932
rect 32508 22194 32564 22204
rect 33180 22372 33236 22382
rect 32396 21700 32452 21710
rect 32284 21588 32340 21598
rect 32284 21494 32340 21532
rect 32060 20916 32116 20926
rect 32060 20822 32116 20860
rect 32396 20580 32452 21644
rect 33180 21698 33236 22316
rect 33180 21646 33182 21698
rect 33234 21646 33236 21698
rect 33180 21634 33236 21646
rect 33292 22260 33348 22270
rect 33068 21364 33124 21374
rect 32396 20486 32452 20524
rect 32508 21362 33124 21364
rect 32508 21310 33070 21362
rect 33122 21310 33124 21362
rect 32508 21308 33124 21310
rect 31948 20078 31950 20130
rect 32002 20078 32004 20130
rect 31388 17442 31444 17454
rect 31388 17390 31390 17442
rect 31442 17390 31444 17442
rect 31388 16994 31444 17390
rect 31388 16942 31390 16994
rect 31442 16942 31444 16994
rect 31388 16884 31444 16942
rect 31724 17442 31780 17454
rect 31724 17390 31726 17442
rect 31778 17390 31780 17442
rect 31724 16884 31780 17390
rect 31836 16884 31892 16894
rect 31388 16882 31892 16884
rect 31388 16830 31838 16882
rect 31890 16830 31892 16882
rect 31388 16828 31892 16830
rect 31388 16436 31444 16446
rect 31388 15428 31444 16380
rect 31836 16098 31892 16828
rect 31836 16046 31838 16098
rect 31890 16046 31892 16098
rect 31836 16034 31892 16046
rect 31388 13074 31444 15372
rect 31948 15148 32004 20078
rect 32284 20130 32340 20142
rect 32284 20078 32286 20130
rect 32338 20078 32340 20130
rect 32284 19460 32340 20078
rect 32284 19394 32340 19404
rect 32060 18676 32116 18686
rect 32060 17554 32116 18620
rect 32396 18676 32452 18686
rect 32396 18582 32452 18620
rect 32508 18562 32564 21308
rect 33068 21298 33124 21308
rect 32620 20802 32676 20814
rect 32620 20750 32622 20802
rect 32674 20750 32676 20802
rect 32620 20020 32676 20750
rect 33292 20802 33348 22204
rect 33292 20750 33294 20802
rect 33346 20750 33348 20802
rect 33292 20692 33348 20750
rect 32620 19954 32676 19964
rect 32956 20636 33348 20692
rect 33404 21812 33460 22876
rect 33516 22838 33572 22876
rect 33628 22260 33684 23886
rect 33740 23940 33796 25228
rect 36428 24948 36484 26460
rect 36764 26402 36820 26852
rect 36764 26350 36766 26402
rect 36818 26350 36820 26402
rect 36764 26338 36820 26350
rect 36876 26740 36932 26750
rect 36876 26290 36932 26684
rect 36876 26238 36878 26290
rect 36930 26238 36932 26290
rect 36876 26068 36932 26238
rect 37100 26292 37156 26302
rect 37212 26292 37268 27580
rect 37436 27188 37492 28364
rect 37436 27122 37492 27132
rect 37548 26908 37604 29036
rect 38556 28868 38612 29148
rect 38668 29110 38724 29148
rect 38556 28812 38948 28868
rect 38444 28756 38500 28766
rect 38444 28662 38500 28700
rect 37996 28644 38052 28654
rect 37660 28642 38052 28644
rect 37660 28590 37998 28642
rect 38050 28590 38052 28642
rect 37660 28588 38052 28590
rect 37660 28082 37716 28588
rect 37996 28578 38052 28588
rect 38892 28642 38948 28812
rect 38892 28590 38894 28642
rect 38946 28590 38948 28642
rect 38892 28578 38948 28590
rect 38108 28530 38164 28542
rect 38108 28478 38110 28530
rect 38162 28478 38164 28530
rect 37660 28030 37662 28082
rect 37714 28030 37716 28082
rect 37660 28018 37716 28030
rect 37996 28084 38052 28094
rect 38108 28084 38164 28478
rect 39004 28420 39060 29260
rect 39116 28756 39172 30158
rect 39228 28868 39284 30268
rect 39452 30994 39508 31006
rect 39452 30942 39454 30994
rect 39506 30942 39508 30994
rect 39452 29988 39508 30942
rect 39564 30884 39620 30894
rect 39788 30884 39844 30894
rect 39564 30882 39788 30884
rect 39564 30830 39566 30882
rect 39618 30830 39788 30882
rect 39564 30828 39788 30830
rect 39564 30818 39620 30828
rect 39788 30210 39844 30828
rect 40012 30436 40068 30446
rect 39788 30158 39790 30210
rect 39842 30158 39844 30210
rect 39788 30146 39844 30158
rect 39900 30380 40012 30436
rect 39452 29932 39620 29988
rect 39564 29428 39620 29932
rect 39228 28802 39284 28812
rect 39452 28868 39508 28878
rect 39116 28690 39172 28700
rect 39452 28530 39508 28812
rect 39452 28478 39454 28530
rect 39506 28478 39508 28530
rect 39452 28466 39508 28478
rect 39564 28530 39620 29372
rect 39676 29426 39732 29438
rect 39676 29374 39678 29426
rect 39730 29374 39732 29426
rect 39676 28756 39732 29374
rect 39676 28690 39732 28700
rect 39788 28644 39844 28654
rect 39900 28644 39956 30380
rect 40012 30370 40068 30380
rect 40124 30322 40180 34862
rect 40348 34242 40404 39788
rect 40460 39060 40516 39070
rect 40460 38966 40516 39004
rect 40684 38276 40740 41244
rect 41132 41234 41188 41244
rect 40908 41076 40964 41086
rect 40796 40962 40852 40974
rect 40796 40910 40798 40962
rect 40850 40910 40852 40962
rect 40796 40516 40852 40910
rect 40796 40450 40852 40460
rect 40908 39844 40964 41020
rect 41244 41076 41300 41468
rect 41244 41010 41300 41020
rect 41356 41074 41412 42588
rect 41468 42532 41524 42542
rect 41468 42438 41524 42476
rect 41468 42084 41524 42094
rect 41468 41748 41524 42028
rect 41468 41682 41524 41692
rect 41580 41972 41636 41982
rect 41356 41022 41358 41074
rect 41410 41022 41412 41074
rect 41356 41010 41412 41022
rect 41468 41074 41524 41086
rect 41468 41022 41470 41074
rect 41522 41022 41524 41074
rect 41020 40964 41076 40974
rect 41020 40626 41076 40908
rect 41020 40574 41022 40626
rect 41074 40574 41076 40626
rect 41020 40562 41076 40574
rect 41132 40962 41188 40974
rect 41132 40910 41134 40962
rect 41186 40910 41188 40962
rect 41020 39844 41076 39854
rect 40908 39842 41076 39844
rect 40908 39790 41022 39842
rect 41074 39790 41076 39842
rect 40908 39788 41076 39790
rect 41020 39778 41076 39788
rect 41132 39618 41188 40910
rect 41468 39844 41524 41022
rect 41468 39778 41524 39788
rect 41132 39566 41134 39618
rect 41186 39566 41188 39618
rect 41132 39554 41188 39566
rect 41244 39730 41300 39742
rect 41244 39678 41246 39730
rect 41298 39678 41300 39730
rect 41020 39172 41076 39182
rect 41020 39058 41076 39116
rect 41020 39006 41022 39058
rect 41074 39006 41076 39058
rect 41020 38994 41076 39006
rect 40572 38164 40628 38174
rect 40684 38164 40740 38220
rect 40572 38162 40740 38164
rect 40572 38110 40574 38162
rect 40626 38110 40740 38162
rect 40572 38108 40740 38110
rect 41132 38836 41188 38846
rect 40572 38098 40628 38108
rect 41132 36820 41188 38780
rect 41244 37044 41300 39678
rect 41356 39284 41412 39294
rect 41356 38946 41412 39228
rect 41356 38894 41358 38946
rect 41410 38894 41412 38946
rect 41356 38882 41412 38894
rect 41468 38948 41524 38958
rect 41580 38948 41636 41916
rect 41804 41970 41860 41982
rect 41804 41918 41806 41970
rect 41858 41918 41860 41970
rect 41804 41300 41860 41918
rect 42028 41970 42084 44492
rect 42252 44482 42308 44492
rect 42476 44322 42532 45612
rect 42812 45602 42868 45612
rect 43260 45602 43316 45612
rect 43148 45332 43204 45342
rect 42812 45330 43204 45332
rect 42812 45278 43150 45330
rect 43202 45278 43204 45330
rect 42812 45276 43204 45278
rect 42812 45106 42868 45276
rect 43148 45266 43204 45276
rect 43484 45330 43540 45612
rect 43484 45278 43486 45330
rect 43538 45278 43540 45330
rect 43372 45220 43428 45230
rect 43036 45108 43092 45118
rect 42812 45054 42814 45106
rect 42866 45054 42868 45106
rect 42812 45042 42868 45054
rect 42924 45106 43092 45108
rect 42924 45054 43038 45106
rect 43090 45054 43092 45106
rect 42924 45052 43092 45054
rect 42476 44270 42478 44322
rect 42530 44270 42532 44322
rect 42476 44212 42532 44270
rect 42476 44146 42532 44156
rect 42924 43876 42980 45052
rect 43036 45042 43092 45052
rect 43260 45106 43316 45118
rect 43260 45054 43262 45106
rect 43314 45054 43316 45106
rect 43036 44772 43092 44782
rect 43036 44434 43092 44716
rect 43260 44548 43316 45054
rect 43260 44482 43316 44492
rect 43036 44382 43038 44434
rect 43090 44382 43092 44434
rect 43036 44370 43092 44382
rect 43372 44434 43428 45164
rect 43372 44382 43374 44434
rect 43426 44382 43428 44434
rect 43372 44370 43428 44382
rect 42924 43810 42980 43820
rect 43036 44212 43092 44222
rect 43036 43650 43092 44156
rect 43484 44210 43540 45278
rect 43484 44158 43486 44210
rect 43538 44158 43540 44210
rect 43484 44146 43540 44158
rect 43036 43598 43038 43650
rect 43090 43598 43092 43650
rect 43036 43586 43092 43598
rect 42476 43540 42532 43550
rect 42476 43446 42532 43484
rect 42812 43540 42868 43550
rect 42812 43446 42868 43484
rect 43484 43540 43540 43550
rect 42924 43426 42980 43438
rect 42924 43374 42926 43426
rect 42978 43374 42980 43426
rect 42924 42980 42980 43374
rect 42924 42924 43204 42980
rect 42476 42868 42532 42878
rect 42532 42812 42756 42868
rect 42476 42774 42532 42812
rect 42364 42644 42420 42654
rect 42364 42550 42420 42588
rect 42028 41918 42030 41970
rect 42082 41918 42084 41970
rect 42028 41906 42084 41918
rect 42140 41972 42196 41982
rect 42364 41972 42420 41982
rect 42140 41970 42420 41972
rect 42140 41918 42142 41970
rect 42194 41918 42366 41970
rect 42418 41918 42420 41970
rect 42140 41916 42420 41918
rect 42140 41906 42196 41916
rect 42364 41906 42420 41916
rect 42700 41748 42756 42812
rect 42812 42756 42868 42766
rect 42812 42662 42868 42700
rect 43148 42754 43204 42924
rect 43148 42702 43150 42754
rect 43202 42702 43204 42754
rect 43148 42690 43204 42702
rect 42924 42644 42980 42654
rect 42924 42550 42980 42588
rect 43484 42308 43540 43484
rect 43596 42980 43652 49532
rect 43820 49364 43876 49374
rect 43708 49308 43820 49364
rect 43708 48244 43764 49308
rect 43820 49298 43876 49308
rect 43820 49026 43876 49038
rect 43820 48974 43822 49026
rect 43874 48974 43876 49026
rect 43820 48916 43876 48974
rect 43932 49028 43988 49038
rect 44156 49028 44212 49646
rect 43932 48934 43988 48972
rect 44044 48972 44212 49028
rect 43820 48850 43876 48860
rect 43820 48244 43876 48254
rect 43708 48242 43876 48244
rect 43708 48190 43822 48242
rect 43874 48190 43876 48242
rect 43708 48188 43876 48190
rect 43820 47570 43876 48188
rect 43820 47518 43822 47570
rect 43874 47518 43876 47570
rect 43708 47348 43764 47358
rect 43708 46562 43764 47292
rect 43708 46510 43710 46562
rect 43762 46510 43764 46562
rect 43708 46498 43764 46510
rect 43820 46452 43876 47518
rect 43820 46004 43876 46396
rect 43932 46004 43988 46014
rect 43820 46002 43988 46004
rect 43820 45950 43934 46002
rect 43986 45950 43988 46002
rect 43820 45948 43988 45950
rect 43932 45938 43988 45948
rect 43708 45668 43764 45678
rect 43708 44660 43764 45612
rect 43932 45556 43988 45566
rect 43708 44594 43764 44604
rect 43820 45332 43876 45342
rect 43820 44210 43876 45276
rect 43932 44996 43988 45500
rect 44044 45220 44100 48972
rect 44156 48802 44212 48814
rect 44156 48750 44158 48802
rect 44210 48750 44212 48802
rect 44156 48242 44212 48750
rect 44156 48190 44158 48242
rect 44210 48190 44212 48242
rect 44156 48178 44212 48190
rect 44268 48020 44324 51660
rect 44380 50428 44436 51884
rect 45276 51716 45332 52332
rect 45276 51650 45332 51660
rect 45276 51380 45332 51390
rect 45332 51324 45444 51380
rect 45276 51286 45332 51324
rect 45388 50482 45444 51324
rect 45388 50430 45390 50482
rect 45442 50430 45444 50482
rect 44380 50372 44884 50428
rect 45388 50418 45444 50430
rect 44604 49924 44660 49934
rect 44828 49924 44884 50372
rect 45500 50148 45556 54348
rect 46284 54404 46340 54414
rect 46284 54310 46340 54348
rect 47068 53732 47124 54462
rect 50988 53842 51044 53854
rect 50988 53790 50990 53842
rect 51042 53790 51044 53842
rect 47740 53732 47796 53742
rect 48188 53732 48244 53742
rect 47068 53730 48244 53732
rect 47068 53678 47742 53730
rect 47794 53678 48190 53730
rect 48242 53678 48244 53730
rect 47068 53676 48244 53678
rect 47740 53666 47796 53676
rect 46956 53618 47012 53630
rect 46956 53566 46958 53618
rect 47010 53566 47012 53618
rect 46620 53284 46676 53294
rect 46620 52162 46676 53228
rect 46620 52110 46622 52162
rect 46674 52110 46676 52162
rect 46620 52098 46676 52110
rect 46732 52274 46788 52286
rect 46732 52222 46734 52274
rect 46786 52222 46788 52274
rect 45836 52050 45892 52062
rect 45836 51998 45838 52050
rect 45890 51998 45892 52050
rect 45724 51380 45780 51390
rect 45724 51286 45780 51324
rect 45388 50092 45556 50148
rect 44492 49922 44884 49924
rect 44492 49870 44606 49922
rect 44658 49870 44884 49922
rect 44492 49868 44884 49870
rect 44940 49924 44996 49934
rect 44380 49026 44436 49038
rect 44380 48974 44382 49026
rect 44434 48974 44436 49026
rect 44380 48804 44436 48974
rect 44380 48738 44436 48748
rect 44380 48468 44436 48506
rect 44380 48402 44436 48412
rect 44380 48244 44436 48254
rect 44492 48244 44548 49868
rect 44604 49858 44660 49868
rect 44940 49364 44996 49868
rect 44716 49308 44996 49364
rect 44380 48242 44548 48244
rect 44380 48190 44382 48242
rect 44434 48190 44548 48242
rect 44380 48188 44548 48190
rect 44380 48178 44436 48188
rect 44156 47964 44324 48020
rect 44380 48020 44436 48030
rect 44156 47572 44212 47964
rect 44156 47478 44212 47516
rect 44268 47460 44324 47470
rect 44268 47366 44324 47404
rect 44380 46900 44436 47964
rect 44380 46806 44436 46844
rect 44492 46676 44548 48188
rect 44604 48242 44660 48254
rect 44604 48190 44606 48242
rect 44658 48190 44660 48242
rect 44604 47012 44660 48190
rect 44716 47124 44772 49308
rect 44828 49140 44884 49150
rect 44828 48244 44884 49084
rect 44940 49026 44996 49308
rect 44940 48974 44942 49026
rect 44994 48974 44996 49026
rect 44940 48962 44996 48974
rect 45276 49922 45332 49934
rect 45276 49870 45278 49922
rect 45330 49870 45332 49922
rect 45276 49028 45332 49870
rect 45276 48962 45332 48972
rect 45164 48916 45220 48926
rect 45052 48914 45220 48916
rect 45052 48862 45166 48914
rect 45218 48862 45220 48914
rect 45052 48860 45220 48862
rect 45052 48580 45108 48860
rect 45164 48850 45220 48860
rect 44828 48178 44884 48188
rect 44940 48524 45108 48580
rect 45276 48804 45332 48814
rect 44940 47460 44996 48524
rect 45164 48468 45220 48478
rect 45276 48468 45332 48748
rect 45164 48466 45332 48468
rect 45164 48414 45166 48466
rect 45218 48414 45332 48466
rect 45164 48412 45332 48414
rect 45388 48468 45444 50092
rect 45612 49924 45668 49934
rect 45836 49924 45892 51998
rect 46396 52050 46452 52062
rect 46396 51998 46398 52050
rect 46450 51998 46452 52050
rect 46396 50484 46452 51998
rect 46508 51380 46564 51390
rect 46508 50594 46564 51324
rect 46732 50706 46788 52222
rect 46844 52164 46900 52174
rect 46844 51602 46900 52108
rect 46844 51550 46846 51602
rect 46898 51550 46900 51602
rect 46844 51538 46900 51550
rect 46732 50654 46734 50706
rect 46786 50654 46788 50706
rect 46732 50642 46788 50654
rect 46508 50542 46510 50594
rect 46562 50542 46564 50594
rect 46508 50530 46564 50542
rect 46844 50596 46900 50634
rect 46844 50530 46900 50540
rect 46956 50428 47012 53566
rect 47516 53508 47572 53518
rect 47068 53172 47124 53182
rect 47068 53078 47124 53116
rect 47516 53170 47572 53452
rect 47516 53118 47518 53170
rect 47570 53118 47572 53170
rect 47516 53106 47572 53118
rect 48076 53172 48132 53182
rect 48076 53078 48132 53116
rect 47964 53058 48020 53070
rect 47964 53006 47966 53058
rect 48018 53006 48020 53058
rect 47740 52162 47796 52174
rect 47740 52110 47742 52162
rect 47794 52110 47796 52162
rect 47180 51828 47236 51838
rect 47180 51492 47236 51772
rect 47404 51716 47460 51726
rect 47292 51492 47348 51502
rect 47180 51490 47348 51492
rect 47180 51438 47294 51490
rect 47346 51438 47348 51490
rect 47180 51436 47348 51438
rect 47180 50596 47236 51436
rect 47292 51426 47348 51436
rect 47180 50530 47236 50540
rect 46284 50036 46340 50046
rect 45612 49922 45892 49924
rect 45612 49870 45614 49922
rect 45666 49870 45892 49922
rect 45612 49868 45892 49870
rect 45612 49858 45668 49868
rect 45836 49700 45892 49868
rect 46172 50034 46340 50036
rect 46172 49982 46286 50034
rect 46338 49982 46340 50034
rect 46172 49980 46340 49982
rect 45836 49634 45892 49644
rect 45948 49810 46004 49822
rect 45948 49758 45950 49810
rect 46002 49758 46004 49810
rect 45500 49476 45556 49486
rect 45500 49250 45556 49420
rect 45724 49364 45780 49374
rect 45500 49198 45502 49250
rect 45554 49198 45556 49250
rect 45500 49186 45556 49198
rect 45612 49308 45724 49364
rect 45612 49026 45668 49308
rect 45724 49298 45780 49308
rect 45836 49140 45892 49150
rect 45612 48974 45614 49026
rect 45666 48974 45668 49026
rect 45612 48962 45668 48974
rect 45724 49084 45836 49140
rect 45724 48802 45780 49084
rect 45836 49074 45892 49084
rect 45724 48750 45726 48802
rect 45778 48750 45780 48802
rect 45724 48738 45780 48750
rect 45164 48402 45220 48412
rect 45388 48402 45444 48412
rect 45724 48468 45780 48478
rect 45948 48468 46004 49758
rect 46172 49476 46228 49980
rect 46284 49970 46340 49980
rect 46284 49812 46340 49822
rect 46284 49718 46340 49756
rect 46172 49410 46228 49420
rect 46284 49028 46340 49038
rect 46284 48934 46340 48972
rect 46172 48916 46228 48926
rect 46172 48822 46228 48860
rect 46060 48804 46116 48814
rect 46060 48710 46116 48748
rect 46396 48692 46452 50428
rect 46620 50372 46676 50382
rect 46620 49810 46676 50316
rect 46620 49758 46622 49810
rect 46674 49758 46676 49810
rect 46620 49746 46676 49758
rect 46732 50372 47012 50428
rect 47404 50482 47460 51660
rect 47740 51380 47796 52110
rect 47964 51604 48020 53006
rect 48188 53060 48244 53676
rect 48860 53618 48916 53630
rect 48860 53566 48862 53618
rect 48914 53566 48916 53618
rect 48860 53172 48916 53566
rect 48860 53106 48916 53116
rect 49420 53508 49476 53518
rect 48748 53060 48804 53070
rect 48188 53004 48468 53060
rect 48188 52836 48244 52846
rect 48188 52742 48244 52780
rect 48300 52500 48356 52510
rect 48076 52164 48132 52174
rect 48076 52070 48132 52108
rect 47964 51538 48020 51548
rect 47740 51314 47796 51324
rect 47404 50430 47406 50482
rect 47458 50430 47460 50482
rect 47404 50418 47460 50430
rect 47964 51266 48020 51278
rect 47964 51214 47966 51266
rect 48018 51214 48020 51266
rect 47964 50428 48020 51214
rect 47180 50372 47236 50382
rect 47964 50372 48132 50428
rect 46732 49140 46788 50372
rect 46844 49810 46900 49822
rect 46844 49758 46846 49810
rect 46898 49758 46900 49810
rect 46844 49252 46900 49758
rect 46956 49812 47012 49822
rect 46956 49718 47012 49756
rect 47068 49810 47124 49822
rect 47068 49758 47070 49810
rect 47122 49758 47124 49810
rect 47068 49252 47124 49758
rect 46844 49186 46900 49196
rect 46956 49196 47124 49252
rect 46732 49074 46788 49084
rect 46620 49026 46676 49038
rect 46620 48974 46622 49026
rect 46674 48974 46676 49026
rect 46620 48916 46676 48974
rect 46956 48916 47012 49196
rect 47180 49138 47236 50316
rect 47964 49922 48020 49934
rect 47964 49870 47966 49922
rect 48018 49870 48020 49922
rect 47516 49810 47572 49822
rect 47516 49758 47518 49810
rect 47570 49758 47572 49810
rect 47292 49588 47348 49598
rect 47292 49250 47348 49532
rect 47292 49198 47294 49250
rect 47346 49198 47348 49250
rect 47292 49186 47348 49198
rect 47180 49086 47182 49138
rect 47234 49086 47236 49138
rect 47180 49074 47236 49086
rect 47516 49028 47572 49758
rect 47964 49812 48020 49870
rect 48076 49924 48132 50372
rect 48076 49858 48132 49868
rect 47964 49746 48020 49756
rect 48076 49698 48132 49710
rect 48076 49646 48078 49698
rect 48130 49646 48132 49698
rect 47964 49028 48020 49038
rect 47516 49026 48020 49028
rect 47516 48974 47966 49026
rect 48018 48974 48020 49026
rect 47516 48972 48020 48974
rect 46620 48860 46900 48916
rect 46172 48636 46676 48692
rect 46060 48468 46116 48478
rect 45948 48466 46116 48468
rect 45948 48414 46062 48466
rect 46114 48414 46116 48466
rect 45948 48412 46116 48414
rect 45724 48374 45780 48412
rect 46060 48402 46116 48412
rect 46172 48466 46228 48636
rect 46172 48414 46174 48466
rect 46226 48414 46228 48466
rect 46172 48402 46228 48414
rect 45052 48356 45108 48366
rect 45052 48262 45108 48300
rect 45164 48244 45220 48254
rect 45948 48244 46004 48254
rect 45220 48188 45332 48244
rect 45164 48178 45220 48188
rect 45276 48130 45332 48188
rect 45276 48078 45278 48130
rect 45330 48078 45332 48130
rect 45276 48066 45332 48078
rect 45612 48242 46004 48244
rect 45612 48190 45950 48242
rect 46002 48190 46004 48242
rect 45612 48188 46004 48190
rect 45500 47796 45556 47806
rect 45500 47572 45556 47740
rect 45388 47570 45556 47572
rect 45388 47518 45502 47570
rect 45554 47518 45556 47570
rect 45388 47516 45556 47518
rect 44996 47404 45108 47460
rect 44940 47394 44996 47404
rect 44828 47348 44884 47358
rect 44828 47236 44884 47292
rect 44940 47236 44996 47246
rect 44828 47234 44996 47236
rect 44828 47182 44942 47234
rect 44994 47182 44996 47234
rect 44828 47180 44996 47182
rect 44940 47170 44996 47180
rect 44716 47068 44884 47124
rect 44660 46956 44772 47012
rect 44604 46946 44660 46956
rect 44604 46676 44660 46686
rect 44492 46674 44660 46676
rect 44492 46622 44606 46674
rect 44658 46622 44660 46674
rect 44492 46620 44660 46622
rect 44604 46610 44660 46620
rect 44604 46228 44660 46238
rect 44492 46172 44604 46228
rect 44268 46004 44324 46014
rect 44268 45668 44324 45948
rect 44268 45574 44324 45612
rect 44492 45444 44548 46172
rect 44604 46162 44660 46172
rect 44716 45556 44772 46956
rect 44268 45388 44548 45444
rect 44604 45500 44772 45556
rect 44268 45330 44324 45388
rect 44268 45278 44270 45330
rect 44322 45278 44324 45330
rect 44268 45266 44324 45278
rect 44044 45154 44100 45164
rect 44156 45106 44212 45118
rect 44156 45054 44158 45106
rect 44210 45054 44212 45106
rect 44156 44996 44212 45054
rect 44492 45106 44548 45118
rect 44492 45054 44494 45106
rect 44546 45054 44548 45106
rect 44380 44996 44436 45006
rect 43932 44940 44100 44996
rect 44156 44940 44380 44996
rect 43820 44158 43822 44210
rect 43874 44158 43876 44210
rect 43820 44146 43876 44158
rect 43932 44322 43988 44334
rect 43932 44270 43934 44322
rect 43986 44270 43988 44322
rect 43596 42914 43652 42924
rect 43820 42980 43876 42990
rect 43932 42980 43988 44270
rect 43820 42978 43988 42980
rect 43820 42926 43822 42978
rect 43874 42926 43988 42978
rect 43820 42924 43988 42926
rect 43820 42914 43876 42924
rect 43596 42756 43652 42766
rect 43932 42756 43988 42766
rect 43596 42754 43988 42756
rect 43596 42702 43598 42754
rect 43650 42702 43934 42754
rect 43986 42702 43988 42754
rect 43596 42700 43988 42702
rect 43596 42690 43652 42700
rect 43932 42690 43988 42700
rect 43484 42252 43764 42308
rect 43708 42194 43764 42252
rect 43708 42142 43710 42194
rect 43762 42142 43764 42194
rect 43148 42028 43428 42084
rect 43036 41972 43092 41982
rect 43148 41972 43204 42028
rect 43036 41970 43204 41972
rect 43036 41918 43038 41970
rect 43090 41918 43204 41970
rect 43036 41916 43204 41918
rect 43036 41906 43092 41916
rect 43260 41860 43316 41870
rect 43148 41858 43316 41860
rect 43148 41806 43262 41858
rect 43314 41806 43316 41858
rect 43148 41804 43316 41806
rect 42812 41748 42868 41758
rect 42700 41746 42868 41748
rect 42700 41694 42814 41746
rect 42866 41694 42868 41746
rect 42700 41692 42868 41694
rect 42812 41682 42868 41692
rect 43036 41748 43092 41758
rect 41804 41234 41860 41244
rect 41916 41412 41972 41422
rect 41916 41298 41972 41356
rect 41916 41246 41918 41298
rect 41970 41246 41972 41298
rect 41916 41234 41972 41246
rect 41804 41076 41860 41086
rect 41804 40626 41860 41020
rect 43036 41074 43092 41692
rect 43036 41022 43038 41074
rect 43090 41022 43092 41074
rect 43036 41010 43092 41022
rect 42700 40964 42756 40974
rect 42588 40962 42756 40964
rect 42588 40910 42702 40962
rect 42754 40910 42756 40962
rect 42588 40908 42756 40910
rect 41804 40574 41806 40626
rect 41858 40574 41860 40626
rect 41804 40562 41860 40574
rect 42028 40628 42084 40638
rect 42028 40534 42084 40572
rect 42252 40402 42308 40414
rect 42252 40350 42254 40402
rect 42306 40350 42308 40402
rect 42140 40290 42196 40302
rect 42140 40238 42142 40290
rect 42194 40238 42196 40290
rect 42140 39508 42196 40238
rect 42140 39442 42196 39452
rect 41524 38892 41636 38948
rect 41916 39172 41972 39182
rect 41468 38882 41524 38892
rect 41692 38834 41748 38846
rect 41692 38782 41694 38834
rect 41746 38782 41748 38834
rect 41468 38722 41524 38734
rect 41468 38670 41470 38722
rect 41522 38670 41524 38722
rect 41468 38164 41524 38670
rect 41468 38098 41524 38108
rect 41692 37268 41748 38782
rect 41916 38834 41972 39116
rect 41916 38782 41918 38834
rect 41970 38782 41972 38834
rect 41916 38770 41972 38782
rect 42252 39060 42308 40350
rect 42588 39844 42644 40908
rect 42700 40898 42756 40908
rect 43036 40740 43092 40750
rect 42588 39778 42644 39788
rect 42700 40628 42756 40638
rect 42252 38836 42308 39004
rect 42476 38948 42532 38958
rect 42364 38836 42420 38846
rect 42252 38834 42420 38836
rect 42252 38782 42366 38834
rect 42418 38782 42420 38834
rect 42252 38780 42420 38782
rect 42364 38770 42420 38780
rect 41804 38724 41860 38734
rect 41804 38610 41860 38668
rect 41804 38558 41806 38610
rect 41858 38558 41860 38610
rect 41804 38546 41860 38558
rect 41916 38612 41972 38622
rect 41692 37202 41748 37212
rect 41244 36978 41300 36988
rect 41132 36764 41300 36820
rect 40908 36372 40964 36382
rect 40908 35922 40964 36316
rect 40908 35870 40910 35922
rect 40962 35870 40964 35922
rect 40908 35364 40964 35870
rect 41132 35810 41188 35822
rect 41132 35758 41134 35810
rect 41186 35758 41188 35810
rect 41132 35588 41188 35758
rect 41244 35810 41300 36764
rect 41244 35758 41246 35810
rect 41298 35758 41300 35810
rect 41244 35746 41300 35758
rect 41580 35812 41636 35822
rect 41580 35718 41636 35756
rect 41132 35522 41188 35532
rect 40908 35298 40964 35308
rect 40460 35140 40516 35150
rect 40460 34914 40516 35084
rect 41356 35026 41412 35038
rect 41356 34974 41358 35026
rect 41410 34974 41412 35026
rect 40460 34862 40462 34914
rect 40514 34862 40516 34914
rect 40460 34850 40516 34862
rect 40684 34916 40740 34926
rect 40684 34802 40740 34860
rect 40684 34750 40686 34802
rect 40738 34750 40740 34802
rect 40684 34738 40740 34750
rect 40796 34804 40852 34814
rect 40796 34710 40852 34748
rect 40348 34190 40350 34242
rect 40402 34190 40404 34242
rect 40348 34178 40404 34190
rect 41132 34132 41188 34142
rect 41356 34132 41412 34974
rect 41804 34916 41860 34926
rect 41132 34130 41412 34132
rect 41132 34078 41134 34130
rect 41186 34078 41412 34130
rect 41132 34076 41412 34078
rect 41692 34860 41804 34916
rect 41692 34130 41748 34860
rect 41804 34822 41860 34860
rect 41692 34078 41694 34130
rect 41746 34078 41748 34130
rect 41132 34020 41188 34076
rect 41692 34066 41748 34078
rect 41132 33954 41188 33964
rect 41916 34020 41972 38556
rect 42476 38500 42532 38892
rect 42700 38834 42756 40572
rect 43036 40626 43092 40684
rect 43036 40574 43038 40626
rect 43090 40574 43092 40626
rect 43036 40562 43092 40574
rect 42924 40404 42980 40414
rect 42924 40310 42980 40348
rect 42924 39732 42980 39742
rect 42924 39618 42980 39676
rect 42924 39566 42926 39618
rect 42978 39566 42980 39618
rect 42924 39554 42980 39566
rect 42700 38782 42702 38834
rect 42754 38782 42756 38834
rect 42700 38770 42756 38782
rect 42812 39508 42868 39518
rect 42812 38836 42868 39452
rect 42924 38836 42980 38846
rect 42812 38834 42980 38836
rect 42812 38782 42926 38834
rect 42978 38782 42980 38834
rect 42812 38780 42980 38782
rect 42924 38770 42980 38780
rect 42588 38724 42644 38762
rect 42588 38658 42644 38668
rect 42476 38444 42644 38500
rect 42476 38052 42532 38062
rect 42252 37604 42308 37614
rect 42028 37042 42084 37054
rect 42028 36990 42030 37042
rect 42082 36990 42084 37042
rect 42028 35924 42084 36990
rect 42140 37042 42196 37054
rect 42140 36990 42142 37042
rect 42194 36990 42196 37042
rect 42140 36820 42196 36990
rect 42140 36754 42196 36764
rect 42028 35868 42196 35924
rect 42028 35698 42084 35710
rect 42028 35646 42030 35698
rect 42082 35646 42084 35698
rect 42028 35588 42084 35646
rect 42028 35522 42084 35532
rect 41916 33954 41972 33964
rect 42028 34132 42084 34142
rect 40236 33908 40292 33918
rect 40236 31948 40292 33852
rect 42028 33460 42084 34076
rect 42140 33572 42196 35868
rect 42252 34914 42308 37548
rect 42364 37268 42420 37278
rect 42364 37174 42420 37212
rect 42476 35698 42532 37996
rect 42588 37266 42644 38444
rect 42700 38164 42756 38174
rect 42700 38070 42756 38108
rect 42700 37940 42756 37950
rect 42700 37378 42756 37884
rect 42700 37326 42702 37378
rect 42754 37326 42756 37378
rect 42700 37314 42756 37326
rect 42588 37214 42590 37266
rect 42642 37214 42644 37266
rect 42588 37202 42644 37214
rect 43036 37044 43092 37054
rect 42476 35646 42478 35698
rect 42530 35646 42532 35698
rect 42476 35634 42532 35646
rect 42812 35812 42868 35822
rect 42252 34862 42254 34914
rect 42306 34862 42308 34914
rect 42252 34850 42308 34862
rect 42700 34916 42756 34926
rect 42700 34822 42756 34860
rect 42812 34914 42868 35756
rect 43036 35700 43092 36988
rect 43148 36820 43204 41804
rect 43260 41794 43316 41804
rect 43372 41636 43428 42028
rect 43596 41972 43652 41982
rect 43596 41636 43652 41916
rect 43372 41580 43652 41636
rect 43372 40964 43428 40974
rect 43372 40740 43428 40908
rect 43372 40674 43428 40684
rect 43148 36754 43204 36764
rect 43260 40402 43316 40414
rect 43260 40350 43262 40402
rect 43314 40350 43316 40402
rect 43148 36372 43204 36382
rect 43148 36278 43204 36316
rect 42812 34862 42814 34914
rect 42866 34862 42868 34914
rect 42812 34850 42868 34862
rect 42924 35698 43092 35700
rect 42924 35646 43038 35698
rect 43090 35646 43092 35698
rect 42924 35644 43092 35646
rect 42588 34690 42644 34702
rect 42924 34692 42980 35644
rect 43036 35634 43092 35644
rect 43260 35698 43316 40350
rect 43372 40402 43428 40414
rect 43372 40350 43374 40402
rect 43426 40350 43428 40402
rect 43372 37604 43428 40350
rect 43484 40404 43540 41580
rect 43596 40628 43652 40638
rect 43596 40534 43652 40572
rect 43484 40348 43652 40404
rect 43484 40180 43540 40190
rect 43484 39844 43540 40124
rect 43484 39730 43540 39788
rect 43484 39678 43486 39730
rect 43538 39678 43540 39730
rect 43484 39666 43540 39678
rect 43596 39508 43652 40348
rect 43484 39452 43652 39508
rect 43484 38836 43540 39452
rect 43596 38948 43652 38958
rect 43708 38948 43764 42142
rect 43820 41076 43876 41086
rect 43820 40964 43876 41020
rect 43820 40962 43988 40964
rect 43820 40910 43822 40962
rect 43874 40910 43988 40962
rect 43820 40908 43988 40910
rect 43820 40898 43876 40908
rect 43820 40404 43876 40414
rect 43820 40310 43876 40348
rect 43932 39732 43988 40908
rect 44044 40514 44100 44940
rect 44380 44930 44436 44940
rect 44492 44212 44548 45054
rect 44492 44146 44548 44156
rect 44380 44098 44436 44110
rect 44380 44046 44382 44098
rect 44434 44046 44436 44098
rect 44380 43540 44436 44046
rect 44380 43474 44436 43484
rect 44268 42756 44324 42766
rect 44268 42662 44324 42700
rect 44156 42530 44212 42542
rect 44156 42478 44158 42530
rect 44210 42478 44212 42530
rect 44156 41972 44212 42478
rect 44156 41906 44212 41916
rect 44044 40462 44046 40514
rect 44098 40462 44100 40514
rect 44044 40450 44100 40462
rect 44380 40404 44436 40414
rect 44380 40310 44436 40348
rect 43932 39666 43988 39676
rect 44492 40290 44548 40302
rect 44492 40238 44494 40290
rect 44546 40238 44548 40290
rect 44044 39396 44100 39406
rect 44044 39394 44212 39396
rect 44044 39342 44046 39394
rect 44098 39342 44212 39394
rect 44044 39340 44212 39342
rect 44044 39330 44100 39340
rect 44156 39172 44212 39340
rect 43820 38948 43876 38958
rect 43708 38946 43876 38948
rect 43708 38894 43822 38946
rect 43874 38894 43876 38946
rect 43708 38892 43876 38894
rect 43596 38854 43652 38892
rect 43484 38770 43540 38780
rect 43372 37538 43428 37548
rect 43484 38050 43540 38062
rect 43484 37998 43486 38050
rect 43538 37998 43540 38050
rect 43484 37156 43540 37998
rect 43820 38052 43876 38892
rect 44156 38834 44212 39116
rect 44380 39060 44436 39070
rect 44380 38966 44436 39004
rect 44156 38782 44158 38834
rect 44210 38782 44212 38834
rect 44156 38770 44212 38782
rect 44156 38612 44212 38622
rect 44492 38612 44548 40238
rect 44604 39284 44660 45500
rect 44716 45108 44772 45118
rect 44716 45014 44772 45052
rect 44828 41524 44884 47068
rect 45052 46898 45108 47404
rect 45052 46846 45054 46898
rect 45106 46846 45108 46898
rect 44940 45108 44996 45118
rect 45052 45108 45108 46846
rect 45276 46900 45332 46910
rect 45388 46900 45444 47516
rect 45500 47506 45556 47516
rect 45612 47124 45668 48188
rect 45948 48178 46004 48188
rect 46620 48242 46676 48636
rect 46620 48190 46622 48242
rect 46674 48190 46676 48242
rect 46620 48178 46676 48190
rect 46844 48468 46900 48860
rect 46956 48850 47012 48860
rect 47068 48802 47124 48814
rect 47068 48750 47070 48802
rect 47122 48750 47124 48802
rect 47068 48692 47124 48750
rect 46172 47572 46228 47582
rect 45836 47458 45892 47470
rect 45836 47406 45838 47458
rect 45890 47406 45892 47458
rect 45276 46898 45444 46900
rect 45276 46846 45278 46898
rect 45330 46846 45444 46898
rect 45276 46844 45444 46846
rect 45500 47068 45668 47124
rect 45724 47236 45780 47246
rect 45276 46834 45332 46844
rect 45164 46562 45220 46574
rect 45164 46510 45166 46562
rect 45218 46510 45220 46562
rect 45164 46228 45220 46510
rect 45164 46162 45220 46172
rect 45388 45892 45444 45902
rect 45164 45666 45220 45678
rect 45164 45614 45166 45666
rect 45218 45614 45220 45666
rect 45164 45332 45220 45614
rect 45164 45266 45220 45276
rect 45388 45220 45444 45836
rect 45164 45108 45220 45118
rect 45052 45106 45220 45108
rect 45052 45054 45166 45106
rect 45218 45054 45220 45106
rect 45052 45052 45220 45054
rect 44940 45014 44996 45052
rect 45164 45042 45220 45052
rect 45388 45106 45444 45164
rect 45388 45054 45390 45106
rect 45442 45054 45444 45106
rect 45388 45042 45444 45054
rect 45500 45108 45556 47068
rect 45612 46900 45668 46910
rect 45612 46674 45668 46844
rect 45612 46622 45614 46674
rect 45666 46622 45668 46674
rect 45612 46610 45668 46622
rect 45612 46452 45668 46462
rect 45612 45890 45668 46396
rect 45612 45838 45614 45890
rect 45666 45838 45668 45890
rect 45612 45826 45668 45838
rect 45724 45890 45780 47180
rect 45836 46004 45892 47406
rect 46172 47458 46228 47516
rect 46172 47406 46174 47458
rect 46226 47406 46228 47458
rect 46172 47394 46228 47406
rect 46284 47460 46340 47470
rect 46284 47458 46564 47460
rect 46284 47406 46286 47458
rect 46338 47406 46564 47458
rect 46284 47404 46564 47406
rect 46284 47394 46340 47404
rect 46396 47234 46452 47246
rect 46396 47182 46398 47234
rect 46450 47182 46452 47234
rect 45836 45938 45892 45948
rect 46284 46900 46340 46910
rect 46284 45892 46340 46844
rect 46396 46340 46452 47182
rect 46508 46900 46564 47404
rect 46508 46834 46564 46844
rect 46452 46284 46564 46340
rect 46396 46274 46452 46284
rect 45724 45838 45726 45890
rect 45778 45838 45780 45890
rect 45724 45826 45780 45838
rect 45948 45890 46340 45892
rect 45948 45838 46286 45890
rect 46338 45838 46340 45890
rect 45948 45836 46340 45838
rect 45836 45778 45892 45790
rect 45836 45726 45838 45778
rect 45890 45726 45892 45778
rect 45500 45052 45668 45108
rect 45276 44996 45332 45034
rect 45276 44930 45332 44940
rect 45500 44884 45556 44894
rect 45276 44772 45332 44782
rect 45276 43764 45332 44716
rect 45164 43204 45220 43214
rect 44940 42868 44996 42878
rect 44940 42754 44996 42812
rect 44940 42702 44942 42754
rect 44994 42702 44996 42754
rect 44940 42690 44996 42702
rect 45164 42756 45220 43148
rect 45164 42642 45220 42700
rect 45164 42590 45166 42642
rect 45218 42590 45220 42642
rect 45164 42578 45220 42590
rect 45276 41972 45332 43708
rect 45500 43762 45556 44828
rect 45500 43710 45502 43762
rect 45554 43710 45556 43762
rect 45500 43698 45556 43710
rect 45500 41972 45556 41982
rect 45276 41970 45556 41972
rect 45276 41918 45278 41970
rect 45330 41918 45502 41970
rect 45554 41918 45556 41970
rect 45276 41916 45556 41918
rect 45276 41906 45332 41916
rect 45500 41906 45556 41916
rect 45612 41748 45668 45052
rect 45724 44212 45780 44222
rect 45836 44212 45892 45726
rect 45948 45330 46004 45836
rect 46284 45826 46340 45836
rect 46396 46116 46452 46126
rect 46396 45668 46452 46060
rect 46284 45612 46452 45668
rect 45948 45278 45950 45330
rect 46002 45278 46004 45330
rect 45948 45266 46004 45278
rect 46060 45332 46116 45342
rect 46060 44322 46116 45276
rect 46060 44270 46062 44322
rect 46114 44270 46116 44322
rect 46060 44258 46116 44270
rect 45948 44212 46004 44222
rect 45836 44156 45948 44212
rect 45724 44118 45780 44156
rect 45948 44146 46004 44156
rect 46172 44098 46228 44110
rect 46172 44046 46174 44098
rect 46226 44046 46228 44098
rect 46172 43652 46228 44046
rect 45836 43540 45892 43550
rect 45836 43426 45892 43484
rect 46172 43538 46228 43596
rect 46172 43486 46174 43538
rect 46226 43486 46228 43538
rect 46172 43474 46228 43486
rect 45836 43374 45838 43426
rect 45890 43374 45892 43426
rect 45836 43362 45892 43374
rect 46284 43204 46340 45612
rect 44828 41458 44884 41468
rect 45164 41692 45668 41748
rect 45724 43148 46340 43204
rect 46396 44996 46452 45006
rect 46508 44996 46564 46284
rect 46396 44994 46564 44996
rect 46396 44942 46398 44994
rect 46450 44942 46564 44994
rect 46396 44940 46564 44942
rect 44940 41186 44996 41198
rect 44940 41134 44942 41186
rect 44994 41134 44996 41186
rect 44940 40964 44996 41134
rect 45164 41076 45220 41692
rect 44940 40898 44996 40908
rect 45052 41074 45220 41076
rect 45052 41022 45166 41074
rect 45218 41022 45220 41074
rect 45052 41020 45220 41022
rect 45052 40740 45108 41020
rect 45164 41010 45220 41020
rect 45276 41524 45332 41534
rect 44716 40684 45108 40740
rect 44716 40516 44772 40684
rect 44716 40402 44772 40460
rect 44716 40350 44718 40402
rect 44770 40350 44772 40402
rect 44716 40338 44772 40350
rect 44940 40402 44996 40414
rect 44940 40350 44942 40402
rect 44994 40350 44996 40402
rect 44828 40180 44884 40190
rect 44716 40178 44884 40180
rect 44716 40126 44830 40178
rect 44882 40126 44884 40178
rect 44716 40124 44884 40126
rect 44716 39284 44772 40124
rect 44828 40114 44884 40124
rect 44940 39730 44996 40350
rect 44940 39678 44942 39730
rect 44994 39678 44996 39730
rect 44940 39666 44996 39678
rect 44828 39508 44884 39518
rect 45052 39508 45108 40684
rect 45164 39620 45220 39630
rect 45164 39526 45220 39564
rect 44828 39506 45108 39508
rect 44828 39454 44830 39506
rect 44882 39454 45108 39506
rect 44828 39452 45108 39454
rect 44828 39442 44884 39452
rect 44716 39228 45108 39284
rect 44604 39060 44660 39228
rect 44604 39004 44884 39060
rect 44604 38948 44660 39004
rect 44604 38882 44660 38892
rect 44716 38836 44772 38846
rect 44716 38722 44772 38780
rect 44716 38670 44718 38722
rect 44770 38670 44772 38722
rect 44716 38658 44772 38670
rect 44156 38610 44548 38612
rect 44156 38558 44158 38610
rect 44210 38558 44548 38610
rect 44156 38556 44548 38558
rect 44156 38546 44212 38556
rect 43932 38276 43988 38286
rect 43932 38162 43988 38220
rect 43932 38110 43934 38162
rect 43986 38110 43988 38162
rect 43932 38098 43988 38110
rect 43820 37986 43876 37996
rect 44828 37938 44884 39004
rect 44828 37886 44830 37938
rect 44882 37886 44884 37938
rect 44828 37874 44884 37886
rect 45052 38052 45108 39228
rect 45276 38388 45332 41468
rect 45500 40404 45556 40414
rect 45500 40310 45556 40348
rect 45388 39956 45444 39966
rect 45388 39618 45444 39900
rect 45388 39566 45390 39618
rect 45442 39566 45444 39618
rect 45388 39554 45444 39566
rect 45724 38668 45780 43148
rect 45836 42868 45892 42878
rect 45836 42774 45892 42812
rect 46284 42754 46340 42766
rect 46284 42702 46286 42754
rect 46338 42702 46340 42754
rect 45836 42082 45892 42094
rect 45836 42030 45838 42082
rect 45890 42030 45892 42082
rect 45836 41748 45892 42030
rect 46284 41972 46340 42702
rect 45892 41692 46116 41748
rect 45836 41682 45892 41692
rect 46060 40402 46116 41692
rect 46172 41300 46228 41310
rect 46284 41300 46340 41916
rect 46172 41298 46340 41300
rect 46172 41246 46174 41298
rect 46226 41246 46340 41298
rect 46172 41244 46340 41246
rect 46172 41234 46228 41244
rect 46060 40350 46062 40402
rect 46114 40350 46116 40402
rect 45836 40178 45892 40190
rect 45836 40126 45838 40178
rect 45890 40126 45892 40178
rect 45836 39956 45892 40126
rect 45836 39890 45892 39900
rect 46060 39620 46116 40350
rect 46060 39554 46116 39564
rect 46172 40292 46228 40302
rect 45276 38322 45332 38332
rect 45612 38612 45780 38668
rect 45500 38052 45556 38062
rect 45052 38050 45556 38052
rect 45052 37998 45054 38050
rect 45106 37998 45502 38050
rect 45554 37998 45556 38050
rect 45052 37996 45556 37998
rect 43820 37826 43876 37838
rect 43820 37774 43822 37826
rect 43874 37774 43876 37826
rect 43820 37268 43876 37774
rect 44604 37492 44660 37502
rect 44604 37398 44660 37436
rect 43820 37202 43876 37212
rect 43708 37156 43764 37166
rect 43484 37100 43708 37156
rect 43708 37062 43764 37100
rect 43372 36932 43428 36942
rect 43372 36484 43428 36876
rect 43372 36418 43428 36428
rect 43484 36820 43540 36830
rect 43260 35646 43262 35698
rect 43314 35646 43316 35698
rect 43260 35634 43316 35646
rect 43484 35812 43540 36764
rect 44156 36596 44212 36606
rect 44156 36502 44212 36540
rect 43820 36484 43876 36494
rect 43820 36482 43988 36484
rect 43820 36430 43822 36482
rect 43874 36430 43988 36482
rect 43820 36428 43988 36430
rect 43820 36418 43876 36428
rect 43036 35364 43092 35374
rect 43036 34802 43092 35308
rect 43036 34750 43038 34802
rect 43090 34750 43092 34802
rect 43036 34738 43092 34750
rect 43484 34804 43540 35756
rect 42588 34638 42590 34690
rect 42642 34638 42644 34690
rect 42588 33908 42644 34638
rect 42700 34636 42980 34692
rect 42700 34242 42756 34636
rect 43372 34356 43428 34366
rect 43484 34356 43540 34748
rect 43372 34354 43540 34356
rect 43372 34302 43374 34354
rect 43426 34302 43540 34354
rect 43372 34300 43540 34302
rect 43596 36258 43652 36270
rect 43596 36206 43598 36258
rect 43650 36206 43652 36258
rect 43372 34290 43428 34300
rect 42700 34190 42702 34242
rect 42754 34190 42756 34242
rect 42700 34178 42756 34190
rect 43036 34132 43092 34142
rect 43036 34038 43092 34076
rect 42588 33842 42644 33852
rect 43596 33908 43652 36206
rect 43932 35810 43988 36428
rect 44940 36482 44996 36494
rect 44940 36430 44942 36482
rect 44994 36430 44996 36482
rect 44380 36372 44436 36382
rect 44268 36036 44324 36046
rect 44268 35922 44324 35980
rect 44268 35870 44270 35922
rect 44322 35870 44324 35922
rect 44268 35858 44324 35870
rect 44380 35922 44436 36316
rect 44380 35870 44382 35922
rect 44434 35870 44436 35922
rect 44380 35858 44436 35870
rect 43932 35758 43934 35810
rect 43986 35758 43988 35810
rect 43932 35746 43988 35758
rect 44492 35812 44548 35822
rect 44716 35812 44772 35822
rect 44492 35718 44548 35756
rect 44604 35810 44772 35812
rect 44604 35758 44718 35810
rect 44770 35758 44772 35810
rect 44604 35756 44772 35758
rect 44604 35140 44660 35756
rect 44716 35746 44772 35756
rect 43932 35084 44660 35140
rect 43932 35026 43988 35084
rect 43932 34974 43934 35026
rect 43986 34974 43988 35026
rect 43932 34580 43988 34974
rect 44940 35028 44996 36430
rect 45052 36372 45108 37996
rect 45500 37490 45556 37996
rect 45500 37438 45502 37490
rect 45554 37438 45556 37490
rect 45500 37426 45556 37438
rect 45164 37268 45220 37278
rect 45164 37174 45220 37212
rect 45500 36932 45556 36942
rect 45164 36372 45220 36382
rect 45500 36372 45556 36876
rect 45052 36370 45220 36372
rect 45052 36318 45166 36370
rect 45218 36318 45220 36370
rect 45052 36316 45220 36318
rect 45164 36306 45220 36316
rect 45388 36370 45556 36372
rect 45388 36318 45502 36370
rect 45554 36318 45556 36370
rect 45388 36316 45556 36318
rect 45388 36036 45444 36316
rect 45500 36306 45556 36316
rect 45388 35922 45444 35980
rect 45388 35870 45390 35922
rect 45442 35870 45444 35922
rect 45388 35858 45444 35870
rect 45052 35028 45108 35038
rect 44940 34972 45052 35028
rect 45052 34914 45108 34972
rect 45052 34862 45054 34914
rect 45106 34862 45108 34914
rect 45052 34850 45108 34862
rect 45388 34692 45444 34702
rect 45388 34598 45444 34636
rect 43932 34514 43988 34524
rect 43596 33842 43652 33852
rect 44604 33908 44660 33918
rect 42140 33516 43652 33572
rect 42028 33404 42532 33460
rect 41468 33122 41524 33134
rect 41468 33070 41470 33122
rect 41522 33070 41524 33122
rect 41020 32676 41076 32686
rect 40908 32674 41076 32676
rect 40908 32622 41022 32674
rect 41074 32622 41076 32674
rect 40908 32620 41076 32622
rect 40236 31892 40404 31948
rect 40348 31890 40404 31892
rect 40348 31838 40350 31890
rect 40402 31838 40404 31890
rect 40348 31826 40404 31838
rect 40236 31780 40292 31790
rect 40236 31686 40292 31724
rect 40796 31666 40852 31678
rect 40796 31614 40798 31666
rect 40850 31614 40852 31666
rect 40124 30270 40126 30322
rect 40178 30270 40180 30322
rect 40124 30258 40180 30270
rect 40236 31220 40292 31230
rect 40236 30210 40292 31164
rect 40796 31108 40852 31614
rect 40796 31042 40852 31052
rect 40348 30994 40404 31006
rect 40348 30942 40350 30994
rect 40402 30942 40404 30994
rect 40348 30884 40404 30942
rect 40348 30818 40404 30828
rect 40908 30436 40964 32620
rect 41020 32610 41076 32620
rect 41132 32562 41188 32574
rect 41132 32510 41134 32562
rect 41186 32510 41188 32562
rect 41020 32338 41076 32350
rect 41020 32286 41022 32338
rect 41074 32286 41076 32338
rect 41020 30994 41076 32286
rect 41132 31220 41188 32510
rect 41468 32564 41524 33070
rect 41356 31892 41412 31902
rect 41356 31556 41412 31836
rect 41356 31490 41412 31500
rect 41132 31154 41188 31164
rect 41244 31444 41300 31454
rect 41020 30942 41022 30994
rect 41074 30942 41076 30994
rect 41020 30930 41076 30942
rect 41244 30994 41300 31388
rect 41244 30942 41246 30994
rect 41298 30942 41300 30994
rect 41244 30930 41300 30942
rect 40908 30370 40964 30380
rect 40236 30158 40238 30210
rect 40290 30158 40292 30210
rect 40236 30146 40292 30158
rect 40348 30324 40404 30334
rect 40348 29538 40404 30268
rect 41244 30324 41300 30334
rect 41244 30230 41300 30268
rect 41468 30100 41524 32508
rect 42140 32564 42196 32602
rect 42140 32498 42196 32508
rect 42476 32450 42532 33404
rect 42476 32398 42478 32450
rect 42530 32398 42532 32450
rect 42476 32386 42532 32398
rect 41804 32338 41860 32350
rect 41804 32286 41806 32338
rect 41858 32286 41860 32338
rect 41468 30006 41524 30044
rect 41692 31108 41748 31118
rect 41804 31108 41860 32286
rect 42140 32338 42196 32350
rect 42140 32286 42142 32338
rect 42194 32286 42196 32338
rect 42140 31948 42196 32286
rect 42140 31892 43092 31948
rect 43036 31780 43092 31892
rect 43596 31892 43652 33516
rect 44604 32674 44660 33852
rect 44604 32622 44606 32674
rect 44658 32622 44660 32674
rect 44604 32610 44660 32622
rect 45612 33572 45668 38612
rect 45948 38500 46004 38510
rect 45948 38162 46004 38444
rect 45948 38110 45950 38162
rect 46002 38110 46004 38162
rect 45948 38098 46004 38110
rect 46060 38388 46116 38398
rect 46060 37828 46116 38332
rect 46060 37266 46116 37772
rect 46060 37214 46062 37266
rect 46114 37214 46116 37266
rect 46060 37202 46116 37214
rect 45836 36708 45892 36718
rect 45724 36652 45836 36708
rect 45724 35698 45780 36652
rect 45836 36642 45892 36652
rect 45836 36260 45892 36270
rect 45836 36166 45892 36204
rect 45724 35646 45726 35698
rect 45778 35646 45780 35698
rect 45724 35634 45780 35646
rect 45612 32676 45668 33516
rect 45836 34692 45892 34702
rect 45836 33346 45892 34636
rect 45836 33294 45838 33346
rect 45890 33294 45892 33346
rect 45836 33282 45892 33294
rect 46172 33458 46228 40236
rect 46396 38668 46452 44940
rect 46508 43538 46564 43550
rect 46508 43486 46510 43538
rect 46562 43486 46564 43538
rect 46508 43316 46564 43486
rect 46508 43250 46564 43260
rect 46732 42644 46788 42654
rect 46732 42550 46788 42588
rect 46620 41860 46676 41870
rect 46620 41766 46676 41804
rect 46844 41636 46900 48412
rect 46956 48636 47124 48692
rect 46956 47124 47012 48636
rect 47180 48244 47236 48254
rect 47180 48150 47236 48188
rect 47964 48132 48020 48972
rect 48076 49028 48132 49646
rect 48076 48962 48132 48972
rect 48188 49586 48244 49598
rect 48188 49534 48190 49586
rect 48242 49534 48244 49586
rect 48076 48132 48132 48142
rect 47964 48130 48132 48132
rect 47964 48078 48078 48130
rect 48130 48078 48132 48130
rect 47964 48076 48132 48078
rect 48076 47684 48132 48076
rect 48188 48020 48244 49534
rect 48188 47954 48244 47964
rect 48188 47684 48244 47694
rect 48076 47628 48188 47684
rect 48188 47618 48244 47628
rect 47740 47572 47796 47582
rect 47068 47458 47124 47470
rect 47068 47406 47070 47458
rect 47122 47406 47124 47458
rect 47068 47348 47124 47406
rect 47068 47282 47124 47292
rect 47740 47346 47796 47516
rect 47740 47294 47742 47346
rect 47794 47294 47796 47346
rect 47740 47282 47796 47294
rect 47964 47570 48020 47582
rect 47964 47518 47966 47570
rect 48018 47518 48020 47570
rect 47964 47348 48020 47518
rect 48076 47460 48132 47470
rect 48076 47366 48132 47404
rect 47964 47282 48020 47292
rect 46956 47068 47124 47124
rect 46956 41972 47012 41982
rect 46956 41878 47012 41916
rect 46620 41580 46900 41636
rect 47068 41636 47124 47068
rect 47964 46562 48020 46574
rect 47964 46510 47966 46562
rect 48018 46510 48020 46562
rect 47180 46228 47236 46238
rect 47180 42754 47236 46172
rect 47516 45332 47572 45342
rect 47292 43652 47348 43662
rect 47292 43538 47348 43596
rect 47292 43486 47294 43538
rect 47346 43486 47348 43538
rect 47292 43474 47348 43486
rect 47404 43316 47460 43326
rect 47404 43222 47460 43260
rect 47180 42702 47182 42754
rect 47234 42702 47236 42754
rect 47180 42690 47236 42702
rect 47292 42644 47348 42654
rect 47292 42550 47348 42588
rect 47516 42420 47572 45276
rect 47628 43540 47684 43550
rect 47628 43446 47684 43484
rect 46396 38612 46564 38668
rect 46396 37828 46452 37838
rect 46284 37826 46452 37828
rect 46284 37774 46398 37826
rect 46450 37774 46452 37826
rect 46284 37772 46452 37774
rect 46284 37492 46340 37772
rect 46396 37762 46452 37772
rect 46284 36482 46340 37436
rect 46396 37380 46452 37390
rect 46396 37044 46452 37324
rect 46396 36978 46452 36988
rect 46508 36932 46564 38612
rect 46620 37268 46676 41580
rect 47068 41570 47124 41580
rect 47180 42364 47572 42420
rect 47628 42644 47684 42654
rect 47068 40852 47124 40862
rect 47180 40852 47236 42364
rect 47292 42196 47348 42206
rect 47292 42102 47348 42140
rect 47628 41972 47684 42588
rect 47852 42196 47908 42234
rect 47852 42130 47908 42140
rect 47124 40796 47236 40852
rect 47292 41970 47684 41972
rect 47292 41918 47630 41970
rect 47682 41918 47684 41970
rect 47292 41916 47684 41918
rect 46732 39732 46788 39742
rect 46732 37938 46788 39676
rect 46844 39060 46900 39070
rect 46844 38946 46900 39004
rect 46844 38894 46846 38946
rect 46898 38894 46900 38946
rect 46844 38882 46900 38894
rect 46732 37886 46734 37938
rect 46786 37886 46788 37938
rect 46732 37874 46788 37886
rect 46620 37202 46676 37212
rect 46732 37268 46788 37278
rect 46732 37266 46900 37268
rect 46732 37214 46734 37266
rect 46786 37214 46900 37266
rect 46732 37212 46900 37214
rect 46732 37202 46788 37212
rect 46508 36866 46564 36876
rect 46844 36484 46900 37212
rect 46284 36430 46286 36482
rect 46338 36430 46340 36482
rect 46284 36418 46340 36430
rect 46508 36482 46900 36484
rect 46508 36430 46846 36482
rect 46898 36430 46900 36482
rect 46508 36428 46900 36430
rect 46508 36370 46564 36428
rect 46844 36418 46900 36428
rect 46508 36318 46510 36370
rect 46562 36318 46564 36370
rect 46284 36260 46340 36270
rect 46284 35924 46340 36204
rect 46508 35924 46564 36318
rect 46284 35922 46564 35924
rect 46284 35870 46286 35922
rect 46338 35870 46564 35922
rect 46284 35868 46564 35870
rect 46284 35858 46340 35868
rect 47068 35700 47124 40796
rect 47292 40626 47348 41916
rect 47628 41906 47684 41916
rect 47852 41972 47908 41982
rect 47292 40574 47294 40626
rect 47346 40574 47348 40626
rect 47180 37044 47236 37054
rect 47180 35922 47236 36988
rect 47292 36484 47348 40574
rect 47740 41858 47796 41870
rect 47740 41806 47742 41858
rect 47794 41806 47796 41858
rect 47628 40516 47684 40526
rect 47740 40516 47796 41806
rect 47852 40626 47908 41916
rect 47964 41300 48020 46510
rect 48076 44322 48132 44334
rect 48076 44270 48078 44322
rect 48130 44270 48132 44322
rect 48076 43764 48132 44270
rect 48300 43988 48356 52444
rect 48412 50428 48468 53004
rect 48524 52948 48580 52958
rect 48524 52162 48580 52892
rect 48748 52500 48804 53004
rect 48972 52948 49028 52958
rect 48972 52854 49028 52892
rect 49420 52946 49476 53452
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 49868 53060 49924 53070
rect 50988 53060 51044 53790
rect 49420 52894 49422 52946
rect 49474 52894 49476 52946
rect 49420 52882 49476 52894
rect 49756 53058 49924 53060
rect 49756 53006 49870 53058
rect 49922 53006 49924 53058
rect 49756 53004 49924 53006
rect 49756 52948 49812 53004
rect 49868 52994 49924 53004
rect 50652 53004 51044 53060
rect 51548 53506 51604 53518
rect 51548 53454 51550 53506
rect 51602 53454 51604 53506
rect 48860 52836 48916 52846
rect 48860 52742 48916 52780
rect 48748 52434 48804 52444
rect 48524 52110 48526 52162
rect 48578 52110 48580 52162
rect 48524 52098 48580 52110
rect 49308 52164 49364 52174
rect 49308 52070 49364 52108
rect 49644 52164 49700 52174
rect 49756 52164 49812 52892
rect 50204 52946 50260 52958
rect 50204 52894 50206 52946
rect 50258 52894 50260 52946
rect 50204 52388 50260 52894
rect 50652 52388 50708 53004
rect 50204 52332 50708 52388
rect 50540 52164 50596 52174
rect 49644 52162 49812 52164
rect 49644 52110 49646 52162
rect 49698 52110 49812 52162
rect 49644 52108 49812 52110
rect 49644 52098 49700 52108
rect 48972 52052 49028 52062
rect 48972 52050 49252 52052
rect 48972 51998 48974 52050
rect 49026 51998 49252 52050
rect 48972 51996 49252 51998
rect 48972 51986 49028 51996
rect 48748 51604 48804 51642
rect 48748 51538 48804 51548
rect 48860 51492 48916 51502
rect 48860 51378 48916 51436
rect 48860 51326 48862 51378
rect 48914 51326 48916 51378
rect 48412 50372 48580 50428
rect 48412 49700 48468 49710
rect 48412 49026 48468 49644
rect 48412 48974 48414 49026
rect 48466 48974 48468 49026
rect 48412 48962 48468 48974
rect 48524 47460 48580 50372
rect 48860 49924 48916 51326
rect 49196 51378 49252 51996
rect 49532 51938 49588 51950
rect 49532 51886 49534 51938
rect 49586 51886 49588 51938
rect 49532 51604 49588 51886
rect 49532 51548 49700 51604
rect 49196 51326 49198 51378
rect 49250 51326 49252 51378
rect 49196 51314 49252 51326
rect 49532 51378 49588 51390
rect 49532 51326 49534 51378
rect 49586 51326 49588 51378
rect 49084 51154 49140 51166
rect 49084 51102 49086 51154
rect 49138 51102 49140 51154
rect 49084 50596 49140 51102
rect 49420 50708 49476 50718
rect 49532 50708 49588 51326
rect 49420 50706 49588 50708
rect 49420 50654 49422 50706
rect 49474 50654 49588 50706
rect 49420 50652 49588 50654
rect 49420 50642 49476 50652
rect 49084 50530 49140 50540
rect 49532 50484 49588 50522
rect 49532 50418 49588 50428
rect 49084 50372 49140 50382
rect 49084 50278 49140 50316
rect 49308 50370 49364 50382
rect 49308 50318 49310 50370
rect 49362 50318 49364 50370
rect 49308 50148 49364 50318
rect 49308 50082 49364 50092
rect 49420 50372 49476 50382
rect 48860 49868 49252 49924
rect 48748 49812 48804 49822
rect 48636 49810 48804 49812
rect 48636 49758 48750 49810
rect 48802 49758 48804 49810
rect 48636 49756 48804 49758
rect 48636 49700 48692 49756
rect 48748 49746 48804 49756
rect 48636 49634 48692 49644
rect 48860 49586 48916 49598
rect 48860 49534 48862 49586
rect 48914 49534 48916 49586
rect 48748 49252 48804 49262
rect 48748 49138 48804 49196
rect 48748 49086 48750 49138
rect 48802 49086 48804 49138
rect 48748 49074 48804 49086
rect 48860 48916 48916 49534
rect 49084 49588 49140 49598
rect 49084 49494 49140 49532
rect 48636 48860 48916 48916
rect 48636 48356 48692 48860
rect 49084 48692 49140 48702
rect 48860 48468 48916 48478
rect 48860 48374 48916 48412
rect 48636 48290 48692 48300
rect 48972 48356 49028 48366
rect 48748 48132 48804 48142
rect 48748 47572 48804 48076
rect 48524 47404 48692 47460
rect 48524 47234 48580 47246
rect 48524 47182 48526 47234
rect 48578 47182 48580 47234
rect 48524 45220 48580 47182
rect 48636 46004 48692 47404
rect 48748 47458 48804 47516
rect 48748 47406 48750 47458
rect 48802 47406 48804 47458
rect 48748 47394 48804 47406
rect 48972 47460 49028 48300
rect 48972 47366 49028 47404
rect 48860 47236 48916 47246
rect 48860 47142 48916 47180
rect 48636 45910 48692 45948
rect 48524 45154 48580 45164
rect 48748 45444 48804 45454
rect 49084 45444 49140 48636
rect 48748 44994 48804 45388
rect 48748 44942 48750 44994
rect 48802 44942 48804 44994
rect 48748 44930 48804 44942
rect 48860 45388 49140 45444
rect 48860 45330 48916 45388
rect 48860 45278 48862 45330
rect 48914 45278 48916 45330
rect 48300 43932 48804 43988
rect 48636 43764 48692 43774
rect 48076 43762 48692 43764
rect 48076 43710 48638 43762
rect 48690 43710 48692 43762
rect 48076 43708 48692 43710
rect 48636 43698 48692 43708
rect 48188 43540 48244 43550
rect 48748 43540 48804 43932
rect 48188 43446 48244 43484
rect 48636 43484 48804 43540
rect 48300 41970 48356 41982
rect 48300 41918 48302 41970
rect 48354 41918 48356 41970
rect 48300 41860 48356 41918
rect 48300 41524 48356 41804
rect 48300 41458 48356 41468
rect 48524 41860 48580 41870
rect 47964 41234 48020 41244
rect 48524 41188 48580 41804
rect 48524 41122 48580 41132
rect 48300 41076 48356 41086
rect 47852 40574 47854 40626
rect 47906 40574 47908 40626
rect 47852 40562 47908 40574
rect 47964 41074 48356 41076
rect 47964 41022 48302 41074
rect 48354 41022 48356 41074
rect 47964 41020 48356 41022
rect 47628 40514 47796 40516
rect 47628 40462 47630 40514
rect 47682 40462 47796 40514
rect 47628 40460 47796 40462
rect 47628 40450 47684 40460
rect 47964 40290 48020 41020
rect 48300 41010 48356 41020
rect 47964 40238 47966 40290
rect 48018 40238 48020 40290
rect 47964 40226 48020 40238
rect 48076 40404 48132 40414
rect 48076 39060 48132 40348
rect 48412 39396 48468 39406
rect 48412 39302 48468 39340
rect 47628 39058 48132 39060
rect 47628 39006 48078 39058
rect 48130 39006 48132 39058
rect 47628 39004 48132 39006
rect 47628 38834 47684 39004
rect 48076 38994 48132 39004
rect 47628 38782 47630 38834
rect 47682 38782 47684 38834
rect 47404 37156 47460 37166
rect 47628 37156 47684 38782
rect 47404 37154 47572 37156
rect 47404 37102 47406 37154
rect 47458 37102 47572 37154
rect 47404 37100 47572 37102
rect 47404 37090 47460 37100
rect 47404 36484 47460 36494
rect 47292 36482 47460 36484
rect 47292 36430 47406 36482
rect 47458 36430 47460 36482
rect 47292 36428 47460 36430
rect 47404 36036 47460 36428
rect 47404 35970 47460 35980
rect 47180 35870 47182 35922
rect 47234 35870 47236 35922
rect 47180 35858 47236 35870
rect 47516 35924 47572 37100
rect 47516 35858 47572 35868
rect 47068 35644 47236 35700
rect 46732 35476 46788 35486
rect 46396 34802 46452 34814
rect 46396 34750 46398 34802
rect 46450 34750 46452 34802
rect 46284 34692 46340 34702
rect 46396 34692 46452 34750
rect 46732 34802 46788 35420
rect 47068 34916 47124 34926
rect 46732 34750 46734 34802
rect 46786 34750 46788 34802
rect 46732 34738 46788 34750
rect 46956 34860 47068 34916
rect 46340 34636 46676 34692
rect 46284 34626 46340 34636
rect 46172 33406 46174 33458
rect 46226 33406 46228 33458
rect 46172 33012 46228 33406
rect 46620 33348 46676 34636
rect 46172 32946 46228 32956
rect 46284 33346 46676 33348
rect 46284 33294 46622 33346
rect 46674 33294 46676 33346
rect 46284 33292 46676 33294
rect 46284 32786 46340 33292
rect 46620 33282 46676 33292
rect 46284 32734 46286 32786
rect 46338 32734 46340 32786
rect 46284 32722 46340 32734
rect 45724 32676 45780 32686
rect 45612 32674 45780 32676
rect 45612 32622 45726 32674
rect 45778 32622 45780 32674
rect 45612 32620 45780 32622
rect 45724 32610 45780 32620
rect 45388 32564 45444 32574
rect 45388 32470 45444 32508
rect 46732 32564 46788 32574
rect 46956 32564 47012 34860
rect 47068 34822 47124 34860
rect 46788 32508 47012 32564
rect 47180 33346 47236 35644
rect 47628 34916 47684 37100
rect 48412 38612 48468 38622
rect 48412 38162 48468 38556
rect 48412 38110 48414 38162
rect 48466 38110 48468 38162
rect 48412 37044 48468 38110
rect 48188 36932 48244 36942
rect 48188 36596 48244 36876
rect 47964 36482 48020 36494
rect 47964 36430 47966 36482
rect 48018 36430 48020 36482
rect 47852 36260 47908 36270
rect 47740 35924 47796 35934
rect 47740 35830 47796 35868
rect 47852 35026 47908 36204
rect 47964 35924 48020 36430
rect 48188 36482 48244 36540
rect 48188 36430 48190 36482
rect 48242 36430 48244 36482
rect 48188 36418 48244 36430
rect 48300 36260 48356 36270
rect 48300 36166 48356 36204
rect 48412 36036 48468 36988
rect 48636 36708 48692 43484
rect 48748 42194 48804 42206
rect 48748 42142 48750 42194
rect 48802 42142 48804 42194
rect 48748 42084 48804 42142
rect 48748 42018 48804 42028
rect 48860 41748 48916 45278
rect 49084 44882 49140 44894
rect 49084 44830 49086 44882
rect 49138 44830 49140 44882
rect 48972 44212 49028 44222
rect 48972 42866 49028 44156
rect 49084 44212 49140 44830
rect 49196 44548 49252 49868
rect 49308 49812 49364 49822
rect 49420 49812 49476 50316
rect 49364 49756 49476 49812
rect 49644 49810 49700 51548
rect 49644 49758 49646 49810
rect 49698 49758 49700 49810
rect 49308 49718 49364 49756
rect 49308 48468 49364 48478
rect 49308 48374 49364 48412
rect 49644 48354 49700 49758
rect 49644 48302 49646 48354
rect 49698 48302 49700 48354
rect 49644 48290 49700 48302
rect 49532 47684 49588 47694
rect 49756 47684 49812 52108
rect 50428 52162 50596 52164
rect 50428 52110 50542 52162
rect 50594 52110 50596 52162
rect 50428 52108 50596 52110
rect 49868 52052 49924 52062
rect 49868 51958 49924 51996
rect 50092 51268 50148 51278
rect 50092 51266 50372 51268
rect 50092 51214 50094 51266
rect 50146 51214 50372 51266
rect 50092 51212 50372 51214
rect 50092 51202 50148 51212
rect 49868 50484 49924 50522
rect 49868 50418 49924 50428
rect 50092 50484 50148 50494
rect 49980 50372 50036 50382
rect 49980 50278 50036 50316
rect 50092 50370 50148 50428
rect 50316 50482 50372 51212
rect 50428 51156 50484 52108
rect 50540 52098 50596 52108
rect 50652 51940 50708 52332
rect 50764 52836 50820 52846
rect 50764 52274 50820 52780
rect 50876 52834 50932 52846
rect 50876 52782 50878 52834
rect 50930 52782 50932 52834
rect 50876 52388 50932 52782
rect 50876 52322 50932 52332
rect 51548 52500 51604 53454
rect 50764 52222 50766 52274
rect 50818 52222 50820 52274
rect 50764 52210 50820 52222
rect 50876 52164 50932 52174
rect 51324 52164 51380 52174
rect 50876 52162 51380 52164
rect 50876 52110 50878 52162
rect 50930 52110 51326 52162
rect 51378 52110 51380 52162
rect 50876 52108 51380 52110
rect 50876 52098 50932 52108
rect 51324 52098 51380 52108
rect 51436 52052 51492 52062
rect 51436 51958 51492 51996
rect 50652 51884 50932 51940
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50876 51604 50932 51884
rect 51212 51938 51268 51950
rect 51212 51886 51214 51938
rect 51266 51886 51268 51938
rect 51212 51716 51268 51886
rect 51548 51716 51604 52444
rect 51884 53508 51940 53518
rect 51884 52276 51940 53452
rect 53788 52946 53844 52958
rect 53788 52894 53790 52946
rect 53842 52894 53844 52946
rect 53004 52836 53060 52846
rect 53004 52742 53060 52780
rect 51884 52162 51940 52220
rect 52780 52276 52836 52286
rect 52780 52182 52836 52220
rect 51884 52110 51886 52162
rect 51938 52110 51940 52162
rect 51884 52098 51940 52110
rect 51212 51660 51604 51716
rect 51996 52052 52052 52062
rect 50764 51548 50932 51604
rect 50764 51380 50820 51548
rect 51660 51492 51716 51502
rect 51660 51398 51716 51436
rect 51996 51490 52052 51996
rect 51996 51438 51998 51490
rect 52050 51438 52052 51490
rect 51996 51426 52052 51438
rect 50764 51286 50820 51324
rect 51884 51380 51940 51390
rect 51884 51286 51940 51324
rect 50876 51268 50932 51278
rect 50876 51174 50932 51212
rect 52556 51266 52612 51278
rect 52556 51214 52558 51266
rect 52610 51214 52612 51266
rect 50428 51100 50820 51156
rect 50764 50818 50820 51100
rect 50764 50766 50766 50818
rect 50818 50766 50820 50818
rect 50764 50754 50820 50766
rect 50316 50430 50318 50482
rect 50370 50430 50372 50482
rect 50316 50418 50372 50430
rect 50876 50594 50932 50606
rect 50876 50542 50878 50594
rect 50930 50542 50932 50594
rect 50876 50484 50932 50542
rect 50876 50418 50932 50428
rect 51100 50594 51156 50606
rect 51100 50542 51102 50594
rect 51154 50542 51156 50594
rect 50092 50318 50094 50370
rect 50146 50318 50148 50370
rect 50092 50306 50148 50318
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50204 49924 50260 49934
rect 50204 49830 50260 49868
rect 51100 49924 51156 50542
rect 51324 50594 51380 50606
rect 51324 50542 51326 50594
rect 51378 50542 51380 50594
rect 51324 50428 51380 50542
rect 51772 50484 51828 50522
rect 51324 50372 51492 50428
rect 51772 50418 51828 50428
rect 52556 50428 52612 51214
rect 52780 51268 52836 51278
rect 53340 51268 53396 51278
rect 52836 51212 52948 51268
rect 52780 51202 52836 51212
rect 52780 50596 52836 50634
rect 52668 50540 52780 50596
rect 52668 50428 52724 50540
rect 52780 50530 52836 50540
rect 52892 50428 52948 51212
rect 53340 51174 53396 51212
rect 53004 51156 53060 51166
rect 53004 50594 53060 51100
rect 53004 50542 53006 50594
rect 53058 50542 53060 50594
rect 53004 50530 53060 50542
rect 51100 49858 51156 49868
rect 50764 49812 50820 49822
rect 50092 49700 50148 49710
rect 50092 49606 50148 49644
rect 49868 49586 49924 49598
rect 49868 49534 49870 49586
rect 49922 49534 49924 49586
rect 49868 48804 49924 49534
rect 50204 49588 50260 49598
rect 49868 48466 49924 48748
rect 49868 48414 49870 48466
rect 49922 48414 49924 48466
rect 49868 48402 49924 48414
rect 50092 49252 50148 49262
rect 49980 48020 50036 48030
rect 49980 47926 50036 47964
rect 50092 47908 50148 49196
rect 50092 47842 50148 47852
rect 49532 47682 49812 47684
rect 49532 47630 49534 47682
rect 49586 47630 49812 47682
rect 49532 47628 49812 47630
rect 50204 47682 50260 49532
rect 50764 49252 50820 49756
rect 50876 49700 50932 49710
rect 50876 49698 51044 49700
rect 50876 49646 50878 49698
rect 50930 49646 51044 49698
rect 50876 49644 51044 49646
rect 50876 49634 50932 49644
rect 50540 49028 50596 49038
rect 50540 48934 50596 48972
rect 50428 48916 50484 48926
rect 50428 48132 50484 48860
rect 50764 48804 50820 49196
rect 50764 48748 50932 48804
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50540 48468 50596 48478
rect 50876 48468 50932 48748
rect 50540 48466 50932 48468
rect 50540 48414 50542 48466
rect 50594 48414 50932 48466
rect 50540 48412 50932 48414
rect 50540 48402 50596 48412
rect 50988 48242 51044 49644
rect 50988 48190 50990 48242
rect 51042 48190 51044 48242
rect 50988 48178 51044 48190
rect 51100 49138 51156 49150
rect 51100 49086 51102 49138
rect 51154 49086 51156 49138
rect 50204 47630 50206 47682
rect 50258 47630 50260 47682
rect 49532 47618 49588 47628
rect 50204 47618 50260 47630
rect 50316 48076 50484 48132
rect 50316 47682 50372 48076
rect 50316 47630 50318 47682
rect 50370 47630 50372 47682
rect 50316 47618 50372 47630
rect 50428 47908 50484 47918
rect 50428 47684 50484 47852
rect 50540 47684 50596 47694
rect 50428 47682 50596 47684
rect 50428 47630 50542 47682
rect 50594 47630 50596 47682
rect 50428 47628 50596 47630
rect 50540 47618 50596 47628
rect 50652 47684 50708 47694
rect 51100 47684 51156 49086
rect 50652 47590 50708 47628
rect 50988 47682 51156 47684
rect 50988 47630 51102 47682
rect 51154 47630 51156 47682
rect 50988 47628 51156 47630
rect 49196 44482 49252 44492
rect 49308 47458 49364 47470
rect 49308 47406 49310 47458
rect 49362 47406 49364 47458
rect 49308 47348 49364 47406
rect 49756 47460 49812 47470
rect 49756 47366 49812 47404
rect 49308 44322 49364 47292
rect 49532 47348 49588 47358
rect 49420 47234 49476 47246
rect 49420 47182 49422 47234
rect 49474 47182 49476 47234
rect 49420 46452 49476 47182
rect 49420 46386 49476 46396
rect 49308 44270 49310 44322
rect 49362 44270 49364 44322
rect 49308 44258 49364 44270
rect 49532 45890 49588 47292
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 49532 45838 49534 45890
rect 49586 45838 49588 45890
rect 49196 44212 49252 44222
rect 49084 44156 49196 44212
rect 49084 43540 49140 44156
rect 49196 44146 49252 44156
rect 49084 43474 49140 43484
rect 49196 43652 49252 43662
rect 49196 43204 49252 43596
rect 49420 43540 49476 43550
rect 49420 43446 49476 43484
rect 49532 43426 49588 45838
rect 49644 46674 49700 46686
rect 49644 46622 49646 46674
rect 49698 46622 49700 46674
rect 49644 44994 49700 46622
rect 50204 46676 50260 46686
rect 50204 46582 50260 46620
rect 49868 46564 49924 46574
rect 49868 46470 49924 46508
rect 50316 46564 50372 46574
rect 50092 46452 50148 46462
rect 50092 45890 50148 46396
rect 50204 46004 50260 46014
rect 50316 46004 50372 46508
rect 50764 46564 50820 46574
rect 50764 46470 50820 46508
rect 50652 46450 50708 46462
rect 50652 46398 50654 46450
rect 50706 46398 50708 46450
rect 50204 46002 50372 46004
rect 50204 45950 50206 46002
rect 50258 45950 50372 46002
rect 50204 45948 50372 45950
rect 50540 46340 50596 46350
rect 50204 45938 50260 45948
rect 50092 45838 50094 45890
rect 50146 45838 50148 45890
rect 50092 45826 50148 45838
rect 50540 45892 50596 46284
rect 50540 45826 50596 45836
rect 50540 45668 50596 45678
rect 50316 45666 50596 45668
rect 50316 45614 50542 45666
rect 50594 45614 50596 45666
rect 50316 45612 50596 45614
rect 50652 45668 50708 46398
rect 50988 46452 51044 47628
rect 51100 47618 51156 47628
rect 51324 48244 51380 48254
rect 51324 47460 51380 48188
rect 51436 47684 51492 50372
rect 51884 50372 51940 50382
rect 52556 50372 52724 50428
rect 51548 49810 51604 49822
rect 51548 49758 51550 49810
rect 51602 49758 51604 49810
rect 51548 49140 51604 49758
rect 51772 49812 51828 49822
rect 51884 49812 51940 50316
rect 51772 49810 52388 49812
rect 51772 49758 51774 49810
rect 51826 49758 52388 49810
rect 51772 49756 52388 49758
rect 51772 49746 51828 49756
rect 51548 48356 51604 49084
rect 51660 49364 51716 49374
rect 51660 49138 51716 49308
rect 51660 49086 51662 49138
rect 51714 49086 51716 49138
rect 51660 49074 51716 49086
rect 51996 49140 52052 49150
rect 51996 49046 52052 49084
rect 52108 49028 52164 49038
rect 52108 48934 52164 48972
rect 51548 48290 51604 48300
rect 52332 48916 52388 49756
rect 52668 49810 52724 50372
rect 52668 49758 52670 49810
rect 52722 49758 52724 49810
rect 52668 49746 52724 49758
rect 52780 50372 52948 50428
rect 53788 50428 53844 52894
rect 53900 51378 53956 51390
rect 53900 51326 53902 51378
rect 53954 51326 53956 51378
rect 53900 51156 53956 51326
rect 53900 51090 53956 51100
rect 54460 51156 54516 51166
rect 54516 51100 54628 51156
rect 54460 51090 54516 51100
rect 54460 50706 54516 50718
rect 54460 50654 54462 50706
rect 54514 50654 54516 50706
rect 54460 50596 54516 50654
rect 54460 50428 54516 50540
rect 54572 50594 54628 51100
rect 54572 50542 54574 50594
rect 54626 50542 54628 50594
rect 54572 50530 54628 50542
rect 54908 50596 54964 50606
rect 54908 50594 55300 50596
rect 54908 50542 54910 50594
rect 54962 50542 55300 50594
rect 54908 50540 55300 50542
rect 54908 50530 54964 50540
rect 53340 50372 53396 50382
rect 53788 50372 53956 50428
rect 54460 50372 54628 50428
rect 52780 49700 52836 50372
rect 53340 50278 53396 50316
rect 53116 49812 53172 49822
rect 53116 49718 53172 49756
rect 53788 49812 53844 49822
rect 53788 49718 53844 49756
rect 52780 49606 52836 49644
rect 53004 49586 53060 49598
rect 53004 49534 53006 49586
rect 53058 49534 53060 49586
rect 52668 49364 52724 49374
rect 52668 49026 52724 49308
rect 52892 49250 52948 49262
rect 52892 49198 52894 49250
rect 52946 49198 52948 49250
rect 52668 48974 52670 49026
rect 52722 48974 52724 49026
rect 52668 48962 52724 48974
rect 52780 49028 52836 49038
rect 52332 48242 52388 48860
rect 52332 48190 52334 48242
rect 52386 48190 52388 48242
rect 52332 48178 52388 48190
rect 52668 48244 52724 48254
rect 51884 48130 51940 48142
rect 51884 48078 51886 48130
rect 51938 48078 51940 48130
rect 51772 47684 51828 47694
rect 51436 47682 51828 47684
rect 51436 47630 51438 47682
rect 51490 47630 51774 47682
rect 51826 47630 51828 47682
rect 51436 47628 51828 47630
rect 51436 47618 51492 47628
rect 51772 47618 51828 47628
rect 51884 47460 51940 48078
rect 51996 47572 52052 47582
rect 51996 47478 52052 47516
rect 52668 47572 52724 48188
rect 52780 48242 52836 48972
rect 52780 48190 52782 48242
rect 52834 48190 52836 48242
rect 52780 48178 52836 48190
rect 51324 47404 51604 47460
rect 51324 47234 51380 47246
rect 51324 47182 51326 47234
rect 51378 47182 51380 47234
rect 51100 47124 51156 47134
rect 51100 46674 51156 47068
rect 51100 46622 51102 46674
rect 51154 46622 51156 46674
rect 51100 46610 51156 46622
rect 50988 46396 51156 46452
rect 50764 46340 50820 46350
rect 50764 45890 50820 46284
rect 50764 45838 50766 45890
rect 50818 45838 50820 45890
rect 50764 45826 50820 45838
rect 50876 45892 50932 45902
rect 50876 45798 50932 45836
rect 51100 45890 51156 46396
rect 51324 46340 51380 47182
rect 51324 46274 51380 46284
rect 51436 47236 51492 47246
rect 51100 45838 51102 45890
rect 51154 45838 51156 45890
rect 50652 45612 50932 45668
rect 49756 45444 49812 45454
rect 49756 45330 49812 45388
rect 50316 45332 50372 45612
rect 50540 45602 50596 45612
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 49756 45278 49758 45330
rect 49810 45278 49812 45330
rect 49756 45266 49812 45278
rect 49980 45276 50372 45332
rect 49980 45218 50036 45276
rect 50764 45220 50820 45230
rect 50876 45220 50932 45612
rect 49980 45166 49982 45218
rect 50034 45166 50036 45218
rect 49980 45154 50036 45166
rect 50540 45218 50932 45220
rect 50540 45166 50766 45218
rect 50818 45166 50932 45218
rect 50540 45164 50932 45166
rect 49644 44942 49646 44994
rect 49698 44942 49700 44994
rect 49644 44930 49700 44942
rect 50316 45108 50372 45118
rect 50204 44212 50260 44222
rect 50092 44100 50148 44110
rect 50092 44006 50148 44044
rect 49532 43374 49534 43426
rect 49586 43374 49588 43426
rect 49532 43362 49588 43374
rect 49644 43540 49700 43550
rect 48972 42814 48974 42866
rect 49026 42814 49028 42866
rect 48972 42802 49028 42814
rect 49084 43148 49252 43204
rect 48860 41682 48916 41692
rect 48972 41972 49028 41982
rect 49084 41972 49140 43148
rect 49644 42196 49700 43484
rect 49644 42130 49700 42140
rect 49868 43316 49924 43326
rect 49532 42084 49588 42094
rect 49532 41990 49588 42028
rect 48972 41970 49140 41972
rect 48972 41918 48974 41970
rect 49026 41918 49140 41970
rect 48972 41916 49140 41918
rect 49196 41970 49252 41982
rect 49196 41918 49198 41970
rect 49250 41918 49252 41970
rect 48972 41524 49028 41916
rect 49084 41748 49140 41758
rect 49084 41654 49140 41692
rect 49196 41636 49252 41918
rect 49196 41570 49252 41580
rect 48860 41468 49028 41524
rect 48748 40964 48804 40974
rect 48748 40626 48804 40908
rect 48748 40574 48750 40626
rect 48802 40574 48804 40626
rect 48748 40562 48804 40574
rect 48860 40404 48916 41468
rect 48972 41300 49028 41310
rect 48972 41186 49028 41244
rect 48972 41134 48974 41186
rect 49026 41134 49028 41186
rect 48972 41122 49028 41134
rect 49532 41300 49588 41310
rect 49532 40626 49588 41244
rect 49756 40964 49812 40974
rect 49756 40870 49812 40908
rect 49532 40574 49534 40626
rect 49586 40574 49588 40626
rect 49084 40516 49140 40526
rect 49084 40422 49140 40460
rect 48748 40348 48916 40404
rect 49532 40404 49588 40574
rect 48748 39396 48804 40348
rect 49532 40338 49588 40348
rect 48748 39330 48804 39340
rect 48860 39620 48916 39630
rect 48860 38834 48916 39564
rect 48860 38782 48862 38834
rect 48914 38782 48916 38834
rect 48860 38612 48916 38782
rect 48860 38546 48916 38556
rect 49084 39396 49140 39406
rect 49084 38724 49140 39340
rect 49196 38724 49252 38734
rect 49084 38722 49252 38724
rect 49084 38670 49198 38722
rect 49250 38670 49252 38722
rect 49084 38668 49252 38670
rect 49084 38276 49140 38668
rect 49196 38658 49252 38668
rect 49868 38668 49924 43260
rect 50204 43204 50260 44156
rect 50316 44210 50372 45052
rect 50428 44324 50484 44334
rect 50540 44324 50596 45164
rect 50764 45154 50820 45164
rect 51100 45108 51156 45838
rect 51324 45892 51380 45902
rect 51436 45892 51492 47180
rect 51324 45890 51492 45892
rect 51324 45838 51326 45890
rect 51378 45838 51492 45890
rect 51324 45836 51492 45838
rect 51324 45826 51380 45836
rect 51100 45014 51156 45052
rect 50428 44322 50596 44324
rect 50428 44270 50430 44322
rect 50482 44270 50596 44322
rect 50428 44268 50596 44270
rect 51212 44994 51268 45006
rect 51212 44942 51214 44994
rect 51266 44942 51268 44994
rect 50428 44258 50484 44268
rect 50316 44158 50318 44210
rect 50370 44158 50372 44210
rect 50316 44146 50372 44158
rect 50764 44210 50820 44222
rect 50764 44158 50766 44210
rect 50818 44158 50820 44210
rect 50764 44100 50820 44158
rect 50876 44212 50932 44222
rect 50876 44118 50932 44156
rect 51100 44212 51156 44222
rect 51100 44118 51156 44156
rect 50764 44034 50820 44044
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50316 43764 50372 43774
rect 50316 43538 50372 43708
rect 50316 43486 50318 43538
rect 50370 43486 50372 43538
rect 50316 43474 50372 43486
rect 50540 43316 50596 43326
rect 50428 43314 50596 43316
rect 50428 43262 50542 43314
rect 50594 43262 50596 43314
rect 50428 43260 50596 43262
rect 50204 43148 50372 43204
rect 50204 41860 50260 41870
rect 49980 41858 50260 41860
rect 49980 41806 50206 41858
rect 50258 41806 50260 41858
rect 49980 41804 50260 41806
rect 49980 41186 50036 41804
rect 50204 41794 50260 41804
rect 49980 41134 49982 41186
rect 50034 41134 50036 41186
rect 49980 40964 50036 41134
rect 50092 41188 50148 41198
rect 50092 41094 50148 41132
rect 50204 41076 50260 41086
rect 50204 40982 50260 41020
rect 49980 40898 50036 40908
rect 50204 40516 50260 40526
rect 50316 40516 50372 43148
rect 50428 42084 50484 43260
rect 50540 43250 50596 43260
rect 50876 43316 50932 43326
rect 50876 43222 50932 43260
rect 50876 42980 50932 42990
rect 50764 42924 50876 42980
rect 50764 42532 50820 42924
rect 50876 42914 50932 42924
rect 50988 42756 51044 42794
rect 50988 42690 51044 42700
rect 50876 42642 50932 42654
rect 50876 42590 50878 42642
rect 50930 42590 50932 42642
rect 50876 42532 50932 42590
rect 50764 42476 50932 42532
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50540 42084 50596 42094
rect 50428 42028 50540 42084
rect 50540 42018 50596 42028
rect 51100 41860 51156 41870
rect 51100 41766 51156 41804
rect 50652 41748 50708 41758
rect 50540 41636 50596 41646
rect 50540 41186 50596 41580
rect 50652 41298 50708 41692
rect 51212 41636 51268 44942
rect 51436 44098 51492 44110
rect 51436 44046 51438 44098
rect 51490 44046 51492 44098
rect 51436 43764 51492 44046
rect 51436 43698 51492 43708
rect 51324 43428 51380 43438
rect 51324 43092 51380 43372
rect 51324 43026 51380 43036
rect 51436 43316 51492 43326
rect 51436 42980 51492 43260
rect 51548 43204 51604 47404
rect 51884 47124 51940 47404
rect 52108 47460 52164 47470
rect 52108 47458 52388 47460
rect 52108 47406 52110 47458
rect 52162 47406 52388 47458
rect 52108 47404 52388 47406
rect 52108 47394 52164 47404
rect 51884 47058 51940 47068
rect 52108 47124 52164 47134
rect 52108 46898 52164 47068
rect 52108 46846 52110 46898
rect 52162 46846 52164 46898
rect 52108 46834 52164 46846
rect 51660 46788 51716 46798
rect 51660 46694 51716 46732
rect 51884 46674 51940 46686
rect 51884 46622 51886 46674
rect 51938 46622 51940 46674
rect 51772 45668 51828 45678
rect 51884 45668 51940 46622
rect 52220 46676 52276 46686
rect 52220 46582 52276 46620
rect 52332 45780 52388 47404
rect 52668 47458 52724 47516
rect 52668 47406 52670 47458
rect 52722 47406 52724 47458
rect 52668 47394 52724 47406
rect 52780 47348 52836 47358
rect 52556 47012 52612 47022
rect 52332 45714 52388 45724
rect 52444 46676 52500 46686
rect 51772 45666 51940 45668
rect 51772 45614 51774 45666
rect 51826 45614 51940 45666
rect 51772 45612 51940 45614
rect 51772 45602 51828 45612
rect 51548 43138 51604 43148
rect 51772 43538 51828 43550
rect 51772 43486 51774 43538
rect 51826 43486 51828 43538
rect 51772 42980 51828 43486
rect 51436 42924 51716 42980
rect 51660 42756 51716 42924
rect 51772 42914 51828 42924
rect 51884 42868 51940 45612
rect 52444 45332 52500 46620
rect 52444 45266 52500 45276
rect 52556 46674 52612 46956
rect 52556 46622 52558 46674
rect 52610 46622 52612 46674
rect 52556 45668 52612 46622
rect 52780 46676 52836 47292
rect 52892 47234 52948 49198
rect 53004 49028 53060 49534
rect 53452 49252 53508 49262
rect 53116 49028 53172 49038
rect 53060 49026 53172 49028
rect 53060 48974 53118 49026
rect 53170 48974 53172 49026
rect 53060 48972 53172 48974
rect 53004 48934 53060 48972
rect 53116 48962 53172 48972
rect 53452 49026 53508 49196
rect 53452 48974 53454 49026
rect 53506 48974 53508 49026
rect 53452 48962 53508 48974
rect 53900 49026 53956 50372
rect 54572 49810 54628 50372
rect 55020 50370 55076 50382
rect 55020 50318 55022 50370
rect 55074 50318 55076 50370
rect 54572 49758 54574 49810
rect 54626 49758 54628 49810
rect 54572 49746 54628 49758
rect 54684 49810 54740 49822
rect 54684 49758 54686 49810
rect 54738 49758 54740 49810
rect 53900 48974 53902 49026
rect 53954 48974 53956 49026
rect 53340 48916 53396 48926
rect 53340 48822 53396 48860
rect 53564 48244 53620 48254
rect 53564 48150 53620 48188
rect 53788 48242 53844 48254
rect 53788 48190 53790 48242
rect 53842 48190 53844 48242
rect 53228 48132 53284 48142
rect 53116 48130 53284 48132
rect 53116 48078 53230 48130
rect 53282 48078 53284 48130
rect 53116 48076 53284 48078
rect 53004 47460 53060 47470
rect 53004 47366 53060 47404
rect 53116 47348 53172 48076
rect 53228 48066 53284 48076
rect 53676 48130 53732 48142
rect 53676 48078 53678 48130
rect 53730 48078 53732 48130
rect 53228 47460 53284 47470
rect 53676 47460 53732 48078
rect 53788 47572 53844 48190
rect 53788 47506 53844 47516
rect 53228 47458 53732 47460
rect 53228 47406 53230 47458
rect 53282 47406 53732 47458
rect 53228 47404 53732 47406
rect 53228 47394 53284 47404
rect 53116 47282 53172 47292
rect 53788 47348 53844 47358
rect 53788 47254 53844 47292
rect 52892 47182 52894 47234
rect 52946 47182 52948 47234
rect 52892 47170 52948 47182
rect 53452 47236 53508 47246
rect 53452 47142 53508 47180
rect 53676 47234 53732 47246
rect 53676 47182 53678 47234
rect 53730 47182 53732 47234
rect 53452 47012 53508 47022
rect 53676 47012 53732 47182
rect 53508 46956 53732 47012
rect 53900 47012 53956 48974
rect 54124 49698 54180 49710
rect 54124 49646 54126 49698
rect 54178 49646 54180 49698
rect 54012 48354 54068 48366
rect 54012 48302 54014 48354
rect 54066 48302 54068 48354
rect 54012 48020 54068 48302
rect 54124 48132 54180 49646
rect 54124 48066 54180 48076
rect 54460 49698 54516 49710
rect 54460 49646 54462 49698
rect 54514 49646 54516 49698
rect 54012 47954 54068 47964
rect 53452 46946 53508 46956
rect 53900 46946 53956 46956
rect 54236 47234 54292 47246
rect 54236 47182 54238 47234
rect 54290 47182 54292 47234
rect 54236 46900 54292 47182
rect 54012 46844 54292 46900
rect 53228 46788 53284 46798
rect 52892 46676 52948 46686
rect 52780 46674 52948 46676
rect 52780 46622 52894 46674
rect 52946 46622 52948 46674
rect 52780 46620 52948 46622
rect 52668 46002 52724 46014
rect 52668 45950 52670 46002
rect 52722 45950 52724 46002
rect 52668 45892 52724 45950
rect 52668 45826 52724 45836
rect 52892 45780 52948 46620
rect 53228 46674 53284 46732
rect 53228 46622 53230 46674
rect 53282 46622 53284 46674
rect 53004 46562 53060 46574
rect 53004 46510 53006 46562
rect 53058 46510 53060 46562
rect 53004 46004 53060 46510
rect 53228 46452 53284 46622
rect 53452 46676 53508 46686
rect 53452 46582 53508 46620
rect 53676 46674 53732 46686
rect 53676 46622 53678 46674
rect 53730 46622 53732 46674
rect 53228 46386 53284 46396
rect 53564 46564 53620 46574
rect 53004 45948 53396 46004
rect 53004 45780 53060 45790
rect 52892 45778 53060 45780
rect 52892 45726 53006 45778
rect 53058 45726 53060 45778
rect 52892 45724 53060 45726
rect 53004 45714 53060 45724
rect 52780 45668 52836 45678
rect 52556 45666 52836 45668
rect 52556 45614 52782 45666
rect 52834 45614 52836 45666
rect 52556 45612 52836 45614
rect 52220 44098 52276 44110
rect 52220 44046 52222 44098
rect 52274 44046 52276 44098
rect 52108 43538 52164 43550
rect 52108 43486 52110 43538
rect 52162 43486 52164 43538
rect 52108 43204 52164 43486
rect 52108 43138 52164 43148
rect 51884 42812 52164 42868
rect 51660 42754 52052 42756
rect 51660 42702 51662 42754
rect 51714 42702 52052 42754
rect 51660 42700 52052 42702
rect 51660 42690 51716 42700
rect 51324 42532 51380 42542
rect 51324 41970 51380 42476
rect 51324 41918 51326 41970
rect 51378 41918 51380 41970
rect 51324 41906 51380 41918
rect 51436 42530 51492 42542
rect 51436 42478 51438 42530
rect 51490 42478 51492 42530
rect 50652 41246 50654 41298
rect 50706 41246 50708 41298
rect 50652 41234 50708 41246
rect 51100 41580 51212 41636
rect 50540 41134 50542 41186
rect 50594 41134 50596 41186
rect 50540 41076 50596 41134
rect 50988 41188 51044 41198
rect 50988 41094 51044 41132
rect 50540 41010 50596 41020
rect 50876 41074 50932 41086
rect 50876 41022 50878 41074
rect 50930 41022 50932 41074
rect 50876 40964 50932 41022
rect 50876 40898 50932 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 51100 40740 51156 41580
rect 51212 41570 51268 41580
rect 51436 41300 51492 42478
rect 51772 42530 51828 42542
rect 51772 42478 51774 42530
rect 51826 42478 51828 42530
rect 51772 41972 51828 42478
rect 51772 41906 51828 41916
rect 51884 42530 51940 42542
rect 51884 42478 51886 42530
rect 51938 42478 51940 42530
rect 51660 41412 51716 41422
rect 51884 41412 51940 42478
rect 51660 41410 51940 41412
rect 51660 41358 51662 41410
rect 51714 41358 51940 41410
rect 51660 41356 51940 41358
rect 51548 41300 51604 41310
rect 51100 40674 51156 40684
rect 51212 41244 51548 41300
rect 50260 40460 50372 40516
rect 50876 40514 50932 40526
rect 50876 40462 50878 40514
rect 50930 40462 50932 40514
rect 50204 40402 50260 40460
rect 50204 40350 50206 40402
rect 50258 40350 50260 40402
rect 50204 40338 50260 40350
rect 50428 39844 50484 39854
rect 50428 39620 50484 39788
rect 50876 39842 50932 40462
rect 50876 39790 50878 39842
rect 50930 39790 50932 39842
rect 50876 39778 50932 39790
rect 50988 40178 51044 40190
rect 50988 40126 50990 40178
rect 51042 40126 51044 40178
rect 50316 39564 50484 39620
rect 50540 39620 50596 39630
rect 50316 39172 50372 39564
rect 50428 39396 50484 39406
rect 50540 39396 50596 39564
rect 50428 39394 50596 39396
rect 50428 39342 50430 39394
rect 50482 39342 50596 39394
rect 50428 39340 50596 39342
rect 50428 39330 50484 39340
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50316 39116 50484 39172
rect 50556 39162 50820 39172
rect 50428 38836 50484 39116
rect 50988 39058 51044 40126
rect 51100 39620 51156 39630
rect 51212 39620 51268 41244
rect 51548 41206 51604 41244
rect 51660 41188 51716 41356
rect 51996 41300 52052 42700
rect 51884 41244 52052 41300
rect 51884 41188 51940 41244
rect 51660 41122 51716 41132
rect 51772 41186 51940 41188
rect 51772 41134 51886 41186
rect 51938 41134 51940 41186
rect 51772 41132 51940 41134
rect 51100 39618 51268 39620
rect 51100 39566 51102 39618
rect 51154 39566 51268 39618
rect 51100 39564 51268 39566
rect 51324 41076 51380 41086
rect 51324 39730 51380 41020
rect 51772 40964 51828 41132
rect 51884 41122 51940 41132
rect 51996 41074 52052 41086
rect 51996 41022 51998 41074
rect 52050 41022 52052 41074
rect 51324 39678 51326 39730
rect 51378 39678 51380 39730
rect 51100 39554 51156 39564
rect 50988 39006 50990 39058
rect 51042 39006 51044 39058
rect 50428 38742 50484 38780
rect 50652 38946 50708 38958
rect 50652 38894 50654 38946
rect 50706 38894 50708 38946
rect 50652 38724 50708 38894
rect 50540 38668 50652 38724
rect 49868 38612 50036 38668
rect 48860 38220 49140 38276
rect 48860 37490 48916 38220
rect 48860 37438 48862 37490
rect 48914 37438 48916 37490
rect 48860 36932 48916 37438
rect 48860 36866 48916 36876
rect 48972 38052 49028 38062
rect 48636 36642 48692 36652
rect 48524 36484 48580 36494
rect 48748 36484 48804 36494
rect 48524 36482 48804 36484
rect 48524 36430 48526 36482
rect 48578 36430 48750 36482
rect 48802 36430 48804 36482
rect 48524 36428 48804 36430
rect 48524 36418 48580 36428
rect 48748 36418 48804 36428
rect 48188 35980 48468 36036
rect 48076 35924 48132 35934
rect 47964 35922 48132 35924
rect 47964 35870 48078 35922
rect 48130 35870 48132 35922
rect 47964 35868 48132 35870
rect 48076 35858 48132 35868
rect 48188 35922 48244 35980
rect 48188 35870 48190 35922
rect 48242 35870 48244 35922
rect 48188 35858 48244 35870
rect 47964 35700 48020 35710
rect 47964 35606 48020 35644
rect 47852 34974 47854 35026
rect 47906 34974 47908 35026
rect 47852 34962 47908 34974
rect 47964 35252 48020 35262
rect 47740 34916 47796 34926
rect 47628 34860 47740 34916
rect 47740 34850 47796 34860
rect 47404 34018 47460 34030
rect 47404 33966 47406 34018
rect 47458 33966 47460 34018
rect 47404 33572 47460 33966
rect 47404 33506 47460 33516
rect 47964 33572 48020 35196
rect 47180 33294 47182 33346
rect 47234 33294 47236 33346
rect 46732 32470 46788 32508
rect 46508 32452 46564 32462
rect 45388 32004 45444 32014
rect 45388 31892 45556 31948
rect 43596 31826 43652 31836
rect 45500 31826 45556 31836
rect 46508 31890 46564 32396
rect 47180 32340 47236 33294
rect 47740 33234 47796 33246
rect 47740 33182 47742 33234
rect 47794 33182 47796 33234
rect 47516 32788 47572 32798
rect 47516 32694 47572 32732
rect 47180 32274 47236 32284
rect 47404 32450 47460 32462
rect 47404 32398 47406 32450
rect 47458 32398 47460 32450
rect 47404 32228 47460 32398
rect 47740 32452 47796 33182
rect 47964 33234 48020 33516
rect 47964 33182 47966 33234
rect 48018 33182 48020 33234
rect 47964 33170 48020 33182
rect 48076 34356 48132 34366
rect 47852 33124 47908 33134
rect 47852 33030 47908 33068
rect 47964 32788 48020 32798
rect 48076 32788 48132 34300
rect 48412 34132 48468 34142
rect 48412 33460 48468 34076
rect 47964 32786 48132 32788
rect 47964 32734 47966 32786
rect 48018 32734 48132 32786
rect 47964 32732 48132 32734
rect 48188 33458 48468 33460
rect 48188 33406 48414 33458
rect 48466 33406 48468 33458
rect 48188 33404 48468 33406
rect 47964 32722 48020 32732
rect 48188 32674 48244 33404
rect 48412 33394 48468 33404
rect 48860 33348 48916 33358
rect 48188 32622 48190 32674
rect 48242 32622 48244 32674
rect 48188 32610 48244 32622
rect 48748 33346 48916 33348
rect 48748 33294 48862 33346
rect 48914 33294 48916 33346
rect 48748 33292 48916 33294
rect 48748 32788 48804 33292
rect 48860 33282 48916 33292
rect 48860 33012 48916 33022
rect 48972 33012 49028 37996
rect 49868 38052 49924 38062
rect 49868 37958 49924 37996
rect 49756 37378 49812 37390
rect 49756 37326 49758 37378
rect 49810 37326 49812 37378
rect 49756 36708 49812 37326
rect 49532 36652 49924 36708
rect 49532 36594 49588 36652
rect 49532 36542 49534 36594
rect 49586 36542 49588 36594
rect 49532 36530 49588 36542
rect 49644 36482 49700 36494
rect 49644 36430 49646 36482
rect 49698 36430 49700 36482
rect 49644 36372 49700 36430
rect 49644 36306 49700 36316
rect 49868 35810 49924 36652
rect 49980 36484 50036 38612
rect 50428 38612 50596 38668
rect 50652 38658 50708 38668
rect 50428 38500 50484 38612
rect 50316 38444 50484 38500
rect 50204 37938 50260 37950
rect 50204 37886 50206 37938
rect 50258 37886 50260 37938
rect 50204 37492 50260 37886
rect 50316 37938 50372 38444
rect 50316 37886 50318 37938
rect 50370 37886 50372 37938
rect 50316 37874 50372 37886
rect 50540 37940 50596 37950
rect 50540 37846 50596 37884
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50204 37426 50260 37436
rect 50988 37380 51044 39006
rect 51324 38946 51380 39678
rect 51436 40908 51828 40964
rect 51884 40964 51940 40974
rect 51436 39618 51492 40908
rect 51660 40740 51716 40750
rect 51660 40402 51716 40684
rect 51660 40350 51662 40402
rect 51714 40350 51716 40402
rect 51660 40338 51716 40350
rect 51884 40402 51940 40908
rect 51884 40350 51886 40402
rect 51938 40350 51940 40402
rect 51884 40338 51940 40350
rect 51996 40292 52052 41022
rect 51996 40226 52052 40236
rect 52108 40068 52164 42812
rect 52220 42308 52276 44046
rect 52444 43652 52500 43662
rect 52556 43652 52612 45612
rect 52780 45602 52836 45612
rect 52668 45106 52724 45118
rect 52668 45054 52670 45106
rect 52722 45054 52724 45106
rect 52668 44884 52724 45054
rect 53340 45108 53396 45948
rect 53452 45892 53508 45902
rect 53564 45892 53620 46508
rect 53676 46004 53732 46622
rect 53900 46564 53956 46574
rect 53900 46470 53956 46508
rect 53676 45948 53844 46004
rect 53452 45890 53620 45892
rect 53452 45838 53454 45890
rect 53506 45838 53620 45890
rect 53452 45836 53620 45838
rect 53452 45826 53508 45836
rect 53676 45778 53732 45790
rect 53676 45726 53678 45778
rect 53730 45726 53732 45778
rect 53564 45108 53620 45118
rect 53340 45052 53564 45108
rect 53564 45014 53620 45052
rect 53676 44996 53732 45726
rect 53788 45220 53844 45948
rect 53900 45892 53956 45902
rect 54012 45892 54068 46844
rect 54460 46788 54516 49646
rect 54684 49700 54740 49758
rect 54684 49634 54740 49644
rect 54572 48916 54628 48926
rect 54572 48822 54628 48860
rect 54572 48130 54628 48142
rect 54572 48078 54574 48130
rect 54626 48078 54628 48130
rect 54572 48020 54628 48078
rect 54572 47954 54628 47964
rect 54460 46722 54516 46732
rect 54796 47458 54852 47470
rect 54796 47406 54798 47458
rect 54850 47406 54852 47458
rect 54796 47012 54852 47406
rect 54124 46676 54180 46686
rect 54124 46674 54292 46676
rect 54124 46622 54126 46674
rect 54178 46622 54292 46674
rect 54124 46620 54292 46622
rect 54124 46610 54180 46620
rect 53900 45890 54068 45892
rect 53900 45838 53902 45890
rect 53954 45838 54068 45890
rect 53900 45836 54068 45838
rect 53900 45826 53956 45836
rect 53788 45106 53844 45164
rect 53788 45054 53790 45106
rect 53842 45054 53844 45106
rect 53788 45042 53844 45054
rect 52892 44884 52948 44894
rect 53116 44884 53172 44894
rect 52668 44882 52948 44884
rect 52668 44830 52894 44882
rect 52946 44830 52948 44882
rect 52668 44828 52948 44830
rect 52444 43650 52612 43652
rect 52444 43598 52446 43650
rect 52498 43598 52612 43650
rect 52444 43596 52612 43598
rect 52780 43650 52836 44828
rect 52892 44818 52948 44828
rect 53004 44828 53116 44884
rect 53004 44212 53060 44828
rect 53116 44818 53172 44828
rect 53340 44884 53396 44894
rect 53340 44882 53508 44884
rect 53340 44830 53342 44882
rect 53394 44830 53508 44882
rect 53340 44828 53508 44830
rect 53340 44818 53396 44828
rect 53340 44548 53396 44558
rect 53228 44546 53396 44548
rect 53228 44494 53342 44546
rect 53394 44494 53396 44546
rect 53228 44492 53396 44494
rect 52780 43598 52782 43650
rect 52834 43598 52836 43650
rect 52444 42532 52500 43596
rect 52780 43586 52836 43598
rect 52892 44098 52948 44110
rect 52892 44046 52894 44098
rect 52946 44046 52948 44098
rect 52444 42466 52500 42476
rect 52556 42754 52612 42766
rect 52556 42702 52558 42754
rect 52610 42702 52612 42754
rect 52556 42308 52612 42702
rect 52892 42644 52948 44046
rect 53004 43650 53060 44156
rect 53004 43598 53006 43650
rect 53058 43598 53060 43650
rect 53004 43586 53060 43598
rect 53116 44322 53172 44334
rect 53116 44270 53118 44322
rect 53170 44270 53172 44322
rect 53116 43652 53172 44270
rect 53116 43586 53172 43596
rect 53116 43428 53172 43438
rect 53228 43428 53284 44492
rect 53340 44482 53396 44492
rect 53452 44324 53508 44828
rect 53564 44324 53620 44334
rect 53452 44268 53564 44324
rect 53564 44258 53620 44268
rect 53676 44322 53732 44940
rect 53676 44270 53678 44322
rect 53730 44270 53732 44322
rect 53676 44258 53732 44270
rect 53900 44324 53956 44334
rect 53900 44230 53956 44268
rect 53564 44098 53620 44110
rect 53564 44046 53566 44098
rect 53618 44046 53620 44098
rect 53564 43652 53620 44046
rect 53788 43652 53844 43662
rect 53564 43650 53844 43652
rect 53564 43598 53790 43650
rect 53842 43598 53844 43650
rect 53564 43596 53844 43598
rect 53788 43586 53844 43596
rect 53116 43426 53284 43428
rect 53116 43374 53118 43426
rect 53170 43374 53284 43426
rect 53116 43372 53284 43374
rect 53116 43362 53172 43372
rect 53564 43316 53620 43326
rect 53228 43314 53620 43316
rect 53228 43262 53566 43314
rect 53618 43262 53620 43314
rect 53228 43260 53620 43262
rect 53116 42868 53172 42878
rect 53228 42868 53284 43260
rect 53564 43250 53620 43260
rect 53900 43316 53956 43326
rect 53900 43222 53956 43260
rect 53676 43204 53732 43214
rect 53116 42866 53284 42868
rect 53116 42814 53118 42866
rect 53170 42814 53284 42866
rect 53116 42812 53284 42814
rect 53564 43092 53620 43102
rect 53116 42802 53172 42812
rect 53004 42756 53060 42766
rect 53004 42662 53060 42700
rect 52892 42578 52948 42588
rect 53228 42644 53284 42654
rect 53228 42550 53284 42588
rect 52220 42252 52612 42308
rect 52220 41970 52276 41982
rect 52220 41918 52222 41970
rect 52274 41918 52276 41970
rect 52220 40180 52276 41918
rect 52444 41972 52500 41982
rect 52444 41878 52500 41916
rect 52220 40114 52276 40124
rect 52556 41524 52612 42252
rect 53116 41972 53172 41982
rect 53452 41972 53508 41982
rect 53116 41970 53508 41972
rect 53116 41918 53118 41970
rect 53170 41918 53454 41970
rect 53506 41918 53508 41970
rect 53116 41916 53508 41918
rect 53116 41906 53172 41916
rect 53452 41906 53508 41916
rect 52892 41858 52948 41870
rect 52892 41806 52894 41858
rect 52946 41806 52948 41858
rect 52668 41748 52724 41758
rect 52668 41654 52724 41692
rect 51436 39566 51438 39618
rect 51490 39566 51492 39618
rect 51436 39554 51492 39566
rect 51996 40012 52164 40068
rect 51996 39508 52052 40012
rect 51996 39442 52052 39452
rect 52220 39508 52276 39518
rect 51436 39396 51492 39406
rect 51436 39058 51492 39340
rect 51436 39006 51438 39058
rect 51490 39006 51492 39058
rect 51436 38994 51492 39006
rect 51324 38894 51326 38946
rect 51378 38894 51380 38946
rect 51324 38882 51380 38894
rect 52220 38834 52276 39452
rect 52220 38782 52222 38834
rect 52274 38782 52276 38834
rect 51436 38724 51492 38734
rect 51324 38162 51380 38174
rect 51324 38110 51326 38162
rect 51378 38110 51380 38162
rect 50988 37314 51044 37324
rect 51100 37490 51156 37502
rect 51100 37438 51102 37490
rect 51154 37438 51156 37490
rect 50876 36596 50932 36606
rect 50092 36484 50148 36494
rect 49980 36482 50148 36484
rect 49980 36430 50094 36482
rect 50146 36430 50148 36482
rect 49980 36428 50148 36430
rect 50092 36418 50148 36428
rect 50876 36482 50932 36540
rect 50876 36430 50878 36482
rect 50930 36430 50932 36482
rect 50428 36370 50484 36382
rect 50428 36318 50430 36370
rect 50482 36318 50484 36370
rect 50316 36260 50372 36270
rect 50316 36166 50372 36204
rect 49868 35758 49870 35810
rect 49922 35758 49924 35810
rect 49868 35746 49924 35758
rect 49196 35700 49252 35710
rect 49196 35606 49252 35644
rect 49980 35700 50036 35710
rect 49532 35588 49588 35598
rect 49532 34130 49588 35532
rect 49980 35028 50036 35644
rect 50428 35140 50484 36318
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50764 35588 50820 35598
rect 50876 35588 50932 36430
rect 50820 35532 50932 35588
rect 50988 35586 51044 35598
rect 50988 35534 50990 35586
rect 51042 35534 51044 35586
rect 50764 35522 50820 35532
rect 50988 35476 51044 35534
rect 50988 35410 51044 35420
rect 50428 35084 50932 35140
rect 49532 34078 49534 34130
rect 49586 34078 49588 34130
rect 49532 34066 49588 34078
rect 49756 35026 50036 35028
rect 49756 34974 49982 35026
rect 50034 34974 50036 35026
rect 49756 34972 50036 34974
rect 49756 34132 49812 34972
rect 49980 34962 50036 34972
rect 50428 34916 50484 34926
rect 50428 34822 50484 34860
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50204 34356 50260 34366
rect 50204 34262 50260 34300
rect 50764 34244 50820 34254
rect 50764 34150 50820 34188
rect 50092 34132 50148 34142
rect 50428 34132 50484 34142
rect 49756 34130 50036 34132
rect 49756 34078 49758 34130
rect 49810 34078 50036 34130
rect 49756 34076 50036 34078
rect 49756 34066 49812 34076
rect 49084 33908 49140 33918
rect 49084 33124 49140 33852
rect 49196 33906 49252 33918
rect 49196 33854 49198 33906
rect 49250 33854 49252 33906
rect 49196 33348 49252 33854
rect 49308 33348 49364 33358
rect 49196 33346 49812 33348
rect 49196 33294 49310 33346
rect 49362 33294 49812 33346
rect 49196 33292 49812 33294
rect 49308 33282 49364 33292
rect 49644 33124 49700 33134
rect 49084 33068 49364 33124
rect 48972 32956 49252 33012
rect 48860 32900 48916 32956
rect 48860 32844 49028 32900
rect 48748 32674 48804 32732
rect 48748 32622 48750 32674
rect 48802 32622 48804 32674
rect 48748 32610 48804 32622
rect 48972 32562 49028 32844
rect 48972 32510 48974 32562
rect 49026 32510 49028 32562
rect 47852 32452 47908 32462
rect 47740 32450 47908 32452
rect 47740 32398 47854 32450
rect 47906 32398 47908 32450
rect 47740 32396 47908 32398
rect 47852 32386 47908 32396
rect 48860 32452 48916 32462
rect 48860 32358 48916 32396
rect 47404 32162 47460 32172
rect 48636 32228 48692 32238
rect 46508 31838 46510 31890
rect 46562 31838 46564 31890
rect 46508 31826 46564 31838
rect 48188 31892 48244 31902
rect 43484 31780 43540 31790
rect 43036 31778 43540 31780
rect 43036 31726 43486 31778
rect 43538 31726 43540 31778
rect 43036 31724 43540 31726
rect 43484 31714 43540 31724
rect 44268 31778 44324 31790
rect 44268 31726 44270 31778
rect 44322 31726 44324 31778
rect 44268 31556 44324 31726
rect 45836 31778 45892 31790
rect 45836 31726 45838 31778
rect 45890 31726 45892 31778
rect 42140 31220 42196 31230
rect 42140 31126 42196 31164
rect 41916 31108 41972 31118
rect 41804 31106 41972 31108
rect 41804 31054 41918 31106
rect 41970 31054 41972 31106
rect 41804 31052 41972 31054
rect 40908 29988 40964 29998
rect 40908 29894 40964 29932
rect 41356 29988 41412 29998
rect 41356 29894 41412 29932
rect 40348 29486 40350 29538
rect 40402 29486 40404 29538
rect 40348 29474 40404 29486
rect 40236 29428 40292 29438
rect 40236 29334 40292 29372
rect 41244 29314 41300 29326
rect 41244 29262 41246 29314
rect 41298 29262 41300 29314
rect 39788 28642 39956 28644
rect 39788 28590 39790 28642
rect 39842 28590 39956 28642
rect 39788 28588 39956 28590
rect 40124 29204 40180 29214
rect 40124 28644 40180 29148
rect 41244 28868 41300 29262
rect 41244 28802 41300 28812
rect 39788 28578 39844 28588
rect 40124 28550 40180 28588
rect 39564 28478 39566 28530
rect 39618 28478 39620 28530
rect 39564 28466 39620 28478
rect 38892 28364 39060 28420
rect 39676 28420 39732 28430
rect 37996 28082 38164 28084
rect 37996 28030 37998 28082
rect 38050 28030 38164 28082
rect 37996 28028 38164 28030
rect 38556 28084 38612 28094
rect 37436 26852 37604 26908
rect 37772 26964 37828 27002
rect 37996 26908 38052 28028
rect 38332 27972 38388 27982
rect 38332 27858 38388 27916
rect 38332 27806 38334 27858
rect 38386 27806 38388 27858
rect 38332 27794 38388 27806
rect 38556 27858 38612 28028
rect 38556 27806 38558 27858
rect 38610 27806 38612 27858
rect 38556 27794 38612 27806
rect 38892 27858 38948 28364
rect 38892 27806 38894 27858
rect 38946 27806 38948 27858
rect 38892 27794 38948 27806
rect 39340 27858 39396 27870
rect 39340 27806 39342 27858
rect 39394 27806 39396 27858
rect 39340 27748 39396 27806
rect 39340 27682 39396 27692
rect 37772 26898 37828 26908
rect 37884 26852 38052 26908
rect 37436 26740 37492 26852
rect 37436 26674 37492 26684
rect 37884 26516 37940 26852
rect 37100 26290 37268 26292
rect 37100 26238 37102 26290
rect 37154 26238 37268 26290
rect 37100 26236 37268 26238
rect 37324 26460 37940 26516
rect 39676 26514 39732 28364
rect 40236 28418 40292 28430
rect 40236 28366 40238 28418
rect 40290 28366 40292 28418
rect 39788 28084 39844 28094
rect 39788 27858 39844 28028
rect 40124 27972 40180 27982
rect 39788 27806 39790 27858
rect 39842 27806 39844 27858
rect 39788 27794 39844 27806
rect 40012 27916 40124 27972
rect 39788 27636 39844 27646
rect 39788 27542 39844 27580
rect 39900 27188 39956 27198
rect 40012 27188 40068 27916
rect 40124 27878 40180 27916
rect 40236 27748 40292 28366
rect 40460 28420 40516 28430
rect 40460 28418 40852 28420
rect 40460 28366 40462 28418
rect 40514 28366 40852 28418
rect 40460 28364 40852 28366
rect 40460 28354 40516 28364
rect 40796 27858 40852 28364
rect 41692 27970 41748 31052
rect 41916 31042 41972 31052
rect 42364 31108 42420 31118
rect 42364 31014 42420 31052
rect 42476 30994 42532 31006
rect 42476 30942 42478 30994
rect 42530 30942 42532 30994
rect 42476 29428 42532 30942
rect 43372 29988 43428 29998
rect 43372 29538 43428 29932
rect 43372 29486 43374 29538
rect 43426 29486 43428 29538
rect 43372 29474 43428 29486
rect 42476 29362 42532 29372
rect 44044 29428 44100 29438
rect 44268 29428 44324 31500
rect 44940 31556 44996 31566
rect 44940 31462 44996 31500
rect 45388 31556 45444 31566
rect 45388 31462 45444 31500
rect 45836 31556 45892 31726
rect 45836 30212 45892 31500
rect 48188 31218 48244 31836
rect 48636 31890 48692 32172
rect 48636 31838 48638 31890
rect 48690 31838 48692 31890
rect 48636 31826 48692 31838
rect 48972 32004 49028 32510
rect 48188 31166 48190 31218
rect 48242 31166 48244 31218
rect 48188 31154 48244 31166
rect 48860 31220 48916 31230
rect 48972 31220 49028 31948
rect 48860 31218 49028 31220
rect 48860 31166 48862 31218
rect 48914 31166 49028 31218
rect 48860 31164 49028 31166
rect 49196 32562 49252 32956
rect 49196 32510 49198 32562
rect 49250 32510 49252 32562
rect 49196 31892 49252 32510
rect 49308 32564 49364 33068
rect 49644 32674 49700 33068
rect 49756 33012 49812 33292
rect 49980 33236 50036 34076
rect 50092 34038 50148 34076
rect 50316 34130 50484 34132
rect 50316 34078 50430 34130
rect 50482 34078 50484 34130
rect 50316 34076 50484 34078
rect 50316 33908 50372 34076
rect 50428 34066 50484 34076
rect 50316 33842 50372 33852
rect 50876 33460 50932 35084
rect 51100 34356 51156 37438
rect 51324 37266 51380 38110
rect 51436 38050 51492 38668
rect 52220 38724 52276 38782
rect 52220 38658 52276 38668
rect 52332 38722 52388 38734
rect 52332 38670 52334 38722
rect 52386 38670 52388 38722
rect 51436 37998 51438 38050
rect 51490 37998 51492 38050
rect 51436 37986 51492 37998
rect 51660 38050 51716 38062
rect 51660 37998 51662 38050
rect 51714 37998 51716 38050
rect 51660 37604 51716 37998
rect 51660 37538 51716 37548
rect 51772 37828 51828 37838
rect 51324 37214 51326 37266
rect 51378 37214 51380 37266
rect 51324 36706 51380 37214
rect 51324 36654 51326 36706
rect 51378 36654 51380 36706
rect 51324 36642 51380 36654
rect 51436 36484 51492 36494
rect 51436 36148 51492 36428
rect 51436 36092 51604 36148
rect 51548 35922 51604 36092
rect 51548 35870 51550 35922
rect 51602 35870 51604 35922
rect 51548 35858 51604 35870
rect 51436 35810 51492 35822
rect 51436 35758 51438 35810
rect 51490 35758 51492 35810
rect 51436 35028 51492 35758
rect 51772 35812 51828 37772
rect 51996 37826 52052 37838
rect 51996 37774 51998 37826
rect 52050 37774 52052 37826
rect 51660 35588 51716 35598
rect 51660 35494 51716 35532
rect 51436 34962 51492 34972
rect 51772 35026 51828 35756
rect 51772 34974 51774 35026
rect 51826 34974 51828 35026
rect 51772 34962 51828 34974
rect 51884 36708 51940 36718
rect 51100 34290 51156 34300
rect 51660 34132 51716 34142
rect 51212 34130 51716 34132
rect 51212 34078 51662 34130
rect 51714 34078 51716 34130
rect 51212 34076 51716 34078
rect 50988 33460 51044 33470
rect 50876 33458 51044 33460
rect 50876 33406 50990 33458
rect 51042 33406 51044 33458
rect 50876 33404 51044 33406
rect 50988 33394 51044 33404
rect 50316 33348 50372 33358
rect 50092 33236 50148 33246
rect 49980 33234 50148 33236
rect 49980 33182 50094 33234
rect 50146 33182 50148 33234
rect 49980 33180 50148 33182
rect 50092 33170 50148 33180
rect 49756 32956 50148 33012
rect 49644 32622 49646 32674
rect 49698 32622 49700 32674
rect 49644 32610 49700 32622
rect 50092 32564 50148 32956
rect 50204 32564 50260 32574
rect 49308 32562 49588 32564
rect 49308 32510 49310 32562
rect 49362 32510 49588 32562
rect 49308 32508 49588 32510
rect 50092 32562 50260 32564
rect 50092 32510 50206 32562
rect 50258 32510 50260 32562
rect 50092 32508 50260 32510
rect 49308 32498 49364 32508
rect 48860 31154 48916 31164
rect 49196 30884 49252 31836
rect 49420 32340 49476 32350
rect 49420 31778 49476 32284
rect 49532 31948 49588 32508
rect 50204 32498 50260 32508
rect 49980 32450 50036 32462
rect 49980 32398 49982 32450
rect 50034 32398 50036 32450
rect 49980 32340 50036 32398
rect 50316 32340 50372 33292
rect 50652 33348 50708 33358
rect 50652 33254 50708 33292
rect 51212 33348 51268 34076
rect 51660 34066 51716 34076
rect 51324 33908 51380 33918
rect 51324 33814 51380 33852
rect 51436 33906 51492 33918
rect 51436 33854 51438 33906
rect 51490 33854 51492 33906
rect 51212 33346 51380 33348
rect 51212 33294 51214 33346
rect 51266 33294 51380 33346
rect 51212 33292 51380 33294
rect 51212 33282 51268 33292
rect 50540 33124 50596 33134
rect 49980 32284 50372 32340
rect 50428 33068 50540 33124
rect 50428 32788 50484 33068
rect 50540 33058 50596 33068
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 51324 32900 51380 33292
rect 51436 33124 51492 33854
rect 51436 33058 51492 33068
rect 51548 33908 51604 33918
rect 50556 32890 50820 32900
rect 51100 32844 51380 32900
rect 50540 32788 50596 32798
rect 50428 32786 50596 32788
rect 50428 32734 50542 32786
rect 50594 32734 50596 32786
rect 50428 32732 50596 32734
rect 49980 32228 50036 32284
rect 49980 32162 50036 32172
rect 49532 31892 49700 31948
rect 49420 31726 49422 31778
rect 49474 31726 49476 31778
rect 49420 31218 49476 31726
rect 49644 31778 49700 31892
rect 50428 31890 50484 32732
rect 50540 32722 50596 32732
rect 50428 31838 50430 31890
rect 50482 31838 50484 31890
rect 50428 31826 50484 31838
rect 49644 31726 49646 31778
rect 49698 31726 49700 31778
rect 49644 31668 49700 31726
rect 49980 31780 50036 31790
rect 49980 31686 50036 31724
rect 50764 31780 50820 31790
rect 50764 31778 50932 31780
rect 50764 31726 50766 31778
rect 50818 31726 50932 31778
rect 50764 31724 50932 31726
rect 50764 31714 50820 31724
rect 49644 31602 49700 31612
rect 49756 31554 49812 31566
rect 50540 31556 50596 31566
rect 49756 31502 49758 31554
rect 49810 31502 49812 31554
rect 49756 31332 49812 31502
rect 50428 31500 50540 31556
rect 49756 31276 50148 31332
rect 49420 31166 49422 31218
rect 49474 31166 49476 31218
rect 49420 31154 49476 31166
rect 50092 30994 50148 31276
rect 50428 31106 50484 31500
rect 50540 31490 50596 31500
rect 50876 31444 50932 31724
rect 51100 31444 51156 32844
rect 51548 32788 51604 33852
rect 51772 33906 51828 33918
rect 51772 33854 51774 33906
rect 51826 33854 51828 33906
rect 51212 32732 51604 32788
rect 51660 33234 51716 33246
rect 51660 33182 51662 33234
rect 51714 33182 51716 33234
rect 51660 32788 51716 33182
rect 51212 32562 51268 32732
rect 51660 32722 51716 32732
rect 51772 32674 51828 33854
rect 51772 32622 51774 32674
rect 51826 32622 51828 32674
rect 51772 32610 51828 32622
rect 51884 33460 51940 36652
rect 51996 36372 52052 37774
rect 52332 37604 52388 38670
rect 52444 38612 52500 38622
rect 52444 38518 52500 38556
rect 52332 37538 52388 37548
rect 52220 37380 52276 37390
rect 52220 37286 52276 37324
rect 52220 36932 52276 36942
rect 52220 36482 52276 36876
rect 52556 36708 52612 41468
rect 52668 41186 52724 41198
rect 52668 41134 52670 41186
rect 52722 41134 52724 41186
rect 52668 40404 52724 41134
rect 52892 41188 52948 41806
rect 53004 41858 53060 41870
rect 53004 41806 53006 41858
rect 53058 41806 53060 41858
rect 53004 41412 53060 41806
rect 53564 41858 53620 43036
rect 53564 41806 53566 41858
rect 53618 41806 53620 41858
rect 53564 41636 53620 41806
rect 53564 41570 53620 41580
rect 53676 42530 53732 43148
rect 54012 43092 54068 45836
rect 54124 46340 54180 46350
rect 54124 45890 54180 46284
rect 54124 45838 54126 45890
rect 54178 45838 54180 45890
rect 54124 45332 54180 45838
rect 54236 45444 54292 46620
rect 54460 46562 54516 46574
rect 54460 46510 54462 46562
rect 54514 46510 54516 46562
rect 54348 46450 54404 46462
rect 54348 46398 54350 46450
rect 54402 46398 54404 46450
rect 54348 45890 54404 46398
rect 54460 46228 54516 46510
rect 54460 46162 54516 46172
rect 54796 46004 54852 46956
rect 54908 46562 54964 46574
rect 54908 46510 54910 46562
rect 54962 46510 54964 46562
rect 54908 46340 54964 46510
rect 54908 46274 54964 46284
rect 54908 46004 54964 46014
rect 54796 45948 54908 46004
rect 54348 45838 54350 45890
rect 54402 45838 54404 45890
rect 54348 45826 54404 45838
rect 54908 45890 54964 45948
rect 54908 45838 54910 45890
rect 54962 45838 54964 45890
rect 54908 45826 54964 45838
rect 54460 45780 54516 45790
rect 54460 45666 54516 45724
rect 54460 45614 54462 45666
rect 54514 45614 54516 45666
rect 54460 45602 54516 45614
rect 55020 45444 55076 50318
rect 55244 49812 55300 50540
rect 55244 49718 55300 49756
rect 56140 50484 56196 50494
rect 55468 47346 55524 47358
rect 55468 47294 55470 47346
rect 55522 47294 55524 47346
rect 55468 47124 55524 47294
rect 55468 47058 55524 47068
rect 55356 46676 55412 46686
rect 55356 46582 55412 46620
rect 55692 45780 55748 45790
rect 55692 45686 55748 45724
rect 54236 45388 54628 45444
rect 54124 45276 54516 45332
rect 54124 45108 54180 45118
rect 54124 45014 54180 45052
rect 54348 44884 54404 44894
rect 54348 44790 54404 44828
rect 54348 44098 54404 44110
rect 54348 44046 54350 44098
rect 54402 44046 54404 44098
rect 54348 43652 54404 44046
rect 54348 43586 54404 43596
rect 54460 43204 54516 45276
rect 54572 44996 54628 45388
rect 54908 45388 55076 45444
rect 55692 45556 55748 45566
rect 54684 45108 54740 45118
rect 54684 44996 54740 45052
rect 54572 44994 54740 44996
rect 54572 44942 54686 44994
rect 54738 44942 54740 44994
rect 54572 44940 54740 44942
rect 54684 44930 54740 44940
rect 54796 44324 54852 44334
rect 54908 44324 54964 45388
rect 55580 45220 55636 45230
rect 55580 45126 55636 45164
rect 55132 45108 55188 45118
rect 55356 45108 55412 45118
rect 55188 45106 55412 45108
rect 55188 45054 55358 45106
rect 55410 45054 55412 45106
rect 55188 45052 55412 45054
rect 55132 45042 55188 45052
rect 55356 45042 55412 45052
rect 55020 44996 55076 45006
rect 55020 44902 55076 44940
rect 55580 44548 55636 44558
rect 55692 44548 55748 45500
rect 55580 44546 55748 44548
rect 55580 44494 55582 44546
rect 55634 44494 55748 44546
rect 55580 44492 55748 44494
rect 55580 44482 55636 44492
rect 54796 44322 54964 44324
rect 54796 44270 54798 44322
rect 54850 44270 54964 44322
rect 54796 44268 54964 44270
rect 54796 44258 54852 44268
rect 54908 43428 54964 44268
rect 55356 44322 55412 44334
rect 55356 44270 55358 44322
rect 55410 44270 55412 44322
rect 55020 44212 55076 44222
rect 55020 44118 55076 44156
rect 54908 43362 54964 43372
rect 55356 44100 55412 44270
rect 54460 43138 54516 43148
rect 53676 42478 53678 42530
rect 53730 42478 53732 42530
rect 53004 41356 53508 41412
rect 53452 41298 53508 41356
rect 53452 41246 53454 41298
rect 53506 41246 53508 41298
rect 53452 41234 53508 41246
rect 52892 41132 53396 41188
rect 52668 40338 52724 40348
rect 53340 41076 53396 41132
rect 53676 41076 53732 42478
rect 53900 43036 54068 43092
rect 53900 41748 53956 43036
rect 54908 42754 54964 42766
rect 54908 42702 54910 42754
rect 54962 42702 54964 42754
rect 54124 42530 54180 42542
rect 54572 42532 54628 42542
rect 54908 42532 54964 42702
rect 55356 42756 55412 44044
rect 55804 44212 55860 44222
rect 55468 43540 55524 43550
rect 55468 43446 55524 43484
rect 55804 43538 55860 44156
rect 55916 44098 55972 44110
rect 55916 44046 55918 44098
rect 55970 44046 55972 44098
rect 55916 43652 55972 44046
rect 56028 43652 56084 43662
rect 55916 43596 56028 43652
rect 56028 43558 56084 43596
rect 55804 43486 55806 43538
rect 55858 43486 55860 43538
rect 55804 43474 55860 43486
rect 55916 43426 55972 43438
rect 55916 43374 55918 43426
rect 55970 43374 55972 43426
rect 55692 43316 55748 43326
rect 55356 42690 55412 42700
rect 55580 42980 55636 42990
rect 54124 42478 54126 42530
rect 54178 42478 54180 42530
rect 53900 41682 53956 41692
rect 54012 41858 54068 41870
rect 54012 41806 54014 41858
rect 54066 41806 54068 41858
rect 54012 41746 54068 41806
rect 54012 41694 54014 41746
rect 54066 41694 54068 41746
rect 54012 41682 54068 41694
rect 53340 41020 53732 41076
rect 52892 40292 52948 40302
rect 52892 39506 52948 40236
rect 53116 39620 53172 39630
rect 52892 39454 52894 39506
rect 52946 39454 52948 39506
rect 52892 39442 52948 39454
rect 53004 39508 53060 39518
rect 53004 39414 53060 39452
rect 53116 39506 53172 39564
rect 53116 39454 53118 39506
rect 53170 39454 53172 39506
rect 53116 39442 53172 39454
rect 52668 39396 52724 39406
rect 52668 39302 52724 39340
rect 52780 39394 52836 39406
rect 52780 39342 52782 39394
rect 52834 39342 52836 39394
rect 52780 39172 52836 39342
rect 53228 39396 53284 39406
rect 52780 39116 53172 39172
rect 53116 38946 53172 39116
rect 53116 38894 53118 38946
rect 53170 38894 53172 38946
rect 53116 38882 53172 38894
rect 53228 38946 53284 39340
rect 53228 38894 53230 38946
rect 53282 38894 53284 38946
rect 53228 38882 53284 38894
rect 52892 38836 52948 38846
rect 52892 38742 52948 38780
rect 53116 38612 53172 38622
rect 53340 38612 53396 41020
rect 54124 40516 54180 42478
rect 54460 42530 54964 42532
rect 54460 42478 54574 42530
rect 54626 42478 54964 42530
rect 54460 42476 54964 42478
rect 54460 41858 54516 42476
rect 54572 42466 54628 42476
rect 55580 42196 55636 42924
rect 55692 42866 55748 43260
rect 55692 42814 55694 42866
rect 55746 42814 55748 42866
rect 55692 42802 55748 42814
rect 54460 41806 54462 41858
rect 54514 41806 54516 41858
rect 53788 40404 53844 40414
rect 53676 40292 53732 40302
rect 53676 40198 53732 40236
rect 53788 39956 53844 40348
rect 54012 40404 54068 40414
rect 54124 40404 54180 40460
rect 54012 40402 54180 40404
rect 54012 40350 54014 40402
rect 54066 40350 54180 40402
rect 54012 40348 54180 40350
rect 54236 41746 54292 41758
rect 54236 41694 54238 41746
rect 54290 41694 54292 41746
rect 54012 40338 54068 40348
rect 53900 40290 53956 40302
rect 53900 40238 53902 40290
rect 53954 40238 53956 40290
rect 53900 40180 53956 40238
rect 53900 40114 53956 40124
rect 53676 39900 53844 39956
rect 53676 39058 53732 39900
rect 54124 39732 54180 39742
rect 54236 39732 54292 41694
rect 54348 40404 54404 40414
rect 54348 40310 54404 40348
rect 54180 39676 54292 39732
rect 54124 39638 54180 39676
rect 54348 39508 54404 39518
rect 54348 39414 54404 39452
rect 53788 39396 53844 39406
rect 53788 39302 53844 39340
rect 53676 39006 53678 39058
rect 53730 39006 53732 39058
rect 53676 38994 53732 39006
rect 54124 38724 54180 38762
rect 54124 38658 54180 38668
rect 53172 38556 53284 38612
rect 53116 38546 53172 38556
rect 53116 38052 53172 38062
rect 53116 37958 53172 37996
rect 52668 37938 52724 37950
rect 52668 37886 52670 37938
rect 52722 37886 52724 37938
rect 52668 37492 52724 37886
rect 52892 37940 52948 37950
rect 52892 37846 52948 37884
rect 52668 37426 52724 37436
rect 52892 37716 52948 37726
rect 52556 36642 52612 36652
rect 52220 36430 52222 36482
rect 52274 36430 52276 36482
rect 52220 36418 52276 36430
rect 52668 36596 52724 36606
rect 52668 36484 52724 36540
rect 52668 36482 52836 36484
rect 52668 36430 52670 36482
rect 52722 36430 52836 36482
rect 52668 36428 52836 36430
rect 52668 36418 52724 36428
rect 51996 35700 52052 36316
rect 52668 36260 52724 36270
rect 52556 36258 52724 36260
rect 52556 36206 52670 36258
rect 52722 36206 52724 36258
rect 52556 36204 52724 36206
rect 52108 35700 52164 35710
rect 51996 35698 52164 35700
rect 51996 35646 52110 35698
rect 52162 35646 52164 35698
rect 51996 35644 52164 35646
rect 52108 35634 52164 35644
rect 52220 35700 52276 35710
rect 52556 35700 52612 36204
rect 52668 36194 52724 36204
rect 52220 35698 52612 35700
rect 52220 35646 52222 35698
rect 52274 35646 52612 35698
rect 52220 35644 52612 35646
rect 52220 35634 52276 35644
rect 52444 35476 52500 35486
rect 52444 35382 52500 35420
rect 52556 35474 52612 35486
rect 52556 35422 52558 35474
rect 52610 35422 52612 35474
rect 52108 35140 52164 35150
rect 52108 35026 52164 35084
rect 52108 34974 52110 35026
rect 52162 34974 52164 35026
rect 52108 34244 52164 34974
rect 52108 34178 52164 34188
rect 52220 34916 52276 34926
rect 52556 34916 52612 35422
rect 52668 35140 52724 35150
rect 52780 35140 52836 36428
rect 52892 35476 52948 37660
rect 53228 37380 53284 38556
rect 53340 38162 53396 38556
rect 53340 38110 53342 38162
rect 53394 38110 53396 38162
rect 53340 38098 53396 38110
rect 54012 38610 54068 38622
rect 54012 38558 54014 38610
rect 54066 38558 54068 38610
rect 53564 38052 53620 38062
rect 53564 37958 53620 37996
rect 54012 38050 54068 38558
rect 54012 37998 54014 38050
rect 54066 37998 54068 38050
rect 54012 37986 54068 37998
rect 54460 38610 54516 41806
rect 54908 41858 54964 41870
rect 54908 41806 54910 41858
rect 54962 41806 54964 41858
rect 54908 41748 54964 41806
rect 54908 41682 54964 41692
rect 55020 41300 55076 41310
rect 54684 40514 54740 40526
rect 54684 40462 54686 40514
rect 54738 40462 54740 40514
rect 54684 39732 54740 40462
rect 55020 40514 55076 41244
rect 55580 41298 55636 42140
rect 55804 42196 55860 42206
rect 55916 42196 55972 43374
rect 55804 42194 55972 42196
rect 55804 42142 55806 42194
rect 55858 42142 55972 42194
rect 55804 42140 55972 42142
rect 55804 42130 55860 42140
rect 56028 42084 56084 42094
rect 56028 41972 56084 42028
rect 55916 41970 56084 41972
rect 55916 41918 56030 41970
rect 56082 41918 56084 41970
rect 55916 41916 56084 41918
rect 55692 41860 55748 41870
rect 55692 41766 55748 41804
rect 55580 41246 55582 41298
rect 55634 41246 55636 41298
rect 55580 41234 55636 41246
rect 55692 41636 55748 41646
rect 55020 40462 55022 40514
rect 55074 40462 55076 40514
rect 55020 40450 55076 40462
rect 55244 40516 55300 40526
rect 55692 40516 55748 41580
rect 55300 40460 55412 40516
rect 55244 40450 55300 40460
rect 55356 40180 55412 40460
rect 55692 40402 55748 40460
rect 55692 40350 55694 40402
rect 55746 40350 55748 40402
rect 55692 40338 55748 40350
rect 55916 40402 55972 41916
rect 56028 41906 56084 41916
rect 55916 40350 55918 40402
rect 55970 40350 55972 40402
rect 55916 40338 55972 40350
rect 55356 40124 55524 40180
rect 54684 39666 54740 39676
rect 55020 39618 55076 39630
rect 55020 39566 55022 39618
rect 55074 39566 55076 39618
rect 55020 39058 55076 39566
rect 55020 39006 55022 39058
rect 55074 39006 55076 39058
rect 55020 38948 55076 39006
rect 54460 38558 54462 38610
rect 54514 38558 54516 38610
rect 53676 37940 53732 37950
rect 53676 37826 53732 37884
rect 53676 37774 53678 37826
rect 53730 37774 53732 37826
rect 53676 37762 53732 37774
rect 53004 36484 53060 36494
rect 53004 36390 53060 36428
rect 53228 36482 53284 37324
rect 53452 37604 53508 37614
rect 53452 37266 53508 37548
rect 54124 37380 54180 37390
rect 54124 37286 54180 37324
rect 53452 37214 53454 37266
rect 53506 37214 53508 37266
rect 53452 37202 53508 37214
rect 53788 37268 53844 37278
rect 53788 37174 53844 37212
rect 54236 37268 54292 37278
rect 54236 37174 54292 37212
rect 54348 37266 54404 37278
rect 54348 37214 54350 37266
rect 54402 37214 54404 37266
rect 53228 36430 53230 36482
rect 53282 36430 53284 36482
rect 53228 36418 53284 36430
rect 53452 36932 53508 36942
rect 53452 36482 53508 36876
rect 54348 36932 54404 37214
rect 54348 36866 54404 36876
rect 53452 36430 53454 36482
rect 53506 36430 53508 36482
rect 53452 36418 53508 36430
rect 54236 36708 54292 36718
rect 53788 36370 53844 36382
rect 53788 36318 53790 36370
rect 53842 36318 53844 36370
rect 53788 35924 53844 36318
rect 54012 36260 54068 36270
rect 54012 36166 54068 36204
rect 53788 35858 53844 35868
rect 53228 35812 53284 35822
rect 53228 35718 53284 35756
rect 54236 35812 54292 36652
rect 54348 36484 54404 36494
rect 54348 36390 54404 36428
rect 53340 35698 53396 35710
rect 53340 35646 53342 35698
rect 53394 35646 53396 35698
rect 52892 35410 52948 35420
rect 53004 35588 53060 35598
rect 52668 35138 52836 35140
rect 52668 35086 52670 35138
rect 52722 35086 52836 35138
rect 52668 35084 52836 35086
rect 53004 35364 53060 35532
rect 53004 35138 53060 35308
rect 53004 35086 53006 35138
rect 53058 35086 53060 35138
rect 52668 35074 52724 35084
rect 53004 35074 53060 35086
rect 53340 35028 53396 35646
rect 53564 35700 53620 35710
rect 53788 35700 53844 35710
rect 53564 35606 53620 35644
rect 53676 35698 53844 35700
rect 53676 35646 53790 35698
rect 53842 35646 53844 35698
rect 53676 35644 53844 35646
rect 53676 35140 53732 35644
rect 53788 35634 53844 35644
rect 54236 35698 54292 35756
rect 54236 35646 54238 35698
rect 54290 35646 54292 35698
rect 54236 35634 54292 35646
rect 54124 35588 54180 35598
rect 53900 35532 54124 35588
rect 53788 35476 53844 35486
rect 53788 35382 53844 35420
rect 53676 35074 53732 35084
rect 53900 35138 53956 35532
rect 54124 35522 54180 35532
rect 53900 35086 53902 35138
rect 53954 35086 53956 35138
rect 53900 35074 53956 35086
rect 53340 34962 53396 34972
rect 53228 34916 53284 34926
rect 52556 34860 53172 34916
rect 52220 34132 52276 34860
rect 53116 34692 53172 34860
rect 53228 34822 53284 34860
rect 53564 34914 53620 34926
rect 54460 34916 54516 38558
rect 54572 38722 54628 38734
rect 54572 38670 54574 38722
rect 54626 38670 54628 38722
rect 54572 37156 54628 38670
rect 55020 38610 55076 38892
rect 55020 38558 55022 38610
rect 55074 38558 55076 38610
rect 55020 38546 55076 38558
rect 55356 39508 55412 39518
rect 55356 39060 55412 39452
rect 54684 37940 54740 37950
rect 54684 37846 54740 37884
rect 54908 37380 54964 37390
rect 54908 37286 54964 37324
rect 54684 37268 54740 37278
rect 54684 37174 54740 37212
rect 55244 37266 55300 37278
rect 55244 37214 55246 37266
rect 55298 37214 55300 37266
rect 54572 37090 54628 37100
rect 55132 37154 55188 37166
rect 55132 37102 55134 37154
rect 55186 37102 55188 37154
rect 54908 37044 54964 37054
rect 54908 36482 54964 36988
rect 54908 36430 54910 36482
rect 54962 36430 54964 36482
rect 54908 36418 54964 36430
rect 54908 36036 54964 36046
rect 54684 35924 54740 35934
rect 53564 34862 53566 34914
rect 53618 34862 53620 34914
rect 53564 34692 53620 34862
rect 54012 34914 54516 34916
rect 54012 34862 54462 34914
rect 54514 34862 54516 34914
rect 54012 34860 54516 34862
rect 53116 34636 53620 34692
rect 53788 34690 53844 34702
rect 53788 34638 53790 34690
rect 53842 34638 53844 34690
rect 53788 34244 53844 34638
rect 53900 34244 53956 34254
rect 53788 34242 53956 34244
rect 53788 34190 53902 34242
rect 53954 34190 53956 34242
rect 53788 34188 53956 34190
rect 53900 34178 53956 34188
rect 52220 34038 52276 34076
rect 52780 34132 52836 34142
rect 52780 34038 52836 34076
rect 53228 34132 53284 34142
rect 53228 34038 53284 34076
rect 54012 34132 54068 34860
rect 54460 34850 54516 34860
rect 54572 35812 54628 35822
rect 54012 33570 54068 34076
rect 54012 33518 54014 33570
rect 54066 33518 54068 33570
rect 51212 32510 51214 32562
rect 51266 32510 51268 32562
rect 51212 32498 51268 32510
rect 51548 32562 51604 32574
rect 51548 32510 51550 32562
rect 51602 32510 51604 32562
rect 51324 32338 51380 32350
rect 51324 32286 51326 32338
rect 51378 32286 51380 32338
rect 51324 31892 51380 32286
rect 51548 32340 51604 32510
rect 51660 32564 51716 32574
rect 51660 32470 51716 32508
rect 51884 32340 51940 33404
rect 52780 33460 52836 33470
rect 52780 33366 52836 33404
rect 54012 33458 54068 33518
rect 54012 33406 54014 33458
rect 54066 33406 54068 33458
rect 54012 33394 54068 33406
rect 54572 33458 54628 35756
rect 54684 35698 54740 35868
rect 54684 35646 54686 35698
rect 54738 35646 54740 35698
rect 54684 34916 54740 35646
rect 54908 35922 54964 35980
rect 54908 35870 54910 35922
rect 54962 35870 54964 35922
rect 54796 35588 54852 35598
rect 54796 35494 54852 35532
rect 54684 34020 54740 34860
rect 54684 33954 54740 33964
rect 54572 33406 54574 33458
rect 54626 33406 54628 33458
rect 54572 33394 54628 33406
rect 54908 33458 54964 35870
rect 55132 35476 55188 37102
rect 55244 36932 55300 37214
rect 55244 35812 55300 36876
rect 55356 36370 55412 39004
rect 55468 39058 55524 40124
rect 55804 39732 55860 39742
rect 55804 39638 55860 39676
rect 55468 39006 55470 39058
rect 55522 39006 55524 39058
rect 55468 37716 55524 39006
rect 55916 38948 55972 38958
rect 55916 38854 55972 38892
rect 56140 38668 56196 50428
rect 56700 49924 56756 49934
rect 56588 49922 56756 49924
rect 56588 49870 56702 49922
rect 56754 49870 56756 49922
rect 56588 49868 56756 49870
rect 56476 49812 56532 49822
rect 56476 49718 56532 49756
rect 56588 48580 56644 49868
rect 56700 49858 56756 49868
rect 56812 49810 56868 49822
rect 56812 49758 56814 49810
rect 56866 49758 56868 49810
rect 56700 49140 56756 49150
rect 56812 49140 56868 49758
rect 57484 49140 57540 49150
rect 56700 49138 57092 49140
rect 56700 49086 56702 49138
rect 56754 49086 57092 49138
rect 56700 49084 57092 49086
rect 56700 49074 56756 49084
rect 57036 49026 57092 49084
rect 57484 49046 57540 49084
rect 57036 48974 57038 49026
rect 57090 48974 57092 49026
rect 57036 48962 57092 48974
rect 56588 48524 57092 48580
rect 57036 48244 57092 48524
rect 57036 48242 57652 48244
rect 57036 48190 57038 48242
rect 57090 48190 57652 48242
rect 57036 48188 57652 48190
rect 57036 48178 57092 48188
rect 56588 48132 56644 48142
rect 56588 48038 56644 48076
rect 57596 47570 57652 48188
rect 57596 47518 57598 47570
rect 57650 47518 57652 47570
rect 57596 47506 57652 47518
rect 57708 46674 57764 46686
rect 57708 46622 57710 46674
rect 57762 46622 57764 46674
rect 57148 46562 57204 46574
rect 57148 46510 57150 46562
rect 57202 46510 57204 46562
rect 57148 46228 57204 46510
rect 56588 45220 56644 45230
rect 56588 45126 56644 45164
rect 57148 45220 57204 46172
rect 57708 46004 57764 46622
rect 57820 46004 57876 46014
rect 57708 46002 57876 46004
rect 57708 45950 57822 46002
rect 57874 45950 57876 46002
rect 57708 45948 57876 45950
rect 57820 45556 57876 45948
rect 57820 45490 57876 45500
rect 57148 45164 57540 45220
rect 57148 45106 57204 45164
rect 57148 45054 57150 45106
rect 57202 45054 57204 45106
rect 57148 45042 57204 45054
rect 57372 44994 57428 45006
rect 57372 44942 57374 44994
rect 57426 44942 57428 44994
rect 57260 44436 57316 44446
rect 57036 44434 57316 44436
rect 57036 44382 57262 44434
rect 57314 44382 57316 44434
rect 57036 44380 57316 44382
rect 56364 44324 56420 44334
rect 56364 44230 56420 44268
rect 56812 44324 56868 44334
rect 57036 44324 57092 44380
rect 57260 44370 57316 44380
rect 56812 44322 57092 44324
rect 56812 44270 56814 44322
rect 56866 44270 57092 44322
rect 56812 44268 57092 44270
rect 56812 44258 56868 44268
rect 56252 44210 56308 44222
rect 56252 44158 56254 44210
rect 56306 44158 56308 44210
rect 56252 43652 56308 44158
rect 56588 44212 56644 44222
rect 56588 44118 56644 44156
rect 57148 44212 57204 44222
rect 57372 44212 57428 44942
rect 57484 44322 57540 45164
rect 57484 44270 57486 44322
rect 57538 44270 57540 44322
rect 57484 44258 57540 44270
rect 57596 44322 57652 44334
rect 57596 44270 57598 44322
rect 57650 44270 57652 44322
rect 57204 44156 57428 44212
rect 57148 44118 57204 44156
rect 57596 44100 57652 44270
rect 57652 44044 57876 44100
rect 57596 44034 57652 44044
rect 56252 43586 56308 43596
rect 57036 43652 57092 43662
rect 57036 43558 57092 43596
rect 56588 43540 56644 43550
rect 56588 43446 56644 43484
rect 56812 43538 56868 43550
rect 56812 43486 56814 43538
rect 56866 43486 56868 43538
rect 56812 43428 56868 43486
rect 56812 43362 56868 43372
rect 57372 43316 57428 43326
rect 57036 43314 57428 43316
rect 57036 43262 57374 43314
rect 57426 43262 57428 43314
rect 57036 43260 57428 43262
rect 56700 42196 56756 42206
rect 56588 42084 56644 42094
rect 56588 40402 56644 42028
rect 56700 42082 56756 42140
rect 56700 42030 56702 42082
rect 56754 42030 56756 42082
rect 56700 42018 56756 42030
rect 57036 42084 57092 43260
rect 57372 43250 57428 43260
rect 57820 42866 57876 44044
rect 57820 42814 57822 42866
rect 57874 42814 57876 42866
rect 57820 42802 57876 42814
rect 57036 41970 57092 42028
rect 57036 41918 57038 41970
rect 57090 41918 57092 41970
rect 57036 41906 57092 41918
rect 57260 41858 57316 41870
rect 57260 41806 57262 41858
rect 57314 41806 57316 41858
rect 57260 41298 57316 41806
rect 57260 41246 57262 41298
rect 57314 41246 57316 41298
rect 56700 41076 56756 41086
rect 56700 40982 56756 41020
rect 56588 40350 56590 40402
rect 56642 40350 56644 40402
rect 56588 40338 56644 40350
rect 56924 40626 56980 40638
rect 56924 40574 56926 40626
rect 56978 40574 56980 40626
rect 56700 38834 56756 38846
rect 56700 38782 56702 38834
rect 56754 38782 56756 38834
rect 55916 38612 56196 38668
rect 56588 38722 56644 38734
rect 56588 38670 56590 38722
rect 56642 38670 56644 38722
rect 55468 37650 55524 37660
rect 55804 37716 55860 37726
rect 55692 37492 55748 37502
rect 55692 37398 55748 37436
rect 55804 37490 55860 37660
rect 55804 37438 55806 37490
rect 55858 37438 55860 37490
rect 55804 37426 55860 37438
rect 55580 37380 55636 37390
rect 55580 37286 55636 37324
rect 55356 36318 55358 36370
rect 55410 36318 55412 36370
rect 55356 36306 55412 36318
rect 55804 37156 55860 37166
rect 55356 35812 55412 35822
rect 55244 35756 55356 35812
rect 55356 35746 55412 35756
rect 55580 35700 55636 35710
rect 55580 35606 55636 35644
rect 55804 35698 55860 37100
rect 55804 35646 55806 35698
rect 55858 35646 55860 35698
rect 55804 35634 55860 35646
rect 55132 35410 55188 35420
rect 55468 35474 55524 35486
rect 55468 35422 55470 35474
rect 55522 35422 55524 35474
rect 55468 35364 55524 35422
rect 55468 35298 55524 35308
rect 55132 35028 55188 35038
rect 55132 34934 55188 34972
rect 54908 33406 54910 33458
rect 54962 33406 54964 33458
rect 54908 33394 54964 33406
rect 55020 33570 55076 33582
rect 55020 33518 55022 33570
rect 55074 33518 55076 33570
rect 52108 32788 52164 32798
rect 52108 32452 52164 32732
rect 54236 32564 54292 32574
rect 54236 32470 54292 32508
rect 55020 32562 55076 33518
rect 55020 32510 55022 32562
rect 55074 32510 55076 32562
rect 55020 32498 55076 32510
rect 52108 32358 52164 32396
rect 52780 32452 52836 32462
rect 51548 32284 51940 32340
rect 51324 31826 51380 31836
rect 51996 32228 52052 32238
rect 51212 31780 51268 31790
rect 51212 31686 51268 31724
rect 51772 31780 51828 31790
rect 51772 31686 51828 31724
rect 51548 31668 51604 31678
rect 51548 31574 51604 31612
rect 50556 31388 50820 31398
rect 50876 31388 51604 31444
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50428 31054 50430 31106
rect 50482 31054 50484 31106
rect 50428 31042 50484 31054
rect 50540 31218 50596 31230
rect 50540 31166 50542 31218
rect 50594 31166 50596 31218
rect 50092 30942 50094 30994
rect 50146 30942 50148 30994
rect 50092 30930 50148 30942
rect 49196 30818 49252 30828
rect 49756 30884 49812 30894
rect 49756 30790 49812 30828
rect 49980 30884 50036 30894
rect 45836 30146 45892 30156
rect 48860 30212 48916 30222
rect 48860 30118 48916 30156
rect 49308 30212 49364 30222
rect 49308 30118 49364 30156
rect 49980 30210 50036 30828
rect 50540 30884 50596 31166
rect 50876 31220 50932 31230
rect 50652 30996 50708 31006
rect 50652 30902 50708 30940
rect 50876 30994 50932 31164
rect 50876 30942 50878 30994
rect 50930 30942 50932 30994
rect 50876 30930 50932 30942
rect 51100 30996 51156 31006
rect 51436 30996 51492 31006
rect 51100 30994 51492 30996
rect 51100 30942 51102 30994
rect 51154 30942 51438 30994
rect 51490 30942 51492 30994
rect 51100 30940 51492 30942
rect 51100 30930 51156 30940
rect 51436 30930 51492 30940
rect 50540 30818 50596 30828
rect 51548 30882 51604 31388
rect 51996 31220 52052 32172
rect 52668 31892 52724 31902
rect 52668 31798 52724 31836
rect 52780 31890 52836 32396
rect 55916 32228 55972 38612
rect 56588 38052 56644 38670
rect 56700 38668 56756 38782
rect 56700 38612 56868 38668
rect 56140 37604 56196 37614
rect 56028 37156 56084 37166
rect 56028 35698 56084 37100
rect 56140 36594 56196 37548
rect 56140 36542 56142 36594
rect 56194 36542 56196 36594
rect 56140 36530 56196 36542
rect 56588 36482 56644 37996
rect 56812 38162 56868 38612
rect 56812 38110 56814 38162
rect 56866 38110 56868 38162
rect 56812 37828 56868 38110
rect 56812 37044 56868 37772
rect 56812 36978 56868 36988
rect 56588 36430 56590 36482
rect 56642 36430 56644 36482
rect 56588 36418 56644 36430
rect 56924 36484 56980 40574
rect 57036 40514 57092 40526
rect 57036 40462 57038 40514
rect 57090 40462 57092 40514
rect 57036 39060 57092 40462
rect 57148 39060 57204 39070
rect 57036 39004 57148 39060
rect 57148 38668 57204 39004
rect 57260 38836 57316 41246
rect 57596 41188 57652 41198
rect 57596 41186 57988 41188
rect 57596 41134 57598 41186
rect 57650 41134 57988 41186
rect 57596 41132 57988 41134
rect 57596 41122 57652 41132
rect 57372 40516 57428 40526
rect 57372 40422 57428 40460
rect 57932 39732 57988 41132
rect 57484 39730 57988 39732
rect 57484 39678 57934 39730
rect 57986 39678 57988 39730
rect 57484 39676 57988 39678
rect 57484 39058 57540 39676
rect 57932 39666 57988 39676
rect 57484 39006 57486 39058
rect 57538 39006 57540 39058
rect 57484 38994 57540 39006
rect 57260 38780 57540 38836
rect 57148 38612 57428 38668
rect 57372 38050 57428 38612
rect 57372 37998 57374 38050
rect 57426 37998 57428 38050
rect 57372 37986 57428 37998
rect 57036 37828 57092 37838
rect 57260 37828 57316 37838
rect 57036 37826 57204 37828
rect 57036 37774 57038 37826
rect 57090 37774 57204 37826
rect 57036 37772 57204 37774
rect 57036 37762 57092 37772
rect 57148 37156 57204 37772
rect 57260 37734 57316 37772
rect 57260 37268 57316 37278
rect 57484 37268 57540 38780
rect 57316 37212 57540 37268
rect 57260 37174 57316 37212
rect 57148 37062 57204 37100
rect 57596 37154 57652 37166
rect 57596 37102 57598 37154
rect 57650 37102 57652 37154
rect 57036 36484 57092 36494
rect 56924 36482 57092 36484
rect 56924 36430 57038 36482
rect 57090 36430 57092 36482
rect 56924 36428 57092 36430
rect 57036 36418 57092 36428
rect 57260 36484 57316 36494
rect 57596 36484 57652 37102
rect 56588 35812 56644 35822
rect 56588 35718 56644 35756
rect 56028 35646 56030 35698
rect 56082 35646 56084 35698
rect 56028 35634 56084 35646
rect 57036 35700 57092 35710
rect 57036 35606 57092 35644
rect 57260 35588 57316 36428
rect 57484 36482 57652 36484
rect 57484 36430 57598 36482
rect 57650 36430 57652 36482
rect 57484 36428 57652 36430
rect 57484 35698 57540 36428
rect 57596 36418 57652 36428
rect 57484 35646 57486 35698
rect 57538 35646 57540 35698
rect 57484 35634 57540 35646
rect 57932 35700 57988 35710
rect 57932 35606 57988 35644
rect 57260 35026 57316 35532
rect 58044 35588 58100 35598
rect 58044 35494 58100 35532
rect 57260 34974 57262 35026
rect 57314 34974 57316 35026
rect 57260 34962 57316 34974
rect 56028 34020 56084 34030
rect 56028 33926 56084 33964
rect 55916 32162 55972 32172
rect 52780 31838 52782 31890
rect 52834 31838 52836 31890
rect 52780 31826 52836 31838
rect 52108 31556 52164 31566
rect 52108 31462 52164 31500
rect 51996 31126 52052 31164
rect 51548 30830 51550 30882
rect 51602 30830 51604 30882
rect 51548 30324 51604 30830
rect 52108 30324 52164 30334
rect 51548 30322 52164 30324
rect 51548 30270 52110 30322
rect 52162 30270 52164 30322
rect 51548 30268 52164 30270
rect 52108 30258 52164 30268
rect 49980 30158 49982 30210
rect 50034 30158 50036 30210
rect 49980 30146 50036 30158
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 44604 29428 44660 29438
rect 44044 29426 44660 29428
rect 44044 29374 44046 29426
rect 44098 29374 44606 29426
rect 44658 29374 44660 29426
rect 44044 29372 44660 29374
rect 42140 28868 42196 28878
rect 42140 28774 42196 28812
rect 42812 28868 42868 28878
rect 41692 27918 41694 27970
rect 41746 27918 41748 27970
rect 41692 27906 41748 27918
rect 41804 28642 41860 28654
rect 41804 28590 41806 28642
rect 41858 28590 41860 28642
rect 41804 27972 41860 28590
rect 41916 28644 41972 28654
rect 41972 28588 42084 28644
rect 41916 28550 41972 28588
rect 42028 28308 42084 28588
rect 42252 28532 42308 28542
rect 42252 28438 42308 28476
rect 42028 28252 42308 28308
rect 41804 27906 41860 27916
rect 40796 27806 40798 27858
rect 40850 27806 40852 27858
rect 40796 27794 40852 27806
rect 41916 27858 41972 27870
rect 41916 27806 41918 27858
rect 41970 27806 41972 27858
rect 40236 27682 40292 27692
rect 40684 27748 40740 27758
rect 39676 26462 39678 26514
rect 39730 26462 39732 26514
rect 37324 26290 37380 26460
rect 39676 26450 39732 26462
rect 39788 27186 40068 27188
rect 39788 27134 39902 27186
rect 39954 27134 40068 27186
rect 39788 27132 40068 27134
rect 40460 27188 40516 27198
rect 37324 26238 37326 26290
rect 37378 26238 37380 26290
rect 37100 26226 37156 26236
rect 37324 26226 37380 26238
rect 39564 26292 39620 26302
rect 39788 26292 39844 27132
rect 39900 27122 39956 27132
rect 39900 26516 39956 26526
rect 39900 26422 39956 26460
rect 40460 26514 40516 27132
rect 40684 27074 40740 27692
rect 41468 27746 41524 27758
rect 41468 27694 41470 27746
rect 41522 27694 41524 27746
rect 41468 27300 41524 27694
rect 41916 27748 41972 27806
rect 41916 27692 42196 27748
rect 41468 27298 41860 27300
rect 41468 27246 41470 27298
rect 41522 27246 41860 27298
rect 41468 27244 41860 27246
rect 40684 27022 40686 27074
rect 40738 27022 40740 27074
rect 40684 27010 40740 27022
rect 40796 27186 40852 27198
rect 40796 27134 40798 27186
rect 40850 27134 40852 27186
rect 40796 26516 40852 27134
rect 40460 26462 40462 26514
rect 40514 26462 40516 26514
rect 40460 26450 40516 26462
rect 40684 26460 40852 26516
rect 40908 27188 40964 27198
rect 39564 26290 39844 26292
rect 39564 26238 39566 26290
rect 39618 26238 39844 26290
rect 39564 26236 39844 26238
rect 40684 26292 40740 26460
rect 39564 26226 39620 26236
rect 36540 26012 36932 26068
rect 36540 25618 36596 26012
rect 36540 25566 36542 25618
rect 36594 25566 36596 25618
rect 36540 25554 36596 25566
rect 39452 25620 39508 25630
rect 39452 25526 39508 25564
rect 40684 25620 40740 26236
rect 40908 26290 40964 27132
rect 40908 26238 40910 26290
rect 40962 26238 40964 26290
rect 40908 26226 40964 26238
rect 41132 27076 41188 27086
rect 41132 26516 41188 27020
rect 41244 26964 41300 26974
rect 41244 26516 41300 26908
rect 41356 26516 41412 26526
rect 41244 26514 41412 26516
rect 41244 26462 41358 26514
rect 41410 26462 41412 26514
rect 41244 26460 41412 26462
rect 41132 26292 41188 26460
rect 41356 26450 41412 26460
rect 41468 26514 41524 27244
rect 41804 27074 41860 27244
rect 41804 27022 41806 27074
rect 41858 27022 41860 27074
rect 41804 27010 41860 27022
rect 42140 27076 42196 27692
rect 42140 26982 42196 27020
rect 42028 26962 42084 26974
rect 42028 26910 42030 26962
rect 42082 26910 42084 26962
rect 42028 26740 42084 26910
rect 41468 26462 41470 26514
rect 41522 26462 41524 26514
rect 41468 26450 41524 26462
rect 41580 26684 42084 26740
rect 41244 26292 41300 26302
rect 41132 26290 41300 26292
rect 41132 26238 41246 26290
rect 41298 26238 41300 26290
rect 41132 26236 41300 26238
rect 41244 26226 41300 26236
rect 40684 25554 40740 25564
rect 41580 25618 41636 26684
rect 42140 26516 42196 26526
rect 42252 26516 42308 28252
rect 42476 26964 42532 26974
rect 42476 26870 42532 26908
rect 42140 26514 42308 26516
rect 42140 26462 42142 26514
rect 42194 26462 42308 26514
rect 42140 26460 42308 26462
rect 42140 26450 42196 26460
rect 41804 26292 41860 26302
rect 41804 26198 41860 26236
rect 42812 25620 42868 28812
rect 44044 28868 44100 29372
rect 44604 29362 44660 29372
rect 44044 28802 44100 28812
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 41580 25566 41582 25618
rect 41634 25566 41636 25618
rect 41580 25554 41636 25566
rect 42364 25618 43428 25620
rect 42364 25566 42814 25618
rect 42866 25566 43428 25618
rect 42364 25564 43428 25566
rect 42364 25506 42420 25564
rect 42812 25554 42868 25564
rect 42364 25454 42366 25506
rect 42418 25454 42420 25506
rect 42364 25442 42420 25454
rect 36876 24948 36932 24958
rect 36092 24946 36932 24948
rect 36092 24894 36430 24946
rect 36482 24894 36878 24946
rect 36930 24894 36932 24946
rect 36092 24892 36932 24894
rect 33852 24836 33908 24846
rect 33852 24742 33908 24780
rect 34860 24612 34916 24622
rect 33852 23940 33908 23950
rect 33740 23884 33852 23940
rect 33740 23492 33796 23502
rect 33740 23266 33796 23436
rect 33740 23214 33742 23266
rect 33794 23214 33796 23266
rect 33740 23202 33796 23214
rect 33852 23044 33908 23884
rect 34860 23828 34916 24556
rect 35980 24612 36036 24622
rect 35980 24518 36036 24556
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 33628 22194 33684 22204
rect 33740 22988 33908 23044
rect 34076 23266 34132 23278
rect 34076 23214 34078 23266
rect 34130 23214 34132 23266
rect 32956 20132 33012 20636
rect 32844 19460 32900 19470
rect 32508 18510 32510 18562
rect 32562 18510 32564 18562
rect 32508 18498 32564 18510
rect 32732 19458 32900 19460
rect 32732 19406 32846 19458
rect 32898 19406 32900 19458
rect 32732 19404 32900 19406
rect 32060 17502 32062 17554
rect 32114 17502 32116 17554
rect 32060 17490 32116 17502
rect 32396 18226 32452 18238
rect 32396 18174 32398 18226
rect 32450 18174 32452 18226
rect 32172 16994 32228 17006
rect 32172 16942 32174 16994
rect 32226 16942 32228 16994
rect 32172 16212 32228 16942
rect 32172 16146 32228 16156
rect 32396 15988 32452 18174
rect 32396 15922 32452 15932
rect 32060 15874 32116 15886
rect 32060 15822 32062 15874
rect 32114 15822 32116 15874
rect 32060 15540 32116 15822
rect 32060 15474 32116 15484
rect 31388 13022 31390 13074
rect 31442 13022 31444 13074
rect 31388 13010 31444 13022
rect 31724 15092 32004 15148
rect 32732 15148 32788 19404
rect 32844 19394 32900 19404
rect 32956 19124 33012 20076
rect 33068 20020 33124 20030
rect 33068 19926 33124 19964
rect 33404 19908 33460 21756
rect 33516 21586 33572 21598
rect 33516 21534 33518 21586
rect 33570 21534 33572 21586
rect 33516 21476 33572 21534
rect 33516 21410 33572 21420
rect 33628 21140 33684 21150
rect 33740 21140 33796 22988
rect 34076 22596 34132 23214
rect 34860 23266 34916 23772
rect 34860 23214 34862 23266
rect 34914 23214 34916 23266
rect 34860 23202 34916 23214
rect 35980 24052 36036 24062
rect 36092 24052 36148 24892
rect 36428 24882 36484 24892
rect 35980 24050 36148 24052
rect 35980 23998 35982 24050
rect 36034 23998 36148 24050
rect 35980 23996 36148 23998
rect 35868 23156 35924 23166
rect 35980 23156 36036 23996
rect 36876 23940 36932 24892
rect 38220 24610 38276 24622
rect 38220 24558 38222 24610
rect 38274 24558 38276 24610
rect 38108 24498 38164 24510
rect 38108 24446 38110 24498
rect 38162 24446 38164 24498
rect 36988 23940 37044 23950
rect 36876 23938 37044 23940
rect 36876 23886 36990 23938
rect 37042 23886 37044 23938
rect 36876 23884 37044 23886
rect 36988 23874 37044 23884
rect 35868 23154 36036 23156
rect 35868 23102 35870 23154
rect 35922 23102 36036 23154
rect 35868 23100 36036 23102
rect 36092 23828 36148 23838
rect 35868 23090 35924 23100
rect 35308 23042 35364 23054
rect 35308 22990 35310 23042
rect 35362 22990 35364 23042
rect 34748 22932 34804 22942
rect 33852 22540 34132 22596
rect 34188 22930 34804 22932
rect 34188 22878 34750 22930
rect 34802 22878 34804 22930
rect 34188 22876 34804 22878
rect 33852 22482 33908 22540
rect 33852 22430 33854 22482
rect 33906 22430 33908 22482
rect 33852 22372 33908 22430
rect 33852 22306 33908 22316
rect 33852 21700 33908 21710
rect 33852 21606 33908 21644
rect 33684 21084 33796 21140
rect 33628 21074 33684 21084
rect 33852 20804 33908 20814
rect 33740 20020 33796 20030
rect 33516 19908 33572 19918
rect 33404 19906 33572 19908
rect 33404 19854 33518 19906
rect 33570 19854 33572 19906
rect 33404 19852 33572 19854
rect 33404 19460 33460 19470
rect 33404 19346 33460 19404
rect 33516 19458 33572 19852
rect 33516 19406 33518 19458
rect 33570 19406 33572 19458
rect 33516 19394 33572 19406
rect 33404 19294 33406 19346
rect 33458 19294 33460 19346
rect 33404 19282 33460 19294
rect 33740 19234 33796 19964
rect 33740 19182 33742 19234
rect 33794 19182 33796 19234
rect 33740 19170 33796 19182
rect 32956 19030 33012 19068
rect 33292 18676 33348 18686
rect 33292 18562 33348 18620
rect 33292 18510 33294 18562
rect 33346 18510 33348 18562
rect 33292 18498 33348 18510
rect 33740 18676 33796 18686
rect 33068 18450 33124 18462
rect 33068 18398 33070 18450
rect 33122 18398 33124 18450
rect 33068 18340 33124 18398
rect 33628 18452 33684 18462
rect 33628 18358 33684 18396
rect 33516 18340 33572 18350
rect 32844 18116 32900 18126
rect 32844 17666 32900 18060
rect 33068 17892 33124 18284
rect 33068 17826 33124 17836
rect 33404 18338 33572 18340
rect 33404 18286 33518 18338
rect 33570 18286 33572 18338
rect 33404 18284 33572 18286
rect 32844 17614 32846 17666
rect 32898 17614 32900 17666
rect 32844 17602 32900 17614
rect 33292 17554 33348 17566
rect 33292 17502 33294 17554
rect 33346 17502 33348 17554
rect 33180 17444 33236 17454
rect 33180 17350 33236 17388
rect 33292 17220 33348 17502
rect 33180 17164 33348 17220
rect 33180 17108 33236 17164
rect 33180 17042 33236 17052
rect 33292 16996 33348 17006
rect 33068 16884 33124 16894
rect 33068 16790 33124 16828
rect 33292 15148 33348 16940
rect 33404 16212 33460 18284
rect 33516 18274 33572 18284
rect 33740 18116 33796 18620
rect 33516 18060 33796 18116
rect 33516 17666 33572 18060
rect 33852 18004 33908 20748
rect 34188 20244 34244 22876
rect 34748 22866 34804 22876
rect 35308 22932 35364 22990
rect 35308 22866 35364 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35084 22484 35140 22494
rect 35084 22390 35140 22428
rect 35980 22484 36036 22494
rect 36092 22484 36148 23772
rect 37772 23828 37828 23838
rect 37772 23734 37828 23772
rect 36540 23044 36596 23054
rect 36540 22950 36596 22988
rect 37436 23044 37492 23054
rect 35980 22482 36148 22484
rect 35980 22430 35982 22482
rect 36034 22430 36148 22482
rect 35980 22428 36148 22430
rect 37436 22482 37492 22988
rect 37436 22430 37438 22482
rect 37490 22430 37492 22482
rect 35980 22418 36036 22428
rect 37436 22418 37492 22430
rect 35644 22372 35700 22382
rect 35644 22278 35700 22316
rect 36988 22372 37044 22382
rect 36988 22278 37044 22316
rect 35308 22260 35364 22270
rect 35196 22204 35308 22260
rect 34300 22146 34356 22158
rect 34300 22094 34302 22146
rect 34354 22094 34356 22146
rect 34300 21588 34356 22094
rect 35084 22036 35140 22046
rect 34300 21522 34356 21532
rect 34636 21700 34692 21710
rect 34636 21586 34692 21644
rect 34636 21534 34638 21586
rect 34690 21534 34692 21586
rect 34636 21522 34692 21534
rect 34076 20188 34244 20244
rect 34412 21474 34468 21486
rect 34412 21422 34414 21474
rect 34466 21422 34468 21474
rect 34412 21364 34468 21422
rect 34972 21476 35028 21486
rect 34860 21364 34916 21374
rect 34412 21362 34916 21364
rect 34412 21310 34862 21362
rect 34914 21310 34916 21362
rect 34412 21308 34916 21310
rect 34076 19236 34132 20188
rect 34188 20018 34244 20030
rect 34188 19966 34190 20018
rect 34242 19966 34244 20018
rect 34188 19460 34244 19966
rect 34412 19908 34468 21308
rect 34860 21298 34916 21308
rect 34412 19842 34468 19852
rect 34636 21140 34692 21150
rect 34636 19906 34692 21084
rect 34636 19854 34638 19906
rect 34690 19854 34692 19906
rect 34636 19684 34692 19854
rect 34188 19394 34244 19404
rect 34412 19628 34692 19684
rect 34076 19180 34244 19236
rect 34076 19012 34132 19022
rect 34076 18918 34132 18956
rect 34188 18788 34244 19180
rect 34412 18900 34468 19628
rect 34972 19460 35028 21420
rect 35084 20188 35140 21980
rect 35196 21810 35252 22204
rect 35308 22166 35364 22204
rect 35868 22260 35924 22270
rect 35868 22166 35924 22204
rect 37548 22260 37604 22270
rect 37884 22260 37940 22270
rect 37604 22258 37940 22260
rect 37604 22206 37886 22258
rect 37938 22206 37940 22258
rect 37604 22204 37940 22206
rect 37548 22166 37604 22204
rect 37884 22194 37940 22204
rect 35420 22148 35476 22158
rect 36092 22148 36148 22158
rect 35420 22146 35588 22148
rect 35420 22094 35422 22146
rect 35474 22094 35588 22146
rect 35420 22092 35588 22094
rect 35420 22082 35476 22092
rect 35196 21758 35198 21810
rect 35250 21758 35252 21810
rect 35196 21746 35252 21758
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 20132 35476 20188
rect 35084 20130 35140 20132
rect 35084 20078 35086 20130
rect 35138 20078 35140 20130
rect 35084 20066 35140 20078
rect 35308 20020 35364 20030
rect 35308 19796 35364 19964
rect 34524 19404 35028 19460
rect 35084 19740 35364 19796
rect 35420 19796 35476 20132
rect 35084 19460 35140 19740
rect 35420 19730 35476 19740
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34524 19122 34580 19404
rect 35084 19234 35140 19404
rect 35084 19182 35086 19234
rect 35138 19182 35140 19234
rect 34524 19070 34526 19122
rect 34578 19070 34580 19122
rect 34524 19012 34580 19070
rect 34748 19122 34804 19134
rect 34748 19070 34750 19122
rect 34802 19070 34804 19122
rect 34524 18946 34580 18956
rect 34636 19010 34692 19022
rect 34636 18958 34638 19010
rect 34690 18958 34692 19010
rect 33516 17614 33518 17666
rect 33570 17614 33572 17666
rect 33516 17602 33572 17614
rect 33628 17948 33908 18004
rect 34076 18732 34244 18788
rect 34300 18844 34468 18900
rect 33404 16156 33572 16212
rect 32732 15092 32900 15148
rect 31724 12516 31780 15092
rect 32620 14980 32676 14990
rect 32508 14924 32620 14980
rect 31948 14644 32004 14654
rect 31948 14550 32004 14588
rect 32284 14420 32340 14430
rect 31948 14306 32004 14318
rect 32172 14308 32228 14318
rect 31948 14254 31950 14306
rect 32002 14254 32004 14306
rect 31948 14196 32004 14254
rect 31948 14130 32004 14140
rect 32060 14306 32228 14308
rect 32060 14254 32174 14306
rect 32226 14254 32228 14306
rect 32060 14252 32228 14254
rect 32060 13970 32116 14252
rect 32172 14242 32228 14252
rect 32060 13918 32062 13970
rect 32114 13918 32116 13970
rect 32060 13906 32116 13918
rect 32172 13972 32228 13982
rect 32284 13972 32340 14364
rect 32172 13970 32340 13972
rect 32172 13918 32174 13970
rect 32226 13918 32340 13970
rect 32172 13916 32340 13918
rect 32396 14418 32452 14430
rect 32396 14366 32398 14418
rect 32450 14366 32452 14418
rect 31948 13746 32004 13758
rect 31948 13694 31950 13746
rect 32002 13694 32004 13746
rect 31836 12740 31892 12750
rect 31836 12646 31892 12684
rect 31724 12460 31892 12516
rect 31388 12180 31444 12190
rect 31724 12180 31780 12190
rect 31388 12178 31780 12180
rect 31388 12126 31390 12178
rect 31442 12126 31726 12178
rect 31778 12126 31780 12178
rect 31388 12124 31780 12126
rect 31388 11956 31444 12124
rect 31724 12114 31780 12124
rect 31388 11890 31444 11900
rect 31836 11394 31892 12460
rect 31836 11342 31838 11394
rect 31890 11342 31892 11394
rect 31836 11330 31892 11342
rect 31500 11170 31556 11182
rect 31500 11118 31502 11170
rect 31554 11118 31556 11170
rect 31164 10610 31332 10612
rect 31164 10558 31166 10610
rect 31218 10558 31332 10610
rect 31164 10556 31332 10558
rect 31388 10722 31444 10734
rect 31388 10670 31390 10722
rect 31442 10670 31444 10722
rect 31164 10546 31220 10556
rect 31388 8932 31444 10670
rect 31388 8866 31444 8876
rect 31276 8148 31332 8158
rect 31276 8054 31332 8092
rect 31500 7588 31556 11118
rect 31948 10276 32004 13694
rect 32060 13748 32116 13758
rect 32060 12404 32116 13692
rect 32172 13300 32228 13916
rect 32396 13636 32452 14366
rect 32508 13746 32564 14924
rect 32620 14914 32676 14924
rect 32620 14308 32676 14318
rect 32620 14214 32676 14252
rect 32732 14306 32788 14318
rect 32732 14254 32734 14306
rect 32786 14254 32788 14306
rect 32732 14196 32788 14254
rect 32732 14130 32788 14140
rect 32844 13860 32900 15092
rect 33068 15092 33348 15148
rect 33404 15988 33460 15998
rect 32956 14308 33012 14318
rect 32956 14214 33012 14252
rect 33068 13972 33124 15092
rect 32508 13694 32510 13746
rect 32562 13694 32564 13746
rect 32508 13682 32564 13694
rect 32620 13804 32900 13860
rect 32956 13916 33124 13972
rect 33180 14418 33236 14430
rect 33180 14366 33182 14418
rect 33234 14366 33236 14418
rect 32396 13570 32452 13580
rect 32620 13524 32676 13804
rect 32172 13234 32228 13244
rect 32508 13468 32676 13524
rect 32172 12852 32228 12862
rect 32396 12852 32452 12862
rect 32172 12850 32396 12852
rect 32172 12798 32174 12850
rect 32226 12798 32396 12850
rect 32172 12796 32396 12798
rect 32172 12786 32228 12796
rect 32396 12786 32452 12796
rect 32060 12310 32116 12348
rect 32508 10836 32564 13468
rect 32956 12850 33012 13916
rect 32956 12798 32958 12850
rect 33010 12798 33012 12850
rect 32956 12786 33012 12798
rect 33068 13746 33124 13758
rect 33068 13694 33070 13746
rect 33122 13694 33124 13746
rect 32508 10770 32564 10780
rect 32620 12738 32676 12750
rect 32620 12686 32622 12738
rect 32674 12686 32676 12738
rect 32620 10500 32676 12686
rect 32844 12738 32900 12750
rect 32844 12686 32846 12738
rect 32898 12686 32900 12738
rect 32844 12404 32900 12686
rect 32844 12338 32900 12348
rect 32172 10444 32676 10500
rect 31948 10220 32116 10276
rect 31948 10050 32004 10062
rect 31948 9998 31950 10050
rect 32002 9998 32004 10050
rect 31948 9938 32004 9998
rect 31948 9886 31950 9938
rect 32002 9886 32004 9938
rect 31948 9874 32004 9886
rect 31948 8148 32004 8158
rect 31948 8054 32004 8092
rect 31500 6692 31556 7532
rect 32060 6804 32116 10220
rect 32172 8260 32228 10444
rect 33068 10276 33124 13694
rect 33180 13076 33236 14366
rect 33292 13860 33348 13898
rect 33292 13794 33348 13804
rect 33404 13858 33460 15932
rect 33516 14980 33572 16156
rect 33628 15148 33684 17948
rect 34076 17666 34132 18732
rect 34300 18676 34356 18844
rect 34076 17614 34078 17666
rect 34130 17614 34132 17666
rect 34076 17602 34132 17614
rect 34188 18620 34356 18676
rect 34636 18676 34692 18958
rect 33964 17556 34020 17566
rect 33740 17442 33796 17454
rect 33740 17390 33742 17442
rect 33794 17390 33796 17442
rect 33740 16996 33796 17390
rect 33740 16930 33796 16940
rect 33852 17444 33908 17454
rect 33852 16994 33908 17388
rect 33964 17442 34020 17500
rect 33964 17390 33966 17442
rect 34018 17390 34020 17442
rect 33964 17378 34020 17390
rect 33852 16942 33854 16994
rect 33906 16942 33908 16994
rect 33852 16930 33908 16942
rect 34188 15148 34244 18620
rect 34636 18610 34692 18620
rect 34748 18564 34804 19070
rect 35084 18676 35140 19182
rect 35420 19124 35476 19134
rect 35532 19124 35588 22092
rect 36092 22054 36148 22092
rect 36316 22148 36372 22158
rect 36316 22054 36372 22092
rect 37324 22146 37380 22158
rect 37324 22094 37326 22146
rect 37378 22094 37380 22146
rect 37324 21924 37380 22094
rect 37324 21858 37380 21868
rect 37996 22146 38052 22158
rect 37996 22094 37998 22146
rect 38050 22094 38052 22146
rect 36428 21700 36484 21710
rect 35084 18610 35140 18620
rect 35308 19122 35588 19124
rect 35308 19070 35422 19122
rect 35474 19070 35588 19122
rect 35308 19068 35588 19070
rect 35644 21588 35700 21598
rect 35756 21588 35812 21598
rect 35700 21586 35812 21588
rect 35700 21534 35758 21586
rect 35810 21534 35812 21586
rect 35700 21532 35812 21534
rect 35644 20914 35700 21532
rect 35756 21522 35812 21532
rect 35644 20862 35646 20914
rect 35698 20862 35700 20914
rect 35644 19908 35700 20862
rect 36428 20804 36484 21644
rect 37996 21588 38052 22094
rect 38108 21924 38164 24446
rect 38220 23044 38276 24558
rect 38668 24612 38724 24622
rect 38668 24610 39956 24612
rect 38668 24558 38670 24610
rect 38722 24558 39956 24610
rect 38668 24556 39956 24558
rect 38668 24546 38724 24556
rect 38220 22978 38276 22988
rect 38556 24498 38612 24510
rect 38556 24446 38558 24498
rect 38610 24446 38612 24498
rect 38220 22148 38276 22158
rect 38220 22054 38276 22092
rect 38556 22036 38612 24446
rect 39900 24050 39956 24556
rect 39900 23998 39902 24050
rect 39954 23998 39956 24050
rect 39900 23986 39956 23998
rect 38668 23044 38724 23054
rect 38668 22950 38724 22988
rect 42476 22484 42532 22494
rect 42924 22484 42980 22494
rect 42476 22482 42980 22484
rect 42476 22430 42478 22482
rect 42530 22430 42926 22482
rect 42978 22430 42980 22482
rect 42476 22428 42980 22430
rect 42476 22418 42532 22428
rect 42924 22418 42980 22428
rect 43372 22482 43428 25564
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 43372 22430 43374 22482
rect 43426 22430 43428 22482
rect 38556 21970 38612 21980
rect 39676 22370 39732 22382
rect 39676 22318 39678 22370
rect 39730 22318 39732 22370
rect 38108 21858 38164 21868
rect 37996 21522 38052 21532
rect 39228 21812 39284 21822
rect 36540 21476 36596 21486
rect 36540 21474 37156 21476
rect 36540 21422 36542 21474
rect 36594 21422 37156 21474
rect 36540 21420 37156 21422
rect 36540 21410 36596 21420
rect 37100 20914 37156 21420
rect 38668 21474 38724 21486
rect 38668 21422 38670 21474
rect 38722 21422 38724 21474
rect 37100 20862 37102 20914
rect 37154 20862 37156 20914
rect 37100 20850 37156 20862
rect 37772 20916 37828 20926
rect 36428 20710 36484 20748
rect 36876 20802 36932 20814
rect 36876 20750 36878 20802
rect 36930 20750 36932 20802
rect 35980 20692 36036 20702
rect 34748 18508 35028 18564
rect 34412 18450 34468 18462
rect 34412 18398 34414 18450
rect 34466 18398 34468 18450
rect 34412 18340 34468 18398
rect 34412 18274 34468 18284
rect 34524 18452 34580 18462
rect 34524 18004 34580 18396
rect 34524 17938 34580 17948
rect 34636 18450 34692 18462
rect 34636 18398 34638 18450
rect 34690 18398 34692 18450
rect 34524 17554 34580 17566
rect 34524 17502 34526 17554
rect 34578 17502 34580 17554
rect 34412 17442 34468 17454
rect 34412 17390 34414 17442
rect 34466 17390 34468 17442
rect 34412 17108 34468 17390
rect 34412 17042 34468 17052
rect 34524 16772 34580 17502
rect 34636 17556 34692 18398
rect 34860 18340 34916 18350
rect 34636 17490 34692 17500
rect 34748 18338 34916 18340
rect 34748 18286 34862 18338
rect 34914 18286 34916 18338
rect 34748 18284 34916 18286
rect 34524 16706 34580 16716
rect 34524 16212 34580 16222
rect 34300 16100 34356 16110
rect 34300 16006 34356 16044
rect 34524 16098 34580 16156
rect 34524 16046 34526 16098
rect 34578 16046 34580 16098
rect 34524 16034 34580 16046
rect 34636 15874 34692 15886
rect 34636 15822 34638 15874
rect 34690 15822 34692 15874
rect 33628 15092 34020 15148
rect 34188 15092 34580 15148
rect 33516 14914 33572 14924
rect 33404 13806 33406 13858
rect 33458 13806 33460 13858
rect 33404 13794 33460 13806
rect 33852 13860 33908 13870
rect 33852 13748 33908 13804
rect 33516 13746 33908 13748
rect 33516 13694 33854 13746
rect 33906 13694 33908 13746
rect 33516 13692 33908 13694
rect 33292 13636 33348 13646
rect 33292 13542 33348 13580
rect 33404 13076 33460 13086
rect 33180 13074 33460 13076
rect 33180 13022 33406 13074
rect 33458 13022 33460 13074
rect 33180 13020 33460 13022
rect 33404 13010 33460 13020
rect 33180 12852 33236 12862
rect 33516 12852 33572 13692
rect 33852 13682 33908 13692
rect 33236 12796 33572 12852
rect 33180 12758 33236 12796
rect 33852 12290 33908 12302
rect 33852 12238 33854 12290
rect 33906 12238 33908 12290
rect 33628 12180 33684 12190
rect 33628 12178 33796 12180
rect 33628 12126 33630 12178
rect 33682 12126 33796 12178
rect 33628 12124 33796 12126
rect 33628 12114 33684 12124
rect 32508 10220 33124 10276
rect 33180 11508 33236 11518
rect 33180 11394 33236 11452
rect 33180 11342 33182 11394
rect 33234 11342 33236 11394
rect 32396 9828 32452 9838
rect 32396 9734 32452 9772
rect 32508 8932 32564 10220
rect 33180 10052 33236 11342
rect 33404 10836 33460 10846
rect 33740 10836 33796 12124
rect 33852 11506 33908 12238
rect 33852 11454 33854 11506
rect 33906 11454 33908 11506
rect 33852 11442 33908 11454
rect 33852 10836 33908 10846
rect 33740 10834 33908 10836
rect 33740 10782 33854 10834
rect 33906 10782 33908 10834
rect 33740 10780 33908 10782
rect 33404 10742 33460 10780
rect 33852 10770 33908 10780
rect 33068 10050 33236 10052
rect 33068 9998 33182 10050
rect 33234 9998 33236 10050
rect 33068 9996 33236 9998
rect 32844 9604 32900 9614
rect 32844 9510 32900 9548
rect 32284 8930 32564 8932
rect 32284 8878 32510 8930
rect 32562 8878 32564 8930
rect 32284 8876 32564 8878
rect 32284 8482 32340 8876
rect 32508 8866 32564 8876
rect 33068 8820 33124 9996
rect 33180 9986 33236 9996
rect 33964 10052 34020 15092
rect 34300 14308 34356 14318
rect 34300 13970 34356 14252
rect 34300 13918 34302 13970
rect 34354 13918 34356 13970
rect 34300 13906 34356 13918
rect 34188 13748 34244 13758
rect 33964 9986 34020 9996
rect 34076 13746 34244 13748
rect 34076 13694 34190 13746
rect 34242 13694 34244 13746
rect 34076 13692 34244 13694
rect 33404 9828 33460 9838
rect 33404 9734 33460 9772
rect 33628 9826 33684 9838
rect 33628 9774 33630 9826
rect 33682 9774 33684 9826
rect 33628 9604 33684 9774
rect 33628 9538 33684 9548
rect 33964 9602 34020 9614
rect 33964 9550 33966 9602
rect 34018 9550 34020 9602
rect 33628 9380 33684 9390
rect 33404 9268 33460 9278
rect 33292 9212 33404 9268
rect 33180 9156 33236 9166
rect 33180 9062 33236 9100
rect 33292 9154 33348 9212
rect 33404 9202 33460 9212
rect 33292 9102 33294 9154
rect 33346 9102 33348 9154
rect 33292 9090 33348 9102
rect 33628 9156 33684 9324
rect 33852 9268 33908 9278
rect 33516 9044 33572 9054
rect 33404 9042 33572 9044
rect 33404 8990 33518 9042
rect 33570 8990 33572 9042
rect 33404 8988 33572 8990
rect 33068 8754 33124 8764
rect 33180 8818 33236 8830
rect 33180 8766 33182 8818
rect 33234 8766 33236 8818
rect 32284 8430 32286 8482
rect 32338 8430 32340 8482
rect 32284 8418 32340 8430
rect 33068 8596 33124 8606
rect 32172 8204 32564 8260
rect 32508 7364 32564 8204
rect 33068 8258 33124 8540
rect 33068 8206 33070 8258
rect 33122 8206 33124 8258
rect 32396 7362 32564 7364
rect 32396 7310 32510 7362
rect 32562 7310 32564 7362
rect 32396 7308 32564 7310
rect 32396 6914 32452 7308
rect 32508 7298 32564 7308
rect 32844 8146 32900 8158
rect 32844 8094 32846 8146
rect 32898 8094 32900 8146
rect 32396 6862 32398 6914
rect 32450 6862 32452 6914
rect 32396 6850 32452 6862
rect 31500 6626 31556 6636
rect 31948 6748 32116 6804
rect 32844 6804 32900 8094
rect 31276 6580 31332 6590
rect 31276 6486 31332 6524
rect 31052 6066 31108 6076
rect 30268 6020 30324 6030
rect 28700 5966 28702 6018
rect 28754 5966 28756 6018
rect 28700 5954 28756 5966
rect 29932 6018 30324 6020
rect 29932 5966 30270 6018
rect 30322 5966 30324 6018
rect 29932 5964 30324 5966
rect 28924 5796 28980 5806
rect 28924 5702 28980 5740
rect 29260 5236 29316 5246
rect 28532 4956 28868 5012
rect 28476 4946 28532 4956
rect 27356 4898 27412 4910
rect 27356 4846 27358 4898
rect 27410 4846 27412 4898
rect 24332 4470 24388 4508
rect 25564 4564 25620 4574
rect 25564 4470 25620 4508
rect 26012 4564 26068 4574
rect 23548 4398 23550 4450
rect 23602 4398 23604 4450
rect 23548 4386 23604 4398
rect 26012 4338 26068 4508
rect 26012 4286 26014 4338
rect 26066 4286 26068 4338
rect 26012 4274 26068 4286
rect 23212 4228 23268 4238
rect 22988 4226 23268 4228
rect 22988 4174 23214 4226
rect 23266 4174 23268 4226
rect 22988 4172 23268 4174
rect 23212 4162 23268 4172
rect 26684 4228 26740 4238
rect 26684 4226 27076 4228
rect 26684 4174 26686 4226
rect 26738 4174 27076 4226
rect 26684 4172 27076 4174
rect 26684 4162 26740 4172
rect 22876 3614 22878 3666
rect 22930 3614 22932 3666
rect 22876 3602 22932 3614
rect 27020 3442 27076 4172
rect 27356 3554 27412 4846
rect 28812 4226 28868 4956
rect 29260 4338 29316 5180
rect 29932 4450 29988 5964
rect 30268 5954 30324 5964
rect 30604 5908 30660 5918
rect 31276 5908 31332 5918
rect 30604 5906 31332 5908
rect 30604 5854 30606 5906
rect 30658 5854 31278 5906
rect 31330 5854 31332 5906
rect 30604 5852 31332 5854
rect 30604 5842 30660 5852
rect 31276 5842 31332 5852
rect 31612 5908 31668 5918
rect 31948 5908 32004 6748
rect 32060 6580 32116 6590
rect 32060 6486 32116 6524
rect 32844 6132 32900 6748
rect 33068 6690 33124 8206
rect 33068 6638 33070 6690
rect 33122 6638 33124 6690
rect 33068 6626 33124 6638
rect 32844 6066 32900 6076
rect 32956 6578 33012 6590
rect 32956 6526 32958 6578
rect 33010 6526 33012 6578
rect 32956 6468 33012 6526
rect 32172 6020 32228 6030
rect 32172 5926 32228 5964
rect 32396 6020 32452 6030
rect 31612 5906 32004 5908
rect 31612 5854 31614 5906
rect 31666 5854 32004 5906
rect 31612 5852 32004 5854
rect 31612 5842 31668 5852
rect 30156 5684 30212 5694
rect 30156 5122 30212 5628
rect 30156 5070 30158 5122
rect 30210 5070 30212 5122
rect 30156 5058 30212 5070
rect 30380 5404 30996 5460
rect 30380 5010 30436 5404
rect 30828 5236 30884 5246
rect 30940 5236 30996 5404
rect 31500 5236 31556 5246
rect 30940 5234 31556 5236
rect 30940 5182 31502 5234
rect 31554 5182 31556 5234
rect 30940 5180 31556 5182
rect 30828 5122 30884 5180
rect 31500 5170 31556 5180
rect 30828 5070 30830 5122
rect 30882 5070 30884 5122
rect 30828 5058 30884 5070
rect 30380 4958 30382 5010
rect 30434 4958 30436 5010
rect 30380 4946 30436 4958
rect 29932 4398 29934 4450
rect 29986 4398 29988 4450
rect 29932 4386 29988 4398
rect 29260 4286 29262 4338
rect 29314 4286 29316 4338
rect 29260 4274 29316 4286
rect 28812 4174 28814 4226
rect 28866 4174 28868 4226
rect 28812 4162 28868 4174
rect 31948 4228 32004 5852
rect 32396 5906 32452 5964
rect 32396 5854 32398 5906
rect 32450 5854 32452 5906
rect 32396 5842 32452 5854
rect 32956 5796 33012 6412
rect 33180 6020 33236 8766
rect 33404 8596 33460 8988
rect 33516 8978 33572 8988
rect 33404 8530 33460 8540
rect 33516 8820 33572 8830
rect 33516 8484 33572 8764
rect 33628 8596 33684 9100
rect 33740 9154 33796 9166
rect 33740 9102 33742 9154
rect 33794 9102 33796 9154
rect 33740 9044 33796 9102
rect 33852 9154 33908 9212
rect 33852 9102 33854 9154
rect 33906 9102 33908 9154
rect 33852 9090 33908 9102
rect 33964 9156 34020 9550
rect 33964 9090 34020 9100
rect 33740 8932 33796 8988
rect 33740 8876 33908 8932
rect 33628 8540 33796 8596
rect 33516 8428 33684 8484
rect 33404 8036 33460 8046
rect 33404 7698 33460 7980
rect 33404 7646 33406 7698
rect 33458 7646 33460 7698
rect 33404 7634 33460 7646
rect 33628 7700 33684 8428
rect 33740 8370 33796 8540
rect 33740 8318 33742 8370
rect 33794 8318 33796 8370
rect 33740 8306 33796 8318
rect 33740 8036 33796 8046
rect 33852 8036 33908 8876
rect 33796 7980 33908 8036
rect 33740 7970 33796 7980
rect 33740 7700 33796 7710
rect 33628 7698 33796 7700
rect 33628 7646 33742 7698
rect 33794 7646 33796 7698
rect 33628 7644 33796 7646
rect 33740 7634 33796 7644
rect 34076 6692 34132 13692
rect 34188 13682 34244 13692
rect 34412 13748 34468 13758
rect 34412 13654 34468 13692
rect 34300 12292 34356 12302
rect 34300 12198 34356 12236
rect 34188 10836 34244 10846
rect 34188 10610 34244 10780
rect 34188 10558 34190 10610
rect 34242 10558 34244 10610
rect 34188 10546 34244 10558
rect 34524 10724 34580 15092
rect 34636 12850 34692 15822
rect 34748 13746 34804 18284
rect 34860 18274 34916 18284
rect 34860 18116 34916 18126
rect 34972 18116 35028 18508
rect 35084 18452 35140 18462
rect 35084 18358 35140 18396
rect 35308 18340 35364 19068
rect 35420 19058 35476 19068
rect 35420 18676 35476 18686
rect 35420 18582 35476 18620
rect 35308 18274 35364 18284
rect 34916 18060 35028 18116
rect 34860 18050 34916 18060
rect 34972 17780 35028 18060
rect 34972 17714 35028 17724
rect 35084 18228 35140 18238
rect 35084 17666 35140 18172
rect 35532 18228 35588 18238
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35084 17614 35086 17666
rect 35138 17614 35140 17666
rect 35084 17602 35140 17614
rect 35532 17666 35588 18172
rect 35532 17614 35534 17666
rect 35586 17614 35588 17666
rect 35532 17602 35588 17614
rect 35196 17556 35252 17566
rect 35196 17462 35252 17500
rect 35308 17442 35364 17454
rect 35308 17390 35310 17442
rect 35362 17390 35364 17442
rect 34972 16996 35028 17006
rect 34860 16940 34972 16996
rect 34860 16098 34916 16940
rect 34972 16930 35028 16940
rect 35308 16660 35364 17390
rect 35532 16884 35588 16894
rect 35644 16884 35700 19852
rect 35756 20580 35812 20590
rect 35756 19234 35812 20524
rect 35868 20020 35924 20030
rect 35868 19926 35924 19964
rect 35756 19182 35758 19234
rect 35810 19182 35812 19234
rect 35756 19170 35812 19182
rect 35868 19796 35924 19806
rect 35868 18674 35924 19740
rect 35980 19346 36036 20636
rect 35980 19294 35982 19346
rect 36034 19294 36036 19346
rect 35980 19282 36036 19294
rect 36092 20578 36148 20590
rect 36092 20526 36094 20578
rect 36146 20526 36148 20578
rect 36092 20188 36148 20526
rect 36316 20578 36372 20590
rect 36316 20526 36318 20578
rect 36370 20526 36372 20578
rect 36316 20468 36372 20526
rect 36316 20402 36372 20412
rect 36876 20188 36932 20750
rect 37324 20690 37380 20702
rect 37324 20638 37326 20690
rect 37378 20638 37380 20690
rect 36092 20132 36932 20188
rect 37212 20468 37268 20478
rect 37212 20244 37268 20412
rect 37212 20178 37268 20188
rect 37324 20468 37380 20638
rect 37548 20692 37604 20702
rect 37548 20598 37604 20636
rect 37772 20692 37828 20860
rect 37996 20916 38052 20926
rect 37996 20822 38052 20860
rect 38668 20916 38724 21422
rect 39116 21362 39172 21374
rect 39116 21310 39118 21362
rect 39170 21310 39172 21362
rect 39116 21028 39172 21310
rect 38668 20850 38724 20860
rect 38892 20972 39172 21028
rect 38444 20804 38500 20814
rect 37772 20626 37828 20636
rect 38332 20692 38388 20702
rect 38332 20598 38388 20636
rect 38444 20690 38500 20748
rect 38444 20638 38446 20690
rect 38498 20638 38500 20690
rect 37884 20578 37940 20590
rect 37884 20526 37886 20578
rect 37938 20526 37940 20578
rect 37884 20468 37940 20526
rect 37324 20412 37940 20468
rect 35868 18622 35870 18674
rect 35922 18622 35924 18674
rect 35868 18610 35924 18622
rect 36092 19122 36148 20132
rect 36764 20130 36820 20132
rect 36764 20078 36766 20130
rect 36818 20078 36820 20130
rect 36764 20066 36820 20078
rect 36092 19070 36094 19122
rect 36146 19070 36148 19122
rect 36092 18450 36148 19070
rect 36092 18398 36094 18450
rect 36146 18398 36148 18450
rect 36092 18386 36148 18398
rect 36204 20018 36260 20030
rect 36204 19966 36206 20018
rect 36258 19966 36260 20018
rect 35980 18338 36036 18350
rect 35980 18286 35982 18338
rect 36034 18286 36036 18338
rect 35980 18228 36036 18286
rect 36204 18228 36260 19966
rect 36540 20018 36596 20030
rect 36540 19966 36542 20018
rect 36594 19966 36596 20018
rect 35980 18172 36260 18228
rect 36316 18340 36372 18350
rect 36092 17892 36148 17902
rect 35980 17890 36148 17892
rect 35980 17838 36094 17890
rect 36146 17838 36148 17890
rect 35980 17836 36148 17838
rect 35980 17780 36036 17836
rect 36092 17826 36148 17836
rect 36316 17892 36372 18284
rect 36540 18340 36596 19966
rect 36652 19906 36708 19918
rect 36652 19854 36654 19906
rect 36706 19854 36708 19906
rect 36652 19348 36708 19854
rect 37212 19908 37268 19918
rect 37212 19814 37268 19852
rect 37324 19572 37380 20412
rect 36652 19282 36708 19292
rect 37212 19516 37380 19572
rect 37660 20244 37716 20254
rect 37660 20130 37716 20188
rect 38444 20188 38500 20638
rect 38668 20692 38724 20702
rect 38892 20692 38948 20972
rect 39004 20804 39060 20814
rect 39004 20710 39060 20748
rect 38668 20690 38892 20692
rect 38668 20638 38670 20690
rect 38722 20638 38892 20690
rect 38668 20636 38892 20638
rect 38668 20626 38724 20636
rect 38892 20598 38948 20636
rect 38892 20356 38948 20366
rect 38444 20132 38724 20188
rect 37660 20078 37662 20130
rect 37714 20078 37716 20130
rect 36540 18274 36596 18284
rect 37100 19234 37156 19246
rect 37100 19182 37102 19234
rect 37154 19182 37156 19234
rect 35980 17714 36036 17724
rect 36204 17780 36260 17790
rect 36204 17686 36260 17724
rect 36316 17554 36372 17836
rect 36316 17502 36318 17554
rect 36370 17502 36372 17554
rect 36316 17490 36372 17502
rect 36428 18004 36484 18014
rect 35588 16828 35700 16884
rect 36204 16884 36260 16894
rect 35532 16818 35588 16828
rect 35980 16772 36036 16782
rect 35980 16678 36036 16716
rect 34860 16046 34862 16098
rect 34914 16046 34916 16098
rect 34860 16034 34916 16046
rect 34972 16604 35364 16660
rect 34860 14420 34916 14430
rect 34972 14420 35028 16604
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 36204 15876 36260 16828
rect 36428 16882 36484 17948
rect 37100 18004 37156 19182
rect 36876 17668 36932 17678
rect 36876 17574 36932 17612
rect 37100 17668 37156 17948
rect 37100 17602 37156 17612
rect 37100 17442 37156 17454
rect 37100 17390 37102 17442
rect 37154 17390 37156 17442
rect 37100 16994 37156 17390
rect 37100 16942 37102 16994
rect 37154 16942 37156 16994
rect 37100 16930 37156 16942
rect 36428 16830 36430 16882
rect 36482 16830 36484 16882
rect 36428 16818 36484 16830
rect 36204 15874 36372 15876
rect 36204 15822 36206 15874
rect 36258 15822 36372 15874
rect 36204 15820 36372 15822
rect 36204 15810 36260 15820
rect 36092 15090 36148 15102
rect 36092 15038 36094 15090
rect 36146 15038 36148 15090
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35980 14756 36036 14766
rect 36092 14756 36148 15038
rect 35308 14700 35812 14756
rect 35308 14530 35364 14700
rect 35308 14478 35310 14530
rect 35362 14478 35364 14530
rect 35308 14466 35364 14478
rect 35644 14530 35700 14542
rect 35644 14478 35646 14530
rect 35698 14478 35700 14530
rect 34860 14418 35028 14420
rect 34860 14366 34862 14418
rect 34914 14366 35028 14418
rect 34860 14364 35028 14366
rect 35084 14420 35140 14430
rect 34860 14354 34916 14364
rect 35084 14326 35140 14364
rect 35196 14306 35252 14318
rect 35196 14254 35198 14306
rect 35250 14254 35252 14306
rect 35196 14084 35252 14254
rect 34972 14028 35252 14084
rect 34748 13694 34750 13746
rect 34802 13694 34804 13746
rect 34748 13682 34804 13694
rect 34860 13748 34916 13758
rect 34860 12962 34916 13692
rect 34972 13188 35028 14028
rect 35308 13972 35364 13982
rect 34972 13122 35028 13132
rect 35084 13970 35364 13972
rect 35084 13918 35310 13970
rect 35362 13918 35364 13970
rect 35084 13916 35364 13918
rect 35084 13076 35140 13916
rect 35308 13906 35364 13916
rect 35644 13860 35700 14478
rect 35420 13804 35700 13860
rect 35420 13746 35476 13804
rect 35420 13694 35422 13746
rect 35474 13694 35476 13746
rect 35420 13524 35476 13694
rect 35420 13458 35476 13468
rect 35644 13524 35700 13534
rect 35644 13430 35700 13468
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35308 13188 35364 13198
rect 35756 13188 35812 14700
rect 35980 14754 36148 14756
rect 35980 14702 35982 14754
rect 36034 14702 36148 14754
rect 35980 14700 36148 14702
rect 35980 14690 36036 14700
rect 36092 14532 36148 14542
rect 35868 14530 36148 14532
rect 35868 14478 36094 14530
rect 36146 14478 36148 14530
rect 35868 14476 36148 14478
rect 35868 13860 35924 14476
rect 36092 14466 36148 14476
rect 35868 13766 35924 13804
rect 35980 14306 36036 14318
rect 35980 14254 35982 14306
rect 36034 14254 36036 14306
rect 35084 13020 35252 13076
rect 34860 12910 34862 12962
rect 34914 12910 34916 12962
rect 34860 12898 34916 12910
rect 34972 12964 35028 12974
rect 34972 12870 35028 12908
rect 34636 12798 34638 12850
rect 34690 12798 34692 12850
rect 34636 12786 34692 12798
rect 34748 12852 34804 12862
rect 34748 12402 34804 12796
rect 34748 12350 34750 12402
rect 34802 12350 34804 12402
rect 34748 12338 34804 12350
rect 35084 12738 35140 12750
rect 35084 12686 35086 12738
rect 35138 12686 35140 12738
rect 34636 12180 34692 12190
rect 34636 12086 34692 12124
rect 34972 12178 35028 12190
rect 34972 12126 34974 12178
rect 35026 12126 35028 12178
rect 34972 11956 35028 12126
rect 34972 11890 35028 11900
rect 34300 10052 34356 10062
rect 34300 9268 34356 9996
rect 34524 10052 34580 10668
rect 34972 10724 35028 10734
rect 34972 10630 35028 10668
rect 34524 9986 34580 9996
rect 34748 10610 34804 10622
rect 34748 10558 34750 10610
rect 34802 10558 34804 10610
rect 34188 8372 34244 8382
rect 34300 8372 34356 9212
rect 34748 9156 34804 10558
rect 34748 9090 34804 9100
rect 35084 9044 35140 12686
rect 35196 12290 35252 13020
rect 35196 12238 35198 12290
rect 35250 12238 35252 12290
rect 35196 12226 35252 12238
rect 35308 12292 35364 13132
rect 35644 13132 35812 13188
rect 35532 13076 35588 13086
rect 35532 12982 35588 13020
rect 35420 12852 35476 12862
rect 35420 12758 35476 12796
rect 35532 12628 35588 12638
rect 35532 12402 35588 12572
rect 35532 12350 35534 12402
rect 35586 12350 35588 12402
rect 35532 12338 35588 12350
rect 35420 12292 35476 12302
rect 35308 12290 35476 12292
rect 35308 12238 35422 12290
rect 35474 12238 35476 12290
rect 35308 12236 35476 12238
rect 35420 12226 35476 12236
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 34972 8988 35140 9044
rect 35196 10052 35252 10062
rect 35196 9492 35252 9996
rect 35644 9828 35700 13132
rect 35756 12964 35812 12974
rect 35756 12870 35812 12908
rect 35980 12962 36036 14254
rect 36092 13748 36148 13758
rect 36092 13654 36148 13692
rect 35980 12910 35982 12962
rect 36034 12910 36036 12962
rect 35980 12898 36036 12910
rect 36204 12404 36260 12414
rect 35868 12402 36260 12404
rect 35868 12350 36206 12402
rect 36258 12350 36260 12402
rect 35868 12348 36260 12350
rect 35868 12178 35924 12348
rect 36204 12338 36260 12348
rect 35868 12126 35870 12178
rect 35922 12126 35924 12178
rect 35868 12114 35924 12126
rect 35980 12178 36036 12190
rect 35980 12126 35982 12178
rect 36034 12126 36036 12178
rect 35980 11732 36036 12126
rect 35868 11676 36036 11732
rect 35868 10834 35924 11676
rect 35868 10782 35870 10834
rect 35922 10782 35924 10834
rect 35868 10770 35924 10782
rect 35980 11506 36036 11518
rect 35980 11454 35982 11506
rect 36034 11454 36036 11506
rect 35980 10724 36036 11454
rect 36316 11508 36372 15820
rect 36540 15540 36596 15550
rect 36428 15538 36596 15540
rect 36428 15486 36542 15538
rect 36594 15486 36596 15538
rect 36428 15484 36596 15486
rect 36428 15090 36484 15484
rect 36540 15474 36596 15484
rect 36988 15540 37044 15550
rect 36428 15038 36430 15090
rect 36482 15038 36484 15090
rect 36428 15026 36484 15038
rect 36540 15316 36596 15326
rect 36428 14420 36484 14430
rect 36428 14326 36484 14364
rect 36428 13970 36484 13982
rect 36428 13918 36430 13970
rect 36482 13918 36484 13970
rect 36428 13524 36484 13918
rect 36540 13746 36596 15260
rect 36988 15314 37044 15484
rect 36988 15262 36990 15314
rect 37042 15262 37044 15314
rect 36876 15204 36932 15214
rect 36876 15090 36932 15148
rect 36876 15038 36878 15090
rect 36930 15038 36932 15090
rect 36876 15026 36932 15038
rect 36988 13858 37044 15262
rect 36988 13806 36990 13858
rect 37042 13806 37044 13858
rect 36988 13794 37044 13806
rect 37212 13858 37268 19516
rect 37548 18340 37604 18350
rect 37436 17780 37492 17790
rect 37436 17666 37492 17724
rect 37436 17614 37438 17666
rect 37490 17614 37492 17666
rect 37436 17602 37492 17614
rect 37324 17554 37380 17566
rect 37324 17502 37326 17554
rect 37378 17502 37380 17554
rect 37324 17444 37380 17502
rect 37324 17388 37492 17444
rect 37436 15876 37492 17388
rect 37436 15810 37492 15820
rect 37324 15428 37380 15438
rect 37548 15428 37604 18284
rect 37324 15426 37604 15428
rect 37324 15374 37326 15426
rect 37378 15374 37604 15426
rect 37324 15372 37604 15374
rect 37324 15362 37380 15372
rect 37660 15148 37716 20078
rect 38668 20130 38724 20132
rect 38668 20078 38670 20130
rect 38722 20078 38724 20130
rect 38668 20066 38724 20078
rect 38780 20130 38836 20142
rect 38780 20078 38782 20130
rect 38834 20078 38836 20130
rect 38332 19908 38388 19918
rect 38780 19908 38836 20078
rect 38332 19906 38836 19908
rect 38332 19854 38334 19906
rect 38386 19854 38836 19906
rect 38332 19852 38836 19854
rect 38892 20020 38948 20300
rect 39116 20132 39172 20142
rect 38332 19842 38388 19852
rect 37772 19348 37828 19358
rect 37772 19254 37828 19292
rect 38108 19348 38164 19358
rect 38108 18450 38164 19292
rect 38108 18398 38110 18450
rect 38162 18398 38164 18450
rect 38108 18386 38164 18398
rect 38444 18788 38500 19852
rect 37996 18340 38052 18350
rect 37996 18246 38052 18284
rect 38220 16772 38276 16782
rect 38220 16210 38276 16716
rect 38220 16158 38222 16210
rect 38274 16158 38276 16210
rect 38220 16146 38276 16158
rect 38108 15876 38164 15886
rect 38108 15782 38164 15820
rect 38444 15148 38500 18732
rect 38780 18676 38836 18686
rect 38892 18676 38948 19964
rect 39004 20076 39116 20132
rect 39004 20018 39060 20076
rect 39004 19966 39006 20018
rect 39058 19966 39060 20018
rect 39004 19954 39060 19966
rect 38780 18674 38948 18676
rect 38780 18622 38782 18674
rect 38834 18622 38948 18674
rect 38780 18620 38948 18622
rect 38780 18610 38836 18620
rect 39116 18564 39172 20076
rect 38892 18562 39172 18564
rect 38892 18510 39118 18562
rect 39170 18510 39172 18562
rect 38892 18508 39172 18510
rect 38892 17666 38948 18508
rect 39116 18498 39172 18508
rect 39228 18116 39284 21756
rect 39340 21698 39396 21710
rect 39340 21646 39342 21698
rect 39394 21646 39396 21698
rect 39340 21588 39396 21646
rect 39676 21700 39732 22318
rect 40348 22260 40404 22270
rect 40236 22258 40404 22260
rect 40236 22206 40350 22258
rect 40402 22206 40404 22258
rect 40236 22204 40404 22206
rect 39676 21634 39732 21644
rect 40124 21812 40180 21822
rect 39340 20244 39396 21532
rect 39788 21586 39844 21598
rect 39788 21534 39790 21586
rect 39842 21534 39844 21586
rect 39452 21476 39508 21486
rect 39788 21476 39844 21534
rect 40124 21586 40180 21756
rect 40236 21810 40292 22204
rect 40348 22194 40404 22204
rect 40236 21758 40238 21810
rect 40290 21758 40292 21810
rect 40236 21746 40292 21758
rect 42812 22146 42868 22158
rect 42812 22094 42814 22146
rect 42866 22094 42868 22146
rect 42812 21812 42868 22094
rect 42812 21746 42868 21756
rect 40908 21700 40964 21710
rect 40348 21588 40404 21598
rect 40124 21534 40126 21586
rect 40178 21534 40180 21586
rect 40124 21522 40180 21534
rect 40236 21586 40404 21588
rect 40236 21534 40350 21586
rect 40402 21534 40404 21586
rect 40236 21532 40404 21534
rect 39452 21474 39844 21476
rect 39452 21422 39454 21474
rect 39506 21422 39844 21474
rect 39452 21420 39844 21422
rect 39452 21410 39508 21420
rect 39676 20916 39732 20926
rect 39676 20914 40180 20916
rect 39676 20862 39678 20914
rect 39730 20862 40180 20914
rect 39676 20860 40180 20862
rect 39676 20850 39732 20860
rect 40124 20802 40180 20860
rect 40124 20750 40126 20802
rect 40178 20750 40180 20802
rect 40124 20738 40180 20750
rect 39788 20692 39844 20702
rect 39788 20598 39844 20636
rect 40236 20692 40292 21532
rect 40348 21522 40404 21532
rect 40908 21586 40964 21644
rect 40908 21534 40910 21586
rect 40962 21534 40964 21586
rect 40572 20916 40628 20926
rect 40796 20916 40852 20926
rect 40572 20914 40796 20916
rect 40572 20862 40574 20914
rect 40626 20862 40796 20914
rect 40572 20860 40796 20862
rect 40572 20850 40628 20860
rect 40796 20850 40852 20860
rect 40236 20626 40292 20636
rect 40460 20802 40516 20814
rect 40460 20750 40462 20802
rect 40514 20750 40516 20802
rect 40460 20692 40516 20750
rect 39564 20578 39620 20590
rect 39564 20526 39566 20578
rect 39618 20526 39620 20578
rect 39564 20188 39620 20526
rect 39340 20178 39396 20188
rect 39452 20132 39620 20188
rect 39676 20356 39732 20366
rect 39452 18452 39508 20132
rect 39676 20130 39732 20300
rect 40236 20244 40292 20282
rect 40236 20178 40292 20188
rect 40012 20132 40068 20142
rect 39676 20078 39678 20130
rect 39730 20078 39732 20130
rect 39676 20066 39732 20078
rect 39788 20076 40012 20132
rect 39788 18562 39844 20076
rect 40012 20038 40068 20076
rect 40236 19906 40292 19918
rect 40236 19854 40238 19906
rect 40290 19854 40292 19906
rect 39900 19348 39956 19358
rect 39900 19254 39956 19292
rect 39788 18510 39790 18562
rect 39842 18510 39844 18562
rect 39788 18498 39844 18510
rect 39228 18050 39284 18060
rect 39340 18450 39508 18452
rect 39340 18398 39454 18450
rect 39506 18398 39508 18450
rect 39340 18396 39508 18398
rect 39340 18004 39396 18396
rect 39452 18386 39508 18396
rect 40012 18450 40068 18462
rect 40012 18398 40014 18450
rect 40066 18398 40068 18450
rect 39900 18340 39956 18350
rect 39900 18246 39956 18284
rect 39340 17938 39396 17948
rect 39452 18226 39508 18238
rect 39452 18174 39454 18226
rect 39506 18174 39508 18226
rect 39004 17780 39060 17790
rect 39004 17686 39060 17724
rect 38892 17614 38894 17666
rect 38946 17614 38948 17666
rect 38892 17602 38948 17614
rect 39116 17666 39172 17678
rect 39116 17614 39118 17666
rect 39170 17614 39172 17666
rect 39116 16884 39172 17614
rect 39452 17666 39508 18174
rect 40012 18228 40068 18398
rect 40236 18452 40292 19854
rect 40348 18452 40404 18462
rect 40236 18450 40404 18452
rect 40236 18398 40350 18450
rect 40402 18398 40404 18450
rect 40236 18396 40404 18398
rect 40348 18386 40404 18396
rect 40460 18452 40516 20636
rect 40684 20690 40740 20702
rect 40684 20638 40686 20690
rect 40738 20638 40740 20690
rect 40684 20580 40740 20638
rect 40684 20514 40740 20524
rect 40460 18386 40516 18396
rect 40908 19908 40964 21534
rect 41692 21474 41748 21486
rect 41692 21422 41694 21474
rect 41746 21422 41748 21474
rect 41692 20916 41748 21422
rect 41692 20850 41748 20860
rect 42364 21476 42420 21486
rect 42364 20914 42420 21420
rect 42364 20862 42366 20914
rect 42418 20862 42420 20914
rect 42364 20850 42420 20862
rect 42252 20692 42308 20702
rect 42252 20598 42308 20636
rect 41244 20578 41300 20590
rect 41244 20526 41246 20578
rect 41298 20526 41300 20578
rect 40908 18450 40964 19852
rect 41132 20020 41188 20030
rect 41020 19236 41076 19246
rect 41132 19236 41188 19964
rect 41244 19348 41300 20526
rect 42252 19908 42308 19918
rect 42252 19814 42308 19852
rect 43372 19908 43428 22430
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 43820 21476 43876 21486
rect 43820 21382 43876 21420
rect 44268 21474 44324 21486
rect 44268 21422 44270 21474
rect 44322 21422 44324 21474
rect 43372 19842 43428 19852
rect 44268 19908 44324 21422
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 41244 19282 41300 19292
rect 42812 19348 42868 19358
rect 41020 19234 41188 19236
rect 41020 19182 41022 19234
rect 41074 19182 41188 19234
rect 41020 19180 41188 19182
rect 41020 19170 41076 19180
rect 40908 18398 40910 18450
rect 40962 18398 40964 18450
rect 40908 18386 40964 18398
rect 41692 18340 41748 18350
rect 41692 18246 41748 18284
rect 40012 18162 40068 18172
rect 40572 17780 40628 17790
rect 42700 17780 42756 17790
rect 40572 17686 40628 17724
rect 42028 17778 42756 17780
rect 42028 17726 42702 17778
rect 42754 17726 42756 17778
rect 42028 17724 42756 17726
rect 39900 17668 39956 17678
rect 39452 17614 39454 17666
rect 39506 17614 39508 17666
rect 39452 17602 39508 17614
rect 39676 17612 39900 17668
rect 39676 17106 39732 17612
rect 39900 17574 39956 17612
rect 39676 17054 39678 17106
rect 39730 17054 39732 17106
rect 39676 17042 39732 17054
rect 42028 16994 42084 17724
rect 42700 17714 42756 17724
rect 42812 17668 42868 19292
rect 43484 19122 43540 19134
rect 43484 19070 43486 19122
rect 43538 19070 43540 19122
rect 43372 19010 43428 19022
rect 43372 18958 43374 19010
rect 43426 18958 43428 19010
rect 43372 18228 43428 18958
rect 43484 18452 43540 19070
rect 44268 18674 44324 19852
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 44268 18622 44270 18674
rect 44322 18622 44324 18674
rect 44268 18610 44324 18622
rect 43484 18396 43876 18452
rect 43820 18338 43876 18396
rect 43820 18286 43822 18338
rect 43874 18286 43876 18338
rect 43820 18274 43876 18286
rect 43372 18162 43428 18172
rect 42812 17444 42868 17612
rect 43148 17444 43204 17454
rect 42812 17442 43204 17444
rect 42812 17390 43150 17442
rect 43202 17390 43204 17442
rect 42812 17388 43204 17390
rect 42028 16942 42030 16994
rect 42082 16942 42084 16994
rect 42028 16930 42084 16942
rect 39116 16818 39172 16828
rect 41916 16884 41972 16894
rect 41916 16790 41972 16828
rect 39228 16772 39284 16782
rect 39228 16678 39284 16716
rect 43148 16212 43204 17388
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 43148 16146 43204 16156
rect 43820 16212 43876 16222
rect 43820 15876 43876 16156
rect 44268 15876 44324 15886
rect 43820 15874 44324 15876
rect 43820 15822 43822 15874
rect 43874 15822 44270 15874
rect 44322 15822 44324 15874
rect 43820 15820 44324 15822
rect 43820 15810 43876 15820
rect 38780 15540 38836 15550
rect 38668 15538 38836 15540
rect 38668 15486 38782 15538
rect 38834 15486 38836 15538
rect 38668 15484 38836 15486
rect 38668 15428 38724 15484
rect 38780 15474 38836 15484
rect 38668 15362 38724 15372
rect 39676 15428 39732 15438
rect 42700 15428 42756 15438
rect 39676 15426 40068 15428
rect 39676 15374 39678 15426
rect 39730 15374 40068 15426
rect 39676 15372 40068 15374
rect 39676 15362 39732 15372
rect 39452 15316 39508 15326
rect 39452 15314 39620 15316
rect 39452 15262 39454 15314
rect 39506 15262 39620 15314
rect 39452 15260 39620 15262
rect 39452 15250 39508 15260
rect 37660 15092 38276 15148
rect 37884 14644 37940 14654
rect 37884 14550 37940 14588
rect 37660 14532 37716 14542
rect 37660 13972 37716 14476
rect 37660 13970 38164 13972
rect 37660 13918 37662 13970
rect 37714 13918 38164 13970
rect 37660 13916 38164 13918
rect 37660 13906 37716 13916
rect 37212 13806 37214 13858
rect 37266 13806 37268 13858
rect 37212 13794 37268 13806
rect 38108 13858 38164 13916
rect 38108 13806 38110 13858
rect 38162 13806 38164 13858
rect 38108 13794 38164 13806
rect 38220 13970 38276 15092
rect 38220 13918 38222 13970
rect 38274 13918 38276 13970
rect 36540 13694 36542 13746
rect 36594 13694 36596 13746
rect 36540 13682 36596 13694
rect 36428 13458 36484 13468
rect 36764 13524 36820 13534
rect 36764 13522 36932 13524
rect 36764 13470 36766 13522
rect 36818 13470 36932 13522
rect 36764 13468 36932 13470
rect 36764 13458 36820 13468
rect 36540 12292 36596 12302
rect 36428 12180 36484 12190
rect 36428 12086 36484 12124
rect 36540 12178 36596 12236
rect 36540 12126 36542 12178
rect 36594 12126 36596 12178
rect 36540 12114 36596 12126
rect 36876 12068 36932 13468
rect 37772 13076 37828 13086
rect 38220 13076 38276 13918
rect 37772 13074 38276 13076
rect 37772 13022 37774 13074
rect 37826 13022 38222 13074
rect 38274 13022 38276 13074
rect 37772 13020 38276 13022
rect 37772 13010 37828 13020
rect 37996 12852 38052 13020
rect 38220 13010 38276 13020
rect 38332 15092 38500 15148
rect 38668 15204 38724 15214
rect 38668 15110 38724 15148
rect 37996 12402 38052 12796
rect 37996 12350 37998 12402
rect 38050 12350 38052 12402
rect 37996 12338 38052 12350
rect 38220 12404 38276 12414
rect 38220 12310 38276 12348
rect 37324 12290 37380 12302
rect 37324 12238 37326 12290
rect 37378 12238 37380 12290
rect 37212 12068 37268 12078
rect 36876 12066 37268 12068
rect 36876 12014 37214 12066
rect 37266 12014 37268 12066
rect 36876 12012 37268 12014
rect 37212 12002 37268 12012
rect 37100 11844 37156 11854
rect 36428 11508 36484 11518
rect 36372 11506 36484 11508
rect 36372 11454 36430 11506
rect 36482 11454 36484 11506
rect 36372 11452 36484 11454
rect 36316 11414 36372 11452
rect 36428 11442 36484 11452
rect 36204 10724 36260 10734
rect 35980 10668 36204 10724
rect 36204 10610 36260 10668
rect 36204 10558 36206 10610
rect 36258 10558 36260 10610
rect 36204 10546 36260 10558
rect 36428 10722 36484 10734
rect 36428 10670 36430 10722
rect 36482 10670 36484 10722
rect 36428 10612 36484 10670
rect 36428 10546 36484 10556
rect 36876 10722 36932 10734
rect 36876 10670 36878 10722
rect 36930 10670 36932 10722
rect 36876 10052 36932 10670
rect 36876 9986 36932 9996
rect 35644 9772 36372 9828
rect 34188 8370 34356 8372
rect 34188 8318 34190 8370
rect 34242 8318 34356 8370
rect 34188 8316 34356 8318
rect 34524 8932 34580 8942
rect 34524 8370 34580 8876
rect 34524 8318 34526 8370
rect 34578 8318 34580 8370
rect 34188 8306 34244 8316
rect 34524 8260 34580 8318
rect 34524 8194 34580 8204
rect 34636 8820 34692 8830
rect 34636 7476 34692 8764
rect 34748 8820 34804 8830
rect 34748 8818 34916 8820
rect 34748 8766 34750 8818
rect 34802 8766 34916 8818
rect 34748 8764 34916 8766
rect 34748 8754 34804 8764
rect 34860 8258 34916 8764
rect 34860 8206 34862 8258
rect 34914 8206 34916 8258
rect 34860 8194 34916 8206
rect 33180 5954 33236 5964
rect 33516 6636 34132 6692
rect 34188 7474 34692 7476
rect 34188 7422 34638 7474
rect 34690 7422 34692 7474
rect 34188 7420 34692 7422
rect 33516 5906 33572 6636
rect 33852 6020 33908 6030
rect 33852 5926 33908 5964
rect 33516 5854 33518 5906
rect 33570 5854 33572 5906
rect 33068 5796 33124 5806
rect 32956 5740 33068 5796
rect 33068 5730 33124 5740
rect 33180 5684 33236 5694
rect 33180 5590 33236 5628
rect 32508 5236 32564 5246
rect 33516 5236 33572 5854
rect 33628 5236 33684 5246
rect 33516 5234 33684 5236
rect 33516 5182 33630 5234
rect 33682 5182 33684 5234
rect 33516 5180 33684 5182
rect 32508 4562 32564 5180
rect 33628 5170 33684 5180
rect 34076 5236 34132 5246
rect 34188 5236 34244 7420
rect 34636 7410 34692 7420
rect 34300 6018 34356 6030
rect 34300 5966 34302 6018
rect 34354 5966 34356 6018
rect 34300 5796 34356 5966
rect 34300 5730 34356 5740
rect 34972 5348 35028 8988
rect 35084 8820 35140 8830
rect 35196 8820 35252 9436
rect 35756 9604 35812 9614
rect 35756 9268 35812 9548
rect 36204 9602 36260 9614
rect 36204 9550 36206 9602
rect 36258 9550 36260 9602
rect 36204 9492 36260 9550
rect 36204 9426 36260 9436
rect 35756 9202 35812 9212
rect 35308 9156 35364 9166
rect 35308 9062 35364 9100
rect 35868 9154 35924 9166
rect 35868 9102 35870 9154
rect 35922 9102 35924 9154
rect 35084 8818 35252 8820
rect 35084 8766 35086 8818
rect 35138 8766 35252 8818
rect 35084 8764 35252 8766
rect 35084 8754 35140 8764
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35868 8372 35924 9102
rect 36204 9044 36260 9054
rect 35868 8306 35924 8316
rect 35980 9042 36260 9044
rect 35980 8990 36206 9042
rect 36258 8990 36260 9042
rect 35980 8988 36260 8990
rect 35196 8036 35252 8046
rect 35196 8034 35364 8036
rect 35196 7982 35198 8034
rect 35250 7982 35364 8034
rect 35196 7980 35364 7982
rect 35196 7970 35252 7980
rect 35308 7586 35364 7980
rect 35308 7534 35310 7586
rect 35362 7534 35364 7586
rect 35308 7522 35364 7534
rect 35756 8034 35812 8046
rect 35756 7982 35758 8034
rect 35810 7982 35812 8034
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35420 6804 35476 6814
rect 35756 6804 35812 7982
rect 35476 6748 35812 6804
rect 35420 6018 35476 6748
rect 35980 6020 36036 8988
rect 36204 8978 36260 8988
rect 36092 8260 36148 8270
rect 36092 8166 36148 8204
rect 35420 5966 35422 6018
rect 35474 5966 35476 6018
rect 35420 5954 35476 5966
rect 35756 6018 36036 6020
rect 35756 5966 35982 6018
rect 36034 5966 36036 6018
rect 35756 5964 36036 5966
rect 35532 5796 35588 5806
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34132 5180 34244 5236
rect 34300 5346 35028 5348
rect 34300 5294 34974 5346
rect 35026 5294 35028 5346
rect 34300 5292 35028 5294
rect 34076 5142 34132 5180
rect 34300 5012 34356 5292
rect 34972 5282 35028 5292
rect 32508 4510 32510 4562
rect 32562 4510 32564 4562
rect 32508 4498 32564 4510
rect 33740 4956 34356 5012
rect 35532 5010 35588 5740
rect 35756 5122 35812 5964
rect 35980 5954 36036 5964
rect 36204 5908 36260 5918
rect 36316 5908 36372 9772
rect 36428 9380 36484 9390
rect 36428 9266 36484 9324
rect 36988 9380 37044 9390
rect 36428 9214 36430 9266
rect 36482 9214 36484 9266
rect 36428 9202 36484 9214
rect 36540 9268 36596 9278
rect 36540 9154 36596 9212
rect 36988 9266 37044 9324
rect 36988 9214 36990 9266
rect 37042 9214 37044 9266
rect 36988 9202 37044 9214
rect 36540 9102 36542 9154
rect 36594 9102 36596 9154
rect 36540 9090 36596 9102
rect 37100 8370 37156 11788
rect 37324 11396 37380 12238
rect 37884 12180 37940 12190
rect 37772 12178 37940 12180
rect 37772 12126 37886 12178
rect 37938 12126 37940 12178
rect 37772 12124 37940 12126
rect 37548 11956 37604 11966
rect 37548 11508 37604 11900
rect 37660 11508 37716 11518
rect 37548 11506 37716 11508
rect 37548 11454 37662 11506
rect 37714 11454 37716 11506
rect 37548 11452 37716 11454
rect 37660 11442 37716 11452
rect 37212 11340 37380 11396
rect 37212 10612 37268 11340
rect 37212 10546 37268 10556
rect 37324 11172 37380 11182
rect 37772 11172 37828 12124
rect 37884 12114 37940 12124
rect 37324 11170 37828 11172
rect 37324 11118 37326 11170
rect 37378 11118 37828 11170
rect 37324 11116 37828 11118
rect 37884 11508 37940 11518
rect 37324 9380 37380 11116
rect 37324 9314 37380 9324
rect 37660 10612 37716 10622
rect 37436 9044 37492 9054
rect 37436 8950 37492 8988
rect 37100 8318 37102 8370
rect 37154 8318 37156 8370
rect 37100 8306 37156 8318
rect 37436 8372 37492 8382
rect 37436 7362 37492 8316
rect 37660 8146 37716 10556
rect 37660 8094 37662 8146
rect 37714 8094 37716 8146
rect 37660 8082 37716 8094
rect 37884 7698 37940 11452
rect 38332 10164 38388 15092
rect 39004 15090 39060 15102
rect 39004 15038 39006 15090
rect 39058 15038 39060 15090
rect 39004 14644 39060 15038
rect 38444 13860 38500 13870
rect 38444 13766 38500 13804
rect 38892 13858 38948 13870
rect 38892 13806 38894 13858
rect 38946 13806 38948 13858
rect 38780 13746 38836 13758
rect 38780 13694 38782 13746
rect 38834 13694 38836 13746
rect 38780 13076 38836 13694
rect 38892 13524 38948 13806
rect 39004 13748 39060 14588
rect 39564 14420 39620 15260
rect 40012 14642 40068 15372
rect 40012 14590 40014 14642
rect 40066 14590 40068 14642
rect 40012 14578 40068 14590
rect 40908 15314 40964 15326
rect 40908 15262 40910 15314
rect 40962 15262 40964 15314
rect 40796 14532 40852 14542
rect 40908 14532 40964 15262
rect 41692 15202 41748 15214
rect 41692 15150 41694 15202
rect 41746 15150 41748 15202
rect 41468 14532 41524 14542
rect 40796 14530 41076 14532
rect 40796 14478 40798 14530
rect 40850 14478 41076 14530
rect 40796 14476 41076 14478
rect 40796 14466 40852 14476
rect 39564 14364 39956 14420
rect 39900 13970 39956 14364
rect 39900 13918 39902 13970
rect 39954 13918 39956 13970
rect 39900 13906 39956 13918
rect 41020 13970 41076 14476
rect 41468 14530 41636 14532
rect 41468 14478 41470 14530
rect 41522 14478 41636 14530
rect 41468 14476 41636 14478
rect 41468 14466 41524 14476
rect 41580 14084 41636 14476
rect 41692 14418 41748 15150
rect 42476 15204 42532 15214
rect 42476 14756 42532 15148
rect 42252 14754 42532 14756
rect 42252 14702 42478 14754
rect 42530 14702 42532 14754
rect 42252 14700 42532 14702
rect 41692 14366 41694 14418
rect 41746 14366 41748 14418
rect 41692 14354 41748 14366
rect 42140 14420 42196 14430
rect 42140 14326 42196 14364
rect 41580 14028 41972 14084
rect 41020 13918 41022 13970
rect 41074 13918 41076 13970
rect 39564 13748 39620 13758
rect 39004 13746 39620 13748
rect 39004 13694 39566 13746
rect 39618 13694 39620 13746
rect 39004 13692 39620 13694
rect 39564 13682 39620 13692
rect 39004 13524 39060 13534
rect 38892 13468 39004 13524
rect 39004 13458 39060 13468
rect 39788 13524 39844 13534
rect 38780 13020 39284 13076
rect 39004 12850 39060 12862
rect 39004 12798 39006 12850
rect 39058 12798 39060 12850
rect 38668 12740 38724 12750
rect 39004 12740 39060 12798
rect 39116 12852 39172 12862
rect 39116 12758 39172 12796
rect 38668 12738 39060 12740
rect 38668 12686 38670 12738
rect 38722 12686 39060 12738
rect 38668 12684 39060 12686
rect 38556 11956 38612 11966
rect 38444 11954 38612 11956
rect 38444 11902 38558 11954
rect 38610 11902 38612 11954
rect 38444 11900 38612 11902
rect 38444 10610 38500 11900
rect 38556 11890 38612 11900
rect 38668 11396 38724 12684
rect 39228 12404 39284 13020
rect 39340 12964 39396 12974
rect 39340 12870 39396 12908
rect 39676 12852 39732 12862
rect 39676 12758 39732 12796
rect 39228 12290 39284 12348
rect 39676 12292 39732 12302
rect 39228 12238 39230 12290
rect 39282 12238 39284 12290
rect 39228 12226 39284 12238
rect 39340 12236 39676 12292
rect 38892 11956 38948 11966
rect 38892 11862 38948 11900
rect 38444 10558 38446 10610
rect 38498 10558 38500 10610
rect 38444 10546 38500 10558
rect 38556 11340 38724 11396
rect 38332 10108 38500 10164
rect 37996 9604 38052 9614
rect 38332 9604 38388 9614
rect 37996 9602 38388 9604
rect 37996 9550 37998 9602
rect 38050 9550 38334 9602
rect 38386 9550 38388 9602
rect 37996 9548 38388 9550
rect 37996 9538 38052 9548
rect 37996 9268 38052 9278
rect 37996 9174 38052 9212
rect 37996 8260 38052 8270
rect 38108 8260 38164 9548
rect 38332 9538 38388 9548
rect 38444 9268 38500 10108
rect 38444 9154 38500 9212
rect 38444 9102 38446 9154
rect 38498 9102 38500 9154
rect 38444 9090 38500 9102
rect 38556 9154 38612 11340
rect 38668 10836 38724 10846
rect 38892 10836 38948 10846
rect 38668 10834 38892 10836
rect 38668 10782 38670 10834
rect 38722 10782 38892 10834
rect 38668 10780 38892 10782
rect 38668 10770 38724 10780
rect 38892 10770 38948 10780
rect 38668 9716 38724 9726
rect 39340 9716 39396 12236
rect 39676 12198 39732 12236
rect 39788 12068 39844 13468
rect 39676 12012 39844 12068
rect 39452 10052 39508 10062
rect 39452 9938 39508 9996
rect 39452 9886 39454 9938
rect 39506 9886 39508 9938
rect 39452 9874 39508 9886
rect 38668 9714 39396 9716
rect 38668 9662 38670 9714
rect 38722 9662 39396 9714
rect 38668 9660 39396 9662
rect 38668 9650 38724 9660
rect 38556 9102 38558 9154
rect 38610 9102 38612 9154
rect 38556 9044 38612 9102
rect 39340 9154 39396 9660
rect 39340 9102 39342 9154
rect 39394 9102 39396 9154
rect 39340 9090 39396 9102
rect 38556 8978 38612 8988
rect 38780 9044 38836 9054
rect 39116 9044 39172 9054
rect 38780 9042 39172 9044
rect 38780 8990 38782 9042
rect 38834 8990 39118 9042
rect 39170 8990 39172 9042
rect 38780 8988 39172 8990
rect 38780 8978 38836 8988
rect 39116 8428 39172 8988
rect 39676 8428 39732 12012
rect 41020 11508 41076 13918
rect 41916 13970 41972 14028
rect 41916 13918 41918 13970
rect 41970 13918 41972 13970
rect 41916 13906 41972 13918
rect 42140 13748 42196 13758
rect 42140 13186 42196 13692
rect 42252 13746 42308 14700
rect 42476 14690 42532 14700
rect 42700 14418 42756 15372
rect 44268 15316 44324 15820
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 44268 15222 44324 15260
rect 45276 15316 45332 15326
rect 43820 15204 43876 15214
rect 44940 15204 44996 15214
rect 43820 15110 43876 15148
rect 44380 15202 44996 15204
rect 44380 15150 44942 15202
rect 44994 15150 44996 15202
rect 44380 15148 44996 15150
rect 44380 14756 44436 15148
rect 44940 15138 44996 15148
rect 44156 14700 44436 14756
rect 43932 14532 43988 14542
rect 43932 14530 44100 14532
rect 43932 14478 43934 14530
rect 43986 14478 44100 14530
rect 43932 14476 44100 14478
rect 43932 14466 43988 14476
rect 42700 14366 42702 14418
rect 42754 14366 42756 14418
rect 42252 13694 42254 13746
rect 42306 13694 42308 13746
rect 42252 13682 42308 13694
rect 42588 13860 42644 13870
rect 42140 13134 42142 13186
rect 42194 13134 42196 13186
rect 42140 13122 42196 13134
rect 42476 12962 42532 12974
rect 42476 12910 42478 12962
rect 42530 12910 42532 12962
rect 42140 11956 42196 11966
rect 42140 11954 42308 11956
rect 42140 11902 42142 11954
rect 42194 11902 42308 11954
rect 42140 11900 42308 11902
rect 42140 11890 42196 11900
rect 40572 11506 41412 11508
rect 40572 11454 41022 11506
rect 41074 11454 41412 11506
rect 40572 11452 41412 11454
rect 40572 11394 40628 11452
rect 41020 11442 41076 11452
rect 40572 11342 40574 11394
rect 40626 11342 40628 11394
rect 40572 11330 40628 11342
rect 41356 11394 41412 11452
rect 41356 11342 41358 11394
rect 41410 11342 41412 11394
rect 39788 11282 39844 11294
rect 39788 11230 39790 11282
rect 39842 11230 39844 11282
rect 39788 10836 39844 11230
rect 39788 10770 39844 10780
rect 40012 10722 40068 10734
rect 40012 10670 40014 10722
rect 40066 10670 40068 10722
rect 39788 10612 39844 10622
rect 39788 10610 39956 10612
rect 39788 10558 39790 10610
rect 39842 10558 39956 10610
rect 39788 10556 39956 10558
rect 39788 10546 39844 10556
rect 39788 10052 39844 10062
rect 39788 9044 39844 9996
rect 39900 9716 39956 10556
rect 40012 9940 40068 10670
rect 40012 9874 40068 9884
rect 41356 10052 41412 11342
rect 42140 11282 42196 11294
rect 42140 11230 42142 11282
rect 42194 11230 42196 11282
rect 42028 10836 42084 10846
rect 42140 10836 42196 11230
rect 42028 10834 42196 10836
rect 42028 10782 42030 10834
rect 42082 10782 42196 10834
rect 42028 10780 42196 10782
rect 42028 10770 42084 10780
rect 42252 10610 42308 11900
rect 42476 11954 42532 12910
rect 42588 12292 42644 13804
rect 42700 12850 42756 14366
rect 43260 14418 43316 14430
rect 43260 14366 43262 14418
rect 43314 14366 43316 14418
rect 42812 13860 42868 13870
rect 42812 13524 42868 13804
rect 42812 13458 42868 13468
rect 43260 13524 43316 14366
rect 44044 14084 44100 14476
rect 44156 14418 44212 14700
rect 44156 14366 44158 14418
rect 44210 14366 44212 14418
rect 44156 14354 44212 14366
rect 44044 14028 44772 14084
rect 44716 13970 44772 14028
rect 44716 13918 44718 13970
rect 44770 13918 44772 13970
rect 44716 13906 44772 13918
rect 43596 13860 43652 13870
rect 43596 13766 43652 13804
rect 43260 13458 43316 13468
rect 43820 13746 43876 13758
rect 43820 13694 43822 13746
rect 43874 13694 43876 13746
rect 43820 12964 43876 13694
rect 44380 13748 44436 13758
rect 44380 13654 44436 13692
rect 45276 13634 45332 15260
rect 47068 15202 47124 15214
rect 47068 15150 47070 15202
rect 47122 15150 47124 15202
rect 47068 13748 47124 15150
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 47068 13682 47124 13692
rect 45276 13582 45278 13634
rect 45330 13582 45332 13634
rect 44604 13076 44660 13086
rect 42700 12798 42702 12850
rect 42754 12798 42756 12850
rect 42700 12786 42756 12798
rect 43260 12850 43316 12862
rect 43260 12798 43262 12850
rect 43314 12798 43316 12850
rect 42700 12292 42756 12302
rect 42588 12290 42756 12292
rect 42588 12238 42702 12290
rect 42754 12238 42756 12290
rect 42588 12236 42756 12238
rect 42700 12226 42756 12236
rect 43148 12292 43204 12302
rect 43148 12198 43204 12236
rect 42476 11902 42478 11954
rect 42530 11902 42532 11954
rect 42476 11620 42532 11902
rect 43260 11956 43316 12798
rect 43820 12178 43876 12908
rect 44044 12962 44100 12974
rect 44044 12910 44046 12962
rect 44098 12910 44100 12962
rect 44044 12404 44100 12910
rect 44268 12852 44324 12862
rect 44268 12758 44324 12796
rect 44044 12338 44100 12348
rect 43932 12292 43988 12302
rect 43932 12198 43988 12236
rect 43820 12126 43822 12178
rect 43874 12126 43876 12178
rect 43820 12114 43876 12126
rect 44604 12178 44660 13020
rect 44604 12126 44606 12178
rect 44658 12126 44660 12178
rect 43260 11890 43316 11900
rect 44604 11956 44660 12126
rect 44604 11890 44660 11900
rect 44828 12964 44884 12974
rect 45276 12964 45332 13582
rect 47740 13076 47796 13086
rect 47740 12982 47796 13020
rect 44828 12962 45332 12964
rect 44828 12910 44830 12962
rect 44882 12910 45332 12962
rect 44828 12908 45332 12910
rect 42476 11554 42532 11564
rect 44268 11620 44324 11630
rect 44268 11506 44324 11564
rect 44268 11454 44270 11506
rect 44322 11454 44324 11506
rect 44268 11442 44324 11454
rect 42252 10558 42254 10610
rect 42306 10558 42308 10610
rect 42252 10546 42308 10558
rect 44828 11172 44884 12908
rect 45612 12852 45668 12862
rect 45612 12758 45668 12796
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 44940 12404 44996 12414
rect 44940 12310 44996 12348
rect 44940 11172 44996 11182
rect 44828 11170 44996 11172
rect 44828 11118 44942 11170
rect 44994 11118 44996 11170
rect 44828 11116 44996 11118
rect 39900 9660 40292 9716
rect 40236 9266 40292 9660
rect 40236 9214 40238 9266
rect 40290 9214 40292 9266
rect 40236 9202 40292 9214
rect 39900 9044 39956 9054
rect 39788 9042 39956 9044
rect 39788 8990 39902 9042
rect 39954 8990 39956 9042
rect 39788 8988 39956 8990
rect 39900 8978 39956 8988
rect 41356 8428 41412 9996
rect 42252 10052 42308 10062
rect 41580 9940 41636 9950
rect 41580 9846 41636 9884
rect 42252 9826 42308 9996
rect 42812 10052 42868 10062
rect 42812 9938 42868 9996
rect 42812 9886 42814 9938
rect 42866 9886 42868 9938
rect 42812 9874 42868 9886
rect 42252 9774 42254 9826
rect 42306 9774 42308 9826
rect 42252 9762 42308 9774
rect 44828 9828 44884 11116
rect 44940 11106 44996 11116
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 44828 9762 44884 9772
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 39116 8372 39620 8428
rect 39676 8372 39956 8428
rect 41356 8372 41636 8428
rect 38052 8204 38164 8260
rect 38220 8260 38276 8270
rect 37996 8194 38052 8204
rect 37884 7646 37886 7698
rect 37938 7646 37940 7698
rect 37884 7634 37940 7646
rect 38220 8146 38276 8204
rect 39340 8260 39396 8270
rect 39340 8166 39396 8204
rect 38220 8094 38222 8146
rect 38274 8094 38276 8146
rect 37436 7310 37438 7362
rect 37490 7310 37492 7362
rect 37436 7298 37492 7310
rect 38220 6802 38276 8094
rect 39564 8146 39620 8372
rect 39564 8094 39566 8146
rect 39618 8094 39620 8146
rect 39564 8082 39620 8094
rect 39900 8146 39956 8372
rect 39900 8094 39902 8146
rect 39954 8094 39956 8146
rect 39004 8036 39060 8046
rect 39900 8036 39956 8094
rect 39004 8034 39508 8036
rect 39004 7982 39006 8034
rect 39058 7982 39508 8034
rect 39004 7980 39508 7982
rect 39004 7970 39060 7980
rect 38444 7588 38500 7598
rect 38444 7364 38500 7532
rect 39116 7588 39172 7598
rect 39116 7586 39396 7588
rect 39116 7534 39118 7586
rect 39170 7534 39396 7586
rect 39116 7532 39396 7534
rect 39116 7522 39172 7532
rect 38780 7474 38836 7486
rect 38780 7422 38782 7474
rect 38834 7422 38836 7474
rect 38780 7364 38836 7422
rect 38444 7308 38836 7364
rect 39340 7364 39396 7532
rect 39452 7586 39508 7980
rect 39452 7534 39454 7586
rect 39506 7534 39508 7586
rect 39452 7522 39508 7534
rect 39676 7980 39956 8036
rect 39676 7364 39732 7980
rect 39340 7308 39732 7364
rect 39788 7586 39844 7598
rect 39788 7534 39790 7586
rect 39842 7534 39844 7586
rect 38220 6750 38222 6802
rect 38274 6750 38276 6802
rect 38220 6738 38276 6750
rect 39788 6580 39844 7534
rect 41132 6692 41188 6702
rect 41580 6692 41636 8372
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 41132 6690 41636 6692
rect 41132 6638 41134 6690
rect 41186 6638 41582 6690
rect 41634 6638 41636 6690
rect 41132 6636 41636 6638
rect 39788 6514 39844 6524
rect 40348 6580 40404 6590
rect 40348 6486 40404 6524
rect 36204 5906 36372 5908
rect 36204 5854 36206 5906
rect 36258 5854 36372 5906
rect 36204 5852 36372 5854
rect 36204 5842 36260 5852
rect 36316 5236 36372 5852
rect 36540 5684 36596 5694
rect 36540 5682 36932 5684
rect 36540 5630 36542 5682
rect 36594 5630 36932 5682
rect 36540 5628 36932 5630
rect 36540 5618 36596 5628
rect 36316 5170 36372 5180
rect 35756 5070 35758 5122
rect 35810 5070 35812 5122
rect 35756 5058 35812 5070
rect 35532 4958 35534 5010
rect 35586 4958 35588 5010
rect 32060 4228 32116 4238
rect 31948 4226 32116 4228
rect 31948 4174 32062 4226
rect 32114 4174 32116 4226
rect 31948 4172 32116 4174
rect 32060 4162 32116 4172
rect 33740 4226 33796 4956
rect 35532 4946 35588 4958
rect 33740 4174 33742 4226
rect 33794 4174 33796 4226
rect 33740 4162 33796 4174
rect 34636 4898 34692 4910
rect 34636 4846 34638 4898
rect 34690 4846 34692 4898
rect 27356 3502 27358 3554
rect 27410 3502 27412 3554
rect 27356 3490 27412 3502
rect 34524 3556 34580 3566
rect 34636 3556 34692 4846
rect 36652 4564 36708 4574
rect 36652 4338 36708 4508
rect 36876 4452 36932 5628
rect 36988 5236 37044 5246
rect 36988 5142 37044 5180
rect 39900 5236 39956 5246
rect 37324 5124 37380 5134
rect 37324 4562 37380 5068
rect 39116 5124 39172 5134
rect 39116 5030 39172 5068
rect 39900 5122 39956 5180
rect 40348 5236 40404 5246
rect 40348 5142 40404 5180
rect 41132 5236 41188 6636
rect 41580 6626 41636 6636
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 41132 5170 41188 5180
rect 39900 5070 39902 5122
rect 39954 5070 39956 5122
rect 37324 4510 37326 4562
rect 37378 4510 37380 4562
rect 37324 4498 37380 4510
rect 37772 4564 37828 4574
rect 37772 4470 37828 4508
rect 39900 4564 39956 5070
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 39900 4498 39956 4508
rect 36988 4452 37044 4462
rect 36876 4450 37044 4452
rect 36876 4398 36990 4450
rect 37042 4398 37044 4450
rect 36876 4396 37044 4398
rect 36988 4386 37044 4396
rect 36652 4286 36654 4338
rect 36706 4286 36708 4338
rect 36652 4274 36708 4286
rect 34524 3554 34692 3556
rect 34524 3502 34526 3554
rect 34578 3502 34692 3554
rect 34524 3500 34692 3502
rect 34748 4228 34804 4238
rect 34524 3490 34580 3500
rect 27020 3390 27022 3442
rect 27074 3390 27076 3442
rect 27020 3378 27076 3390
rect 34748 3442 34804 4172
rect 35868 4228 35924 4238
rect 35868 4134 35924 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34748 3390 34750 3442
rect 34802 3390 34804 3442
rect 34748 3378 34804 3390
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
<< via2 >>
rect 1596 53788 1652 53844
rect 2380 53506 2436 53508
rect 2380 53454 2382 53506
rect 2382 53454 2434 53506
rect 2434 53454 2436 53506
rect 2380 53452 2436 53454
rect 3500 54236 3556 54292
rect 3164 53452 3220 53508
rect 2492 52668 2548 52724
rect 4620 56306 4676 56308
rect 4620 56254 4622 56306
rect 4622 56254 4674 56306
rect 4674 56254 4676 56306
rect 4620 56252 4676 56254
rect 5516 56306 5572 56308
rect 5516 56254 5518 56306
rect 5518 56254 5570 56306
rect 5570 56254 5572 56306
rect 5516 56252 5572 56254
rect 5852 56194 5908 56196
rect 5852 56142 5854 56194
rect 5854 56142 5906 56194
rect 5906 56142 5908 56194
rect 5852 56140 5908 56142
rect 9100 56140 9156 56196
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4060 53788 4116 53844
rect 3836 53730 3892 53732
rect 3836 53678 3838 53730
rect 3838 53678 3890 53730
rect 3890 53678 3892 53730
rect 3836 53676 3892 53678
rect 5516 54290 5572 54292
rect 5516 54238 5518 54290
rect 5518 54238 5570 54290
rect 5570 54238 5572 54290
rect 5516 54236 5572 54238
rect 4844 53676 4900 53732
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 3724 52332 3780 52388
rect 4620 52108 4676 52164
rect 6076 53058 6132 53060
rect 6076 53006 6078 53058
rect 6078 53006 6130 53058
rect 6130 53006 6132 53058
rect 6076 53004 6132 53006
rect 5180 52834 5236 52836
rect 5180 52782 5182 52834
rect 5182 52782 5234 52834
rect 5234 52782 5236 52834
rect 5180 52780 5236 52782
rect 6972 54290 7028 54292
rect 6972 54238 6974 54290
rect 6974 54238 7026 54290
rect 7026 54238 7028 54290
rect 6972 54236 7028 54238
rect 6300 52892 6356 52948
rect 6188 52780 6244 52836
rect 4844 52220 4900 52276
rect 5180 52332 5236 52388
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 2044 50034 2100 50036
rect 2044 49982 2046 50034
rect 2046 49982 2098 50034
rect 2098 49982 2100 50034
rect 2044 49980 2100 49982
rect 2716 49980 2772 50036
rect 3500 49810 3556 49812
rect 3500 49758 3502 49810
rect 3502 49758 3554 49810
rect 3554 49758 3556 49810
rect 3500 49756 3556 49758
rect 4620 49756 4676 49812
rect 5516 52722 5572 52724
rect 5516 52670 5518 52722
rect 5518 52670 5570 52722
rect 5570 52670 5572 52722
rect 5516 52668 5572 52670
rect 5740 52332 5796 52388
rect 5628 52220 5684 52276
rect 5852 52162 5908 52164
rect 5852 52110 5854 52162
rect 5854 52110 5906 52162
rect 5906 52110 5908 52162
rect 5852 52108 5908 52110
rect 5404 51324 5460 51380
rect 2716 49250 2772 49252
rect 2716 49198 2718 49250
rect 2718 49198 2770 49250
rect 2770 49198 2772 49250
rect 2716 49196 2772 49198
rect 2940 48914 2996 48916
rect 2940 48862 2942 48914
rect 2942 48862 2994 48914
rect 2994 48862 2996 48914
rect 2940 48860 2996 48862
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 3388 48860 3444 48916
rect 3500 49196 3556 49252
rect 4732 49026 4788 49028
rect 4732 48974 4734 49026
rect 4734 48974 4786 49026
rect 4786 48974 4788 49026
rect 4732 48972 4788 48974
rect 4396 48914 4452 48916
rect 4396 48862 4398 48914
rect 4398 48862 4450 48914
rect 4450 48862 4452 48914
rect 4396 48860 4452 48862
rect 3836 48412 3892 48468
rect 5740 50428 5796 50484
rect 6076 51378 6132 51380
rect 6076 51326 6078 51378
rect 6078 51326 6130 51378
rect 6130 51326 6132 51378
rect 6076 51324 6132 51326
rect 6972 53004 7028 53060
rect 6860 52780 6916 52836
rect 7420 53004 7476 53060
rect 7308 52946 7364 52948
rect 7308 52894 7310 52946
rect 7310 52894 7362 52946
rect 7362 52894 7364 52946
rect 7308 52892 7364 52894
rect 7868 52162 7924 52164
rect 7868 52110 7870 52162
rect 7870 52110 7922 52162
rect 7922 52110 7924 52162
rect 7868 52108 7924 52110
rect 6972 51100 7028 51156
rect 5852 50092 5908 50148
rect 6860 50428 6916 50484
rect 5964 49756 6020 49812
rect 5628 48914 5684 48916
rect 5628 48862 5630 48914
rect 5630 48862 5682 48914
rect 5682 48862 5684 48914
rect 5628 48860 5684 48862
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 6300 50034 6356 50036
rect 6300 49982 6302 50034
rect 6302 49982 6354 50034
rect 6354 49982 6356 50034
rect 6300 49980 6356 49982
rect 6412 49756 6468 49812
rect 6188 49644 6244 49700
rect 5740 47570 5796 47572
rect 5740 47518 5742 47570
rect 5742 47518 5794 47570
rect 5794 47518 5796 47570
rect 5740 47516 5796 47518
rect 4956 47458 5012 47460
rect 4956 47406 4958 47458
rect 4958 47406 5010 47458
rect 5010 47406 5012 47458
rect 4956 47404 5012 47406
rect 5628 47346 5684 47348
rect 5628 47294 5630 47346
rect 5630 47294 5682 47346
rect 5682 47294 5684 47346
rect 5628 47292 5684 47294
rect 2940 47068 2996 47124
rect 4844 46620 4900 46676
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 2268 45948 2324 46004
rect 4396 45948 4452 46004
rect 5964 47458 6020 47460
rect 5964 47406 5966 47458
rect 5966 47406 6018 47458
rect 6018 47406 6020 47458
rect 5964 47404 6020 47406
rect 6636 47516 6692 47572
rect 5964 46732 6020 46788
rect 4956 46396 5012 46452
rect 5068 46114 5124 46116
rect 5068 46062 5070 46114
rect 5070 46062 5122 46114
rect 5122 46062 5124 46114
rect 5068 46060 5124 46062
rect 5740 46450 5796 46452
rect 5740 46398 5742 46450
rect 5742 46398 5794 46450
rect 5794 46398 5796 46450
rect 5740 46396 5796 46398
rect 6972 49810 7028 49812
rect 6972 49758 6974 49810
rect 6974 49758 7026 49810
rect 7026 49758 7028 49810
rect 6972 49756 7028 49758
rect 7196 49810 7252 49812
rect 7196 49758 7198 49810
rect 7198 49758 7250 49810
rect 7250 49758 7252 49810
rect 7196 49756 7252 49758
rect 7084 48972 7140 49028
rect 6972 48466 7028 48468
rect 6972 48414 6974 48466
rect 6974 48414 7026 48466
rect 7026 48414 7028 48466
rect 6972 48412 7028 48414
rect 6972 47852 7028 47908
rect 6860 46786 6916 46788
rect 6860 46734 6862 46786
rect 6862 46734 6914 46786
rect 6914 46734 6916 46786
rect 6860 46732 6916 46734
rect 6300 46674 6356 46676
rect 6300 46622 6302 46674
rect 6302 46622 6354 46674
rect 6354 46622 6356 46674
rect 6300 46620 6356 46622
rect 6076 46060 6132 46116
rect 6412 46060 6468 46116
rect 7644 50092 7700 50148
rect 8876 54236 8932 54292
rect 8876 51324 8932 51380
rect 8428 51100 8484 51156
rect 8204 49756 8260 49812
rect 7756 47964 7812 48020
rect 6972 46002 7028 46004
rect 6972 45950 6974 46002
rect 6974 45950 7026 46002
rect 7026 45950 7028 46002
rect 6972 45948 7028 45950
rect 7196 46620 7252 46676
rect 6972 45388 7028 45444
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 7644 46674 7700 46676
rect 7644 46622 7646 46674
rect 7646 46622 7698 46674
rect 7698 46622 7700 46674
rect 7644 46620 7700 46622
rect 8092 45388 8148 45444
rect 7644 45276 7700 45332
rect 8988 48972 9044 49028
rect 8876 48130 8932 48132
rect 8876 48078 8878 48130
rect 8878 48078 8930 48130
rect 8930 48078 8932 48130
rect 8876 48076 8932 48078
rect 8764 46956 8820 47012
rect 8988 47404 9044 47460
rect 8652 46732 8708 46788
rect 8428 46674 8484 46676
rect 8428 46622 8430 46674
rect 8430 46622 8482 46674
rect 8482 46622 8484 46674
rect 8428 46620 8484 46622
rect 8092 45164 8148 45220
rect 7420 44434 7476 44436
rect 7420 44382 7422 44434
rect 7422 44382 7474 44434
rect 7474 44382 7476 44434
rect 7420 44380 7476 44382
rect 7980 44380 8036 44436
rect 7308 44322 7364 44324
rect 7308 44270 7310 44322
rect 7310 44270 7362 44322
rect 7362 44270 7364 44322
rect 7308 44268 7364 44270
rect 7196 44210 7252 44212
rect 7196 44158 7198 44210
rect 7198 44158 7250 44210
rect 7250 44158 7252 44210
rect 7196 44156 7252 44158
rect 7868 43932 7924 43988
rect 7644 43708 7700 43764
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 6748 42754 6804 42756
rect 6748 42702 6750 42754
rect 6750 42702 6802 42754
rect 6802 42702 6804 42754
rect 6748 42700 6804 42702
rect 7532 42700 7588 42756
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5068 40962 5124 40964
rect 5068 40910 5070 40962
rect 5070 40910 5122 40962
rect 5122 40910 5124 40962
rect 5068 40908 5124 40910
rect 1820 40348 1876 40404
rect 4060 40402 4116 40404
rect 4060 40350 4062 40402
rect 4062 40350 4114 40402
rect 4114 40350 4116 40402
rect 4060 40348 4116 40350
rect 3276 40290 3332 40292
rect 3276 40238 3278 40290
rect 3278 40238 3330 40290
rect 3330 40238 3332 40290
rect 3276 40236 3332 40238
rect 3052 40178 3108 40180
rect 3052 40126 3054 40178
rect 3054 40126 3106 40178
rect 3106 40126 3108 40178
rect 3052 40124 3108 40126
rect 3948 40124 4004 40180
rect 3612 39228 3668 39284
rect 2940 38946 2996 38948
rect 2940 38894 2942 38946
rect 2942 38894 2994 38946
rect 2994 38894 2996 38946
rect 2940 38892 2996 38894
rect 3052 38834 3108 38836
rect 3052 38782 3054 38834
rect 3054 38782 3106 38834
rect 3106 38782 3108 38834
rect 3052 38780 3108 38782
rect 3388 38780 3444 38836
rect 2716 37884 2772 37940
rect 2380 37490 2436 37492
rect 2380 37438 2382 37490
rect 2382 37438 2434 37490
rect 2434 37438 2436 37490
rect 2380 37436 2436 37438
rect 2492 36988 2548 37044
rect 2156 35980 2212 36036
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 6860 41858 6916 41860
rect 6860 41806 6862 41858
rect 6862 41806 6914 41858
rect 6914 41806 6916 41858
rect 6860 41804 6916 41806
rect 6076 40908 6132 40964
rect 5068 40348 5124 40404
rect 7420 40348 7476 40404
rect 7868 40796 7924 40852
rect 4844 39676 4900 39732
rect 5740 39730 5796 39732
rect 5740 39678 5742 39730
rect 5742 39678 5794 39730
rect 5794 39678 5796 39730
rect 5740 39676 5796 39678
rect 6076 39618 6132 39620
rect 6076 39566 6078 39618
rect 6078 39566 6130 39618
rect 6130 39566 6132 39618
rect 6076 39564 6132 39566
rect 4060 39452 4116 39508
rect 3836 38892 3892 38948
rect 3724 38834 3780 38836
rect 3724 38782 3726 38834
rect 3726 38782 3778 38834
rect 3778 38782 3780 38834
rect 3724 38780 3780 38782
rect 5628 39506 5684 39508
rect 5628 39454 5630 39506
rect 5630 39454 5682 39506
rect 5682 39454 5684 39506
rect 5628 39452 5684 39454
rect 4284 38892 4340 38948
rect 6412 39228 6468 39284
rect 5180 38892 5236 38948
rect 4732 38834 4788 38836
rect 4732 38782 4734 38834
rect 4734 38782 4786 38834
rect 4786 38782 4788 38834
rect 4732 38780 4788 38782
rect 4620 38556 4676 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 3948 37938 4004 37940
rect 3948 37886 3950 37938
rect 3950 37886 4002 37938
rect 4002 37886 4004 37938
rect 3948 37884 4004 37886
rect 4844 38332 4900 38388
rect 3724 37826 3780 37828
rect 3724 37774 3726 37826
rect 3726 37774 3778 37826
rect 3778 37774 3780 37826
rect 3724 37772 3780 37774
rect 3500 37436 3556 37492
rect 3724 37212 3780 37268
rect 3052 37100 3108 37156
rect 4620 37266 4676 37268
rect 4620 37214 4622 37266
rect 4622 37214 4674 37266
rect 4674 37214 4676 37266
rect 4620 37212 4676 37214
rect 5068 37826 5124 37828
rect 5068 37774 5070 37826
rect 5070 37774 5122 37826
rect 5122 37774 5124 37826
rect 5068 37772 5124 37774
rect 5404 38610 5460 38612
rect 5404 38558 5406 38610
rect 5406 38558 5458 38610
rect 5458 38558 5460 38610
rect 5404 38556 5460 38558
rect 5740 38610 5796 38612
rect 5740 38558 5742 38610
rect 5742 38558 5794 38610
rect 5794 38558 5796 38610
rect 5740 38556 5796 38558
rect 5180 37266 5236 37268
rect 5180 37214 5182 37266
rect 5182 37214 5234 37266
rect 5234 37214 5236 37266
rect 5180 37212 5236 37214
rect 5852 37212 5908 37268
rect 6300 38556 6356 38612
rect 6076 37100 6132 37156
rect 3948 37042 4004 37044
rect 3948 36990 3950 37042
rect 3950 36990 4002 37042
rect 4002 36990 4004 37042
rect 3948 36988 4004 36990
rect 3052 35980 3108 36036
rect 3948 35586 4004 35588
rect 3948 35534 3950 35586
rect 3950 35534 4002 35586
rect 4002 35534 4004 35586
rect 3948 35532 4004 35534
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 5068 36988 5124 37044
rect 5292 36652 5348 36708
rect 4620 36316 4676 36372
rect 4956 36370 5012 36372
rect 4956 36318 4958 36370
rect 4958 36318 5010 36370
rect 5010 36318 5012 36370
rect 4956 36316 5012 36318
rect 5292 35980 5348 36036
rect 5740 36428 5796 36484
rect 4284 35532 4340 35588
rect 6076 36428 6132 36484
rect 6188 37324 6244 37380
rect 6300 37100 6356 37156
rect 6188 36988 6244 37044
rect 6860 38556 6916 38612
rect 7084 39676 7140 39732
rect 6412 36652 6468 36708
rect 5964 36204 6020 36260
rect 5404 35420 5460 35476
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4620 35084 4676 35140
rect 1820 34972 1876 35028
rect 3276 34972 3332 35028
rect 2940 33852 2996 33908
rect 4844 35026 4900 35028
rect 4844 34974 4846 35026
rect 4846 34974 4898 35026
rect 4898 34974 4900 35026
rect 4844 34972 4900 34974
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5292 34636 5348 34692
rect 5068 34524 5124 34580
rect 6748 35644 6804 35700
rect 6076 35308 6132 35364
rect 6076 34860 6132 34916
rect 5964 34076 6020 34132
rect 5068 33852 5124 33908
rect 4844 32732 4900 32788
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 6748 34914 6804 34916
rect 6748 34862 6750 34914
rect 6750 34862 6802 34914
rect 6802 34862 6804 34914
rect 6748 34860 6804 34862
rect 7196 39564 7252 39620
rect 7308 36316 7364 36372
rect 7196 34914 7252 34916
rect 7196 34862 7198 34914
rect 7198 34862 7250 34914
rect 7250 34862 7252 34914
rect 7196 34860 7252 34862
rect 6972 34802 7028 34804
rect 6972 34750 6974 34802
rect 6974 34750 7026 34802
rect 7026 34750 7028 34802
rect 6972 34748 7028 34750
rect 8764 45388 8820 45444
rect 8988 45724 9044 45780
rect 9884 54236 9940 54292
rect 9996 54572 10052 54628
rect 14364 56306 14420 56308
rect 14364 56254 14366 56306
rect 14366 56254 14418 56306
rect 14418 56254 14420 56306
rect 14364 56252 14420 56254
rect 15036 56194 15092 56196
rect 15036 56142 15038 56194
rect 15038 56142 15090 56194
rect 15090 56142 15092 56194
rect 15036 56140 15092 56142
rect 13916 55970 13972 55972
rect 13916 55918 13918 55970
rect 13918 55918 13970 55970
rect 13970 55918 13972 55970
rect 13916 55916 13972 55918
rect 14812 55356 14868 55412
rect 15372 56140 15428 56196
rect 15372 55468 15428 55524
rect 15932 56082 15988 56084
rect 15932 56030 15934 56082
rect 15934 56030 15986 56082
rect 15986 56030 15988 56082
rect 15932 56028 15988 56030
rect 16604 56252 16660 56308
rect 16156 55916 16212 55972
rect 16492 55580 16548 55636
rect 16716 55916 16772 55972
rect 16380 55468 16436 55524
rect 15932 55298 15988 55300
rect 15932 55246 15934 55298
rect 15934 55246 15986 55298
rect 15986 55246 15988 55298
rect 15932 55244 15988 55246
rect 16828 55468 16884 55524
rect 16940 55356 16996 55412
rect 17500 55244 17556 55300
rect 15596 54684 15652 54740
rect 16604 54684 16660 54740
rect 10668 54626 10724 54628
rect 10668 54574 10670 54626
rect 10670 54574 10722 54626
rect 10722 54574 10724 54626
rect 10668 54572 10724 54574
rect 11452 54572 11508 54628
rect 17612 55020 17668 55076
rect 16380 54514 16436 54516
rect 16380 54462 16382 54514
rect 16382 54462 16434 54514
rect 16434 54462 16436 54514
rect 16380 54460 16436 54462
rect 12796 53564 12852 53620
rect 13580 53564 13636 53620
rect 14252 53116 14308 53172
rect 15148 53564 15204 53620
rect 9660 51548 9716 51604
rect 9548 49980 9604 50036
rect 11004 51602 11060 51604
rect 11004 51550 11006 51602
rect 11006 51550 11058 51602
rect 11058 51550 11060 51602
rect 11004 51548 11060 51550
rect 11676 52332 11732 52388
rect 11340 51548 11396 51604
rect 11452 51996 11508 52052
rect 9772 51324 9828 51380
rect 10220 51378 10276 51380
rect 10220 51326 10222 51378
rect 10222 51326 10274 51378
rect 10274 51326 10276 51378
rect 10220 51324 10276 51326
rect 11340 51324 11396 51380
rect 11900 52050 11956 52052
rect 11900 51998 11902 52050
rect 11902 51998 11954 52050
rect 11954 51998 11956 52050
rect 11900 51996 11956 51998
rect 10444 50764 10500 50820
rect 11340 50764 11396 50820
rect 9884 50652 9940 50708
rect 11228 50652 11284 50708
rect 10892 50594 10948 50596
rect 10892 50542 10894 50594
rect 10894 50542 10946 50594
rect 10946 50542 10948 50594
rect 10892 50540 10948 50542
rect 10108 50482 10164 50484
rect 10108 50430 10110 50482
rect 10110 50430 10162 50482
rect 10162 50430 10164 50482
rect 10108 50428 10164 50430
rect 10780 50482 10836 50484
rect 10780 50430 10782 50482
rect 10782 50430 10834 50482
rect 10834 50430 10836 50482
rect 10780 50428 10836 50430
rect 11452 50428 11508 50484
rect 10108 49084 10164 49140
rect 9100 45612 9156 45668
rect 9548 48018 9604 48020
rect 9548 47966 9550 48018
rect 9550 47966 9602 48018
rect 9602 47966 9604 48018
rect 9548 47964 9604 47966
rect 9660 47852 9716 47908
rect 9996 49026 10052 49028
rect 9996 48974 9998 49026
rect 9998 48974 10050 49026
rect 10050 48974 10052 49026
rect 9996 48972 10052 48974
rect 9884 48130 9940 48132
rect 9884 48078 9886 48130
rect 9886 48078 9938 48130
rect 9938 48078 9940 48130
rect 9884 48076 9940 48078
rect 10668 49756 10724 49812
rect 10332 49138 10388 49140
rect 10332 49086 10334 49138
rect 10334 49086 10386 49138
rect 10386 49086 10388 49138
rect 10332 49084 10388 49086
rect 10108 47852 10164 47908
rect 9884 46956 9940 47012
rect 10220 46674 10276 46676
rect 10220 46622 10222 46674
rect 10222 46622 10274 46674
rect 10274 46622 10276 46674
rect 10220 46620 10276 46622
rect 9660 45778 9716 45780
rect 9660 45726 9662 45778
rect 9662 45726 9714 45778
rect 9714 45726 9716 45778
rect 9660 45724 9716 45726
rect 9660 45388 9716 45444
rect 9436 43932 9492 43988
rect 9548 44268 9604 44324
rect 10220 45218 10276 45220
rect 10220 45166 10222 45218
rect 10222 45166 10274 45218
rect 10274 45166 10276 45218
rect 10220 45164 10276 45166
rect 9772 44156 9828 44212
rect 10556 46844 10612 46900
rect 11564 49810 11620 49812
rect 11564 49758 11566 49810
rect 11566 49758 11618 49810
rect 11618 49758 11620 49810
rect 11564 49756 11620 49758
rect 11228 49532 11284 49588
rect 11228 48972 11284 49028
rect 12348 51548 12404 51604
rect 11900 50594 11956 50596
rect 11900 50542 11902 50594
rect 11902 50542 11954 50594
rect 11954 50542 11956 50594
rect 11900 50540 11956 50542
rect 12572 50652 12628 50708
rect 12460 50482 12516 50484
rect 12460 50430 12462 50482
rect 12462 50430 12514 50482
rect 12514 50430 12516 50482
rect 12460 50428 12516 50430
rect 11900 49810 11956 49812
rect 11900 49758 11902 49810
rect 11902 49758 11954 49810
rect 11954 49758 11956 49810
rect 11900 49756 11956 49758
rect 12460 49810 12516 49812
rect 12460 49758 12462 49810
rect 12462 49758 12514 49810
rect 12514 49758 12516 49810
rect 12460 49756 12516 49758
rect 12348 49644 12404 49700
rect 11788 49586 11844 49588
rect 11788 49534 11790 49586
rect 11790 49534 11842 49586
rect 11842 49534 11844 49586
rect 11788 49532 11844 49534
rect 11676 49196 11732 49252
rect 12012 49308 12068 49364
rect 11116 48860 11172 48916
rect 11564 48300 11620 48356
rect 12684 49644 12740 49700
rect 11900 48914 11956 48916
rect 11900 48862 11902 48914
rect 11902 48862 11954 48914
rect 11954 48862 11956 48914
rect 11900 48860 11956 48862
rect 13132 51378 13188 51380
rect 13132 51326 13134 51378
rect 13134 51326 13186 51378
rect 13186 51326 13188 51378
rect 13132 51324 13188 51326
rect 17836 55244 17892 55300
rect 15820 53564 15876 53620
rect 18060 55580 18116 55636
rect 18060 55020 18116 55076
rect 18172 53788 18228 53844
rect 16380 53452 16436 53508
rect 16044 53170 16100 53172
rect 16044 53118 16046 53170
rect 16046 53118 16098 53170
rect 16098 53118 16100 53170
rect 16044 53116 16100 53118
rect 15820 52332 15876 52388
rect 16604 52946 16660 52948
rect 16604 52894 16606 52946
rect 16606 52894 16658 52946
rect 16658 52894 16660 52946
rect 16604 52892 16660 52894
rect 17052 53506 17108 53508
rect 17052 53454 17054 53506
rect 17054 53454 17106 53506
rect 17106 53454 17108 53506
rect 17052 53452 17108 53454
rect 16268 52332 16324 52388
rect 15484 52050 15540 52052
rect 15484 51998 15486 52050
rect 15486 51998 15538 52050
rect 15538 51998 15540 52050
rect 15484 51996 15540 51998
rect 15148 51324 15204 51380
rect 17052 52162 17108 52164
rect 17052 52110 17054 52162
rect 17054 52110 17106 52162
rect 17106 52110 17108 52162
rect 17052 52108 17108 52110
rect 16604 51996 16660 52052
rect 16940 51884 16996 51940
rect 15932 51324 15988 51380
rect 16156 51324 16212 51380
rect 15932 50706 15988 50708
rect 15932 50654 15934 50706
rect 15934 50654 15986 50706
rect 15986 50654 15988 50706
rect 15932 50652 15988 50654
rect 16716 51490 16772 51492
rect 16716 51438 16718 51490
rect 16718 51438 16770 51490
rect 16770 51438 16772 51490
rect 16716 51436 16772 51438
rect 19068 55970 19124 55972
rect 19068 55918 19070 55970
rect 19070 55918 19122 55970
rect 19122 55918 19124 55970
rect 19068 55916 19124 55918
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 19852 55916 19908 55972
rect 18844 55356 18900 55412
rect 18396 55298 18452 55300
rect 18396 55246 18398 55298
rect 18398 55246 18450 55298
rect 18450 55246 18452 55298
rect 18396 55244 18452 55246
rect 18844 55186 18900 55188
rect 18844 55134 18846 55186
rect 18846 55134 18898 55186
rect 18898 55134 18900 55186
rect 18844 55132 18900 55134
rect 18956 55020 19012 55076
rect 18732 54460 18788 54516
rect 19292 55356 19348 55412
rect 19628 55244 19684 55300
rect 19964 55356 20020 55412
rect 20524 55356 20580 55412
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19404 54572 19460 54628
rect 19292 54514 19348 54516
rect 19292 54462 19294 54514
rect 19294 54462 19346 54514
rect 19346 54462 19348 54514
rect 19292 54460 19348 54462
rect 19404 54402 19460 54404
rect 19404 54350 19406 54402
rect 19406 54350 19458 54402
rect 19458 54350 19460 54402
rect 19404 54348 19460 54350
rect 18844 53842 18900 53844
rect 18844 53790 18846 53842
rect 18846 53790 18898 53842
rect 18898 53790 18900 53842
rect 18844 53788 18900 53790
rect 20300 54460 20356 54516
rect 19852 53788 19908 53844
rect 20748 54626 20804 54628
rect 20748 54574 20750 54626
rect 20750 54574 20802 54626
rect 20802 54574 20804 54626
rect 20748 54572 20804 54574
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 17500 52332 17556 52388
rect 17612 52108 17668 52164
rect 16716 50428 16772 50484
rect 13916 50316 13972 50372
rect 16380 50370 16436 50372
rect 16380 50318 16382 50370
rect 16382 50318 16434 50370
rect 16434 50318 16436 50370
rect 16380 50316 16436 50318
rect 12796 49308 12852 49364
rect 12796 48860 12852 48916
rect 11004 47458 11060 47460
rect 11004 47406 11006 47458
rect 11006 47406 11058 47458
rect 11058 47406 11060 47458
rect 11004 47404 11060 47406
rect 11228 47570 11284 47572
rect 11228 47518 11230 47570
rect 11230 47518 11282 47570
rect 11282 47518 11284 47570
rect 11228 47516 11284 47518
rect 11228 47180 11284 47236
rect 10668 46732 10724 46788
rect 11676 46732 11732 46788
rect 11788 47180 11844 47236
rect 13580 48354 13636 48356
rect 13580 48302 13582 48354
rect 13582 48302 13634 48354
rect 13634 48302 13636 48354
rect 13580 48300 13636 48302
rect 15036 48300 15092 48356
rect 16044 48354 16100 48356
rect 16044 48302 16046 48354
rect 16046 48302 16098 48354
rect 16098 48302 16100 48354
rect 16044 48300 16100 48302
rect 16156 48242 16212 48244
rect 16156 48190 16158 48242
rect 16158 48190 16210 48242
rect 16210 48190 16212 48242
rect 16156 48188 16212 48190
rect 14812 47516 14868 47572
rect 12572 47458 12628 47460
rect 12572 47406 12574 47458
rect 12574 47406 12626 47458
rect 12626 47406 12628 47458
rect 12572 47404 12628 47406
rect 11340 46060 11396 46116
rect 10556 45276 10612 45332
rect 11900 46844 11956 46900
rect 12796 46844 12852 46900
rect 14028 46786 14084 46788
rect 14028 46734 14030 46786
rect 14030 46734 14082 46786
rect 14082 46734 14084 46786
rect 14028 46732 14084 46734
rect 16604 49420 16660 49476
rect 16828 49810 16884 49812
rect 16828 49758 16830 49810
rect 16830 49758 16882 49810
rect 16882 49758 16884 49810
rect 16828 49756 16884 49758
rect 17948 52050 18004 52052
rect 17948 51998 17950 52050
rect 17950 51998 18002 52050
rect 18002 51998 18004 52050
rect 17948 51996 18004 51998
rect 18060 51436 18116 51492
rect 18732 52834 18788 52836
rect 18732 52782 18734 52834
rect 18734 52782 18786 52834
rect 18786 52782 18788 52834
rect 18732 52780 18788 52782
rect 18284 52332 18340 52388
rect 18508 52274 18564 52276
rect 18508 52222 18510 52274
rect 18510 52222 18562 52274
rect 18562 52222 18564 52274
rect 18508 52220 18564 52222
rect 18396 51938 18452 51940
rect 18396 51886 18398 51938
rect 18398 51886 18450 51938
rect 18450 51886 18452 51938
rect 18396 51884 18452 51886
rect 17388 50482 17444 50484
rect 17388 50430 17390 50482
rect 17390 50430 17442 50482
rect 17442 50430 17444 50482
rect 17388 50428 17444 50430
rect 18284 51548 18340 51604
rect 19628 52892 19684 52948
rect 19404 52780 19460 52836
rect 19740 52162 19796 52164
rect 19740 52110 19742 52162
rect 19742 52110 19794 52162
rect 19794 52110 19796 52162
rect 19740 52108 19796 52110
rect 19292 51548 19348 51604
rect 18172 50706 18228 50708
rect 18172 50654 18174 50706
rect 18174 50654 18226 50706
rect 18226 50654 18228 50706
rect 18172 50652 18228 50654
rect 19180 51212 19236 51268
rect 18956 50594 19012 50596
rect 18956 50542 18958 50594
rect 18958 50542 19010 50594
rect 19010 50542 19012 50594
rect 18956 50540 19012 50542
rect 18844 50482 18900 50484
rect 18844 50430 18846 50482
rect 18846 50430 18898 50482
rect 18898 50430 18900 50482
rect 18844 50428 18900 50430
rect 17724 49810 17780 49812
rect 17724 49758 17726 49810
rect 17726 49758 17778 49810
rect 17778 49758 17780 49810
rect 17724 49756 17780 49758
rect 17052 49532 17108 49588
rect 17164 49420 17220 49476
rect 17948 49420 18004 49476
rect 17276 48860 17332 48916
rect 15260 47516 15316 47572
rect 16604 47516 16660 47572
rect 16268 47404 16324 47460
rect 17836 48802 17892 48804
rect 17836 48750 17838 48802
rect 17838 48750 17890 48802
rect 17890 48750 17892 48802
rect 17836 48748 17892 48750
rect 17500 48188 17556 48244
rect 13356 46060 13412 46116
rect 13244 45612 13300 45668
rect 12796 45276 12852 45332
rect 12124 44434 12180 44436
rect 12124 44382 12126 44434
rect 12126 44382 12178 44434
rect 12178 44382 12180 44434
rect 12124 44380 12180 44382
rect 17948 46674 18004 46676
rect 17948 46622 17950 46674
rect 17950 46622 18002 46674
rect 18002 46622 18004 46674
rect 17948 46620 18004 46622
rect 16940 46002 16996 46004
rect 16940 45950 16942 46002
rect 16942 45950 16994 46002
rect 16994 45950 16996 46002
rect 16940 45948 16996 45950
rect 17612 46002 17668 46004
rect 17612 45950 17614 46002
rect 17614 45950 17666 46002
rect 17666 45950 17668 46002
rect 17612 45948 17668 45950
rect 17836 46002 17892 46004
rect 17836 45950 17838 46002
rect 17838 45950 17890 46002
rect 17890 45950 17892 46002
rect 17836 45948 17892 45950
rect 14812 45778 14868 45780
rect 14812 45726 14814 45778
rect 14814 45726 14866 45778
rect 14866 45726 14868 45778
rect 14812 45724 14868 45726
rect 15372 45724 15428 45780
rect 14140 45106 14196 45108
rect 14140 45054 14142 45106
rect 14142 45054 14194 45106
rect 14194 45054 14196 45106
rect 14140 45052 14196 45054
rect 14588 45106 14644 45108
rect 14588 45054 14590 45106
rect 14590 45054 14642 45106
rect 14642 45054 14644 45106
rect 14588 45052 14644 45054
rect 13244 44380 13300 44436
rect 11676 44044 11732 44100
rect 10556 43932 10612 43988
rect 10108 43762 10164 43764
rect 10108 43710 10110 43762
rect 10110 43710 10162 43762
rect 10162 43710 10164 43762
rect 10108 43708 10164 43710
rect 11452 43650 11508 43652
rect 11452 43598 11454 43650
rect 11454 43598 11506 43650
rect 11506 43598 11508 43650
rect 11452 43596 11508 43598
rect 8988 41916 9044 41972
rect 8876 41804 8932 41860
rect 8092 40908 8148 40964
rect 9996 42530 10052 42532
rect 9996 42478 9998 42530
rect 9998 42478 10050 42530
rect 10050 42478 10052 42530
rect 9996 42476 10052 42478
rect 9212 40962 9268 40964
rect 9212 40910 9214 40962
rect 9214 40910 9266 40962
rect 9266 40910 9268 40962
rect 9212 40908 9268 40910
rect 10780 42530 10836 42532
rect 10780 42478 10782 42530
rect 10782 42478 10834 42530
rect 10834 42478 10836 42530
rect 10780 42476 10836 42478
rect 12348 44044 12404 44100
rect 9996 40908 10052 40964
rect 10108 41916 10164 41972
rect 8316 40348 8372 40404
rect 7980 39788 8036 39844
rect 8316 39618 8372 39620
rect 8316 39566 8318 39618
rect 8318 39566 8370 39618
rect 8370 39566 8372 39618
rect 8316 39564 8372 39566
rect 9772 40290 9828 40292
rect 9772 40238 9774 40290
rect 9774 40238 9826 40290
rect 9826 40238 9828 40290
rect 9772 40236 9828 40238
rect 8764 39676 8820 39732
rect 9660 39618 9716 39620
rect 9660 39566 9662 39618
rect 9662 39566 9714 39618
rect 9714 39566 9716 39618
rect 9660 39564 9716 39566
rect 10108 40514 10164 40516
rect 10108 40462 10110 40514
rect 10110 40462 10162 40514
rect 10162 40462 10164 40514
rect 10108 40460 10164 40462
rect 10220 40402 10276 40404
rect 10220 40350 10222 40402
rect 10222 40350 10274 40402
rect 10274 40350 10276 40402
rect 10220 40348 10276 40350
rect 10556 41970 10612 41972
rect 10556 41918 10558 41970
rect 10558 41918 10610 41970
rect 10610 41918 10612 41970
rect 10556 41916 10612 41918
rect 11116 42476 11172 42532
rect 11788 42530 11844 42532
rect 11788 42478 11790 42530
rect 11790 42478 11842 42530
rect 11842 42478 11844 42530
rect 11788 42476 11844 42478
rect 12236 42476 12292 42532
rect 10668 40572 10724 40628
rect 11452 40572 11508 40628
rect 10332 40124 10388 40180
rect 10892 40348 10948 40404
rect 10108 39842 10164 39844
rect 10108 39790 10110 39842
rect 10110 39790 10162 39842
rect 10162 39790 10164 39842
rect 10108 39788 10164 39790
rect 7644 38668 7700 38724
rect 9212 39394 9268 39396
rect 9212 39342 9214 39394
rect 9214 39342 9266 39394
rect 9266 39342 9268 39394
rect 9212 39340 9268 39342
rect 8764 38834 8820 38836
rect 8764 38782 8766 38834
rect 8766 38782 8818 38834
rect 8818 38782 8820 38834
rect 8764 38780 8820 38782
rect 7532 38556 7588 38612
rect 8316 38332 8372 38388
rect 7532 37996 7588 38052
rect 7756 37378 7812 37380
rect 7756 37326 7758 37378
rect 7758 37326 7810 37378
rect 7810 37326 7812 37378
rect 7756 37324 7812 37326
rect 8428 37772 8484 37828
rect 9212 37826 9268 37828
rect 9212 37774 9214 37826
rect 9214 37774 9266 37826
rect 9266 37774 9268 37826
rect 9212 37772 9268 37774
rect 8316 36706 8372 36708
rect 8316 36654 8318 36706
rect 8318 36654 8370 36706
rect 8370 36654 8372 36706
rect 8316 36652 8372 36654
rect 8204 36540 8260 36596
rect 7532 36370 7588 36372
rect 7532 36318 7534 36370
rect 7534 36318 7586 36370
rect 7586 36318 7588 36370
rect 7532 36316 7588 36318
rect 8204 36258 8260 36260
rect 8204 36206 8206 36258
rect 8206 36206 8258 36258
rect 8258 36206 8260 36258
rect 8204 36204 8260 36206
rect 7420 35474 7476 35476
rect 7420 35422 7422 35474
rect 7422 35422 7474 35474
rect 7474 35422 7476 35474
rect 7420 35420 7476 35422
rect 7420 34690 7476 34692
rect 7420 34638 7422 34690
rect 7422 34638 7474 34690
rect 7474 34638 7476 34690
rect 7420 34636 7476 34638
rect 7756 34860 7812 34916
rect 7868 34802 7924 34804
rect 7868 34750 7870 34802
rect 7870 34750 7922 34802
rect 7922 34750 7924 34802
rect 7868 34748 7924 34750
rect 8876 36428 8932 36484
rect 9100 36764 9156 36820
rect 8652 35586 8708 35588
rect 8652 35534 8654 35586
rect 8654 35534 8706 35586
rect 8706 35534 8708 35586
rect 8652 35532 8708 35534
rect 8652 35196 8708 35252
rect 8428 34914 8484 34916
rect 8428 34862 8430 34914
rect 8430 34862 8482 34914
rect 8482 34862 8484 34914
rect 8428 34860 8484 34862
rect 9772 38220 9828 38276
rect 9884 39340 9940 39396
rect 9884 39004 9940 39060
rect 9660 38108 9716 38164
rect 9996 38834 10052 38836
rect 9996 38782 9998 38834
rect 9998 38782 10050 38834
rect 10050 38782 10052 38834
rect 9996 38780 10052 38782
rect 9660 36764 9716 36820
rect 9436 36482 9492 36484
rect 9436 36430 9438 36482
rect 9438 36430 9490 36482
rect 9490 36430 9492 36482
rect 9436 36428 9492 36430
rect 8204 34748 8260 34804
rect 9324 35532 9380 35588
rect 7196 34130 7252 34132
rect 7196 34078 7198 34130
rect 7198 34078 7250 34130
rect 7250 34078 7252 34130
rect 7196 34076 7252 34078
rect 9884 37100 9940 37156
rect 10556 39394 10612 39396
rect 10556 39342 10558 39394
rect 10558 39342 10610 39394
rect 10610 39342 10612 39394
rect 10556 39340 10612 39342
rect 10780 39228 10836 39284
rect 11116 39788 11172 39844
rect 11004 39618 11060 39620
rect 11004 39566 11006 39618
rect 11006 39566 11058 39618
rect 11058 39566 11060 39618
rect 11004 39564 11060 39566
rect 11340 39116 11396 39172
rect 10220 38946 10276 38948
rect 10220 38894 10222 38946
rect 10222 38894 10274 38946
rect 10274 38894 10276 38946
rect 10220 38892 10276 38894
rect 10444 38444 10500 38500
rect 10332 38332 10388 38388
rect 10220 38220 10276 38276
rect 10668 38332 10724 38388
rect 10668 38108 10724 38164
rect 10444 37938 10500 37940
rect 10444 37886 10446 37938
rect 10446 37886 10498 37938
rect 10498 37886 10500 37938
rect 10444 37884 10500 37886
rect 10556 37660 10612 37716
rect 10108 36652 10164 36708
rect 10108 36482 10164 36484
rect 10108 36430 10110 36482
rect 10110 36430 10162 36482
rect 10162 36430 10164 36482
rect 10108 36428 10164 36430
rect 9660 35196 9716 35252
rect 10332 35084 10388 35140
rect 9884 34972 9940 35028
rect 9996 34802 10052 34804
rect 9996 34750 9998 34802
rect 9998 34750 10050 34802
rect 10050 34750 10052 34802
rect 9996 34748 10052 34750
rect 12460 40684 12516 40740
rect 11564 40460 11620 40516
rect 12908 40460 12964 40516
rect 12012 40236 12068 40292
rect 11900 39340 11956 39396
rect 11564 39058 11620 39060
rect 11564 39006 11566 39058
rect 11566 39006 11618 39058
rect 11618 39006 11620 39058
rect 11564 39004 11620 39006
rect 12012 38892 12068 38948
rect 12348 39676 12404 39732
rect 12796 39564 12852 39620
rect 12684 39116 12740 39172
rect 12460 38780 12516 38836
rect 11564 38444 11620 38500
rect 11116 37660 11172 37716
rect 10780 36428 10836 36484
rect 10668 36316 10724 36372
rect 10892 35868 10948 35924
rect 11340 37042 11396 37044
rect 11340 36990 11342 37042
rect 11342 36990 11394 37042
rect 11394 36990 11396 37042
rect 11340 36988 11396 36990
rect 11564 36652 11620 36708
rect 11228 36092 11284 36148
rect 11564 35868 11620 35924
rect 11788 37100 11844 37156
rect 11676 36428 11732 36484
rect 12124 36540 12180 36596
rect 12124 36204 12180 36260
rect 11116 35084 11172 35140
rect 11452 35196 11508 35252
rect 9884 33964 9940 34020
rect 10444 34412 10500 34468
rect 10892 34802 10948 34804
rect 10892 34750 10894 34802
rect 10894 34750 10946 34802
rect 10946 34750 10948 34802
rect 10892 34748 10948 34750
rect 12572 38610 12628 38612
rect 12572 38558 12574 38610
rect 12574 38558 12626 38610
rect 12626 38558 12628 38610
rect 12572 38556 12628 38558
rect 12796 38946 12852 38948
rect 12796 38894 12798 38946
rect 12798 38894 12850 38946
rect 12850 38894 12852 38946
rect 12796 38892 12852 38894
rect 12796 38220 12852 38276
rect 13132 39340 13188 39396
rect 13020 38668 13076 38724
rect 12908 38108 12964 38164
rect 13020 37324 13076 37380
rect 14812 44434 14868 44436
rect 14812 44382 14814 44434
rect 14814 44382 14866 44434
rect 14866 44382 14868 44434
rect 14812 44380 14868 44382
rect 15148 44380 15204 44436
rect 14364 41970 14420 41972
rect 14364 41918 14366 41970
rect 14366 41918 14418 41970
rect 14418 41918 14420 41970
rect 14364 41916 14420 41918
rect 14252 41692 14308 41748
rect 13468 40626 13524 40628
rect 13468 40574 13470 40626
rect 13470 40574 13522 40626
rect 13522 40574 13524 40626
rect 13468 40572 13524 40574
rect 14812 41020 14868 41076
rect 13580 40402 13636 40404
rect 13580 40350 13582 40402
rect 13582 40350 13634 40402
rect 13634 40350 13636 40402
rect 13580 40348 13636 40350
rect 13468 40178 13524 40180
rect 13468 40126 13470 40178
rect 13470 40126 13522 40178
rect 13522 40126 13524 40178
rect 13468 40124 13524 40126
rect 13468 39788 13524 39844
rect 13580 39730 13636 39732
rect 13580 39678 13582 39730
rect 13582 39678 13634 39730
rect 13634 39678 13636 39730
rect 13580 39676 13636 39678
rect 13468 39618 13524 39620
rect 13468 39566 13470 39618
rect 13470 39566 13522 39618
rect 13522 39566 13524 39618
rect 13468 39564 13524 39566
rect 14252 40908 14308 40964
rect 15260 41186 15316 41188
rect 15260 41134 15262 41186
rect 15262 41134 15314 41186
rect 15314 41134 15316 41186
rect 15260 41132 15316 41134
rect 13580 38946 13636 38948
rect 13580 38894 13582 38946
rect 13582 38894 13634 38946
rect 13634 38894 13636 38946
rect 13580 38892 13636 38894
rect 15260 40908 15316 40964
rect 15148 40796 15204 40852
rect 14812 40626 14868 40628
rect 14812 40574 14814 40626
rect 14814 40574 14866 40626
rect 14866 40574 14868 40626
rect 14812 40572 14868 40574
rect 14588 40460 14644 40516
rect 14476 40402 14532 40404
rect 14476 40350 14478 40402
rect 14478 40350 14530 40402
rect 14530 40350 14532 40402
rect 14476 40348 14532 40350
rect 14364 38892 14420 38948
rect 13356 38668 13412 38724
rect 13468 38444 13524 38500
rect 13804 38050 13860 38052
rect 13804 37998 13806 38050
rect 13806 37998 13858 38050
rect 13858 37998 13860 38050
rect 13804 37996 13860 37998
rect 14252 38834 14308 38836
rect 14252 38782 14254 38834
rect 14254 38782 14306 38834
rect 14306 38782 14308 38834
rect 14252 38780 14308 38782
rect 15148 40236 15204 40292
rect 14924 39452 14980 39508
rect 16268 45164 16324 45220
rect 17948 45388 18004 45444
rect 17836 45164 17892 45220
rect 16716 45052 16772 45108
rect 15484 44098 15540 44100
rect 15484 44046 15486 44098
rect 15486 44046 15538 44098
rect 15538 44046 15540 44098
rect 15484 44044 15540 44046
rect 16716 43932 16772 43988
rect 17052 43596 17108 43652
rect 16716 42924 16772 42980
rect 16044 41970 16100 41972
rect 16044 41918 16046 41970
rect 16046 41918 16098 41970
rect 16098 41918 16100 41970
rect 16044 41916 16100 41918
rect 15820 41132 15876 41188
rect 16268 41186 16324 41188
rect 16268 41134 16270 41186
rect 16270 41134 16322 41186
rect 16322 41134 16324 41186
rect 16268 41132 16324 41134
rect 16044 41020 16100 41076
rect 15372 40012 15428 40068
rect 16380 41020 16436 41076
rect 16156 40796 16212 40852
rect 16044 40460 16100 40516
rect 15820 40236 15876 40292
rect 16268 40012 16324 40068
rect 15820 39618 15876 39620
rect 15820 39566 15822 39618
rect 15822 39566 15874 39618
rect 15874 39566 15876 39618
rect 15820 39564 15876 39566
rect 15932 39452 15988 39508
rect 15148 38668 15204 38724
rect 14476 38444 14532 38500
rect 13468 37884 13524 37940
rect 13468 36540 13524 36596
rect 12796 36370 12852 36372
rect 12796 36318 12798 36370
rect 12798 36318 12850 36370
rect 12850 36318 12852 36370
rect 12796 36316 12852 36318
rect 12684 35980 12740 36036
rect 11564 34748 11620 34804
rect 11004 34636 11060 34692
rect 10444 34130 10500 34132
rect 10444 34078 10446 34130
rect 10446 34078 10498 34130
rect 10498 34078 10500 34130
rect 10444 34076 10500 34078
rect 11564 34412 11620 34468
rect 11004 34130 11060 34132
rect 11004 34078 11006 34130
rect 11006 34078 11058 34130
rect 11058 34078 11060 34130
rect 11004 34076 11060 34078
rect 9324 33516 9380 33572
rect 8540 33068 8596 33124
rect 6524 32786 6580 32788
rect 6524 32734 6526 32786
rect 6526 32734 6578 32786
rect 6578 32734 6580 32786
rect 6524 32732 6580 32734
rect 6524 31836 6580 31892
rect 6748 32396 6804 32452
rect 7756 31836 7812 31892
rect 8204 31836 8260 31892
rect 7868 31276 7924 31332
rect 7308 30716 7364 30772
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 1596 29932 1652 29988
rect 8764 31948 8820 32004
rect 9100 32732 9156 32788
rect 9660 31948 9716 32004
rect 11788 34690 11844 34692
rect 11788 34638 11790 34690
rect 11790 34638 11842 34690
rect 11842 34638 11844 34690
rect 11788 34636 11844 34638
rect 12796 34076 12852 34132
rect 10892 31948 10948 32004
rect 10556 31836 10612 31892
rect 10556 31388 10612 31444
rect 10332 31218 10388 31220
rect 10332 31166 10334 31218
rect 10334 31166 10386 31218
rect 10386 31166 10388 31218
rect 10332 31164 10388 31166
rect 11116 31388 11172 31444
rect 11228 31948 11284 32004
rect 11116 30994 11172 30996
rect 11116 30942 11118 30994
rect 11118 30942 11170 30994
rect 11170 30942 11172 30994
rect 11116 30940 11172 30942
rect 8988 30828 9044 30884
rect 10220 30770 10276 30772
rect 10220 30718 10222 30770
rect 10222 30718 10274 30770
rect 10274 30718 10276 30770
rect 10220 30716 10276 30718
rect 9212 30268 9268 30324
rect 5180 29260 5236 29316
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 6188 29260 6244 29316
rect 6748 29260 6804 29316
rect 6524 29036 6580 29092
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3500 26290 3556 26292
rect 3500 26238 3502 26290
rect 3502 26238 3554 26290
rect 3554 26238 3556 26290
rect 3500 26236 3556 26238
rect 6524 27356 6580 27412
rect 4956 26236 5012 26292
rect 4172 26178 4228 26180
rect 4172 26126 4174 26178
rect 4174 26126 4226 26178
rect 4226 26126 4228 26178
rect 4172 26124 4228 26126
rect 5628 26124 5684 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 5964 26124 6020 26180
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 6300 25452 6356 25508
rect 6972 29036 7028 29092
rect 8204 29260 8260 29316
rect 12012 31948 12068 32004
rect 11452 31836 11508 31892
rect 11340 31276 11396 31332
rect 12236 31724 12292 31780
rect 12460 31164 12516 31220
rect 12012 30994 12068 30996
rect 12012 30942 12014 30994
rect 12014 30942 12066 30994
rect 12066 30942 12068 30994
rect 12012 30940 12068 30942
rect 12572 30994 12628 30996
rect 12572 30942 12574 30994
rect 12574 30942 12626 30994
rect 12626 30942 12628 30994
rect 12572 30940 12628 30942
rect 12348 30716 12404 30772
rect 12796 30604 12852 30660
rect 13468 35698 13524 35700
rect 13468 35646 13470 35698
rect 13470 35646 13522 35698
rect 13522 35646 13524 35698
rect 13468 35644 13524 35646
rect 13468 34524 13524 34580
rect 13580 34412 13636 34468
rect 13468 34354 13524 34356
rect 13468 34302 13470 34354
rect 13470 34302 13522 34354
rect 13522 34302 13524 34354
rect 13468 34300 13524 34302
rect 13020 31724 13076 31780
rect 13244 34130 13300 34132
rect 13244 34078 13246 34130
rect 13246 34078 13298 34130
rect 13298 34078 13300 34130
rect 13244 34076 13300 34078
rect 11452 30268 11508 30324
rect 12796 30210 12852 30212
rect 12796 30158 12798 30210
rect 12798 30158 12850 30210
rect 12850 30158 12852 30210
rect 12796 30156 12852 30158
rect 11564 30044 11620 30100
rect 9772 29314 9828 29316
rect 9772 29262 9774 29314
rect 9774 29262 9826 29314
rect 9826 29262 9828 29314
rect 9772 29260 9828 29262
rect 12012 29650 12068 29652
rect 12012 29598 12014 29650
rect 12014 29598 12066 29650
rect 12066 29598 12068 29650
rect 12012 29596 12068 29598
rect 12796 29372 12852 29428
rect 12460 29202 12516 29204
rect 12460 29150 12462 29202
rect 12462 29150 12514 29202
rect 12514 29150 12516 29202
rect 12460 29148 12516 29150
rect 12908 28028 12964 28084
rect 13132 30492 13188 30548
rect 9660 27916 9716 27972
rect 7756 27804 7812 27860
rect 8428 27804 8484 27860
rect 7980 27580 8036 27636
rect 7644 26962 7700 26964
rect 7644 26910 7646 26962
rect 7646 26910 7698 26962
rect 7698 26910 7700 26962
rect 7644 26908 7700 26910
rect 3948 23660 4004 23716
rect 3276 23154 3332 23156
rect 3276 23102 3278 23154
rect 3278 23102 3330 23154
rect 3330 23102 3332 23154
rect 3276 23100 3332 23102
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 5852 23714 5908 23716
rect 5852 23662 5854 23714
rect 5854 23662 5906 23714
rect 5906 23662 5908 23714
rect 5852 23660 5908 23662
rect 5740 23100 5796 23156
rect 5740 22428 5796 22484
rect 5964 23324 6020 23380
rect 6524 23436 6580 23492
rect 6076 23042 6132 23044
rect 6076 22990 6078 23042
rect 6078 22990 6130 23042
rect 6130 22990 6132 23042
rect 6076 22988 6132 22990
rect 6748 22428 6804 22484
rect 7308 26290 7364 26292
rect 7308 26238 7310 26290
rect 7310 26238 7362 26290
rect 7362 26238 7364 26290
rect 7308 26236 7364 26238
rect 6972 26012 7028 26068
rect 7308 25506 7364 25508
rect 7308 25454 7310 25506
rect 7310 25454 7362 25506
rect 7362 25454 7364 25506
rect 7308 25452 7364 25454
rect 7420 25340 7476 25396
rect 7756 26236 7812 26292
rect 7644 25618 7700 25620
rect 7644 25566 7646 25618
rect 7646 25566 7698 25618
rect 7698 25566 7700 25618
rect 7644 25564 7700 25566
rect 8540 26962 8596 26964
rect 8540 26910 8542 26962
rect 8542 26910 8594 26962
rect 8594 26910 8596 26962
rect 8540 26908 8596 26910
rect 7644 25004 7700 25060
rect 7980 25340 8036 25396
rect 8764 26290 8820 26292
rect 8764 26238 8766 26290
rect 8766 26238 8818 26290
rect 8818 26238 8820 26290
rect 8764 26236 8820 26238
rect 8764 25394 8820 25396
rect 8764 25342 8766 25394
rect 8766 25342 8818 25394
rect 8818 25342 8820 25394
rect 8764 25340 8820 25342
rect 8428 24892 8484 24948
rect 9548 27356 9604 27412
rect 10220 27970 10276 27972
rect 10220 27918 10222 27970
rect 10222 27918 10274 27970
rect 10274 27918 10276 27970
rect 10220 27916 10276 27918
rect 9884 27858 9940 27860
rect 9884 27806 9886 27858
rect 9886 27806 9938 27858
rect 9938 27806 9940 27858
rect 9884 27804 9940 27806
rect 10556 27858 10612 27860
rect 10556 27806 10558 27858
rect 10558 27806 10610 27858
rect 10610 27806 10612 27858
rect 10556 27804 10612 27806
rect 9436 26236 9492 26292
rect 9996 26908 10052 26964
rect 9660 26178 9716 26180
rect 9660 26126 9662 26178
rect 9662 26126 9714 26178
rect 9714 26126 9716 26178
rect 9660 26124 9716 26126
rect 9548 26012 9604 26068
rect 10108 26236 10164 26292
rect 9324 25452 9380 25508
rect 9548 25004 9604 25060
rect 9212 24892 9268 24948
rect 7084 23826 7140 23828
rect 7084 23774 7086 23826
rect 7086 23774 7138 23826
rect 7138 23774 7140 23826
rect 7084 23772 7140 23774
rect 7308 23548 7364 23604
rect 7532 23378 7588 23380
rect 7532 23326 7534 23378
rect 7534 23326 7586 23378
rect 7586 23326 7588 23378
rect 7532 23324 7588 23326
rect 7420 23212 7476 23268
rect 7420 22988 7476 23044
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 7868 23436 7924 23492
rect 10332 25618 10388 25620
rect 10332 25566 10334 25618
rect 10334 25566 10386 25618
rect 10386 25566 10388 25618
rect 10332 25564 10388 25566
rect 10332 24834 10388 24836
rect 10332 24782 10334 24834
rect 10334 24782 10386 24834
rect 10386 24782 10388 24834
rect 10332 24780 10388 24782
rect 7980 23324 8036 23380
rect 8652 24498 8708 24500
rect 8652 24446 8654 24498
rect 8654 24446 8706 24498
rect 8706 24446 8708 24498
rect 8652 24444 8708 24446
rect 8540 24108 8596 24164
rect 9324 24162 9380 24164
rect 9324 24110 9326 24162
rect 9326 24110 9378 24162
rect 9378 24110 9380 24162
rect 9324 24108 9380 24110
rect 8428 23772 8484 23828
rect 7980 22428 8036 22484
rect 9212 23826 9268 23828
rect 9212 23774 9214 23826
rect 9214 23774 9266 23826
rect 9266 23774 9268 23826
rect 9212 23772 9268 23774
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 6076 18450 6132 18452
rect 6076 18398 6078 18450
rect 6078 18398 6130 18450
rect 6130 18398 6132 18450
rect 6076 18396 6132 18398
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 6076 15148 6132 15204
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 8988 22482 9044 22484
rect 8988 22430 8990 22482
rect 8990 22430 9042 22482
rect 9042 22430 9044 22482
rect 8988 22428 9044 22430
rect 10332 23436 10388 23492
rect 11116 26962 11172 26964
rect 11116 26910 11118 26962
rect 11118 26910 11170 26962
rect 11170 26910 11172 26962
rect 11116 26908 11172 26910
rect 14028 36482 14084 36484
rect 14028 36430 14030 36482
rect 14030 36430 14082 36482
rect 14082 36430 14084 36482
rect 14028 36428 14084 36430
rect 13916 36204 13972 36260
rect 14140 36204 14196 36260
rect 13804 35644 13860 35700
rect 13916 35586 13972 35588
rect 13916 35534 13918 35586
rect 13918 35534 13970 35586
rect 13970 35534 13972 35586
rect 13916 35532 13972 35534
rect 13804 35196 13860 35252
rect 14028 34636 14084 34692
rect 14476 36764 14532 36820
rect 15036 38220 15092 38276
rect 14812 37212 14868 37268
rect 14364 36316 14420 36372
rect 14700 36988 14756 37044
rect 14252 35196 14308 35252
rect 14588 36258 14644 36260
rect 14588 36206 14590 36258
rect 14590 36206 14642 36258
rect 14642 36206 14644 36258
rect 14588 36204 14644 36206
rect 15036 36652 15092 36708
rect 14812 36482 14868 36484
rect 14812 36430 14814 36482
rect 14814 36430 14866 36482
rect 14866 36430 14868 36482
rect 14812 36428 14868 36430
rect 14700 35868 14756 35924
rect 14924 35980 14980 36036
rect 15148 36316 15204 36372
rect 14812 35810 14868 35812
rect 14812 35758 14814 35810
rect 14814 35758 14866 35810
rect 14866 35758 14868 35810
rect 14812 35756 14868 35758
rect 14252 34412 14308 34468
rect 14588 34412 14644 34468
rect 13916 33122 13972 33124
rect 13916 33070 13918 33122
rect 13918 33070 13970 33122
rect 13970 33070 13972 33122
rect 13916 33068 13972 33070
rect 13916 32732 13972 32788
rect 13468 31778 13524 31780
rect 13468 31726 13470 31778
rect 13470 31726 13522 31778
rect 13522 31726 13524 31778
rect 13468 31724 13524 31726
rect 14700 34076 14756 34132
rect 14812 33852 14868 33908
rect 14140 33346 14196 33348
rect 14140 33294 14142 33346
rect 14142 33294 14194 33346
rect 14194 33294 14196 33346
rect 14140 33292 14196 33294
rect 14028 31612 14084 31668
rect 13916 31554 13972 31556
rect 13916 31502 13918 31554
rect 13918 31502 13970 31554
rect 13970 31502 13972 31554
rect 13916 31500 13972 31502
rect 14700 32956 14756 33012
rect 15484 38332 15540 38388
rect 15708 38162 15764 38164
rect 15708 38110 15710 38162
rect 15710 38110 15762 38162
rect 15762 38110 15764 38162
rect 15708 38108 15764 38110
rect 15372 36876 15428 36932
rect 15932 37436 15988 37492
rect 15596 37042 15652 37044
rect 15596 36990 15598 37042
rect 15598 36990 15650 37042
rect 15650 36990 15652 37042
rect 15596 36988 15652 36990
rect 18060 43932 18116 43988
rect 18172 44156 18228 44212
rect 17836 43596 17892 43652
rect 19516 50428 19572 50484
rect 18956 49810 19012 49812
rect 18956 49758 18958 49810
rect 18958 49758 19010 49810
rect 19010 49758 19012 49810
rect 18956 49756 19012 49758
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19964 51266 20020 51268
rect 19964 51214 19966 51266
rect 19966 51214 20018 51266
rect 20018 51214 20020 51266
rect 19964 51212 20020 51214
rect 19964 50876 20020 50932
rect 21084 55356 21140 55412
rect 21420 54684 21476 54740
rect 21980 54738 22036 54740
rect 21980 54686 21982 54738
rect 21982 54686 22034 54738
rect 22034 54686 22036 54738
rect 21980 54684 22036 54686
rect 22652 54738 22708 54740
rect 22652 54686 22654 54738
rect 22654 54686 22706 54738
rect 22706 54686 22708 54738
rect 22652 54684 22708 54686
rect 21532 52108 21588 52164
rect 21868 52556 21924 52612
rect 21980 52220 22036 52276
rect 21756 51548 21812 51604
rect 21532 50652 21588 50708
rect 19628 50316 19684 50372
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 18732 49532 18788 49588
rect 19068 49532 19124 49588
rect 18732 49308 18788 49364
rect 18620 49026 18676 49028
rect 18620 48974 18622 49026
rect 18622 48974 18674 49026
rect 18674 48974 18676 49026
rect 18620 48972 18676 48974
rect 18508 48914 18564 48916
rect 18508 48862 18510 48914
rect 18510 48862 18562 48914
rect 18562 48862 18564 48914
rect 18508 48860 18564 48862
rect 18620 47404 18676 47460
rect 19180 49308 19236 49364
rect 19068 49084 19124 49140
rect 19964 49532 20020 49588
rect 20076 49308 20132 49364
rect 20188 49250 20244 49252
rect 20188 49198 20190 49250
rect 20190 49198 20242 49250
rect 20242 49198 20244 49250
rect 20188 49196 20244 49198
rect 20412 50316 20468 50372
rect 19628 49026 19684 49028
rect 19628 48974 19630 49026
rect 19630 48974 19682 49026
rect 19682 48974 19684 49026
rect 19628 48972 19684 48974
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19740 48412 19796 48468
rect 20636 49810 20692 49812
rect 20636 49758 20638 49810
rect 20638 49758 20690 49810
rect 20690 49758 20692 49810
rect 20636 49756 20692 49758
rect 20412 48748 20468 48804
rect 20524 49308 20580 49364
rect 21308 49308 21364 49364
rect 20524 48860 20580 48916
rect 20860 48972 20916 49028
rect 20748 48636 20804 48692
rect 19852 47570 19908 47572
rect 19852 47518 19854 47570
rect 19854 47518 19906 47570
rect 19906 47518 19908 47570
rect 19852 47516 19908 47518
rect 19404 47292 19460 47348
rect 19180 45666 19236 45668
rect 19180 45614 19182 45666
rect 19182 45614 19234 45666
rect 19234 45614 19236 45666
rect 19180 45612 19236 45614
rect 18956 44380 19012 44436
rect 18396 43596 18452 43652
rect 17052 42866 17108 42868
rect 17052 42814 17054 42866
rect 17054 42814 17106 42866
rect 17106 42814 17108 42866
rect 17052 42812 17108 42814
rect 17276 42700 17332 42756
rect 16940 40572 16996 40628
rect 16828 40348 16884 40404
rect 17388 41692 17444 41748
rect 17276 41410 17332 41412
rect 17276 41358 17278 41410
rect 17278 41358 17330 41410
rect 17330 41358 17332 41410
rect 17276 41356 17332 41358
rect 17836 42866 17892 42868
rect 17836 42814 17838 42866
rect 17838 42814 17890 42866
rect 17890 42814 17892 42866
rect 17836 42812 17892 42814
rect 18060 42924 18116 42980
rect 17724 41970 17780 41972
rect 17724 41918 17726 41970
rect 17726 41918 17778 41970
rect 17778 41918 17780 41970
rect 17724 41916 17780 41918
rect 17948 42364 18004 42420
rect 17948 41692 18004 41748
rect 16604 39676 16660 39732
rect 16828 39900 16884 39956
rect 16828 39004 16884 39060
rect 16828 38834 16884 38836
rect 16828 38782 16830 38834
rect 16830 38782 16882 38834
rect 16882 38782 16884 38834
rect 16828 38780 16884 38782
rect 16604 38108 16660 38164
rect 16156 36316 16212 36372
rect 16044 36258 16100 36260
rect 16044 36206 16046 36258
rect 16046 36206 16098 36258
rect 16098 36206 16100 36258
rect 16044 36204 16100 36206
rect 16268 36204 16324 36260
rect 15372 35922 15428 35924
rect 15372 35870 15374 35922
rect 15374 35870 15426 35922
rect 15426 35870 15428 35922
rect 15372 35868 15428 35870
rect 15596 35698 15652 35700
rect 15596 35646 15598 35698
rect 15598 35646 15650 35698
rect 15650 35646 15652 35698
rect 15596 35644 15652 35646
rect 15260 35084 15316 35140
rect 16492 35698 16548 35700
rect 16492 35646 16494 35698
rect 16494 35646 16546 35698
rect 16546 35646 16548 35698
rect 16492 35644 16548 35646
rect 16044 35474 16100 35476
rect 16044 35422 16046 35474
rect 16046 35422 16098 35474
rect 16098 35422 16100 35474
rect 16044 35420 16100 35422
rect 15932 35308 15988 35364
rect 15484 34972 15540 35028
rect 15596 34524 15652 34580
rect 15036 33292 15092 33348
rect 15148 34076 15204 34132
rect 15484 33964 15540 34020
rect 15260 33068 15316 33124
rect 15596 33122 15652 33124
rect 15596 33070 15598 33122
rect 15598 33070 15650 33122
rect 15650 33070 15652 33122
rect 15596 33068 15652 33070
rect 15596 32674 15652 32676
rect 15596 32622 15598 32674
rect 15598 32622 15650 32674
rect 15650 32622 15652 32674
rect 15596 32620 15652 32622
rect 15372 32450 15428 32452
rect 15372 32398 15374 32450
rect 15374 32398 15426 32450
rect 15426 32398 15428 32450
rect 15372 32396 15428 32398
rect 15820 32732 15876 32788
rect 15820 32396 15876 32452
rect 15372 32060 15428 32116
rect 14812 31666 14868 31668
rect 14812 31614 14814 31666
rect 14814 31614 14866 31666
rect 14866 31614 14868 31666
rect 14812 31612 14868 31614
rect 13916 30940 13972 30996
rect 14028 30882 14084 30884
rect 14028 30830 14030 30882
rect 14030 30830 14082 30882
rect 14082 30830 14084 30882
rect 14028 30828 14084 30830
rect 13692 30492 13748 30548
rect 13804 30604 13860 30660
rect 13468 30098 13524 30100
rect 13468 30046 13470 30098
rect 13470 30046 13522 30098
rect 13522 30046 13524 30098
rect 13468 30044 13524 30046
rect 13356 29596 13412 29652
rect 13468 28924 13524 28980
rect 13244 28588 13300 28644
rect 13020 27634 13076 27636
rect 13020 27582 13022 27634
rect 13022 27582 13074 27634
rect 13074 27582 13076 27634
rect 13020 27580 13076 27582
rect 12236 27074 12292 27076
rect 12236 27022 12238 27074
rect 12238 27022 12290 27074
rect 12290 27022 12292 27074
rect 12236 27020 12292 27022
rect 13132 27020 13188 27076
rect 11340 26348 11396 26404
rect 10780 24946 10836 24948
rect 10780 24894 10782 24946
rect 10782 24894 10834 24946
rect 10834 24894 10836 24946
rect 10780 24892 10836 24894
rect 10668 24834 10724 24836
rect 10668 24782 10670 24834
rect 10670 24782 10722 24834
rect 10722 24782 10724 24834
rect 10668 24780 10724 24782
rect 10780 23826 10836 23828
rect 10780 23774 10782 23826
rect 10782 23774 10834 23826
rect 10834 23774 10836 23826
rect 10780 23772 10836 23774
rect 12236 26402 12292 26404
rect 12236 26350 12238 26402
rect 12238 26350 12290 26402
rect 12290 26350 12292 26402
rect 12236 26348 12292 26350
rect 13356 28812 13412 28868
rect 14252 30380 14308 30436
rect 15036 31724 15092 31780
rect 15260 31500 15316 31556
rect 15036 30604 15092 30660
rect 15148 31052 15204 31108
rect 14924 30434 14980 30436
rect 14924 30382 14926 30434
rect 14926 30382 14978 30434
rect 14978 30382 14980 30434
rect 14924 30380 14980 30382
rect 15036 30268 15092 30324
rect 14140 30156 14196 30212
rect 13804 29426 13860 29428
rect 13804 29374 13806 29426
rect 13806 29374 13858 29426
rect 13858 29374 13860 29426
rect 13804 29372 13860 29374
rect 14700 30044 14756 30100
rect 16268 34860 16324 34916
rect 16380 34524 16436 34580
rect 16268 34242 16324 34244
rect 16268 34190 16270 34242
rect 16270 34190 16322 34242
rect 16322 34190 16324 34242
rect 16268 34188 16324 34190
rect 16492 34130 16548 34132
rect 16492 34078 16494 34130
rect 16494 34078 16546 34130
rect 16546 34078 16548 34130
rect 16492 34076 16548 34078
rect 16828 37100 16884 37156
rect 17612 41074 17668 41076
rect 17612 41022 17614 41074
rect 17614 41022 17666 41074
rect 17666 41022 17668 41074
rect 17612 41020 17668 41022
rect 17164 40012 17220 40068
rect 17164 38108 17220 38164
rect 16940 36988 16996 37044
rect 16828 35868 16884 35924
rect 16716 35532 16772 35588
rect 16604 33852 16660 33908
rect 16156 32620 16212 32676
rect 16044 31778 16100 31780
rect 16044 31726 16046 31778
rect 16046 31726 16098 31778
rect 16098 31726 16100 31778
rect 16044 31724 16100 31726
rect 16044 31276 16100 31332
rect 16604 31724 16660 31780
rect 15708 31106 15764 31108
rect 15708 31054 15710 31106
rect 15710 31054 15762 31106
rect 15762 31054 15764 31106
rect 15708 31052 15764 31054
rect 15596 30492 15652 30548
rect 15260 30268 15316 30324
rect 15708 30322 15764 30324
rect 15708 30270 15710 30322
rect 15710 30270 15762 30322
rect 15762 30270 15764 30322
rect 15708 30268 15764 30270
rect 14476 29820 14532 29876
rect 14252 29260 14308 29316
rect 13804 28924 13860 28980
rect 13468 28642 13524 28644
rect 13468 28590 13470 28642
rect 13470 28590 13522 28642
rect 13522 28590 13524 28642
rect 13468 28588 13524 28590
rect 14812 29708 14868 29764
rect 14476 28812 14532 28868
rect 14700 28812 14756 28868
rect 15932 29708 15988 29764
rect 16268 31500 16324 31556
rect 16268 30994 16324 30996
rect 16268 30942 16270 30994
rect 16270 30942 16322 30994
rect 16322 30942 16324 30994
rect 16268 30940 16324 30942
rect 16604 31106 16660 31108
rect 16604 31054 16606 31106
rect 16606 31054 16658 31106
rect 16658 31054 16660 31106
rect 16604 31052 16660 31054
rect 15148 29596 15204 29652
rect 15036 29538 15092 29540
rect 15036 29486 15038 29538
rect 15038 29486 15090 29538
rect 15090 29486 15092 29538
rect 15036 29484 15092 29486
rect 16156 29484 16212 29540
rect 15820 29426 15876 29428
rect 15820 29374 15822 29426
rect 15822 29374 15874 29426
rect 15874 29374 15876 29426
rect 15820 29372 15876 29374
rect 14364 28476 14420 28532
rect 14028 28418 14084 28420
rect 14028 28366 14030 28418
rect 14030 28366 14082 28418
rect 14082 28366 14084 28418
rect 14028 28364 14084 28366
rect 13580 27858 13636 27860
rect 13580 27806 13582 27858
rect 13582 27806 13634 27858
rect 13634 27806 13636 27858
rect 13580 27804 13636 27806
rect 14700 27804 14756 27860
rect 14364 27580 14420 27636
rect 14252 27020 14308 27076
rect 11900 25116 11956 25172
rect 11452 25004 11508 25060
rect 12236 24332 12292 24388
rect 12348 24444 12404 24500
rect 12348 23660 12404 23716
rect 10892 23324 10948 23380
rect 13020 24780 13076 24836
rect 14140 26236 14196 26292
rect 14140 25452 14196 25508
rect 13356 25116 13412 25172
rect 13692 25228 13748 25284
rect 13804 25004 13860 25060
rect 15036 27074 15092 27076
rect 15036 27022 15038 27074
rect 15038 27022 15090 27074
rect 15090 27022 15092 27074
rect 15036 27020 15092 27022
rect 15148 26348 15204 26404
rect 14476 26236 14532 26292
rect 14924 26012 14980 26068
rect 14700 25506 14756 25508
rect 14700 25454 14702 25506
rect 14702 25454 14754 25506
rect 14754 25454 14756 25506
rect 14700 25452 14756 25454
rect 14588 25282 14644 25284
rect 14588 25230 14590 25282
rect 14590 25230 14642 25282
rect 14642 25230 14644 25282
rect 14588 25228 14644 25230
rect 14588 24834 14644 24836
rect 14588 24782 14590 24834
rect 14590 24782 14642 24834
rect 14642 24782 14644 24834
rect 14588 24780 14644 24782
rect 12908 24332 12964 24388
rect 13468 23660 13524 23716
rect 10220 22428 10276 22484
rect 8092 20524 8148 20580
rect 8652 19404 8708 19460
rect 11004 22428 11060 22484
rect 12908 22482 12964 22484
rect 12908 22430 12910 22482
rect 12910 22430 12962 22482
rect 12962 22430 12964 22482
rect 12908 22428 12964 22430
rect 15260 26290 15316 26292
rect 15260 26238 15262 26290
rect 15262 26238 15314 26290
rect 15314 26238 15316 26290
rect 15260 26236 15316 26238
rect 15708 29148 15764 29204
rect 15596 27746 15652 27748
rect 15596 27694 15598 27746
rect 15598 27694 15650 27746
rect 15650 27694 15652 27746
rect 15596 27692 15652 27694
rect 15484 26066 15540 26068
rect 15484 26014 15486 26066
rect 15486 26014 15538 26066
rect 15538 26014 15540 26066
rect 15484 26012 15540 26014
rect 16044 28530 16100 28532
rect 16044 28478 16046 28530
rect 16046 28478 16098 28530
rect 16098 28478 16100 28530
rect 16044 28476 16100 28478
rect 16044 28252 16100 28308
rect 16156 28140 16212 28196
rect 15820 27186 15876 27188
rect 15820 27134 15822 27186
rect 15822 27134 15874 27186
rect 15874 27134 15876 27186
rect 15820 27132 15876 27134
rect 15820 26514 15876 26516
rect 15820 26462 15822 26514
rect 15822 26462 15874 26514
rect 15874 26462 15876 26514
rect 15820 26460 15876 26462
rect 16716 29372 16772 29428
rect 16492 28364 16548 28420
rect 17164 37884 17220 37940
rect 17164 37548 17220 37604
rect 17836 40908 17892 40964
rect 18844 42476 18900 42532
rect 18620 42252 18676 42308
rect 18172 41692 18228 41748
rect 18396 41804 18452 41860
rect 18060 41580 18116 41636
rect 18396 41244 18452 41300
rect 18508 40684 18564 40740
rect 17500 39730 17556 39732
rect 17500 39678 17502 39730
rect 17502 39678 17554 39730
rect 17554 39678 17556 39730
rect 17500 39676 17556 39678
rect 17724 39676 17780 39732
rect 17836 40348 17892 40404
rect 18284 40348 18340 40404
rect 18284 39900 18340 39956
rect 17500 38668 17556 38724
rect 17388 37772 17444 37828
rect 17388 37490 17444 37492
rect 17388 37438 17390 37490
rect 17390 37438 17442 37490
rect 17442 37438 17444 37490
rect 17388 37436 17444 37438
rect 17612 37100 17668 37156
rect 17836 38780 17892 38836
rect 17836 37548 17892 37604
rect 18284 38780 18340 38836
rect 18172 38722 18228 38724
rect 18172 38670 18174 38722
rect 18174 38670 18226 38722
rect 18226 38670 18228 38722
rect 18172 38668 18228 38670
rect 17948 37436 18004 37492
rect 18508 39618 18564 39620
rect 18508 39566 18510 39618
rect 18510 39566 18562 39618
rect 18562 39566 18564 39618
rect 18508 39564 18564 39566
rect 18508 38108 18564 38164
rect 17388 35586 17444 35588
rect 17388 35534 17390 35586
rect 17390 35534 17442 35586
rect 17442 35534 17444 35586
rect 17388 35532 17444 35534
rect 17500 34860 17556 34916
rect 17500 34076 17556 34132
rect 17612 34412 17668 34468
rect 17612 33852 17668 33908
rect 17724 35420 17780 35476
rect 17052 32732 17108 32788
rect 17164 33068 17220 33124
rect 16940 32620 16996 32676
rect 17388 32786 17444 32788
rect 17388 32734 17390 32786
rect 17390 32734 17442 32786
rect 17442 32734 17444 32786
rect 17388 32732 17444 32734
rect 17388 31500 17444 31556
rect 17388 31218 17444 31220
rect 17388 31166 17390 31218
rect 17390 31166 17442 31218
rect 17442 31166 17444 31218
rect 17388 31164 17444 31166
rect 17612 31106 17668 31108
rect 17612 31054 17614 31106
rect 17614 31054 17666 31106
rect 17666 31054 17668 31106
rect 17612 31052 17668 31054
rect 17164 30716 17220 30772
rect 17948 36316 18004 36372
rect 18284 35420 18340 35476
rect 17948 33122 18004 33124
rect 17948 33070 17950 33122
rect 17950 33070 18002 33122
rect 18002 33070 18004 33122
rect 17948 33068 18004 33070
rect 18844 41970 18900 41972
rect 18844 41918 18846 41970
rect 18846 41918 18898 41970
rect 18898 41918 18900 41970
rect 18844 41916 18900 41918
rect 18732 41356 18788 41412
rect 19068 41692 19124 41748
rect 19068 40908 19124 40964
rect 18844 40402 18900 40404
rect 18844 40350 18846 40402
rect 18846 40350 18898 40402
rect 18898 40350 18900 40402
rect 18844 40348 18900 40350
rect 19068 40348 19124 40404
rect 18844 39730 18900 39732
rect 18844 39678 18846 39730
rect 18846 39678 18898 39730
rect 18898 39678 18900 39730
rect 18844 39676 18900 39678
rect 18844 39116 18900 39172
rect 19292 41804 19348 41860
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20524 47682 20580 47684
rect 20524 47630 20526 47682
rect 20526 47630 20578 47682
rect 20578 47630 20580 47682
rect 20524 47628 20580 47630
rect 20412 46956 20468 47012
rect 21644 49196 21700 49252
rect 21420 48972 21476 49028
rect 21532 48860 21588 48916
rect 21084 48748 21140 48804
rect 20972 48466 21028 48468
rect 20972 48414 20974 48466
rect 20974 48414 21026 48466
rect 21026 48414 21028 48466
rect 20972 48412 21028 48414
rect 20748 47292 20804 47348
rect 20412 46620 20468 46676
rect 19628 45612 19684 45668
rect 19516 45164 19572 45220
rect 19516 44434 19572 44436
rect 19516 44382 19518 44434
rect 19518 44382 19570 44434
rect 19570 44382 19572 44434
rect 19516 44380 19572 44382
rect 20076 45724 20132 45780
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 20076 44828 20132 44884
rect 19852 44210 19908 44212
rect 19852 44158 19854 44210
rect 19854 44158 19906 44210
rect 19906 44158 19908 44210
rect 19852 44156 19908 44158
rect 19628 43932 19684 43988
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19516 42476 19572 42532
rect 21420 47628 21476 47684
rect 21420 47458 21476 47460
rect 21420 47406 21422 47458
rect 21422 47406 21474 47458
rect 21474 47406 21476 47458
rect 21420 47404 21476 47406
rect 23548 55020 23604 55076
rect 23324 53788 23380 53844
rect 22876 53730 22932 53732
rect 22876 53678 22878 53730
rect 22878 53678 22930 53730
rect 22930 53678 22932 53730
rect 22876 53676 22932 53678
rect 22540 51602 22596 51604
rect 22540 51550 22542 51602
rect 22542 51550 22594 51602
rect 22594 51550 22596 51602
rect 22540 51548 22596 51550
rect 22652 51324 22708 51380
rect 22092 50876 22148 50932
rect 22988 51212 23044 51268
rect 22652 50594 22708 50596
rect 22652 50542 22654 50594
rect 22654 50542 22706 50594
rect 22706 50542 22708 50594
rect 22652 50540 22708 50542
rect 22428 50482 22484 50484
rect 22428 50430 22430 50482
rect 22430 50430 22482 50482
rect 22482 50430 22484 50482
rect 22428 50428 22484 50430
rect 21868 49308 21924 49364
rect 22092 49196 22148 49252
rect 21868 49026 21924 49028
rect 21868 48974 21870 49026
rect 21870 48974 21922 49026
rect 21922 48974 21924 49026
rect 21868 48972 21924 48974
rect 21756 48636 21812 48692
rect 22540 48412 22596 48468
rect 22540 47682 22596 47684
rect 22540 47630 22542 47682
rect 22542 47630 22594 47682
rect 22594 47630 22596 47682
rect 22540 47628 22596 47630
rect 22316 47346 22372 47348
rect 22316 47294 22318 47346
rect 22318 47294 22370 47346
rect 22370 47294 22372 47346
rect 22316 47292 22372 47294
rect 20860 45164 20916 45220
rect 21308 46562 21364 46564
rect 21308 46510 21310 46562
rect 21310 46510 21362 46562
rect 21362 46510 21364 46562
rect 21308 46508 21364 46510
rect 22988 47234 23044 47236
rect 22988 47182 22990 47234
rect 22990 47182 23042 47234
rect 23042 47182 23044 47234
rect 22988 47180 23044 47182
rect 21756 46732 21812 46788
rect 21196 45612 21252 45668
rect 20412 44322 20468 44324
rect 20412 44270 20414 44322
rect 20414 44270 20466 44322
rect 20466 44270 20468 44322
rect 20412 44268 20468 44270
rect 20412 43260 20468 43316
rect 20188 42700 20244 42756
rect 19628 42252 19684 42308
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19852 42028 19908 42084
rect 19292 41186 19348 41188
rect 19292 41134 19294 41186
rect 19294 41134 19346 41186
rect 19346 41134 19348 41186
rect 19292 41132 19348 41134
rect 19516 41020 19572 41076
rect 19292 40626 19348 40628
rect 19292 40574 19294 40626
rect 19294 40574 19346 40626
rect 19346 40574 19348 40626
rect 19292 40572 19348 40574
rect 19292 39900 19348 39956
rect 19180 39564 19236 39620
rect 19180 38946 19236 38948
rect 19180 38894 19182 38946
rect 19182 38894 19234 38946
rect 19234 38894 19236 38946
rect 19180 38892 19236 38894
rect 18732 36428 18788 36484
rect 18956 37436 19012 37492
rect 19180 37436 19236 37492
rect 18396 34636 18452 34692
rect 18396 34076 18452 34132
rect 18284 33964 18340 34020
rect 18620 33180 18676 33236
rect 19404 38668 19460 38724
rect 19964 41804 20020 41860
rect 19964 41580 20020 41636
rect 19740 41186 19796 41188
rect 19740 41134 19742 41186
rect 19742 41134 19794 41186
rect 19794 41134 19796 41186
rect 19740 41132 19796 41134
rect 20636 41074 20692 41076
rect 20636 41022 20638 41074
rect 20638 41022 20690 41074
rect 20690 41022 20692 41074
rect 20636 41020 20692 41022
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 20300 40962 20356 40964
rect 20300 40910 20302 40962
rect 20302 40910 20354 40962
rect 20354 40910 20356 40962
rect 20300 40908 20356 40910
rect 20636 40626 20692 40628
rect 20636 40574 20638 40626
rect 20638 40574 20690 40626
rect 20690 40574 20692 40626
rect 20636 40572 20692 40574
rect 19628 39900 19684 39956
rect 20076 39506 20132 39508
rect 20076 39454 20078 39506
rect 20078 39454 20130 39506
rect 20130 39454 20132 39506
rect 20076 39452 20132 39454
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19628 38162 19684 38164
rect 19628 38110 19630 38162
rect 19630 38110 19682 38162
rect 19682 38110 19684 38162
rect 19628 38108 19684 38110
rect 20076 38722 20132 38724
rect 20076 38670 20078 38722
rect 20078 38670 20130 38722
rect 20130 38670 20132 38722
rect 20076 38668 20132 38670
rect 21756 45164 21812 45220
rect 21308 44156 21364 44212
rect 21196 43596 21252 43652
rect 21532 43708 21588 43764
rect 23212 52108 23268 52164
rect 23436 53452 23492 53508
rect 23436 52668 23492 52724
rect 23324 51884 23380 51940
rect 23660 53842 23716 53844
rect 23660 53790 23662 53842
rect 23662 53790 23714 53842
rect 23714 53790 23716 53842
rect 23660 53788 23716 53790
rect 23884 52556 23940 52612
rect 24668 55244 24724 55300
rect 24668 54738 24724 54740
rect 24668 54686 24670 54738
rect 24670 54686 24722 54738
rect 24722 54686 24724 54738
rect 24668 54684 24724 54686
rect 25676 55298 25732 55300
rect 25676 55246 25678 55298
rect 25678 55246 25730 55298
rect 25730 55246 25732 55298
rect 25676 55244 25732 55246
rect 26460 55186 26516 55188
rect 26460 55134 26462 55186
rect 26462 55134 26514 55186
rect 26514 55134 26516 55186
rect 26460 55132 26516 55134
rect 24332 53730 24388 53732
rect 24332 53678 24334 53730
rect 24334 53678 24386 53730
rect 24386 53678 24388 53730
rect 24332 53676 24388 53678
rect 24220 52722 24276 52724
rect 24220 52670 24222 52722
rect 24222 52670 24274 52722
rect 24274 52670 24276 52722
rect 24220 52668 24276 52670
rect 23660 51996 23716 52052
rect 23772 51884 23828 51940
rect 23324 50876 23380 50932
rect 23100 45164 23156 45220
rect 23884 51490 23940 51492
rect 23884 51438 23886 51490
rect 23886 51438 23938 51490
rect 23938 51438 23940 51490
rect 23884 51436 23940 51438
rect 23772 51212 23828 51268
rect 23660 50540 23716 50596
rect 23772 50428 23828 50484
rect 24108 50594 24164 50596
rect 24108 50542 24110 50594
rect 24110 50542 24162 50594
rect 24162 50542 24164 50594
rect 24108 50540 24164 50542
rect 24556 52722 24612 52724
rect 24556 52670 24558 52722
rect 24558 52670 24610 52722
rect 24610 52670 24612 52722
rect 24556 52668 24612 52670
rect 25564 53676 25620 53732
rect 24892 52556 24948 52612
rect 24444 52162 24500 52164
rect 24444 52110 24446 52162
rect 24446 52110 24498 52162
rect 24498 52110 24500 52162
rect 24444 52108 24500 52110
rect 24668 52050 24724 52052
rect 24668 51998 24670 52050
rect 24670 51998 24722 52050
rect 24722 51998 24724 52050
rect 24668 51996 24724 51998
rect 26124 52108 26180 52164
rect 24668 50652 24724 50708
rect 24444 50540 24500 50596
rect 23660 49420 23716 49476
rect 23996 48914 24052 48916
rect 23996 48862 23998 48914
rect 23998 48862 24050 48914
rect 24050 48862 24052 48914
rect 23996 48860 24052 48862
rect 23660 46786 23716 46788
rect 23660 46734 23662 46786
rect 23662 46734 23714 46786
rect 23714 46734 23716 46786
rect 23660 46732 23716 46734
rect 24556 50482 24612 50484
rect 24556 50430 24558 50482
rect 24558 50430 24610 50482
rect 24610 50430 24612 50482
rect 24556 50428 24612 50430
rect 24332 46508 24388 46564
rect 22092 44210 22148 44212
rect 22092 44158 22094 44210
rect 22094 44158 22146 44210
rect 22146 44158 22148 44210
rect 22092 44156 22148 44158
rect 22988 43708 23044 43764
rect 22428 43484 22484 43540
rect 21308 42642 21364 42644
rect 21308 42590 21310 42642
rect 21310 42590 21362 42642
rect 21362 42590 21364 42642
rect 21308 42588 21364 42590
rect 21196 42476 21252 42532
rect 20860 42028 20916 42084
rect 20972 41970 21028 41972
rect 20972 41918 20974 41970
rect 20974 41918 21026 41970
rect 21026 41918 21028 41970
rect 20972 41916 21028 41918
rect 21532 42252 21588 42308
rect 21532 41970 21588 41972
rect 21532 41918 21534 41970
rect 21534 41918 21586 41970
rect 21586 41918 21588 41970
rect 21532 41916 21588 41918
rect 22652 43372 22708 43428
rect 23324 43484 23380 43540
rect 23884 43426 23940 43428
rect 23884 43374 23886 43426
rect 23886 43374 23938 43426
rect 23938 43374 23940 43426
rect 23884 43372 23940 43374
rect 23100 42812 23156 42868
rect 23548 42754 23604 42756
rect 23548 42702 23550 42754
rect 23550 42702 23602 42754
rect 23602 42702 23604 42754
rect 23548 42700 23604 42702
rect 21868 42530 21924 42532
rect 21868 42478 21870 42530
rect 21870 42478 21922 42530
rect 21922 42478 21924 42530
rect 21868 42476 21924 42478
rect 22092 42194 22148 42196
rect 22092 42142 22094 42194
rect 22094 42142 22146 42194
rect 22146 42142 22148 42194
rect 22092 42140 22148 42142
rect 23212 42140 23268 42196
rect 21756 41916 21812 41972
rect 22092 41244 22148 41300
rect 21980 41132 22036 41188
rect 21084 39788 21140 39844
rect 21084 39004 21140 39060
rect 20300 38834 20356 38836
rect 20300 38782 20302 38834
rect 20302 38782 20354 38834
rect 20354 38782 20356 38834
rect 20300 38780 20356 38782
rect 20188 38444 20244 38500
rect 20636 38610 20692 38612
rect 20636 38558 20638 38610
rect 20638 38558 20690 38610
rect 20690 38558 20692 38610
rect 20636 38556 20692 38558
rect 20412 38444 20468 38500
rect 21196 38444 21252 38500
rect 20524 38332 20580 38388
rect 20636 38274 20692 38276
rect 20636 38222 20638 38274
rect 20638 38222 20690 38274
rect 20690 38222 20692 38274
rect 20636 38220 20692 38222
rect 21756 40572 21812 40628
rect 21644 40460 21700 40516
rect 21532 39506 21588 39508
rect 21532 39454 21534 39506
rect 21534 39454 21586 39506
rect 21586 39454 21588 39506
rect 21532 39452 21588 39454
rect 21756 39788 21812 39844
rect 21868 39452 21924 39508
rect 21532 38668 21588 38724
rect 22428 41298 22484 41300
rect 22428 41246 22430 41298
rect 22430 41246 22482 41298
rect 22482 41246 22484 41298
rect 22428 41244 22484 41246
rect 23212 41244 23268 41300
rect 22316 40684 22372 40740
rect 23212 40626 23268 40628
rect 23212 40574 23214 40626
rect 23214 40574 23266 40626
rect 23266 40574 23268 40626
rect 23212 40572 23268 40574
rect 23324 40684 23380 40740
rect 22540 40402 22596 40404
rect 22540 40350 22542 40402
rect 22542 40350 22594 40402
rect 22594 40350 22596 40402
rect 22540 40348 22596 40350
rect 22988 39788 23044 39844
rect 22092 39618 22148 39620
rect 22092 39566 22094 39618
rect 22094 39566 22146 39618
rect 22146 39566 22148 39618
rect 22092 39564 22148 39566
rect 22092 38892 22148 38948
rect 21532 38444 21588 38500
rect 20636 37884 20692 37940
rect 20188 37826 20244 37828
rect 20188 37774 20190 37826
rect 20190 37774 20242 37826
rect 20242 37774 20244 37826
rect 20188 37772 20244 37774
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20524 37548 20580 37604
rect 19852 37436 19908 37492
rect 20748 37436 20804 37492
rect 19628 36876 19684 36932
rect 20300 37266 20356 37268
rect 20300 37214 20302 37266
rect 20302 37214 20354 37266
rect 20354 37214 20356 37266
rect 20300 37212 20356 37214
rect 19964 36764 20020 36820
rect 19292 35308 19348 35364
rect 19628 35980 19684 36036
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19516 35922 19572 35924
rect 19516 35870 19518 35922
rect 19518 35870 19570 35922
rect 19570 35870 19572 35922
rect 19516 35868 19572 35870
rect 20412 36988 20468 37044
rect 20860 36988 20916 37044
rect 20636 36370 20692 36372
rect 20636 36318 20638 36370
rect 20638 36318 20690 36370
rect 20690 36318 20692 36370
rect 20636 36316 20692 36318
rect 20636 35644 20692 35700
rect 20860 35532 20916 35588
rect 20748 35308 20804 35364
rect 19516 34914 19572 34916
rect 19516 34862 19518 34914
rect 19518 34862 19570 34914
rect 19570 34862 19572 34914
rect 19516 34860 19572 34862
rect 18284 32956 18340 33012
rect 18172 32620 18228 32676
rect 17948 32450 18004 32452
rect 17948 32398 17950 32450
rect 17950 32398 18002 32450
rect 18002 32398 18004 32450
rect 17948 32396 18004 32398
rect 18396 31724 18452 31780
rect 18284 31388 18340 31444
rect 18060 31164 18116 31220
rect 18396 30940 18452 30996
rect 18396 30492 18452 30548
rect 19964 34860 20020 34916
rect 20188 34636 20244 34692
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 20188 34300 20244 34356
rect 19740 33852 19796 33908
rect 19292 33404 19348 33460
rect 19068 33180 19124 33236
rect 18620 32674 18676 32676
rect 18620 32622 18622 32674
rect 18622 32622 18674 32674
rect 18674 32622 18676 32674
rect 18620 32620 18676 32622
rect 18620 32396 18676 32452
rect 18620 31948 18676 32004
rect 18508 30268 18564 30324
rect 17500 30210 17556 30212
rect 17500 30158 17502 30210
rect 17502 30158 17554 30210
rect 17554 30158 17556 30210
rect 17500 30156 17556 30158
rect 17500 29426 17556 29428
rect 17500 29374 17502 29426
rect 17502 29374 17554 29426
rect 17554 29374 17556 29426
rect 17500 29372 17556 29374
rect 19180 33068 19236 33124
rect 19292 32956 19348 33012
rect 19516 32732 19572 32788
rect 19068 32620 19124 32676
rect 18844 32284 18900 32340
rect 18172 30210 18228 30212
rect 18172 30158 18174 30210
rect 18174 30158 18226 30210
rect 18226 30158 18228 30210
rect 18172 30156 18228 30158
rect 17836 29820 17892 29876
rect 17948 29596 18004 29652
rect 18284 29596 18340 29652
rect 17052 28642 17108 28644
rect 17052 28590 17054 28642
rect 17054 28590 17106 28642
rect 17106 28590 17108 28642
rect 17052 28588 17108 28590
rect 17276 28476 17332 28532
rect 16380 27692 16436 27748
rect 17724 28588 17780 28644
rect 17724 28418 17780 28420
rect 17724 28366 17726 28418
rect 17726 28366 17778 28418
rect 17778 28366 17780 28418
rect 17724 28364 17780 28366
rect 17948 28418 18004 28420
rect 17948 28366 17950 28418
rect 17950 28366 18002 28418
rect 18002 28366 18004 28418
rect 17948 28364 18004 28366
rect 18172 28588 18228 28644
rect 18620 30210 18676 30212
rect 18620 30158 18622 30210
rect 18622 30158 18674 30210
rect 18674 30158 18676 30210
rect 18620 30156 18676 30158
rect 18620 29650 18676 29652
rect 18620 29598 18622 29650
rect 18622 29598 18674 29650
rect 18674 29598 18676 29650
rect 18620 29596 18676 29598
rect 18732 28700 18788 28756
rect 20300 33906 20356 33908
rect 20300 33854 20302 33906
rect 20302 33854 20354 33906
rect 20354 33854 20356 33906
rect 20300 33852 20356 33854
rect 19964 33404 20020 33460
rect 20300 33458 20356 33460
rect 20300 33406 20302 33458
rect 20302 33406 20354 33458
rect 20354 33406 20356 33458
rect 20300 33404 20356 33406
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20636 34636 20692 34692
rect 20748 34018 20804 34020
rect 20748 33966 20750 34018
rect 20750 33966 20802 34018
rect 20802 33966 20804 34018
rect 20748 33964 20804 33966
rect 21308 37826 21364 37828
rect 21308 37774 21310 37826
rect 21310 37774 21362 37826
rect 21362 37774 21364 37826
rect 21308 37772 21364 37774
rect 21308 37266 21364 37268
rect 21308 37214 21310 37266
rect 21310 37214 21362 37266
rect 21362 37214 21364 37266
rect 21308 37212 21364 37214
rect 21644 37826 21700 37828
rect 21644 37774 21646 37826
rect 21646 37774 21698 37826
rect 21698 37774 21700 37826
rect 21644 37772 21700 37774
rect 21532 36652 21588 36708
rect 21420 36594 21476 36596
rect 21420 36542 21422 36594
rect 21422 36542 21474 36594
rect 21474 36542 21476 36594
rect 21420 36540 21476 36542
rect 21308 36258 21364 36260
rect 21308 36206 21310 36258
rect 21310 36206 21362 36258
rect 21362 36206 21364 36258
rect 21308 36204 21364 36206
rect 21196 35586 21252 35588
rect 21196 35534 21198 35586
rect 21198 35534 21250 35586
rect 21250 35534 21252 35586
rect 21196 35532 21252 35534
rect 20748 33516 20804 33572
rect 20748 33068 20804 33124
rect 20412 31778 20468 31780
rect 20412 31726 20414 31778
rect 20414 31726 20466 31778
rect 20466 31726 20468 31778
rect 20412 31724 20468 31726
rect 19628 31612 19684 31668
rect 20188 31554 20244 31556
rect 20188 31502 20190 31554
rect 20190 31502 20242 31554
rect 20242 31502 20244 31554
rect 20188 31500 20244 31502
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 18956 30268 19012 30324
rect 19068 30156 19124 30212
rect 18620 28530 18676 28532
rect 18620 28478 18622 28530
rect 18622 28478 18674 28530
rect 18674 28478 18676 28530
rect 18620 28476 18676 28478
rect 18956 29596 19012 29652
rect 19628 30994 19684 30996
rect 19628 30942 19630 30994
rect 19630 30942 19682 30994
rect 19682 30942 19684 30994
rect 19628 30940 19684 30942
rect 19404 30882 19460 30884
rect 19404 30830 19406 30882
rect 19406 30830 19458 30882
rect 19458 30830 19460 30882
rect 19404 30828 19460 30830
rect 20524 30716 20580 30772
rect 20188 30604 20244 30660
rect 21084 34748 21140 34804
rect 21420 34802 21476 34804
rect 21420 34750 21422 34802
rect 21422 34750 21474 34802
rect 21474 34750 21476 34802
rect 21420 34748 21476 34750
rect 21644 35586 21700 35588
rect 21644 35534 21646 35586
rect 21646 35534 21698 35586
rect 21698 35534 21700 35586
rect 21644 35532 21700 35534
rect 21644 34524 21700 34580
rect 21644 34354 21700 34356
rect 21644 34302 21646 34354
rect 21646 34302 21698 34354
rect 21698 34302 21700 34354
rect 21644 34300 21700 34302
rect 20972 32508 21028 32564
rect 21196 33516 21252 33572
rect 21980 37266 22036 37268
rect 21980 37214 21982 37266
rect 21982 37214 22034 37266
rect 22034 37214 22036 37266
rect 21980 37212 22036 37214
rect 22204 37938 22260 37940
rect 22204 37886 22206 37938
rect 22206 37886 22258 37938
rect 22258 37886 22260 37938
rect 22204 37884 22260 37886
rect 22540 37938 22596 37940
rect 22540 37886 22542 37938
rect 22542 37886 22594 37938
rect 22594 37886 22596 37938
rect 22540 37884 22596 37886
rect 22316 37772 22372 37828
rect 22764 37660 22820 37716
rect 22540 37378 22596 37380
rect 22540 37326 22542 37378
rect 22542 37326 22594 37378
rect 22594 37326 22596 37378
rect 22540 37324 22596 37326
rect 23212 38780 23268 38836
rect 23436 40124 23492 40180
rect 23548 38946 23604 38948
rect 23548 38894 23550 38946
rect 23550 38894 23602 38946
rect 23602 38894 23604 38946
rect 23548 38892 23604 38894
rect 23660 38556 23716 38612
rect 22764 36540 22820 36596
rect 22540 35922 22596 35924
rect 22540 35870 22542 35922
rect 22542 35870 22594 35922
rect 22594 35870 22596 35922
rect 22540 35868 22596 35870
rect 22428 35756 22484 35812
rect 22764 36370 22820 36372
rect 22764 36318 22766 36370
rect 22766 36318 22818 36370
rect 22818 36318 22820 36370
rect 22764 36316 22820 36318
rect 22652 35644 22708 35700
rect 22204 35532 22260 35588
rect 22540 35532 22596 35588
rect 22428 35308 22484 35364
rect 21980 34524 22036 34580
rect 21420 33122 21476 33124
rect 21420 33070 21422 33122
rect 21422 33070 21474 33122
rect 21474 33070 21476 33122
rect 21420 33068 21476 33070
rect 21308 32396 21364 32452
rect 20748 32284 20804 32340
rect 21196 31836 21252 31892
rect 20748 31778 20804 31780
rect 20748 31726 20750 31778
rect 20750 31726 20802 31778
rect 20802 31726 20804 31778
rect 20748 31724 20804 31726
rect 21084 31612 21140 31668
rect 21084 31218 21140 31220
rect 21084 31166 21086 31218
rect 21086 31166 21138 31218
rect 21138 31166 21140 31218
rect 21084 31164 21140 31166
rect 21196 31052 21252 31108
rect 20972 30994 21028 30996
rect 20972 30942 20974 30994
rect 20974 30942 21026 30994
rect 21026 30942 21028 30994
rect 20972 30940 21028 30942
rect 19852 30044 19908 30100
rect 19292 29820 19348 29876
rect 19068 28642 19124 28644
rect 19068 28590 19070 28642
rect 19070 28590 19122 28642
rect 19122 28590 19124 28642
rect 19068 28588 19124 28590
rect 19516 28700 19572 28756
rect 19404 28642 19460 28644
rect 19404 28590 19406 28642
rect 19406 28590 19458 28642
rect 19458 28590 19460 28642
rect 19404 28588 19460 28590
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 21196 30268 21252 30324
rect 21308 31164 21364 31220
rect 19964 29484 20020 29540
rect 21644 33292 21700 33348
rect 22204 34300 22260 34356
rect 22092 33516 22148 33572
rect 21756 33234 21812 33236
rect 21756 33182 21758 33234
rect 21758 33182 21810 33234
rect 21810 33182 21812 33234
rect 21756 33180 21812 33182
rect 22652 35196 22708 35252
rect 22652 34130 22708 34132
rect 22652 34078 22654 34130
rect 22654 34078 22706 34130
rect 22706 34078 22708 34130
rect 22652 34076 22708 34078
rect 22652 33740 22708 33796
rect 22092 33068 22148 33124
rect 21644 32060 21700 32116
rect 21980 32450 22036 32452
rect 21980 32398 21982 32450
rect 21982 32398 22034 32450
rect 22034 32398 22036 32450
rect 21980 32396 22036 32398
rect 21868 31836 21924 31892
rect 21980 32060 22036 32116
rect 22204 32508 22260 32564
rect 21868 30716 21924 30772
rect 21532 30210 21588 30212
rect 21532 30158 21534 30210
rect 21534 30158 21586 30210
rect 21586 30158 21588 30210
rect 21532 30156 21588 30158
rect 21308 29596 21364 29652
rect 20524 29484 20580 29540
rect 20860 29538 20916 29540
rect 20860 29486 20862 29538
rect 20862 29486 20914 29538
rect 20914 29486 20916 29538
rect 20860 29484 20916 29486
rect 19964 28588 20020 28644
rect 20300 29260 20356 29316
rect 20636 28700 20692 28756
rect 20188 28476 20244 28532
rect 19628 28140 19684 28196
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 21532 28700 21588 28756
rect 22428 31836 22484 31892
rect 22540 31778 22596 31780
rect 22540 31726 22542 31778
rect 22542 31726 22594 31778
rect 22594 31726 22596 31778
rect 22540 31724 22596 31726
rect 22652 31666 22708 31668
rect 22652 31614 22654 31666
rect 22654 31614 22706 31666
rect 22706 31614 22708 31666
rect 22652 31612 22708 31614
rect 22988 36764 23044 36820
rect 23436 37884 23492 37940
rect 23436 36482 23492 36484
rect 23436 36430 23438 36482
rect 23438 36430 23490 36482
rect 23490 36430 23492 36482
rect 23436 36428 23492 36430
rect 25564 51324 25620 51380
rect 25564 51154 25620 51156
rect 25564 51102 25566 51154
rect 25566 51102 25618 51154
rect 25618 51102 25620 51154
rect 25564 51100 25620 51102
rect 25452 49868 25508 49924
rect 25340 49532 25396 49588
rect 27468 56028 27524 56084
rect 28700 56082 28756 56084
rect 28700 56030 28702 56082
rect 28702 56030 28754 56082
rect 28754 56030 28756 56082
rect 28700 56028 28756 56030
rect 30044 56252 30100 56308
rect 28588 55692 28644 55748
rect 27356 55356 27412 55412
rect 27804 55132 27860 55188
rect 28028 52946 28084 52948
rect 28028 52894 28030 52946
rect 28030 52894 28082 52946
rect 28082 52894 28084 52946
rect 28028 52892 28084 52894
rect 26908 52668 26964 52724
rect 27468 52444 27524 52500
rect 26348 51772 26404 51828
rect 26460 51660 26516 51716
rect 26236 50482 26292 50484
rect 26236 50430 26238 50482
rect 26238 50430 26290 50482
rect 26290 50430 26292 50482
rect 26236 50428 26292 50430
rect 26236 49026 26292 49028
rect 26236 48974 26238 49026
rect 26238 48974 26290 49026
rect 26290 48974 26292 49026
rect 26236 48972 26292 48974
rect 26124 48860 26180 48916
rect 25228 47292 25284 47348
rect 25788 46508 25844 46564
rect 24444 44268 24500 44324
rect 25788 45612 25844 45668
rect 24108 43596 24164 43652
rect 24332 42866 24388 42868
rect 24332 42814 24334 42866
rect 24334 42814 24386 42866
rect 24386 42814 24388 42866
rect 24332 42812 24388 42814
rect 24556 42700 24612 42756
rect 24780 43260 24836 43316
rect 24220 39452 24276 39508
rect 24556 40572 24612 40628
rect 24556 39058 24612 39060
rect 24556 39006 24558 39058
rect 24558 39006 24610 39058
rect 24610 39006 24612 39058
rect 24556 39004 24612 39006
rect 24108 38892 24164 38948
rect 24332 38834 24388 38836
rect 24332 38782 24334 38834
rect 24334 38782 24386 38834
rect 24386 38782 24388 38834
rect 24332 38780 24388 38782
rect 23772 37884 23828 37940
rect 23996 37660 24052 37716
rect 24332 38556 24388 38612
rect 24220 38220 24276 38276
rect 24220 37100 24276 37156
rect 23324 35868 23380 35924
rect 22988 35196 23044 35252
rect 23548 35698 23604 35700
rect 23548 35646 23550 35698
rect 23550 35646 23602 35698
rect 23602 35646 23604 35698
rect 23548 35644 23604 35646
rect 23772 35698 23828 35700
rect 23772 35646 23774 35698
rect 23774 35646 23826 35698
rect 23826 35646 23828 35698
rect 23772 35644 23828 35646
rect 24108 36482 24164 36484
rect 24108 36430 24110 36482
rect 24110 36430 24162 36482
rect 24162 36430 24164 36482
rect 24108 36428 24164 36430
rect 23996 35922 24052 35924
rect 23996 35870 23998 35922
rect 23998 35870 24050 35922
rect 24050 35870 24052 35922
rect 23996 35868 24052 35870
rect 24556 36370 24612 36372
rect 24556 36318 24558 36370
rect 24558 36318 24610 36370
rect 24610 36318 24612 36370
rect 24556 36316 24612 36318
rect 24444 36258 24500 36260
rect 24444 36206 24446 36258
rect 24446 36206 24498 36258
rect 24498 36206 24500 36258
rect 24444 36204 24500 36206
rect 23436 35196 23492 35252
rect 23100 33180 23156 33236
rect 22876 31612 22932 31668
rect 22764 31052 22820 31108
rect 24332 35084 24388 35140
rect 23884 34748 23940 34804
rect 23884 34188 23940 34244
rect 24332 34914 24388 34916
rect 24332 34862 24334 34914
rect 24334 34862 24386 34914
rect 24386 34862 24388 34914
rect 24332 34860 24388 34862
rect 24108 34690 24164 34692
rect 24108 34638 24110 34690
rect 24110 34638 24162 34690
rect 24162 34638 24164 34690
rect 24108 34636 24164 34638
rect 24220 34412 24276 34468
rect 24668 35084 24724 35140
rect 24220 33906 24276 33908
rect 24220 33854 24222 33906
rect 24222 33854 24274 33906
rect 24274 33854 24276 33906
rect 24220 33852 24276 33854
rect 23996 33628 24052 33684
rect 23772 32060 23828 32116
rect 24220 32732 24276 32788
rect 23548 31836 23604 31892
rect 23212 31778 23268 31780
rect 23212 31726 23214 31778
rect 23214 31726 23266 31778
rect 23266 31726 23268 31778
rect 23212 31724 23268 31726
rect 23324 31276 23380 31332
rect 23100 30716 23156 30772
rect 23324 30716 23380 30772
rect 22428 30044 22484 30100
rect 22652 30098 22708 30100
rect 22652 30046 22654 30098
rect 22654 30046 22706 30098
rect 22706 30046 22708 30098
rect 22652 30044 22708 30046
rect 24332 32562 24388 32564
rect 24332 32510 24334 32562
rect 24334 32510 24386 32562
rect 24386 32510 24388 32562
rect 24332 32508 24388 32510
rect 24556 32956 24612 33012
rect 24668 32844 24724 32900
rect 25340 45388 25396 45444
rect 26236 45666 26292 45668
rect 26236 45614 26238 45666
rect 26238 45614 26290 45666
rect 26290 45614 26292 45666
rect 26236 45612 26292 45614
rect 26348 45388 26404 45444
rect 25676 44882 25732 44884
rect 25676 44830 25678 44882
rect 25678 44830 25730 44882
rect 25730 44830 25732 44882
rect 25676 44828 25732 44830
rect 26012 44882 26068 44884
rect 26012 44830 26014 44882
rect 26014 44830 26066 44882
rect 26066 44830 26068 44882
rect 26012 44828 26068 44830
rect 25452 44268 25508 44324
rect 25340 42700 25396 42756
rect 27132 52162 27188 52164
rect 27132 52110 27134 52162
rect 27134 52110 27186 52162
rect 27186 52110 27188 52162
rect 27132 52108 27188 52110
rect 27468 52220 27524 52276
rect 27132 51324 27188 51380
rect 27916 52668 27972 52724
rect 30268 55692 30324 55748
rect 29596 55410 29652 55412
rect 29596 55358 29598 55410
rect 29598 55358 29650 55410
rect 29650 55358 29652 55410
rect 29596 55356 29652 55358
rect 31052 56306 31108 56308
rect 31052 56254 31054 56306
rect 31054 56254 31106 56306
rect 31106 56254 31108 56306
rect 31052 56252 31108 56254
rect 31388 56252 31444 56308
rect 32620 56252 32676 56308
rect 30380 55074 30436 55076
rect 30380 55022 30382 55074
rect 30382 55022 30434 55074
rect 30434 55022 30436 55074
rect 30380 55020 30436 55022
rect 31276 54460 31332 54516
rect 28924 54402 28980 54404
rect 28924 54350 28926 54402
rect 28926 54350 28978 54402
rect 28978 54350 28980 54402
rect 28924 54348 28980 54350
rect 29372 53676 29428 53732
rect 28364 53004 28420 53060
rect 29596 53004 29652 53060
rect 28140 52332 28196 52388
rect 28812 52834 28868 52836
rect 28812 52782 28814 52834
rect 28814 52782 28866 52834
rect 28866 52782 28868 52834
rect 28812 52780 28868 52782
rect 28588 52220 28644 52276
rect 28924 52444 28980 52500
rect 29148 52946 29204 52948
rect 29148 52894 29150 52946
rect 29150 52894 29202 52946
rect 29202 52894 29204 52946
rect 29148 52892 29204 52894
rect 33180 57036 33236 57092
rect 33628 56252 33684 56308
rect 34636 57036 34692 57092
rect 34076 55580 34132 55636
rect 35308 56306 35364 56308
rect 35308 56254 35310 56306
rect 35310 56254 35362 56306
rect 35362 56254 35364 56306
rect 35308 56252 35364 56254
rect 36764 57036 36820 57092
rect 36316 56252 36372 56308
rect 37436 56140 37492 56196
rect 32396 54514 32452 54516
rect 32396 54462 32398 54514
rect 32398 54462 32450 54514
rect 32450 54462 32452 54514
rect 32396 54460 32452 54462
rect 32284 54348 32340 54404
rect 34188 53900 34244 53956
rect 31948 53730 32004 53732
rect 31948 53678 31950 53730
rect 31950 53678 32002 53730
rect 32002 53678 32004 53730
rect 31948 53676 32004 53678
rect 33180 53676 33236 53732
rect 29932 53004 29988 53060
rect 30716 53058 30772 53060
rect 30716 53006 30718 53058
rect 30718 53006 30770 53058
rect 30770 53006 30772 53058
rect 30716 53004 30772 53006
rect 30268 52780 30324 52836
rect 29820 52722 29876 52724
rect 29820 52670 29822 52722
rect 29822 52670 29874 52722
rect 29874 52670 29876 52722
rect 29820 52668 29876 52670
rect 28924 52220 28980 52276
rect 30044 52386 30100 52388
rect 30044 52334 30046 52386
rect 30046 52334 30098 52386
rect 30098 52334 30100 52386
rect 30044 52332 30100 52334
rect 27804 52108 27860 52164
rect 28924 51602 28980 51604
rect 28924 51550 28926 51602
rect 28926 51550 28978 51602
rect 28978 51550 28980 51602
rect 28924 51548 28980 51550
rect 28700 51490 28756 51492
rect 28700 51438 28702 51490
rect 28702 51438 28754 51490
rect 28754 51438 28756 51490
rect 28700 51436 28756 51438
rect 27916 51324 27972 51380
rect 26796 50594 26852 50596
rect 26796 50542 26798 50594
rect 26798 50542 26850 50594
rect 26850 50542 26852 50594
rect 26796 50540 26852 50542
rect 27132 50428 27188 50484
rect 26684 49868 26740 49924
rect 26796 49756 26852 49812
rect 26572 49420 26628 49476
rect 26572 49250 26628 49252
rect 26572 49198 26574 49250
rect 26574 49198 26626 49250
rect 26626 49198 26628 49250
rect 26572 49196 26628 49198
rect 27468 51100 27524 51156
rect 27468 50818 27524 50820
rect 27468 50766 27470 50818
rect 27470 50766 27522 50818
rect 27522 50766 27524 50818
rect 27468 50764 27524 50766
rect 27356 50316 27412 50372
rect 27692 50540 27748 50596
rect 27580 49922 27636 49924
rect 27580 49870 27582 49922
rect 27582 49870 27634 49922
rect 27634 49870 27636 49922
rect 27580 49868 27636 49870
rect 27132 49196 27188 49252
rect 27356 49532 27412 49588
rect 27356 49308 27412 49364
rect 26908 48860 26964 48916
rect 27244 48748 27300 48804
rect 27020 48354 27076 48356
rect 27020 48302 27022 48354
rect 27022 48302 27074 48354
rect 27074 48302 27076 48354
rect 27020 48300 27076 48302
rect 27468 48972 27524 49028
rect 27804 49532 27860 49588
rect 28140 50818 28196 50820
rect 28140 50766 28142 50818
rect 28142 50766 28194 50818
rect 28194 50766 28196 50818
rect 28140 50764 28196 50766
rect 28252 50594 28308 50596
rect 28252 50542 28254 50594
rect 28254 50542 28306 50594
rect 28306 50542 28308 50594
rect 28252 50540 28308 50542
rect 28028 49922 28084 49924
rect 28028 49870 28030 49922
rect 28030 49870 28082 49922
rect 28082 49870 28084 49922
rect 28028 49868 28084 49870
rect 28140 49756 28196 49812
rect 27692 48412 27748 48468
rect 27468 48300 27524 48356
rect 29148 52162 29204 52164
rect 29148 52110 29150 52162
rect 29150 52110 29202 52162
rect 29202 52110 29204 52162
rect 29148 52108 29204 52110
rect 28476 50706 28532 50708
rect 28476 50654 28478 50706
rect 28478 50654 28530 50706
rect 28530 50654 28532 50706
rect 28476 50652 28532 50654
rect 28364 50316 28420 50372
rect 28812 50540 28868 50596
rect 28924 49810 28980 49812
rect 28924 49758 28926 49810
rect 28926 49758 28978 49810
rect 28978 49758 28980 49810
rect 28924 49756 28980 49758
rect 28700 49308 28756 49364
rect 28812 49420 28868 49476
rect 28364 49196 28420 49252
rect 28588 49138 28644 49140
rect 28588 49086 28590 49138
rect 28590 49086 28642 49138
rect 28642 49086 28644 49138
rect 28588 49084 28644 49086
rect 28252 49026 28308 49028
rect 28252 48974 28254 49026
rect 28254 48974 28306 49026
rect 28306 48974 28308 49026
rect 28252 48972 28308 48974
rect 28812 48860 28868 48916
rect 29036 49308 29092 49364
rect 28476 48802 28532 48804
rect 28476 48750 28478 48802
rect 28478 48750 28530 48802
rect 28530 48750 28532 48802
rect 28476 48748 28532 48750
rect 28252 48354 28308 48356
rect 28252 48302 28254 48354
rect 28254 48302 28306 48354
rect 28306 48302 28308 48354
rect 28252 48300 28308 48302
rect 28588 48300 28644 48356
rect 29372 49980 29428 50036
rect 31276 52668 31332 52724
rect 29596 51212 29652 51268
rect 29708 51548 29764 51604
rect 30604 51548 30660 51604
rect 30268 51212 30324 51268
rect 30268 50764 30324 50820
rect 29932 50652 29988 50708
rect 29820 50428 29876 50484
rect 29372 49810 29428 49812
rect 29372 49758 29374 49810
rect 29374 49758 29426 49810
rect 29426 49758 29428 49810
rect 29372 49756 29428 49758
rect 29596 49420 29652 49476
rect 29260 49250 29316 49252
rect 29260 49198 29262 49250
rect 29262 49198 29314 49250
rect 29314 49198 29316 49250
rect 29260 49196 29316 49198
rect 29148 49084 29204 49140
rect 29932 49980 29988 50036
rect 29372 48972 29428 49028
rect 30044 49644 30100 49700
rect 29260 48802 29316 48804
rect 29260 48750 29262 48802
rect 29262 48750 29314 48802
rect 29314 48750 29316 48802
rect 29260 48748 29316 48750
rect 30492 50482 30548 50484
rect 30492 50430 30494 50482
rect 30494 50430 30546 50482
rect 30546 50430 30548 50482
rect 30492 50428 30548 50430
rect 30380 49756 30436 49812
rect 31276 50652 31332 50708
rect 30716 49756 30772 49812
rect 33292 52220 33348 52276
rect 33404 52108 33460 52164
rect 32284 51938 32340 51940
rect 32284 51886 32286 51938
rect 32286 51886 32338 51938
rect 32338 51886 32340 51938
rect 32284 51884 32340 51886
rect 33180 51884 33236 51940
rect 31948 50764 32004 50820
rect 31836 50706 31892 50708
rect 31836 50654 31838 50706
rect 31838 50654 31890 50706
rect 31890 50654 31892 50706
rect 31836 50652 31892 50654
rect 32172 50594 32228 50596
rect 32172 50542 32174 50594
rect 32174 50542 32226 50594
rect 32226 50542 32228 50594
rect 32172 50540 32228 50542
rect 31164 49868 31220 49924
rect 31052 49644 31108 49700
rect 31164 49532 31220 49588
rect 31052 49420 31108 49476
rect 30268 49196 30324 49252
rect 30940 49196 30996 49252
rect 30828 49138 30884 49140
rect 30828 49086 30830 49138
rect 30830 49086 30882 49138
rect 30882 49086 30884 49138
rect 30828 49084 30884 49086
rect 29708 48802 29764 48804
rect 29708 48750 29710 48802
rect 29710 48750 29762 48802
rect 29762 48750 29764 48802
rect 29708 48748 29764 48750
rect 30604 48802 30660 48804
rect 30604 48750 30606 48802
rect 30606 48750 30658 48802
rect 30658 48750 30660 48802
rect 30604 48748 30660 48750
rect 30156 48636 30212 48692
rect 30828 48636 30884 48692
rect 29820 48188 29876 48244
rect 31052 48412 31108 48468
rect 31276 49308 31332 49364
rect 31388 50092 31444 50148
rect 31836 50370 31892 50372
rect 31836 50318 31838 50370
rect 31838 50318 31890 50370
rect 31890 50318 31892 50370
rect 31836 50316 31892 50318
rect 31612 49868 31668 49924
rect 31724 49420 31780 49476
rect 31836 49756 31892 49812
rect 31612 49308 31668 49364
rect 31612 48972 31668 49028
rect 31612 48242 31668 48244
rect 31612 48190 31614 48242
rect 31614 48190 31666 48242
rect 31666 48190 31668 48242
rect 31612 48188 31668 48190
rect 32284 50204 32340 50260
rect 34076 52274 34132 52276
rect 34076 52222 34078 52274
rect 34078 52222 34130 52274
rect 34130 52222 34132 52274
rect 34076 52220 34132 52222
rect 33852 52108 33908 52164
rect 33068 50652 33124 50708
rect 33404 50764 33460 50820
rect 32508 50370 32564 50372
rect 32508 50318 32510 50370
rect 32510 50318 32562 50370
rect 32562 50318 32564 50370
rect 32508 50316 32564 50318
rect 32396 50092 32452 50148
rect 33180 50316 33236 50372
rect 33292 50428 33348 50484
rect 32284 49868 32340 49924
rect 32060 49420 32116 49476
rect 32172 49644 32228 49700
rect 32732 49644 32788 49700
rect 32732 49026 32788 49028
rect 32732 48974 32734 49026
rect 32734 48974 32786 49026
rect 32786 48974 32788 49026
rect 32732 48972 32788 48974
rect 33852 51602 33908 51604
rect 33852 51550 33854 51602
rect 33854 51550 33906 51602
rect 33906 51550 33908 51602
rect 33852 51548 33908 51550
rect 35196 55690 35252 55692
rect 34972 55580 35028 55636
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 34860 55132 34916 55188
rect 35756 54514 35812 54516
rect 35756 54462 35758 54514
rect 35758 54462 35810 54514
rect 35810 54462 35812 54514
rect 35756 54460 35812 54462
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35756 53788 35812 53844
rect 35980 53788 36036 53844
rect 34300 52556 34356 52612
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34972 52274 35028 52276
rect 34972 52222 34974 52274
rect 34974 52222 35026 52274
rect 35026 52222 35028 52274
rect 34972 52220 35028 52222
rect 36204 55186 36260 55188
rect 36204 55134 36206 55186
rect 36206 55134 36258 55186
rect 36258 55134 36260 55186
rect 36204 55132 36260 55134
rect 37100 54460 37156 54516
rect 37100 53842 37156 53844
rect 37100 53790 37102 53842
rect 37102 53790 37154 53842
rect 37154 53790 37156 53842
rect 37100 53788 37156 53790
rect 36428 53004 36484 53060
rect 35644 52220 35700 52276
rect 34300 50482 34356 50484
rect 34300 50430 34302 50482
rect 34302 50430 34354 50482
rect 34354 50430 34356 50482
rect 34300 50428 34356 50430
rect 35084 51324 35140 51380
rect 34188 49698 34244 49700
rect 34188 49646 34190 49698
rect 34190 49646 34242 49698
rect 34242 49646 34244 49698
rect 34188 49644 34244 49646
rect 31948 48354 32004 48356
rect 31948 48302 31950 48354
rect 31950 48302 32002 48354
rect 32002 48302 32004 48354
rect 31948 48300 32004 48302
rect 32956 48076 33012 48132
rect 32956 47180 33012 47236
rect 27356 46562 27412 46564
rect 27356 46510 27358 46562
rect 27358 46510 27410 46562
rect 27410 46510 27412 46562
rect 27356 46508 27412 46510
rect 30156 46620 30212 46676
rect 27916 45948 27972 46004
rect 26684 45666 26740 45668
rect 26684 45614 26686 45666
rect 26686 45614 26738 45666
rect 26738 45614 26740 45666
rect 26684 45612 26740 45614
rect 27580 44828 27636 44884
rect 27244 43650 27300 43652
rect 27244 43598 27246 43650
rect 27246 43598 27298 43650
rect 27298 43598 27300 43650
rect 27244 43596 27300 43598
rect 29820 45948 29876 46004
rect 28924 45612 28980 45668
rect 28700 44044 28756 44100
rect 29260 44994 29316 44996
rect 29260 44942 29262 44994
rect 29262 44942 29314 44994
rect 29314 44942 29316 44994
rect 29260 44940 29316 44942
rect 29260 44098 29316 44100
rect 29260 44046 29262 44098
rect 29262 44046 29314 44098
rect 29314 44046 29316 44098
rect 29260 44044 29316 44046
rect 27132 43484 27188 43540
rect 26460 42252 26516 42308
rect 28700 43650 28756 43652
rect 28700 43598 28702 43650
rect 28702 43598 28754 43650
rect 28754 43598 28756 43650
rect 28700 43596 28756 43598
rect 28588 43484 28644 43540
rect 25676 40460 25732 40516
rect 26348 39900 26404 39956
rect 26460 40348 26516 40404
rect 26572 40236 26628 40292
rect 26572 39900 26628 39956
rect 25228 39452 25284 39508
rect 26236 39228 26292 39284
rect 25228 39116 25284 39172
rect 25340 38834 25396 38836
rect 25340 38782 25342 38834
rect 25342 38782 25394 38834
rect 25394 38782 25396 38834
rect 25340 38780 25396 38782
rect 25228 38668 25284 38724
rect 24892 38220 24948 38276
rect 24892 35644 24948 35700
rect 24892 35308 24948 35364
rect 24892 34748 24948 34804
rect 24780 32732 24836 32788
rect 25676 37548 25732 37604
rect 27580 40236 27636 40292
rect 27916 41804 27972 41860
rect 28812 41858 28868 41860
rect 28812 41806 28814 41858
rect 28814 41806 28866 41858
rect 28866 41806 28868 41858
rect 28812 41804 28868 41806
rect 28588 41186 28644 41188
rect 28588 41134 28590 41186
rect 28590 41134 28642 41186
rect 28642 41134 28644 41186
rect 28588 41132 28644 41134
rect 29148 41916 29204 41972
rect 30828 46620 30884 46676
rect 30380 44380 30436 44436
rect 30492 43650 30548 43652
rect 30492 43598 30494 43650
rect 30494 43598 30546 43650
rect 30546 43598 30548 43650
rect 30492 43596 30548 43598
rect 31388 46674 31444 46676
rect 31388 46622 31390 46674
rect 31390 46622 31442 46674
rect 31442 46622 31444 46674
rect 31388 46620 31444 46622
rect 31052 46562 31108 46564
rect 31052 46510 31054 46562
rect 31054 46510 31106 46562
rect 31106 46510 31108 46562
rect 31052 46508 31108 46510
rect 32060 46508 32116 46564
rect 31724 46060 31780 46116
rect 32396 46450 32452 46452
rect 32396 46398 32398 46450
rect 32398 46398 32450 46450
rect 32450 46398 32452 46450
rect 32396 46396 32452 46398
rect 31948 45890 32004 45892
rect 31948 45838 31950 45890
rect 31950 45838 32002 45890
rect 32002 45838 32004 45890
rect 31948 45836 32004 45838
rect 31052 45612 31108 45668
rect 31388 44940 31444 44996
rect 31388 44322 31444 44324
rect 31388 44270 31390 44322
rect 31390 44270 31442 44322
rect 31442 44270 31444 44322
rect 31388 44268 31444 44270
rect 32172 44322 32228 44324
rect 32172 44270 32174 44322
rect 32174 44270 32226 44322
rect 32226 44270 32228 44322
rect 32172 44268 32228 44270
rect 32508 44268 32564 44324
rect 31052 44156 31108 44212
rect 31948 43596 32004 43652
rect 30716 42700 30772 42756
rect 30828 41916 30884 41972
rect 29260 41186 29316 41188
rect 29260 41134 29262 41186
rect 29262 41134 29314 41186
rect 29314 41134 29316 41186
rect 29260 41132 29316 41134
rect 27804 40348 27860 40404
rect 26684 39004 26740 39060
rect 26796 39228 26852 39284
rect 26572 38892 26628 38948
rect 26348 38780 26404 38836
rect 26236 38668 26292 38724
rect 27692 39116 27748 39172
rect 27132 38892 27188 38948
rect 27468 38834 27524 38836
rect 27468 38782 27470 38834
rect 27470 38782 27522 38834
rect 27522 38782 27524 38834
rect 27468 38780 27524 38782
rect 27580 38556 27636 38612
rect 26348 37548 26404 37604
rect 26684 37772 26740 37828
rect 26236 36764 26292 36820
rect 25676 36316 25732 36372
rect 25340 34690 25396 34692
rect 25340 34638 25342 34690
rect 25342 34638 25394 34690
rect 25394 34638 25396 34690
rect 25340 34636 25396 34638
rect 27804 37938 27860 37940
rect 27804 37886 27806 37938
rect 27806 37886 27858 37938
rect 27858 37886 27860 37938
rect 27804 37884 27860 37886
rect 26796 36652 26852 36708
rect 26908 36764 26964 36820
rect 26460 36482 26516 36484
rect 26460 36430 26462 36482
rect 26462 36430 26514 36482
rect 26514 36430 26516 36482
rect 26460 36428 26516 36430
rect 26796 36370 26852 36372
rect 26796 36318 26798 36370
rect 26798 36318 26850 36370
rect 26850 36318 26852 36370
rect 26796 36316 26852 36318
rect 26684 36092 26740 36148
rect 25676 35084 25732 35140
rect 26236 35868 26292 35924
rect 25900 35084 25956 35140
rect 25676 34914 25732 34916
rect 25676 34862 25678 34914
rect 25678 34862 25730 34914
rect 25730 34862 25732 34914
rect 25676 34860 25732 34862
rect 26012 34860 26068 34916
rect 26012 34636 26068 34692
rect 25676 34188 25732 34244
rect 25116 33346 25172 33348
rect 25116 33294 25118 33346
rect 25118 33294 25170 33346
rect 25170 33294 25172 33346
rect 25116 33292 25172 33294
rect 26796 35810 26852 35812
rect 26796 35758 26798 35810
rect 26798 35758 26850 35810
rect 26850 35758 26852 35810
rect 26796 35756 26852 35758
rect 26460 34914 26516 34916
rect 26460 34862 26462 34914
rect 26462 34862 26514 34914
rect 26514 34862 26516 34914
rect 26460 34860 26516 34862
rect 26012 33852 26068 33908
rect 24556 31948 24612 32004
rect 24780 32508 24836 32564
rect 23548 30156 23604 30212
rect 22540 29260 22596 29316
rect 24556 31388 24612 31444
rect 23996 30940 24052 30996
rect 24444 31276 24500 31332
rect 24332 30770 24388 30772
rect 24332 30718 24334 30770
rect 24334 30718 24386 30770
rect 24386 30718 24388 30770
rect 24332 30716 24388 30718
rect 24220 30604 24276 30660
rect 25452 33068 25508 33124
rect 25116 32508 25172 32564
rect 25228 32844 25284 32900
rect 25004 32396 25060 32452
rect 24892 31164 24948 31220
rect 25004 31388 25060 31444
rect 24892 30716 24948 30772
rect 24892 30268 24948 30324
rect 26236 33180 26292 33236
rect 25676 33068 25732 33124
rect 25452 32620 25508 32676
rect 25340 31724 25396 31780
rect 25340 31164 25396 31220
rect 25788 32562 25844 32564
rect 25788 32510 25790 32562
rect 25790 32510 25842 32562
rect 25842 32510 25844 32562
rect 25788 32508 25844 32510
rect 25900 31948 25956 32004
rect 25900 31724 25956 31780
rect 25788 31388 25844 31444
rect 26124 32508 26180 32564
rect 25228 30210 25284 30212
rect 25228 30158 25230 30210
rect 25230 30158 25282 30210
rect 25282 30158 25284 30210
rect 25228 30156 25284 30158
rect 27020 36092 27076 36148
rect 27244 37100 27300 37156
rect 26796 34860 26852 34916
rect 27132 34914 27188 34916
rect 27132 34862 27134 34914
rect 27134 34862 27186 34914
rect 27186 34862 27188 34914
rect 27132 34860 27188 34862
rect 27580 37378 27636 37380
rect 27580 37326 27582 37378
rect 27582 37326 27634 37378
rect 27634 37326 27636 37378
rect 27580 37324 27636 37326
rect 27804 37324 27860 37380
rect 27580 36428 27636 36484
rect 27804 36258 27860 36260
rect 27804 36206 27806 36258
rect 27806 36206 27858 36258
rect 27858 36206 27860 36258
rect 27804 36204 27860 36206
rect 27804 35980 27860 36036
rect 26908 34690 26964 34692
rect 26908 34638 26910 34690
rect 26910 34638 26962 34690
rect 26962 34638 26964 34690
rect 26908 34636 26964 34638
rect 26908 34242 26964 34244
rect 26908 34190 26910 34242
rect 26910 34190 26962 34242
rect 26962 34190 26964 34242
rect 26908 34188 26964 34190
rect 26796 33740 26852 33796
rect 27020 33852 27076 33908
rect 26908 33628 26964 33684
rect 27804 35532 27860 35588
rect 28028 39788 28084 39844
rect 28028 39618 28084 39620
rect 28028 39566 28030 39618
rect 28030 39566 28082 39618
rect 28082 39566 28084 39618
rect 28028 39564 28084 39566
rect 28028 39116 28084 39172
rect 28924 38946 28980 38948
rect 28924 38894 28926 38946
rect 28926 38894 28978 38946
rect 28978 38894 28980 38946
rect 28924 38892 28980 38894
rect 28364 38556 28420 38612
rect 28588 37996 28644 38052
rect 28364 37938 28420 37940
rect 28364 37886 28366 37938
rect 28366 37886 28418 37938
rect 28418 37886 28420 37938
rect 28364 37884 28420 37886
rect 28252 37490 28308 37492
rect 28252 37438 28254 37490
rect 28254 37438 28306 37490
rect 28306 37438 28308 37490
rect 28252 37436 28308 37438
rect 29260 37938 29316 37940
rect 29260 37886 29262 37938
rect 29262 37886 29314 37938
rect 29314 37886 29316 37938
rect 29260 37884 29316 37886
rect 29148 37436 29204 37492
rect 28588 36428 28644 36484
rect 28588 35698 28644 35700
rect 28588 35646 28590 35698
rect 28590 35646 28642 35698
rect 28642 35646 28644 35698
rect 28588 35644 28644 35646
rect 28252 35308 28308 35364
rect 27804 34690 27860 34692
rect 27804 34638 27806 34690
rect 27806 34638 27858 34690
rect 27858 34638 27860 34690
rect 27804 34636 27860 34638
rect 27580 33852 27636 33908
rect 27468 33346 27524 33348
rect 27468 33294 27470 33346
rect 27470 33294 27522 33346
rect 27522 33294 27524 33346
rect 27468 33292 27524 33294
rect 27356 33234 27412 33236
rect 27356 33182 27358 33234
rect 27358 33182 27410 33234
rect 27410 33182 27412 33234
rect 27356 33180 27412 33182
rect 27804 33516 27860 33572
rect 27692 33404 27748 33460
rect 27692 33180 27748 33236
rect 26236 31666 26292 31668
rect 26236 31614 26238 31666
rect 26238 31614 26290 31666
rect 26290 31614 26292 31666
rect 26236 31612 26292 31614
rect 23660 29538 23716 29540
rect 23660 29486 23662 29538
rect 23662 29486 23714 29538
rect 23714 29486 23716 29538
rect 23660 29484 23716 29486
rect 25228 29260 25284 29316
rect 26572 31554 26628 31556
rect 26572 31502 26574 31554
rect 26574 31502 26626 31554
rect 26626 31502 26628 31554
rect 26572 31500 26628 31502
rect 26460 31164 26516 31220
rect 26348 30156 26404 30212
rect 27020 32732 27076 32788
rect 27020 31724 27076 31780
rect 27356 31724 27412 31780
rect 27804 32732 27860 32788
rect 28028 33404 28084 33460
rect 27692 32674 27748 32676
rect 27692 32622 27694 32674
rect 27694 32622 27746 32674
rect 27746 32622 27748 32674
rect 27692 32620 27748 32622
rect 27132 31276 27188 31332
rect 26684 30268 26740 30324
rect 25340 29484 25396 29540
rect 24444 29148 24500 29204
rect 21420 28476 21476 28532
rect 22428 28530 22484 28532
rect 22428 28478 22430 28530
rect 22430 28478 22482 28530
rect 22482 28478 22484 28530
rect 22428 28476 22484 28478
rect 23324 28530 23380 28532
rect 23324 28478 23326 28530
rect 23326 28478 23378 28530
rect 23378 28478 23380 28530
rect 23324 28476 23380 28478
rect 21868 28418 21924 28420
rect 21868 28366 21870 28418
rect 21870 28366 21922 28418
rect 21922 28366 21924 28418
rect 21868 28364 21924 28366
rect 22540 28252 22596 28308
rect 23324 28252 23380 28308
rect 22876 27804 22932 27860
rect 17836 27020 17892 27076
rect 18060 26908 18116 26964
rect 17836 26796 17892 26852
rect 14812 24556 14868 24612
rect 16716 26290 16772 26292
rect 16716 26238 16718 26290
rect 16718 26238 16770 26290
rect 16770 26238 16772 26290
rect 16716 26236 16772 26238
rect 17388 26236 17444 26292
rect 16604 26178 16660 26180
rect 16604 26126 16606 26178
rect 16606 26126 16658 26178
rect 16658 26126 16660 26178
rect 16604 26124 16660 26126
rect 16044 25282 16100 25284
rect 16044 25230 16046 25282
rect 16046 25230 16098 25282
rect 16098 25230 16100 25282
rect 16044 25228 16100 25230
rect 16044 24668 16100 24724
rect 14028 24050 14084 24052
rect 14028 23998 14030 24050
rect 14030 23998 14082 24050
rect 14082 23998 14084 24050
rect 14028 23996 14084 23998
rect 13804 22482 13860 22484
rect 13804 22430 13806 22482
rect 13806 22430 13858 22482
rect 13858 22430 13860 22482
rect 13804 22428 13860 22430
rect 14140 23324 14196 23380
rect 14476 23826 14532 23828
rect 14476 23774 14478 23826
rect 14478 23774 14530 23826
rect 14530 23774 14532 23826
rect 14476 23772 14532 23774
rect 14140 22316 14196 22372
rect 14252 22540 14308 22596
rect 11676 21868 11732 21924
rect 14028 21868 14084 21924
rect 11340 21756 11396 21812
rect 12124 21756 12180 21812
rect 12012 21420 12068 21476
rect 11340 20578 11396 20580
rect 11340 20526 11342 20578
rect 11342 20526 11394 20578
rect 11394 20526 11396 20578
rect 11340 20524 11396 20526
rect 11228 20412 11284 20468
rect 12460 20914 12516 20916
rect 12460 20862 12462 20914
rect 12462 20862 12514 20914
rect 12514 20862 12516 20914
rect 12460 20860 12516 20862
rect 13020 21474 13076 21476
rect 13020 21422 13022 21474
rect 13022 21422 13074 21474
rect 13074 21422 13076 21474
rect 13020 21420 13076 21422
rect 13468 21308 13524 21364
rect 13468 20860 13524 20916
rect 12012 20412 12068 20468
rect 7420 18396 7476 18452
rect 8428 18396 8484 18452
rect 7868 18172 7924 18228
rect 9660 18450 9716 18452
rect 9660 18398 9662 18450
rect 9662 18398 9714 18450
rect 9714 18398 9716 18450
rect 9660 18396 9716 18398
rect 13356 20076 13412 20132
rect 14028 20802 14084 20804
rect 14028 20750 14030 20802
rect 14030 20750 14082 20802
rect 14082 20750 14084 20802
rect 14028 20748 14084 20750
rect 14252 21420 14308 21476
rect 15820 23938 15876 23940
rect 15820 23886 15822 23938
rect 15822 23886 15874 23938
rect 15874 23886 15876 23938
rect 15820 23884 15876 23886
rect 16156 24332 16212 24388
rect 16492 24332 16548 24388
rect 16044 23996 16100 24052
rect 16268 24108 16324 24164
rect 15932 23772 15988 23828
rect 15148 22540 15204 22596
rect 15708 22370 15764 22372
rect 15708 22318 15710 22370
rect 15710 22318 15762 22370
rect 15762 22318 15764 22370
rect 15708 22316 15764 22318
rect 15484 22092 15540 22148
rect 14812 21532 14868 21588
rect 14588 21308 14644 21364
rect 16268 21644 16324 21700
rect 15820 21532 15876 21588
rect 15148 21196 15204 21252
rect 14924 20914 14980 20916
rect 14924 20862 14926 20914
rect 14926 20862 14978 20914
rect 14978 20862 14980 20914
rect 14924 20860 14980 20862
rect 13580 20412 13636 20468
rect 15372 20412 15428 20468
rect 14924 20076 14980 20132
rect 12348 20018 12404 20020
rect 12348 19966 12350 20018
rect 12350 19966 12402 20018
rect 12402 19966 12404 20018
rect 12348 19964 12404 19966
rect 12124 19458 12180 19460
rect 12124 19406 12126 19458
rect 12126 19406 12178 19458
rect 12178 19406 12180 19458
rect 12124 19404 12180 19406
rect 15148 19516 15204 19572
rect 12124 18956 12180 19012
rect 10668 18396 10724 18452
rect 10780 18226 10836 18228
rect 10780 18174 10782 18226
rect 10782 18174 10834 18226
rect 10834 18174 10836 18226
rect 10780 18172 10836 18174
rect 8876 18060 8932 18116
rect 11116 17836 11172 17892
rect 9884 16268 9940 16324
rect 11564 17052 11620 17108
rect 11228 16322 11284 16324
rect 11228 16270 11230 16322
rect 11230 16270 11282 16322
rect 11282 16270 11284 16322
rect 11228 16268 11284 16270
rect 11788 16268 11844 16324
rect 8876 15484 8932 15540
rect 7980 15148 8036 15204
rect 8540 15148 8596 15204
rect 11900 17164 11956 17220
rect 12012 18396 12068 18452
rect 12348 18450 12404 18452
rect 12348 18398 12350 18450
rect 12350 18398 12402 18450
rect 12402 18398 12404 18450
rect 12348 18396 12404 18398
rect 12460 17778 12516 17780
rect 12460 17726 12462 17778
rect 12462 17726 12514 17778
rect 12514 17726 12516 17778
rect 12460 17724 12516 17726
rect 14476 18956 14532 19012
rect 14476 17890 14532 17892
rect 14476 17838 14478 17890
rect 14478 17838 14530 17890
rect 14530 17838 14532 17890
rect 14476 17836 14532 17838
rect 14588 17442 14644 17444
rect 14588 17390 14590 17442
rect 14590 17390 14642 17442
rect 14642 17390 14644 17442
rect 14588 17388 14644 17390
rect 13132 16882 13188 16884
rect 13132 16830 13134 16882
rect 13134 16830 13186 16882
rect 13186 16830 13188 16882
rect 13132 16828 13188 16830
rect 9660 15202 9716 15204
rect 9660 15150 9662 15202
rect 9662 15150 9714 15202
rect 9714 15150 9716 15202
rect 9660 15148 9716 15150
rect 10444 15148 10500 15204
rect 11900 15148 11956 15204
rect 9884 13746 9940 13748
rect 9884 13694 9886 13746
rect 9886 13694 9938 13746
rect 9938 13694 9940 13746
rect 9884 13692 9940 13694
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 8988 13468 9044 13524
rect 11116 13746 11172 13748
rect 11116 13694 11118 13746
rect 11118 13694 11170 13746
rect 11170 13694 11172 13746
rect 11116 13692 11172 13694
rect 10220 13468 10276 13524
rect 12796 16716 12852 16772
rect 14700 16322 14756 16324
rect 14700 16270 14702 16322
rect 14702 16270 14754 16322
rect 14754 16270 14756 16322
rect 14700 16268 14756 16270
rect 13804 15932 13860 15988
rect 12796 15148 12852 15204
rect 15036 17276 15092 17332
rect 14924 16770 14980 16772
rect 14924 16718 14926 16770
rect 14926 16718 14978 16770
rect 14978 16718 14980 16770
rect 14924 16716 14980 16718
rect 15036 16268 15092 16324
rect 16380 21474 16436 21476
rect 16380 21422 16382 21474
rect 16382 21422 16434 21474
rect 16434 21422 16436 21474
rect 16380 21420 16436 21422
rect 16268 21196 16324 21252
rect 16828 24834 16884 24836
rect 16828 24782 16830 24834
rect 16830 24782 16882 24834
rect 16882 24782 16884 24834
rect 16828 24780 16884 24782
rect 23436 27858 23492 27860
rect 23436 27806 23438 27858
rect 23438 27806 23490 27858
rect 23490 27806 23492 27858
rect 23436 27804 23492 27806
rect 25452 29314 25508 29316
rect 25452 29262 25454 29314
rect 25454 29262 25506 29314
rect 25506 29262 25508 29314
rect 25452 29260 25508 29262
rect 25900 29314 25956 29316
rect 25900 29262 25902 29314
rect 25902 29262 25954 29314
rect 25954 29262 25956 29314
rect 25900 29260 25956 29262
rect 26908 29426 26964 29428
rect 26908 29374 26910 29426
rect 26910 29374 26962 29426
rect 26962 29374 26964 29426
rect 26908 29372 26964 29374
rect 26460 29260 26516 29316
rect 27244 29596 27300 29652
rect 27468 31388 27524 31444
rect 27916 31778 27972 31780
rect 27916 31726 27918 31778
rect 27918 31726 27970 31778
rect 27970 31726 27972 31778
rect 27916 31724 27972 31726
rect 28028 31388 28084 31444
rect 28588 35084 28644 35140
rect 29260 36652 29316 36708
rect 29148 35980 29204 36036
rect 29260 35644 29316 35700
rect 28924 35308 28980 35364
rect 28812 34860 28868 34916
rect 30044 39058 30100 39060
rect 30044 39006 30046 39058
rect 30046 39006 30098 39058
rect 30098 39006 30100 39058
rect 30044 39004 30100 39006
rect 29708 38946 29764 38948
rect 29708 38894 29710 38946
rect 29710 38894 29762 38946
rect 29762 38894 29764 38946
rect 29708 38892 29764 38894
rect 30044 38050 30100 38052
rect 30044 37998 30046 38050
rect 30046 37998 30098 38050
rect 30098 37998 30100 38050
rect 30044 37996 30100 37998
rect 29596 36482 29652 36484
rect 29596 36430 29598 36482
rect 29598 36430 29650 36482
rect 29650 36430 29652 36482
rect 29596 36428 29652 36430
rect 29820 35698 29876 35700
rect 29820 35646 29822 35698
rect 29822 35646 29874 35698
rect 29874 35646 29876 35698
rect 29820 35644 29876 35646
rect 30492 40460 30548 40516
rect 30268 39676 30324 39732
rect 30044 36482 30100 36484
rect 30044 36430 30046 36482
rect 30046 36430 30098 36482
rect 30098 36430 30100 36482
rect 30044 36428 30100 36430
rect 30716 39618 30772 39620
rect 30716 39566 30718 39618
rect 30718 39566 30770 39618
rect 30770 39566 30772 39618
rect 30716 39564 30772 39566
rect 30828 39340 30884 39396
rect 32844 43484 32900 43540
rect 31276 42476 31332 42532
rect 31164 41916 31220 41972
rect 31052 40348 31108 40404
rect 31164 40236 31220 40292
rect 31164 39676 31220 39732
rect 31052 39394 31108 39396
rect 31052 39342 31054 39394
rect 31054 39342 31106 39394
rect 31106 39342 31108 39394
rect 31052 39340 31108 39342
rect 30940 39058 30996 39060
rect 30940 39006 30942 39058
rect 30942 39006 30994 39058
rect 30994 39006 30996 39058
rect 30940 39004 30996 39006
rect 32508 42140 32564 42196
rect 31724 41186 31780 41188
rect 31724 41134 31726 41186
rect 31726 41134 31778 41186
rect 31778 41134 31780 41186
rect 31724 41132 31780 41134
rect 31612 39340 31668 39396
rect 31612 39116 31668 39172
rect 30380 38556 30436 38612
rect 30940 37996 30996 38052
rect 30268 36258 30324 36260
rect 30268 36206 30270 36258
rect 30270 36206 30322 36258
rect 30322 36206 30324 36258
rect 30268 36204 30324 36206
rect 29932 35532 29988 35588
rect 29484 35084 29540 35140
rect 28588 33964 28644 34020
rect 28364 33852 28420 33908
rect 28252 33180 28308 33236
rect 28476 33628 28532 33684
rect 28812 33516 28868 33572
rect 28588 32562 28644 32564
rect 28588 32510 28590 32562
rect 28590 32510 28642 32562
rect 28642 32510 28644 32562
rect 28588 32508 28644 32510
rect 28252 31724 28308 31780
rect 29148 34914 29204 34916
rect 29148 34862 29150 34914
rect 29150 34862 29202 34914
rect 29202 34862 29204 34914
rect 29148 34860 29204 34862
rect 29372 34914 29428 34916
rect 29372 34862 29374 34914
rect 29374 34862 29426 34914
rect 29426 34862 29428 34914
rect 29372 34860 29428 34862
rect 29708 35196 29764 35252
rect 29148 33234 29204 33236
rect 29148 33182 29150 33234
rect 29150 33182 29202 33234
rect 29202 33182 29204 33234
rect 29148 33180 29204 33182
rect 30268 35196 30324 35252
rect 30044 34412 30100 34468
rect 29372 32732 29428 32788
rect 29260 32562 29316 32564
rect 29260 32510 29262 32562
rect 29262 32510 29314 32562
rect 29314 32510 29316 32562
rect 29260 32508 29316 32510
rect 29820 32396 29876 32452
rect 29260 31724 29316 31780
rect 29820 32172 29876 32228
rect 29148 31666 29204 31668
rect 29148 31614 29150 31666
rect 29150 31614 29202 31666
rect 29202 31614 29204 31666
rect 29148 31612 29204 31614
rect 29484 31554 29540 31556
rect 29484 31502 29486 31554
rect 29486 31502 29538 31554
rect 29538 31502 29540 31554
rect 29484 31500 29540 31502
rect 29484 30994 29540 30996
rect 29484 30942 29486 30994
rect 29486 30942 29538 30994
rect 29538 30942 29540 30994
rect 29484 30940 29540 30942
rect 30044 31778 30100 31780
rect 30044 31726 30046 31778
rect 30046 31726 30098 31778
rect 30098 31726 30100 31778
rect 30044 31724 30100 31726
rect 28700 29932 28756 29988
rect 27804 29426 27860 29428
rect 27804 29374 27806 29426
rect 27806 29374 27858 29426
rect 27858 29374 27860 29426
rect 27804 29372 27860 29374
rect 24444 28364 24500 28420
rect 24780 28082 24836 28084
rect 24780 28030 24782 28082
rect 24782 28030 24834 28082
rect 24834 28030 24836 28082
rect 24780 28028 24836 28030
rect 25452 28082 25508 28084
rect 25452 28030 25454 28082
rect 25454 28030 25506 28082
rect 25506 28030 25508 28082
rect 25452 28028 25508 28030
rect 24108 27804 24164 27860
rect 24668 27804 24724 27860
rect 24332 27356 24388 27412
rect 22428 26908 22484 26964
rect 20524 26850 20580 26852
rect 20524 26798 20526 26850
rect 20526 26798 20578 26850
rect 20578 26798 20580 26850
rect 20524 26796 20580 26798
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19180 26348 19236 26404
rect 18284 26290 18340 26292
rect 18284 26238 18286 26290
rect 18286 26238 18338 26290
rect 18338 26238 18340 26290
rect 18284 26236 18340 26238
rect 18844 26290 18900 26292
rect 18844 26238 18846 26290
rect 18846 26238 18898 26290
rect 18898 26238 18900 26290
rect 18844 26236 18900 26238
rect 17500 25394 17556 25396
rect 17500 25342 17502 25394
rect 17502 25342 17554 25394
rect 17554 25342 17556 25394
rect 17500 25340 17556 25342
rect 17612 24722 17668 24724
rect 17612 24670 17614 24722
rect 17614 24670 17666 24722
rect 17666 24670 17668 24722
rect 17612 24668 17668 24670
rect 17836 24444 17892 24500
rect 18284 26066 18340 26068
rect 18284 26014 18286 26066
rect 18286 26014 18338 26066
rect 18338 26014 18340 26066
rect 18284 26012 18340 26014
rect 19852 26402 19908 26404
rect 19852 26350 19854 26402
rect 19854 26350 19906 26402
rect 19906 26350 19908 26402
rect 19852 26348 19908 26350
rect 19068 26066 19124 26068
rect 19068 26014 19070 26066
rect 19070 26014 19122 26066
rect 19122 26014 19124 26066
rect 19068 26012 19124 26014
rect 20300 25340 20356 25396
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 22092 26460 22148 26516
rect 25228 27356 25284 27412
rect 27468 28754 27524 28756
rect 27468 28702 27470 28754
rect 27470 28702 27522 28754
rect 27522 28702 27524 28754
rect 27468 28700 27524 28702
rect 28700 29484 28756 29540
rect 29820 30828 29876 30884
rect 30604 33964 30660 34020
rect 30828 34914 30884 34916
rect 30828 34862 30830 34914
rect 30830 34862 30882 34914
rect 30882 34862 30884 34914
rect 30828 34860 30884 34862
rect 32508 41074 32564 41076
rect 32508 41022 32510 41074
rect 32510 41022 32562 41074
rect 32562 41022 32564 41074
rect 32508 41020 32564 41022
rect 32060 40402 32116 40404
rect 32060 40350 32062 40402
rect 32062 40350 32114 40402
rect 32114 40350 32116 40402
rect 32060 40348 32116 40350
rect 32508 40236 32564 40292
rect 31836 39116 31892 39172
rect 32284 38892 32340 38948
rect 31612 37996 31668 38052
rect 31276 37436 31332 37492
rect 31836 37436 31892 37492
rect 31388 36204 31444 36260
rect 31052 36092 31108 36148
rect 31500 35868 31556 35924
rect 31276 35084 31332 35140
rect 30716 33740 30772 33796
rect 31052 34690 31108 34692
rect 31052 34638 31054 34690
rect 31054 34638 31106 34690
rect 31106 34638 31108 34690
rect 31052 34636 31108 34638
rect 30604 33346 30660 33348
rect 30604 33294 30606 33346
rect 30606 33294 30658 33346
rect 30658 33294 30660 33346
rect 30604 33292 30660 33294
rect 31948 37212 32004 37268
rect 32172 35308 32228 35364
rect 32284 34972 32340 35028
rect 32732 35644 32788 35700
rect 32508 35474 32564 35476
rect 32508 35422 32510 35474
rect 32510 35422 32562 35474
rect 32562 35422 32564 35474
rect 32508 35420 32564 35422
rect 31836 34802 31892 34804
rect 31836 34750 31838 34802
rect 31838 34750 31890 34802
rect 31890 34750 31892 34802
rect 31836 34748 31892 34750
rect 30940 34076 30996 34132
rect 30940 33852 30996 33908
rect 30828 32562 30884 32564
rect 30828 32510 30830 32562
rect 30830 32510 30882 32562
rect 30882 32510 30884 32562
rect 30828 32508 30884 32510
rect 30716 32172 30772 32228
rect 30492 31724 30548 31780
rect 31724 34242 31780 34244
rect 31724 34190 31726 34242
rect 31726 34190 31778 34242
rect 31778 34190 31780 34242
rect 31724 34188 31780 34190
rect 31948 34130 32004 34132
rect 31948 34078 31950 34130
rect 31950 34078 32002 34130
rect 32002 34078 32004 34130
rect 31948 34076 32004 34078
rect 31500 33740 31556 33796
rect 32620 34802 32676 34804
rect 32620 34750 32622 34802
rect 32622 34750 32674 34802
rect 32674 34750 32676 34802
rect 32620 34748 32676 34750
rect 32172 33852 32228 33908
rect 32844 35532 32900 35588
rect 31836 32562 31892 32564
rect 31836 32510 31838 32562
rect 31838 32510 31890 32562
rect 31890 32510 31892 32562
rect 31836 32508 31892 32510
rect 31612 32450 31668 32452
rect 31612 32398 31614 32450
rect 31614 32398 31666 32450
rect 31666 32398 31668 32450
rect 31612 32396 31668 32398
rect 31388 32338 31444 32340
rect 31388 32286 31390 32338
rect 31390 32286 31442 32338
rect 31442 32286 31444 32338
rect 31388 32284 31444 32286
rect 31164 32172 31220 32228
rect 30604 31948 30660 32004
rect 30380 30156 30436 30212
rect 29596 29538 29652 29540
rect 29596 29486 29598 29538
rect 29598 29486 29650 29538
rect 29650 29486 29652 29538
rect 29596 29484 29652 29486
rect 28364 29036 28420 29092
rect 32060 32732 32116 32788
rect 34188 46956 34244 47012
rect 33516 46844 33572 46900
rect 34748 46002 34804 46004
rect 34748 45950 34750 46002
rect 34750 45950 34802 46002
rect 34802 45950 34804 46002
rect 34748 45948 34804 45950
rect 33180 45836 33236 45892
rect 33292 44322 33348 44324
rect 33292 44270 33294 44322
rect 33294 44270 33346 44322
rect 33346 44270 33348 44322
rect 33292 44268 33348 44270
rect 34524 45106 34580 45108
rect 34524 45054 34526 45106
rect 34526 45054 34578 45106
rect 34578 45054 34580 45106
rect 34524 45052 34580 45054
rect 33964 44268 34020 44324
rect 33516 44098 33572 44100
rect 33516 44046 33518 44098
rect 33518 44046 33570 44098
rect 33570 44046 33572 44098
rect 33516 44044 33572 44046
rect 34188 44156 34244 44212
rect 33628 43538 33684 43540
rect 33628 43486 33630 43538
rect 33630 43486 33682 43538
rect 33682 43486 33684 43538
rect 33628 43484 33684 43486
rect 33740 42866 33796 42868
rect 33740 42814 33742 42866
rect 33742 42814 33794 42866
rect 33794 42814 33796 42866
rect 33740 42812 33796 42814
rect 33740 41692 33796 41748
rect 33516 41020 33572 41076
rect 33404 40908 33460 40964
rect 33516 40348 33572 40404
rect 33068 40236 33124 40292
rect 33516 37324 33572 37380
rect 33964 39564 34020 39620
rect 33628 36204 33684 36260
rect 33852 35810 33908 35812
rect 33852 35758 33854 35810
rect 33854 35758 33906 35810
rect 33906 35758 33908 35810
rect 33852 35756 33908 35758
rect 33740 35586 33796 35588
rect 33740 35534 33742 35586
rect 33742 35534 33794 35586
rect 33794 35534 33796 35586
rect 33740 35532 33796 35534
rect 34076 36540 34132 36596
rect 34636 44044 34692 44100
rect 35868 51378 35924 51380
rect 35868 51326 35870 51378
rect 35870 51326 35922 51378
rect 35922 51326 35924 51378
rect 35868 51324 35924 51326
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 37100 51660 37156 51716
rect 36540 51100 36596 51156
rect 36316 50428 36372 50484
rect 36316 49586 36372 49588
rect 36316 49534 36318 49586
rect 36318 49534 36370 49586
rect 36370 49534 36372 49586
rect 36316 49532 36372 49534
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 36652 49698 36708 49700
rect 36652 49646 36654 49698
rect 36654 49646 36706 49698
rect 36706 49646 36708 49698
rect 36652 49644 36708 49646
rect 36764 49532 36820 49588
rect 35644 48130 35700 48132
rect 35644 48078 35646 48130
rect 35646 48078 35698 48130
rect 35698 48078 35700 48130
rect 35644 48076 35700 48078
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35532 46844 35588 46900
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 36316 48914 36372 48916
rect 36316 48862 36318 48914
rect 36318 48862 36370 48914
rect 36370 48862 36372 48914
rect 36316 48860 36372 48862
rect 36204 46844 36260 46900
rect 36764 47404 36820 47460
rect 36428 46844 36484 46900
rect 36204 46620 36260 46676
rect 36428 46284 36484 46340
rect 37436 53900 37492 53956
rect 37996 57036 38052 57092
rect 38108 56924 38164 56980
rect 38556 56028 38612 56084
rect 37660 54684 37716 54740
rect 38892 54738 38948 54740
rect 38892 54686 38894 54738
rect 38894 54686 38946 54738
rect 38946 54686 38948 54738
rect 38892 54684 38948 54686
rect 39116 56306 39172 56308
rect 39116 56254 39118 56306
rect 39118 56254 39170 56306
rect 39170 56254 39172 56306
rect 39116 56252 39172 56254
rect 39900 56252 39956 56308
rect 39788 56082 39844 56084
rect 39788 56030 39790 56082
rect 39790 56030 39842 56082
rect 39842 56030 39844 56082
rect 39788 56028 39844 56030
rect 40572 56924 40628 56980
rect 41132 56306 41188 56308
rect 41132 56254 41134 56306
rect 41134 56254 41186 56306
rect 41186 56254 41188 56306
rect 41132 56252 41188 56254
rect 41580 56252 41636 56308
rect 41356 56194 41412 56196
rect 41356 56142 41358 56194
rect 41358 56142 41410 56194
rect 41410 56142 41412 56194
rect 41356 56140 41412 56142
rect 40348 55916 40404 55972
rect 39452 55356 39508 55412
rect 40684 55410 40740 55412
rect 40684 55358 40686 55410
rect 40686 55358 40738 55410
rect 40738 55358 40740 55410
rect 40684 55356 40740 55358
rect 41244 56028 41300 56084
rect 41580 56028 41636 56084
rect 42028 56082 42084 56084
rect 42028 56030 42030 56082
rect 42030 56030 42082 56082
rect 42082 56030 42084 56082
rect 42028 56028 42084 56030
rect 38780 54460 38836 54516
rect 37772 53788 37828 53844
rect 40908 54514 40964 54516
rect 40908 54462 40910 54514
rect 40910 54462 40962 54514
rect 40962 54462 40964 54514
rect 40908 54460 40964 54462
rect 37548 53004 37604 53060
rect 38892 52220 38948 52276
rect 37884 52108 37940 52164
rect 37436 51378 37492 51380
rect 37436 51326 37438 51378
rect 37438 51326 37490 51378
rect 37490 51326 37492 51378
rect 37436 51324 37492 51326
rect 39452 52834 39508 52836
rect 39452 52782 39454 52834
rect 39454 52782 39506 52834
rect 39506 52782 39508 52834
rect 39452 52780 39508 52782
rect 38108 51772 38164 51828
rect 37660 51154 37716 51156
rect 37660 51102 37662 51154
rect 37662 51102 37714 51154
rect 37714 51102 37716 51154
rect 37660 51100 37716 51102
rect 38668 51660 38724 51716
rect 38108 51436 38164 51492
rect 38556 51154 38612 51156
rect 38556 51102 38558 51154
rect 38558 51102 38610 51154
rect 38610 51102 38612 51154
rect 38556 51100 38612 51102
rect 39676 51996 39732 52052
rect 39116 51772 39172 51828
rect 37548 50482 37604 50484
rect 37548 50430 37550 50482
rect 37550 50430 37602 50482
rect 37602 50430 37604 50482
rect 37548 50428 37604 50430
rect 38444 50482 38500 50484
rect 38444 50430 38446 50482
rect 38446 50430 38498 50482
rect 38498 50430 38500 50482
rect 38444 50428 38500 50430
rect 37884 50204 37940 50260
rect 42700 55970 42756 55972
rect 42700 55918 42702 55970
rect 42702 55918 42754 55970
rect 42754 55918 42756 55970
rect 42700 55916 42756 55918
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 41580 53788 41636 53844
rect 40796 52892 40852 52948
rect 42476 53842 42532 53844
rect 42476 53790 42478 53842
rect 42478 53790 42530 53842
rect 42530 53790 42532 53842
rect 42476 53788 42532 53790
rect 42364 53730 42420 53732
rect 42364 53678 42366 53730
rect 42366 53678 42418 53730
rect 42418 53678 42420 53730
rect 42364 53676 42420 53678
rect 42588 53506 42644 53508
rect 42588 53454 42590 53506
rect 42590 53454 42642 53506
rect 42642 53454 42644 53506
rect 42588 53452 42644 53454
rect 43036 53564 43092 53620
rect 43484 53730 43540 53732
rect 43484 53678 43486 53730
rect 43486 53678 43538 53730
rect 43538 53678 43540 53730
rect 43484 53676 43540 53678
rect 41692 52892 41748 52948
rect 40796 52274 40852 52276
rect 40796 52222 40798 52274
rect 40798 52222 40850 52274
rect 40850 52222 40852 52274
rect 40796 52220 40852 52222
rect 40124 51548 40180 51604
rect 40348 52050 40404 52052
rect 40348 51998 40350 52050
rect 40350 51998 40402 52050
rect 40402 51998 40404 52050
rect 40348 51996 40404 51998
rect 41020 51884 41076 51940
rect 40908 51548 40964 51604
rect 38668 49810 38724 49812
rect 38668 49758 38670 49810
rect 38670 49758 38722 49810
rect 38722 49758 38724 49810
rect 38668 49756 38724 49758
rect 37324 48860 37380 48916
rect 37996 48076 38052 48132
rect 38556 48188 38612 48244
rect 38892 47964 38948 48020
rect 39116 48242 39172 48244
rect 39116 48190 39118 48242
rect 39118 48190 39170 48242
rect 39170 48190 39172 48242
rect 39116 48188 39172 48190
rect 37100 47458 37156 47460
rect 37100 47406 37102 47458
rect 37102 47406 37154 47458
rect 37154 47406 37156 47458
rect 37100 47404 37156 47406
rect 37100 46898 37156 46900
rect 37100 46846 37102 46898
rect 37102 46846 37154 46898
rect 37154 46846 37156 46898
rect 37100 46844 37156 46846
rect 36876 46620 36932 46676
rect 36764 46172 36820 46228
rect 37212 46396 37268 46452
rect 35308 45106 35364 45108
rect 35308 45054 35310 45106
rect 35310 45054 35362 45106
rect 35362 45054 35364 45106
rect 35308 45052 35364 45054
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35308 44210 35364 44212
rect 35308 44158 35310 44210
rect 35310 44158 35362 44210
rect 35362 44158 35364 44210
rect 35308 44156 35364 44158
rect 35644 44156 35700 44212
rect 34748 43596 34804 43652
rect 34412 43538 34468 43540
rect 34412 43486 34414 43538
rect 34414 43486 34466 43538
rect 34466 43486 34468 43538
rect 34412 43484 34468 43486
rect 34636 42924 34692 42980
rect 34860 43538 34916 43540
rect 34860 43486 34862 43538
rect 34862 43486 34914 43538
rect 34914 43486 34916 43538
rect 34860 43484 34916 43486
rect 35308 43426 35364 43428
rect 35308 43374 35310 43426
rect 35310 43374 35362 43426
rect 35362 43374 35364 43426
rect 35308 43372 35364 43374
rect 35644 43650 35700 43652
rect 35644 43598 35646 43650
rect 35646 43598 35698 43650
rect 35698 43598 35700 43650
rect 35644 43596 35700 43598
rect 35420 43260 35476 43316
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 34300 40012 34356 40068
rect 34300 39676 34356 39732
rect 34412 39564 34468 39620
rect 34300 39058 34356 39060
rect 34300 39006 34302 39058
rect 34302 39006 34354 39058
rect 34354 39006 34356 39058
rect 34300 39004 34356 39006
rect 34188 36428 34244 36484
rect 34412 37772 34468 37828
rect 34188 36204 34244 36260
rect 34076 35532 34132 35588
rect 33964 34972 34020 35028
rect 32508 33404 32564 33460
rect 33068 34748 33124 34804
rect 32732 33234 32788 33236
rect 32732 33182 32734 33234
rect 32734 33182 32786 33234
rect 32786 33182 32788 33234
rect 32732 33180 32788 33182
rect 31948 32396 32004 32452
rect 32060 31948 32116 32004
rect 30940 30940 30996 30996
rect 32396 32396 32452 32452
rect 32396 31052 32452 31108
rect 30940 30268 30996 30324
rect 32620 29820 32676 29876
rect 31948 29596 32004 29652
rect 32284 29538 32340 29540
rect 32284 29486 32286 29538
rect 32286 29486 32338 29538
rect 32338 29486 32340 29538
rect 32284 29484 32340 29486
rect 32508 29426 32564 29428
rect 32508 29374 32510 29426
rect 32510 29374 32562 29426
rect 32562 29374 32564 29426
rect 32508 29372 32564 29374
rect 30828 29148 30884 29204
rect 29932 28700 29988 28756
rect 30604 28588 30660 28644
rect 30156 27970 30212 27972
rect 30156 27918 30158 27970
rect 30158 27918 30210 27970
rect 30210 27918 30212 27970
rect 30156 27916 30212 27918
rect 30716 27916 30772 27972
rect 29260 27074 29316 27076
rect 29260 27022 29262 27074
rect 29262 27022 29314 27074
rect 29314 27022 29316 27074
rect 29260 27020 29316 27022
rect 32620 28588 32676 28644
rect 32508 28418 32564 28420
rect 32508 28366 32510 28418
rect 32510 28366 32562 28418
rect 32562 28366 32564 28418
rect 32508 28364 32564 28366
rect 32060 27916 32116 27972
rect 32284 27858 32340 27860
rect 32284 27806 32286 27858
rect 32286 27806 32338 27858
rect 32338 27806 32340 27858
rect 32284 27804 32340 27806
rect 16604 22092 16660 22148
rect 16828 22258 16884 22260
rect 16828 22206 16830 22258
rect 16830 22206 16882 22258
rect 16882 22206 16884 22258
rect 16828 22204 16884 22206
rect 16716 21532 16772 21588
rect 16716 21362 16772 21364
rect 16716 21310 16718 21362
rect 16718 21310 16770 21362
rect 16770 21310 16772 21362
rect 16716 21308 16772 21310
rect 16492 20748 16548 20804
rect 16604 21084 16660 21140
rect 17388 22540 17444 22596
rect 17388 22204 17444 22260
rect 17500 21698 17556 21700
rect 17500 21646 17502 21698
rect 17502 21646 17554 21698
rect 17554 21646 17556 21698
rect 17500 21644 17556 21646
rect 16716 20690 16772 20692
rect 16716 20638 16718 20690
rect 16718 20638 16770 20690
rect 16770 20638 16772 20690
rect 16716 20636 16772 20638
rect 16828 20524 16884 20580
rect 16716 20018 16772 20020
rect 16716 19966 16718 20018
rect 16718 19966 16770 20018
rect 16770 19966 16772 20018
rect 16716 19964 16772 19966
rect 17388 20018 17444 20020
rect 17388 19966 17390 20018
rect 17390 19966 17442 20018
rect 17442 19966 17444 20018
rect 17388 19964 17444 19966
rect 16156 19346 16212 19348
rect 16156 19294 16158 19346
rect 16158 19294 16210 19346
rect 16210 19294 16212 19346
rect 16156 19292 16212 19294
rect 15484 17666 15540 17668
rect 15484 17614 15486 17666
rect 15486 17614 15538 17666
rect 15538 17614 15540 17666
rect 15484 17612 15540 17614
rect 16044 16882 16100 16884
rect 16044 16830 16046 16882
rect 16046 16830 16098 16882
rect 16098 16830 16100 16882
rect 16044 16828 16100 16830
rect 15820 16716 15876 16772
rect 14812 15932 14868 15988
rect 15932 15986 15988 15988
rect 15932 15934 15934 15986
rect 15934 15934 15986 15986
rect 15986 15934 15988 15986
rect 15932 15932 15988 15934
rect 16268 16322 16324 16324
rect 16268 16270 16270 16322
rect 16270 16270 16322 16322
rect 16322 16270 16324 16322
rect 16268 16268 16324 16270
rect 15596 15202 15652 15204
rect 15596 15150 15598 15202
rect 15598 15150 15650 15202
rect 15650 15150 15652 15202
rect 15596 15148 15652 15150
rect 11452 13804 11508 13860
rect 11340 13580 11396 13636
rect 11004 13020 11060 13076
rect 8540 12684 8596 12740
rect 11900 14364 11956 14420
rect 12236 14364 12292 14420
rect 18284 24610 18340 24612
rect 18284 24558 18286 24610
rect 18286 24558 18338 24610
rect 18338 24558 18340 24610
rect 18284 24556 18340 24558
rect 18508 24220 18564 24276
rect 19068 24722 19124 24724
rect 19068 24670 19070 24722
rect 19070 24670 19122 24722
rect 19122 24670 19124 24722
rect 19068 24668 19124 24670
rect 19292 24722 19348 24724
rect 19292 24670 19294 24722
rect 19294 24670 19346 24722
rect 19346 24670 19348 24722
rect 19292 24668 19348 24670
rect 19628 24668 19684 24724
rect 18732 24444 18788 24500
rect 18060 23884 18116 23940
rect 18732 23884 18788 23940
rect 18172 21868 18228 21924
rect 18172 21644 18228 21700
rect 20748 24722 20804 24724
rect 20748 24670 20750 24722
rect 20750 24670 20802 24722
rect 20802 24670 20804 24722
rect 20748 24668 20804 24670
rect 20076 24220 20132 24276
rect 20412 23938 20468 23940
rect 20412 23886 20414 23938
rect 20414 23886 20466 23938
rect 20466 23886 20468 23938
rect 20412 23884 20468 23886
rect 20188 23772 20244 23828
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19068 22876 19124 22932
rect 18956 22540 19012 22596
rect 19740 23042 19796 23044
rect 19740 22990 19742 23042
rect 19742 22990 19794 23042
rect 19794 22990 19796 23042
rect 19740 22988 19796 22990
rect 17724 19516 17780 19572
rect 18396 21532 18452 21588
rect 19068 20860 19124 20916
rect 19180 21644 19236 21700
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19628 21532 19684 21588
rect 18508 20636 18564 20692
rect 18844 19292 18900 19348
rect 18508 18284 18564 18340
rect 18956 18172 19012 18228
rect 18284 17948 18340 18004
rect 18396 17836 18452 17892
rect 17836 17724 17892 17780
rect 17500 17276 17556 17332
rect 16828 16994 16884 16996
rect 16828 16942 16830 16994
rect 16830 16942 16882 16994
rect 16882 16942 16884 16994
rect 16828 16940 16884 16942
rect 17500 16994 17556 16996
rect 17500 16942 17502 16994
rect 17502 16942 17554 16994
rect 17554 16942 17556 16994
rect 17500 16940 17556 16942
rect 16716 16828 16772 16884
rect 18284 17388 18340 17444
rect 18396 17276 18452 17332
rect 18284 16716 18340 16772
rect 16380 14418 16436 14420
rect 16380 14366 16382 14418
rect 16382 14366 16434 14418
rect 16434 14366 16436 14418
rect 16380 14364 16436 14366
rect 13692 13858 13748 13860
rect 13692 13806 13694 13858
rect 13694 13806 13746 13858
rect 13746 13806 13748 13858
rect 13692 13804 13748 13806
rect 11564 13074 11620 13076
rect 11564 13022 11566 13074
rect 11566 13022 11618 13074
rect 11618 13022 11620 13074
rect 11564 13020 11620 13022
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 12460 11900 12516 11956
rect 14028 13020 14084 13076
rect 14364 13020 14420 13076
rect 14700 13522 14756 13524
rect 14700 13470 14702 13522
rect 14702 13470 14754 13522
rect 14754 13470 14756 13522
rect 14700 13468 14756 13470
rect 15372 13132 15428 13188
rect 14252 11954 14308 11956
rect 14252 11902 14254 11954
rect 14254 11902 14306 11954
rect 14306 11902 14308 11954
rect 14252 11900 14308 11902
rect 13468 10668 13524 10724
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 13244 10498 13300 10500
rect 13244 10446 13246 10498
rect 13246 10446 13298 10498
rect 13298 10446 13300 10498
rect 13244 10444 13300 10446
rect 15148 11788 15204 11844
rect 11676 9714 11732 9716
rect 11676 9662 11678 9714
rect 11678 9662 11730 9714
rect 11730 9662 11732 9714
rect 11676 9660 11732 9662
rect 14028 9714 14084 9716
rect 14028 9662 14030 9714
rect 14030 9662 14082 9714
rect 14082 9662 14084 9714
rect 14028 9660 14084 9662
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 11900 8764 11956 8820
rect 14476 10722 14532 10724
rect 14476 10670 14478 10722
rect 14478 10670 14530 10722
rect 14530 10670 14532 10722
rect 14476 10668 14532 10670
rect 14364 10444 14420 10500
rect 14700 10498 14756 10500
rect 14700 10446 14702 10498
rect 14702 10446 14754 10498
rect 14754 10446 14756 10498
rect 14700 10444 14756 10446
rect 16940 15372 16996 15428
rect 17388 15202 17444 15204
rect 17388 15150 17390 15202
rect 17390 15150 17442 15202
rect 17442 15150 17444 15202
rect 17388 15148 17444 15150
rect 17388 14700 17444 14756
rect 16492 13580 16548 13636
rect 16716 13132 16772 13188
rect 15820 12908 15876 12964
rect 16044 11676 16100 11732
rect 15708 10668 15764 10724
rect 15260 9996 15316 10052
rect 14812 9660 14868 9716
rect 15932 9548 15988 9604
rect 14924 9154 14980 9156
rect 14924 9102 14926 9154
rect 14926 9102 14978 9154
rect 14978 9102 14980 9154
rect 14924 9100 14980 9102
rect 15036 9042 15092 9044
rect 15036 8990 15038 9042
rect 15038 8990 15090 9042
rect 15090 8990 15092 9042
rect 15036 8988 15092 8990
rect 13916 8818 13972 8820
rect 13916 8766 13918 8818
rect 13918 8766 13970 8818
rect 13970 8766 13972 8818
rect 13916 8764 13972 8766
rect 15148 8370 15204 8372
rect 15148 8318 15150 8370
rect 15150 8318 15202 8370
rect 15202 8318 15204 8370
rect 15148 8316 15204 8318
rect 12236 7474 12292 7476
rect 12236 7422 12238 7474
rect 12238 7422 12290 7474
rect 12290 7422 12292 7474
rect 12236 7420 12292 7422
rect 13580 7420 13636 7476
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 16716 11228 16772 11284
rect 16268 11170 16324 11172
rect 16268 11118 16270 11170
rect 16270 11118 16322 11170
rect 16322 11118 16324 11170
rect 16268 11116 16324 11118
rect 17724 15090 17780 15092
rect 17724 15038 17726 15090
rect 17726 15038 17778 15090
rect 17778 15038 17780 15090
rect 17724 15036 17780 15038
rect 17612 13858 17668 13860
rect 17612 13806 17614 13858
rect 17614 13806 17666 13858
rect 17666 13806 17668 13858
rect 17612 13804 17668 13806
rect 17276 13244 17332 13300
rect 17500 13020 17556 13076
rect 17164 12124 17220 12180
rect 18844 17778 18900 17780
rect 18844 17726 18846 17778
rect 18846 17726 18898 17778
rect 18898 17726 18900 17778
rect 18844 17724 18900 17726
rect 18620 17500 18676 17556
rect 19068 20524 19124 20580
rect 19180 20412 19236 20468
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19740 20242 19796 20244
rect 19740 20190 19742 20242
rect 19742 20190 19794 20242
rect 19794 20190 19796 20242
rect 19740 20188 19796 20190
rect 20188 18956 20244 19012
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18620 19684 18676
rect 19628 18338 19684 18340
rect 19628 18286 19630 18338
rect 19630 18286 19682 18338
rect 19682 18286 19684 18338
rect 19628 18284 19684 18286
rect 19292 17948 19348 18004
rect 19180 17164 19236 17220
rect 19628 17666 19684 17668
rect 19628 17614 19630 17666
rect 19630 17614 19682 17666
rect 19682 17614 19684 17666
rect 19628 17612 19684 17614
rect 19852 17554 19908 17556
rect 19852 17502 19854 17554
rect 19854 17502 19906 17554
rect 19906 17502 19908 17554
rect 19852 17500 19908 17502
rect 19628 17388 19684 17444
rect 20412 23548 20468 23604
rect 20860 24220 20916 24276
rect 20636 23324 20692 23380
rect 20748 23548 20804 23604
rect 20972 23772 21028 23828
rect 20972 23154 21028 23156
rect 20972 23102 20974 23154
rect 20974 23102 21026 23154
rect 21026 23102 21028 23154
rect 20972 23100 21028 23102
rect 20412 22594 20468 22596
rect 20412 22542 20414 22594
rect 20414 22542 20466 22594
rect 20466 22542 20468 22594
rect 20412 22540 20468 22542
rect 20524 20914 20580 20916
rect 20524 20862 20526 20914
rect 20526 20862 20578 20914
rect 20578 20862 20580 20914
rect 20524 20860 20580 20862
rect 20412 20802 20468 20804
rect 20412 20750 20414 20802
rect 20414 20750 20466 20802
rect 20466 20750 20468 20802
rect 20412 20748 20468 20750
rect 20412 20412 20468 20468
rect 20412 19292 20468 19348
rect 20524 18732 20580 18788
rect 21308 23826 21364 23828
rect 21308 23774 21310 23826
rect 21310 23774 21362 23826
rect 21362 23774 21364 23826
rect 21308 23772 21364 23774
rect 21756 23772 21812 23828
rect 21532 23548 21588 23604
rect 21420 23436 21476 23492
rect 21644 23324 21700 23380
rect 23548 23826 23604 23828
rect 23548 23774 23550 23826
rect 23550 23774 23602 23826
rect 23602 23774 23604 23826
rect 23548 23772 23604 23774
rect 23212 23714 23268 23716
rect 23212 23662 23214 23714
rect 23214 23662 23266 23714
rect 23266 23662 23268 23714
rect 23212 23660 23268 23662
rect 23996 23660 24052 23716
rect 22204 23100 22260 23156
rect 22764 22988 22820 23044
rect 21980 22876 22036 22932
rect 21420 22146 21476 22148
rect 21420 22094 21422 22146
rect 21422 22094 21474 22146
rect 21474 22094 21476 22146
rect 21420 22092 21476 22094
rect 22652 22092 22708 22148
rect 21980 21980 22036 22036
rect 21980 21586 22036 21588
rect 21980 21534 21982 21586
rect 21982 21534 22034 21586
rect 22034 21534 22036 21586
rect 21980 21532 22036 21534
rect 22652 21420 22708 21476
rect 21084 20748 21140 20804
rect 21084 19906 21140 19908
rect 21084 19854 21086 19906
rect 21086 19854 21138 19906
rect 21138 19854 21140 19906
rect 21084 19852 21140 19854
rect 21308 19010 21364 19012
rect 21308 18958 21310 19010
rect 21310 18958 21362 19010
rect 21362 18958 21364 19010
rect 21308 18956 21364 18958
rect 20524 17724 20580 17780
rect 20300 17388 20356 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20188 16940 20244 16996
rect 20188 16268 20244 16324
rect 20300 16492 20356 16548
rect 20076 16156 20132 16212
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19292 15426 19348 15428
rect 19292 15374 19294 15426
rect 19294 15374 19346 15426
rect 19346 15374 19348 15426
rect 19292 15372 19348 15374
rect 19628 15314 19684 15316
rect 19628 15262 19630 15314
rect 19630 15262 19682 15314
rect 19682 15262 19684 15314
rect 19628 15260 19684 15262
rect 19180 14476 19236 14532
rect 18620 13746 18676 13748
rect 18620 13694 18622 13746
rect 18622 13694 18674 13746
rect 18674 13694 18676 13746
rect 18620 13692 18676 13694
rect 20076 14700 20132 14756
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20972 18172 21028 18228
rect 20972 17164 21028 17220
rect 21980 20690 22036 20692
rect 21980 20638 21982 20690
rect 21982 20638 22034 20690
rect 22034 20638 22036 20690
rect 21980 20636 22036 20638
rect 21756 20524 21812 20580
rect 22204 20578 22260 20580
rect 22204 20526 22206 20578
rect 22206 20526 22258 20578
rect 22258 20526 22260 20578
rect 22204 20524 22260 20526
rect 21532 20412 21588 20468
rect 22428 20412 22484 20468
rect 21644 19234 21700 19236
rect 21644 19182 21646 19234
rect 21646 19182 21698 19234
rect 21698 19182 21700 19234
rect 21644 19180 21700 19182
rect 22092 19852 22148 19908
rect 22316 19740 22372 19796
rect 22428 19292 22484 19348
rect 22540 20188 22596 20244
rect 23660 22540 23716 22596
rect 22876 20860 22932 20916
rect 24220 22988 24276 23044
rect 24108 22316 24164 22372
rect 22988 20636 23044 20692
rect 23660 20524 23716 20580
rect 23772 20188 23828 20244
rect 23100 20076 23156 20132
rect 23100 19852 23156 19908
rect 23548 19794 23604 19796
rect 23548 19742 23550 19794
rect 23550 19742 23602 19794
rect 23602 19742 23604 19794
rect 23548 19740 23604 19742
rect 23996 20524 24052 20580
rect 24220 20130 24276 20132
rect 24220 20078 24222 20130
rect 24222 20078 24274 20130
rect 24274 20078 24276 20130
rect 24220 20076 24276 20078
rect 24444 20018 24500 20020
rect 24444 19966 24446 20018
rect 24446 19966 24498 20018
rect 24498 19966 24500 20018
rect 24444 19964 24500 19966
rect 23996 19346 24052 19348
rect 23996 19294 23998 19346
rect 23998 19294 24050 19346
rect 24050 19294 24052 19346
rect 23996 19292 24052 19294
rect 23884 19068 23940 19124
rect 23436 19010 23492 19012
rect 23436 18958 23438 19010
rect 23438 18958 23490 19010
rect 23490 18958 23492 19010
rect 23436 18956 23492 18958
rect 21756 17612 21812 17668
rect 22428 17948 22484 18004
rect 22092 17388 22148 17444
rect 21308 15260 21364 15316
rect 20748 14700 20804 14756
rect 20636 14476 20692 14532
rect 20860 14364 20916 14420
rect 19180 13634 19236 13636
rect 19180 13582 19182 13634
rect 19182 13582 19234 13634
rect 19234 13582 19236 13634
rect 19180 13580 19236 13582
rect 18060 13244 18116 13300
rect 18508 13132 18564 13188
rect 17724 12962 17780 12964
rect 17724 12910 17726 12962
rect 17726 12910 17778 12962
rect 17778 12910 17780 12962
rect 17724 12908 17780 12910
rect 17500 11676 17556 11732
rect 17612 10780 17668 10836
rect 18508 11004 18564 11060
rect 17836 10610 17892 10612
rect 17836 10558 17838 10610
rect 17838 10558 17890 10610
rect 17890 10558 17892 10610
rect 17836 10556 17892 10558
rect 18620 10556 18676 10612
rect 17388 10444 17444 10500
rect 18284 10498 18340 10500
rect 18284 10446 18286 10498
rect 18286 10446 18338 10498
rect 18338 10446 18340 10498
rect 18284 10444 18340 10446
rect 16940 9660 16996 9716
rect 17500 9884 17556 9940
rect 18060 9884 18116 9940
rect 17948 9714 18004 9716
rect 17948 9662 17950 9714
rect 17950 9662 18002 9714
rect 18002 9662 18004 9714
rect 17948 9660 18004 9662
rect 17164 9602 17220 9604
rect 17164 9550 17166 9602
rect 17166 9550 17218 9602
rect 17218 9550 17220 9602
rect 17164 9548 17220 9550
rect 16156 8988 16212 9044
rect 15484 6914 15540 6916
rect 15484 6862 15486 6914
rect 15486 6862 15538 6914
rect 15538 6862 15540 6914
rect 15484 6860 15540 6862
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 13468 4956 13524 5012
rect 14028 4956 14084 5012
rect 14476 5122 14532 5124
rect 14476 5070 14478 5122
rect 14478 5070 14530 5122
rect 14530 5070 14532 5122
rect 14476 5068 14532 5070
rect 15148 5068 15204 5124
rect 15932 6860 15988 6916
rect 16044 5964 16100 6020
rect 16380 8316 16436 8372
rect 16716 8316 16772 8372
rect 17724 8988 17780 9044
rect 17836 8316 17892 8372
rect 15484 5068 15540 5124
rect 16940 5740 16996 5796
rect 16828 4956 16884 5012
rect 17164 4956 17220 5012
rect 14700 4450 14756 4452
rect 14700 4398 14702 4450
rect 14702 4398 14754 4450
rect 14754 4398 14756 4450
rect 14700 4396 14756 4398
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 17388 4450 17444 4452
rect 17388 4398 17390 4450
rect 17390 4398 17442 4450
rect 17442 4398 17444 4450
rect 17388 4396 17444 4398
rect 18172 8204 18228 8260
rect 18620 9436 18676 9492
rect 18732 9826 18788 9828
rect 18732 9774 18734 9826
rect 18734 9774 18786 9826
rect 18786 9774 18788 9826
rect 18732 9772 18788 9774
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19852 12178 19908 12180
rect 19852 12126 19854 12178
rect 19854 12126 19906 12178
rect 19906 12126 19908 12178
rect 19852 12124 19908 12126
rect 19852 11676 19908 11732
rect 19180 11004 19236 11060
rect 20188 11506 20244 11508
rect 20188 11454 20190 11506
rect 20190 11454 20242 11506
rect 20242 11454 20244 11506
rect 20188 11452 20244 11454
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 18956 10610 19012 10612
rect 18956 10558 18958 10610
rect 18958 10558 19010 10610
rect 19010 10558 19012 10610
rect 18956 10556 19012 10558
rect 19628 10610 19684 10612
rect 19628 10558 19630 10610
rect 19630 10558 19682 10610
rect 19682 10558 19684 10610
rect 19628 10556 19684 10558
rect 21756 15148 21812 15204
rect 22428 17164 22484 17220
rect 22988 17948 23044 18004
rect 23324 17500 23380 17556
rect 23996 18060 24052 18116
rect 23772 17500 23828 17556
rect 21980 14418 22036 14420
rect 21980 14366 21982 14418
rect 21982 14366 22034 14418
rect 22034 14366 22036 14418
rect 21980 14364 22036 14366
rect 21756 13804 21812 13860
rect 19180 9714 19236 9716
rect 19180 9662 19182 9714
rect 19182 9662 19234 9714
rect 19234 9662 19236 9714
rect 19180 9660 19236 9662
rect 19628 9996 19684 10052
rect 19292 9548 19348 9604
rect 19516 9660 19572 9716
rect 19516 9436 19572 9492
rect 20524 9996 20580 10052
rect 20636 11676 20692 11732
rect 19740 9714 19796 9716
rect 19740 9662 19742 9714
rect 19742 9662 19794 9714
rect 19794 9662 19796 9714
rect 19740 9660 19796 9662
rect 20188 9602 20244 9604
rect 20188 9550 20190 9602
rect 20190 9550 20242 9602
rect 20242 9550 20244 9602
rect 20188 9548 20244 9550
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 18844 7586 18900 7588
rect 18844 7534 18846 7586
rect 18846 7534 18898 7586
rect 18898 7534 18900 7586
rect 18844 7532 18900 7534
rect 19964 8764 20020 8820
rect 19404 8316 19460 8372
rect 19516 8204 19572 8260
rect 20524 8818 20580 8820
rect 20524 8766 20526 8818
rect 20526 8766 20578 8818
rect 20578 8766 20580 8818
rect 20524 8764 20580 8766
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 21756 12012 21812 12068
rect 21644 11452 21700 11508
rect 20748 10610 20804 10612
rect 20748 10558 20750 10610
rect 20750 10558 20802 10610
rect 20802 10558 20804 10610
rect 20748 10556 20804 10558
rect 21196 9996 21252 10052
rect 21980 11340 22036 11396
rect 21980 10556 22036 10612
rect 22204 14364 22260 14420
rect 22092 10668 22148 10724
rect 22316 10722 22372 10724
rect 22316 10670 22318 10722
rect 22318 10670 22370 10722
rect 22370 10670 22372 10722
rect 22316 10668 22372 10670
rect 22092 9826 22148 9828
rect 22092 9774 22094 9826
rect 22094 9774 22146 9826
rect 22146 9774 22148 9826
rect 22092 9772 22148 9774
rect 21868 9154 21924 9156
rect 21868 9102 21870 9154
rect 21870 9102 21922 9154
rect 21922 9102 21924 9154
rect 21868 9100 21924 9102
rect 21532 8876 21588 8932
rect 20636 8370 20692 8372
rect 20636 8318 20638 8370
rect 20638 8318 20690 8370
rect 20690 8318 20692 8370
rect 20636 8316 20692 8318
rect 20412 7308 20468 7364
rect 21756 6636 21812 6692
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 18396 6018 18452 6020
rect 18396 5966 18398 6018
rect 18398 5966 18450 6018
rect 18450 5966 18452 6018
rect 18396 5964 18452 5966
rect 17836 5794 17892 5796
rect 17836 5742 17838 5794
rect 17838 5742 17890 5794
rect 17890 5742 17892 5794
rect 17836 5740 17892 5742
rect 19292 5292 19348 5348
rect 18732 4450 18788 4452
rect 18732 4398 18734 4450
rect 18734 4398 18786 4450
rect 18786 4398 18788 4450
rect 18732 4396 18788 4398
rect 20636 5292 20692 5348
rect 20412 4956 20468 5012
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20972 4956 21028 5012
rect 21756 5964 21812 6020
rect 21420 5682 21476 5684
rect 21420 5630 21422 5682
rect 21422 5630 21474 5682
rect 21474 5630 21476 5682
rect 21420 5628 21476 5630
rect 22204 8876 22260 8932
rect 21980 8146 22036 8148
rect 21980 8094 21982 8146
rect 21982 8094 22034 8146
rect 22034 8094 22036 8146
rect 21980 8092 22036 8094
rect 22988 16770 23044 16772
rect 22988 16718 22990 16770
rect 22990 16718 23042 16770
rect 23042 16718 23044 16770
rect 22988 16716 23044 16718
rect 23324 16604 23380 16660
rect 22876 16380 22932 16436
rect 22764 16210 22820 16212
rect 22764 16158 22766 16210
rect 22766 16158 22818 16210
rect 22818 16158 22820 16210
rect 22764 16156 22820 16158
rect 23324 16156 23380 16212
rect 22876 15202 22932 15204
rect 22876 15150 22878 15202
rect 22878 15150 22930 15202
rect 22930 15150 22932 15202
rect 22876 15148 22932 15150
rect 22540 13746 22596 13748
rect 22540 13694 22542 13746
rect 22542 13694 22594 13746
rect 22594 13694 22596 13746
rect 22540 13692 22596 13694
rect 23324 13970 23380 13972
rect 23324 13918 23326 13970
rect 23326 13918 23378 13970
rect 23378 13918 23380 13970
rect 23324 13916 23380 13918
rect 23324 13746 23380 13748
rect 23324 13694 23326 13746
rect 23326 13694 23378 13746
rect 23378 13694 23380 13746
rect 23324 13692 23380 13694
rect 22988 12738 23044 12740
rect 22988 12686 22990 12738
rect 22990 12686 23042 12738
rect 23042 12686 23044 12738
rect 22988 12684 23044 12686
rect 22764 12348 22820 12404
rect 22988 12460 23044 12516
rect 22764 12066 22820 12068
rect 22764 12014 22766 12066
rect 22766 12014 22818 12066
rect 22818 12014 22820 12066
rect 22764 12012 22820 12014
rect 22540 11676 22596 11732
rect 23212 12402 23268 12404
rect 23212 12350 23214 12402
rect 23214 12350 23266 12402
rect 23266 12350 23268 12402
rect 23212 12348 23268 12350
rect 23660 16940 23716 16996
rect 23884 16828 23940 16884
rect 24444 19122 24500 19124
rect 24444 19070 24446 19122
rect 24446 19070 24498 19122
rect 24498 19070 24500 19122
rect 24444 19068 24500 19070
rect 24332 18060 24388 18116
rect 24668 25282 24724 25284
rect 24668 25230 24670 25282
rect 24670 25230 24722 25282
rect 24722 25230 24724 25282
rect 24668 25228 24724 25230
rect 25340 25282 25396 25284
rect 25340 25230 25342 25282
rect 25342 25230 25394 25282
rect 25394 25230 25396 25282
rect 25340 25228 25396 25230
rect 25788 25228 25844 25284
rect 26460 23996 26516 24052
rect 24668 23660 24724 23716
rect 24780 23324 24836 23380
rect 25564 23378 25620 23380
rect 25564 23326 25566 23378
rect 25566 23326 25618 23378
rect 25618 23326 25620 23378
rect 25564 23324 25620 23326
rect 24780 22594 24836 22596
rect 24780 22542 24782 22594
rect 24782 22542 24834 22594
rect 24834 22542 24836 22594
rect 24780 22540 24836 22542
rect 25452 22428 25508 22484
rect 25116 22370 25172 22372
rect 25116 22318 25118 22370
rect 25118 22318 25170 22370
rect 25170 22318 25172 22370
rect 25116 22316 25172 22318
rect 24668 22092 24724 22148
rect 26460 23154 26516 23156
rect 26460 23102 26462 23154
rect 26462 23102 26514 23154
rect 26514 23102 26516 23154
rect 26460 23100 26516 23102
rect 26236 23042 26292 23044
rect 26236 22990 26238 23042
rect 26238 22990 26290 23042
rect 26290 22990 26292 23042
rect 26236 22988 26292 22990
rect 25900 22540 25956 22596
rect 27804 23996 27860 24052
rect 25564 22146 25620 22148
rect 25564 22094 25566 22146
rect 25566 22094 25618 22146
rect 25618 22094 25620 22146
rect 25564 22092 25620 22094
rect 24668 21868 24724 21924
rect 26460 20076 26516 20132
rect 25116 19292 25172 19348
rect 25452 20018 25508 20020
rect 25452 19966 25454 20018
rect 25454 19966 25506 20018
rect 25506 19966 25508 20018
rect 25452 19964 25508 19966
rect 24668 18562 24724 18564
rect 24668 18510 24670 18562
rect 24670 18510 24722 18562
rect 24722 18510 24724 18562
rect 24668 18508 24724 18510
rect 26348 19906 26404 19908
rect 26348 19854 26350 19906
rect 26350 19854 26402 19906
rect 26402 19854 26404 19906
rect 26348 19852 26404 19854
rect 26124 19010 26180 19012
rect 26124 18958 26126 19010
rect 26126 18958 26178 19010
rect 26178 18958 26180 19010
rect 26124 18956 26180 18958
rect 26684 18956 26740 19012
rect 24780 18172 24836 18228
rect 24556 17276 24612 17332
rect 24444 17052 24500 17108
rect 23996 16658 24052 16660
rect 23996 16606 23998 16658
rect 23998 16606 24050 16658
rect 24050 16606 24052 16658
rect 23996 16604 24052 16606
rect 24220 16044 24276 16100
rect 24220 15260 24276 15316
rect 23884 14418 23940 14420
rect 23884 14366 23886 14418
rect 23886 14366 23938 14418
rect 23938 14366 23940 14418
rect 23884 14364 23940 14366
rect 23548 12684 23604 12740
rect 23436 11900 23492 11956
rect 22428 10108 22484 10164
rect 23100 11340 23156 11396
rect 22764 10668 22820 10724
rect 23212 11116 23268 11172
rect 23212 10610 23268 10612
rect 23212 10558 23214 10610
rect 23214 10558 23266 10610
rect 23266 10558 23268 10610
rect 23212 10556 23268 10558
rect 23548 10780 23604 10836
rect 22652 9996 22708 10052
rect 22540 9772 22596 9828
rect 22764 9212 22820 9268
rect 22316 7532 22372 7588
rect 22316 7362 22372 7364
rect 22316 7310 22318 7362
rect 22318 7310 22370 7362
rect 22370 7310 22372 7362
rect 22316 7308 22372 7310
rect 22988 9714 23044 9716
rect 22988 9662 22990 9714
rect 22990 9662 23042 9714
rect 23042 9662 23044 9714
rect 22988 9660 23044 9662
rect 23660 9266 23716 9268
rect 23660 9214 23662 9266
rect 23662 9214 23714 9266
rect 23714 9214 23716 9266
rect 23660 9212 23716 9214
rect 22988 9100 23044 9156
rect 23212 8930 23268 8932
rect 23212 8878 23214 8930
rect 23214 8878 23266 8930
rect 23266 8878 23268 8930
rect 23212 8876 23268 8878
rect 22540 8316 22596 8372
rect 23884 13580 23940 13636
rect 24668 16380 24724 16436
rect 24444 16268 24500 16324
rect 24780 16156 24836 16212
rect 24444 16098 24500 16100
rect 24444 16046 24446 16098
rect 24446 16046 24498 16098
rect 24498 16046 24500 16098
rect 24444 16044 24500 16046
rect 24332 14364 24388 14420
rect 23996 13356 24052 13412
rect 24220 13522 24276 13524
rect 24220 13470 24222 13522
rect 24222 13470 24274 13522
rect 24274 13470 24276 13522
rect 24220 13468 24276 13470
rect 24108 13244 24164 13300
rect 24220 12348 24276 12404
rect 24444 13746 24500 13748
rect 24444 13694 24446 13746
rect 24446 13694 24498 13746
rect 24498 13694 24500 13746
rect 24444 13692 24500 13694
rect 24556 13468 24612 13524
rect 24556 13186 24612 13188
rect 24556 13134 24558 13186
rect 24558 13134 24610 13186
rect 24610 13134 24612 13186
rect 24556 13132 24612 13134
rect 24444 12178 24500 12180
rect 24444 12126 24446 12178
rect 24446 12126 24498 12178
rect 24498 12126 24500 12178
rect 24444 12124 24500 12126
rect 23884 11788 23940 11844
rect 23884 11452 23940 11508
rect 24332 11394 24388 11396
rect 24332 11342 24334 11394
rect 24334 11342 24386 11394
rect 24386 11342 24388 11394
rect 24332 11340 24388 11342
rect 24220 11282 24276 11284
rect 24220 11230 24222 11282
rect 24222 11230 24274 11282
rect 24274 11230 24276 11282
rect 24220 11228 24276 11230
rect 24332 10556 24388 10612
rect 23548 8370 23604 8372
rect 23548 8318 23550 8370
rect 23550 8318 23602 8370
rect 23602 8318 23604 8370
rect 23548 8316 23604 8318
rect 23212 8092 23268 8148
rect 22652 6636 22708 6692
rect 23436 7474 23492 7476
rect 23436 7422 23438 7474
rect 23438 7422 23490 7474
rect 23490 7422 23492 7474
rect 23436 7420 23492 7422
rect 23212 6578 23268 6580
rect 23212 6526 23214 6578
rect 23214 6526 23266 6578
rect 23266 6526 23268 6578
rect 23212 6524 23268 6526
rect 22540 6300 22596 6356
rect 23212 6300 23268 6356
rect 22988 5628 23044 5684
rect 22316 5234 22372 5236
rect 22316 5182 22318 5234
rect 22318 5182 22370 5234
rect 22370 5182 22372 5234
rect 22316 5180 22372 5182
rect 22876 4956 22932 5012
rect 22652 4898 22708 4900
rect 22652 4846 22654 4898
rect 22654 4846 22706 4898
rect 22706 4846 22708 4898
rect 22652 4844 22708 4846
rect 21868 4396 21924 4452
rect 23548 7308 23604 7364
rect 23772 8316 23828 8372
rect 25676 18226 25732 18228
rect 25676 18174 25678 18226
rect 25678 18174 25730 18226
rect 25730 18174 25732 18226
rect 25676 18172 25732 18174
rect 26012 18060 26068 18116
rect 26348 18172 26404 18228
rect 25564 17948 25620 18004
rect 25900 17666 25956 17668
rect 25900 17614 25902 17666
rect 25902 17614 25954 17666
rect 25954 17614 25956 17666
rect 25900 17612 25956 17614
rect 26348 17554 26404 17556
rect 26348 17502 26350 17554
rect 26350 17502 26402 17554
rect 26402 17502 26404 17554
rect 26348 17500 26404 17502
rect 25564 17276 25620 17332
rect 25788 17388 25844 17444
rect 25004 16716 25060 16772
rect 24780 12796 24836 12852
rect 25452 16882 25508 16884
rect 25452 16830 25454 16882
rect 25454 16830 25506 16882
rect 25506 16830 25508 16882
rect 25452 16828 25508 16830
rect 25116 13804 25172 13860
rect 26124 17276 26180 17332
rect 26572 17276 26628 17332
rect 26572 16994 26628 16996
rect 26572 16942 26574 16994
rect 26574 16942 26626 16994
rect 26626 16942 26628 16994
rect 26572 16940 26628 16942
rect 26124 16828 26180 16884
rect 25900 15372 25956 15428
rect 25788 15314 25844 15316
rect 25788 15262 25790 15314
rect 25790 15262 25842 15314
rect 25842 15262 25844 15314
rect 25788 15260 25844 15262
rect 26684 16492 26740 16548
rect 26684 15484 26740 15540
rect 26124 15426 26180 15428
rect 26124 15374 26126 15426
rect 26126 15374 26178 15426
rect 26178 15374 26180 15426
rect 26124 15372 26180 15374
rect 25676 14364 25732 14420
rect 25340 13916 25396 13972
rect 25228 13580 25284 13636
rect 25340 13356 25396 13412
rect 25452 13132 25508 13188
rect 25788 14306 25844 14308
rect 25788 14254 25790 14306
rect 25790 14254 25842 14306
rect 25842 14254 25844 14306
rect 25788 14252 25844 14254
rect 25676 13692 25732 13748
rect 25788 14028 25844 14084
rect 25676 13522 25732 13524
rect 25676 13470 25678 13522
rect 25678 13470 25730 13522
rect 25730 13470 25732 13522
rect 25676 13468 25732 13470
rect 25564 13020 25620 13076
rect 26124 14028 26180 14084
rect 27132 23772 27188 23828
rect 27020 22930 27076 22932
rect 27020 22878 27022 22930
rect 27022 22878 27074 22930
rect 27074 22878 27076 22930
rect 27020 22876 27076 22878
rect 27020 21980 27076 22036
rect 26908 19906 26964 19908
rect 26908 19854 26910 19906
rect 26910 19854 26962 19906
rect 26962 19854 26964 19906
rect 26908 19852 26964 19854
rect 27244 23100 27300 23156
rect 27692 23826 27748 23828
rect 27692 23774 27694 23826
rect 27694 23774 27746 23826
rect 27746 23774 27748 23826
rect 27692 23772 27748 23774
rect 28028 22876 28084 22932
rect 27356 22482 27412 22484
rect 27356 22430 27358 22482
rect 27358 22430 27410 22482
rect 27410 22430 27412 22482
rect 27356 22428 27412 22430
rect 28028 21810 28084 21812
rect 28028 21758 28030 21810
rect 28030 21758 28082 21810
rect 28082 21758 28084 21810
rect 28028 21756 28084 21758
rect 27244 21644 27300 21700
rect 27692 20130 27748 20132
rect 27692 20078 27694 20130
rect 27694 20078 27746 20130
rect 27746 20078 27748 20130
rect 27692 20076 27748 20078
rect 27916 20076 27972 20132
rect 27132 19628 27188 19684
rect 27804 19740 27860 19796
rect 27020 19404 27076 19460
rect 27020 18732 27076 18788
rect 27356 19010 27412 19012
rect 27356 18958 27358 19010
rect 27358 18958 27410 19010
rect 27410 18958 27412 19010
rect 27356 18956 27412 18958
rect 27244 18508 27300 18564
rect 28028 19628 28084 19684
rect 27580 18732 27636 18788
rect 27356 18396 27412 18452
rect 27020 18284 27076 18340
rect 27356 18226 27412 18228
rect 27356 18174 27358 18226
rect 27358 18174 27410 18226
rect 27410 18174 27412 18226
rect 27356 18172 27412 18174
rect 27020 17666 27076 17668
rect 27020 17614 27022 17666
rect 27022 17614 27074 17666
rect 27074 17614 27076 17666
rect 27020 17612 27076 17614
rect 27580 17612 27636 17668
rect 27468 17554 27524 17556
rect 27468 17502 27470 17554
rect 27470 17502 27522 17554
rect 27522 17502 27524 17554
rect 27468 17500 27524 17502
rect 27132 17276 27188 17332
rect 27132 17052 27188 17108
rect 26796 15372 26852 15428
rect 27132 16882 27188 16884
rect 27132 16830 27134 16882
rect 27134 16830 27186 16882
rect 27186 16830 27188 16882
rect 27132 16828 27188 16830
rect 26908 15148 26964 15204
rect 27468 17276 27524 17332
rect 28140 18956 28196 19012
rect 28140 18732 28196 18788
rect 28028 18450 28084 18452
rect 28028 18398 28030 18450
rect 28030 18398 28082 18450
rect 28082 18398 28084 18450
rect 28028 18396 28084 18398
rect 34860 40962 34916 40964
rect 34860 40910 34862 40962
rect 34862 40910 34914 40962
rect 34914 40910 34916 40962
rect 34860 40908 34916 40910
rect 35196 40908 35252 40964
rect 35868 45948 35924 46004
rect 36540 46060 36596 46116
rect 37548 46956 37604 47012
rect 37996 46956 38052 47012
rect 38332 46844 38388 46900
rect 37884 46562 37940 46564
rect 37884 46510 37886 46562
rect 37886 46510 37938 46562
rect 37938 46510 37940 46562
rect 37884 46508 37940 46510
rect 37548 46396 37604 46452
rect 37996 46284 38052 46340
rect 40236 51324 40292 51380
rect 40012 50652 40068 50708
rect 40124 50540 40180 50596
rect 40348 50482 40404 50484
rect 40348 50430 40350 50482
rect 40350 50430 40402 50482
rect 40402 50430 40404 50482
rect 40348 50428 40404 50430
rect 39676 48972 39732 49028
rect 40012 50204 40068 50260
rect 40796 50428 40852 50484
rect 41020 50764 41076 50820
rect 41244 50540 41300 50596
rect 41356 50428 41412 50484
rect 40124 49756 40180 49812
rect 40012 49026 40068 49028
rect 40012 48974 40014 49026
rect 40014 48974 40066 49026
rect 40066 48974 40068 49026
rect 40012 48972 40068 48974
rect 37548 46060 37604 46116
rect 37324 45948 37380 46004
rect 37548 45724 37604 45780
rect 37100 45666 37156 45668
rect 37100 45614 37102 45666
rect 37102 45614 37154 45666
rect 37154 45614 37156 45666
rect 37100 45612 37156 45614
rect 37660 45612 37716 45668
rect 36876 44604 36932 44660
rect 38108 45778 38164 45780
rect 38108 45726 38110 45778
rect 38110 45726 38162 45778
rect 38162 45726 38164 45778
rect 38108 45724 38164 45726
rect 37996 45330 38052 45332
rect 37996 45278 37998 45330
rect 37998 45278 38050 45330
rect 38050 45278 38052 45330
rect 37996 45276 38052 45278
rect 38892 46956 38948 47012
rect 38780 46562 38836 46564
rect 38780 46510 38782 46562
rect 38782 46510 38834 46562
rect 38834 46510 38836 46562
rect 38780 46508 38836 46510
rect 41580 51772 41636 51828
rect 41804 51548 41860 51604
rect 42140 52946 42196 52948
rect 42140 52894 42142 52946
rect 42142 52894 42194 52946
rect 42194 52894 42196 52946
rect 42140 52892 42196 52894
rect 42364 52780 42420 52836
rect 42140 52162 42196 52164
rect 42140 52110 42142 52162
rect 42142 52110 42194 52162
rect 42194 52110 42196 52162
rect 42140 52108 42196 52110
rect 42364 52108 42420 52164
rect 41804 51266 41860 51268
rect 41804 51214 41806 51266
rect 41806 51214 41858 51266
rect 41858 51214 41860 51266
rect 41804 51212 41860 51214
rect 41916 50988 41972 51044
rect 42140 51884 42196 51940
rect 41692 50652 41748 50708
rect 42140 51378 42196 51380
rect 42140 51326 42142 51378
rect 42142 51326 42194 51378
rect 42194 51326 42196 51378
rect 42140 51324 42196 51326
rect 41692 50092 41748 50148
rect 40012 46844 40068 46900
rect 39004 45778 39060 45780
rect 39004 45726 39006 45778
rect 39006 45726 39058 45778
rect 39058 45726 39060 45778
rect 39004 45724 39060 45726
rect 39228 45388 39284 45444
rect 38780 45330 38836 45332
rect 38780 45278 38782 45330
rect 38782 45278 38834 45330
rect 38834 45278 38836 45330
rect 38780 45276 38836 45278
rect 38444 45106 38500 45108
rect 38444 45054 38446 45106
rect 38446 45054 38498 45106
rect 38498 45054 38500 45106
rect 38444 45052 38500 45054
rect 35980 44322 36036 44324
rect 35980 44270 35982 44322
rect 35982 44270 36034 44322
rect 36034 44270 36036 44322
rect 35980 44268 36036 44270
rect 37660 44322 37716 44324
rect 37660 44270 37662 44322
rect 37662 44270 37714 44322
rect 37714 44270 37716 44322
rect 37660 44268 37716 44270
rect 39452 44994 39508 44996
rect 39452 44942 39454 44994
rect 39454 44942 39506 44994
rect 39506 44942 39508 44994
rect 39452 44940 39508 44942
rect 39004 44828 39060 44884
rect 38220 44434 38276 44436
rect 38220 44382 38222 44434
rect 38222 44382 38274 44434
rect 38274 44382 38276 44434
rect 38220 44380 38276 44382
rect 36652 44044 36708 44100
rect 36092 43538 36148 43540
rect 36092 43486 36094 43538
rect 36094 43486 36146 43538
rect 36146 43486 36148 43538
rect 36092 43484 36148 43486
rect 35868 42812 35924 42868
rect 36204 43260 36260 43316
rect 36540 42924 36596 42980
rect 36316 42866 36372 42868
rect 36316 42814 36318 42866
rect 36318 42814 36370 42866
rect 36370 42814 36372 42866
rect 36316 42812 36372 42814
rect 36204 42754 36260 42756
rect 36204 42702 36206 42754
rect 36206 42702 36258 42754
rect 36258 42702 36260 42754
rect 36204 42700 36260 42702
rect 36092 40962 36148 40964
rect 36092 40910 36094 40962
rect 36094 40910 36146 40962
rect 36146 40910 36148 40962
rect 36092 40908 36148 40910
rect 35644 40460 35700 40516
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34636 39058 34692 39060
rect 34636 39006 34638 39058
rect 34638 39006 34690 39058
rect 34690 39006 34692 39058
rect 34636 39004 34692 39006
rect 35196 38834 35252 38836
rect 35196 38782 35198 38834
rect 35198 38782 35250 38834
rect 35250 38782 35252 38834
rect 35196 38780 35252 38782
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34748 37996 34804 38052
rect 35420 38050 35476 38052
rect 35420 37998 35422 38050
rect 35422 37998 35474 38050
rect 35474 37998 35476 38050
rect 35420 37996 35476 37998
rect 36540 40908 36596 40964
rect 36092 40348 36148 40404
rect 36092 39618 36148 39620
rect 36092 39566 36094 39618
rect 36094 39566 36146 39618
rect 36146 39566 36148 39618
rect 36092 39564 36148 39566
rect 35980 39228 36036 39284
rect 35756 37996 35812 38052
rect 35980 38780 36036 38836
rect 35084 37826 35140 37828
rect 35084 37774 35086 37826
rect 35086 37774 35138 37826
rect 35138 37774 35140 37826
rect 35084 37772 35140 37774
rect 34524 36652 34580 36708
rect 34412 35756 34468 35812
rect 34636 35586 34692 35588
rect 34636 35534 34638 35586
rect 34638 35534 34690 35586
rect 34690 35534 34692 35586
rect 34636 35532 34692 35534
rect 36652 39564 36708 39620
rect 36540 38892 36596 38948
rect 36316 38780 36372 38836
rect 36652 38444 36708 38500
rect 36316 37826 36372 37828
rect 36316 37774 36318 37826
rect 36318 37774 36370 37826
rect 36370 37774 36372 37826
rect 36316 37772 36372 37774
rect 35532 37266 35588 37268
rect 35532 37214 35534 37266
rect 35534 37214 35586 37266
rect 35586 37214 35588 37266
rect 35532 37212 35588 37214
rect 34860 36428 34916 36484
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35084 36428 35140 36484
rect 35308 36652 35364 36708
rect 34860 36258 34916 36260
rect 34860 36206 34862 36258
rect 34862 36206 34914 36258
rect 34914 36206 34916 36258
rect 34860 36204 34916 36206
rect 35420 36428 35476 36484
rect 34972 35420 35028 35476
rect 35084 35980 35140 36036
rect 35308 35810 35364 35812
rect 35308 35758 35310 35810
rect 35310 35758 35362 35810
rect 35362 35758 35364 35810
rect 35308 35756 35364 35758
rect 36316 37436 36372 37492
rect 35980 36482 36036 36484
rect 35980 36430 35982 36482
rect 35982 36430 36034 36482
rect 36034 36430 36036 36482
rect 35980 36428 36036 36430
rect 35084 35532 35140 35588
rect 34412 35026 34468 35028
rect 34412 34974 34414 35026
rect 34414 34974 34466 35026
rect 34466 34974 34468 35026
rect 34412 34972 34468 34974
rect 34860 34972 34916 35028
rect 33180 33964 33236 34020
rect 34300 34018 34356 34020
rect 34300 33966 34302 34018
rect 34302 33966 34354 34018
rect 34354 33966 34356 34018
rect 34300 33964 34356 33966
rect 34300 33234 34356 33236
rect 34300 33182 34302 33234
rect 34302 33182 34354 33234
rect 34354 33182 34356 33234
rect 34300 33180 34356 33182
rect 33628 33068 33684 33124
rect 33180 32956 33236 33012
rect 33740 32956 33796 33012
rect 33068 32562 33124 32564
rect 33068 32510 33070 32562
rect 33070 32510 33122 32562
rect 33122 32510 33124 32562
rect 33068 32508 33124 32510
rect 33628 32284 33684 32340
rect 33068 31724 33124 31780
rect 34188 31778 34244 31780
rect 34188 31726 34190 31778
rect 34190 31726 34242 31778
rect 34242 31726 34244 31778
rect 34188 31724 34244 31726
rect 34524 33068 34580 33124
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35644 34972 35700 35028
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34636 32956 34692 33012
rect 35196 32732 35252 32788
rect 34412 31612 34468 31668
rect 33292 31500 33348 31556
rect 33964 31106 34020 31108
rect 33964 31054 33966 31106
rect 33966 31054 34018 31106
rect 34018 31054 34020 31106
rect 33964 31052 34020 31054
rect 33404 30380 33460 30436
rect 33180 30268 33236 30324
rect 33068 30156 33124 30212
rect 32844 29372 32900 29428
rect 32844 27804 32900 27860
rect 30716 26124 30772 26180
rect 31612 26178 31668 26180
rect 31612 26126 31614 26178
rect 31614 26126 31666 26178
rect 31666 26126 31668 26178
rect 31612 26124 31668 26126
rect 28812 23772 28868 23828
rect 28476 23042 28532 23044
rect 28476 22990 28478 23042
rect 28478 22990 28530 23042
rect 28530 22990 28532 23042
rect 28476 22988 28532 22990
rect 29036 22876 29092 22932
rect 29260 22988 29316 23044
rect 29484 22428 29540 22484
rect 29372 22370 29428 22372
rect 29372 22318 29374 22370
rect 29374 22318 29426 22370
rect 29426 22318 29428 22370
rect 29372 22316 29428 22318
rect 30940 22316 30996 22372
rect 29484 21980 29540 22036
rect 30268 22092 30324 22148
rect 28588 21810 28644 21812
rect 28588 21758 28590 21810
rect 28590 21758 28642 21810
rect 28642 21758 28644 21810
rect 28588 21756 28644 21758
rect 28364 19740 28420 19796
rect 29036 18620 29092 18676
rect 28364 18450 28420 18452
rect 28364 18398 28366 18450
rect 28366 18398 28418 18450
rect 28418 18398 28420 18450
rect 28364 18396 28420 18398
rect 28812 18450 28868 18452
rect 28812 18398 28814 18450
rect 28814 18398 28866 18450
rect 28866 18398 28868 18450
rect 28812 18396 28868 18398
rect 29260 21532 29316 21588
rect 29484 21084 29540 21140
rect 30044 21084 30100 21140
rect 29372 20076 29428 20132
rect 29596 20018 29652 20020
rect 29596 19966 29598 20018
rect 29598 19966 29650 20018
rect 29650 19966 29652 20018
rect 29596 19964 29652 19966
rect 29932 19964 29988 20020
rect 29596 19010 29652 19012
rect 29596 18958 29598 19010
rect 29598 18958 29650 19010
rect 29650 18958 29652 19010
rect 29596 18956 29652 18958
rect 29820 18620 29876 18676
rect 30156 18844 30212 18900
rect 29484 18508 29540 18564
rect 28028 18172 28084 18228
rect 27916 17388 27972 17444
rect 28028 17106 28084 17108
rect 28028 17054 28030 17106
rect 28030 17054 28082 17106
rect 28082 17054 28084 17106
rect 28028 17052 28084 17054
rect 27916 15484 27972 15540
rect 28028 15426 28084 15428
rect 28028 15374 28030 15426
rect 28030 15374 28082 15426
rect 28082 15374 28084 15426
rect 28028 15372 28084 15374
rect 26796 14476 26852 14532
rect 26572 13746 26628 13748
rect 26572 13694 26574 13746
rect 26574 13694 26626 13746
rect 26626 13694 26628 13746
rect 26572 13692 26628 13694
rect 26460 13468 26516 13524
rect 26012 13356 26068 13412
rect 26348 13244 26404 13300
rect 25900 12962 25956 12964
rect 25900 12910 25902 12962
rect 25902 12910 25954 12962
rect 25954 12910 25956 12962
rect 25900 12908 25956 12910
rect 26908 14418 26964 14420
rect 26908 14366 26910 14418
rect 26910 14366 26962 14418
rect 26962 14366 26964 14418
rect 26908 14364 26964 14366
rect 26572 12908 26628 12964
rect 25564 12850 25620 12852
rect 25564 12798 25566 12850
rect 25566 12798 25618 12850
rect 25618 12798 25620 12850
rect 25564 12796 25620 12798
rect 24780 12124 24836 12180
rect 25228 12684 25284 12740
rect 25900 12684 25956 12740
rect 25900 12402 25956 12404
rect 25900 12350 25902 12402
rect 25902 12350 25954 12402
rect 25954 12350 25956 12402
rect 25900 12348 25956 12350
rect 25340 12178 25396 12180
rect 25340 12126 25342 12178
rect 25342 12126 25394 12178
rect 25394 12126 25396 12178
rect 25340 12124 25396 12126
rect 25228 11900 25284 11956
rect 27468 14252 27524 14308
rect 27244 12348 27300 12404
rect 27692 14700 27748 14756
rect 27468 12460 27524 12516
rect 27580 12850 27636 12852
rect 27580 12798 27582 12850
rect 27582 12798 27634 12850
rect 27634 12798 27636 12850
rect 27580 12796 27636 12798
rect 27580 12348 27636 12404
rect 28252 16994 28308 16996
rect 28252 16942 28254 16994
rect 28254 16942 28306 16994
rect 28306 16942 28308 16994
rect 28252 16940 28308 16942
rect 28364 16156 28420 16212
rect 28252 13916 28308 13972
rect 28364 14252 28420 14308
rect 27916 13858 27972 13860
rect 27916 13806 27918 13858
rect 27918 13806 27970 13858
rect 27970 13806 27972 13858
rect 27916 13804 27972 13806
rect 28252 12850 28308 12852
rect 28252 12798 28254 12850
rect 28254 12798 28306 12850
rect 28306 12798 28308 12850
rect 28252 12796 28308 12798
rect 28364 12348 28420 12404
rect 27244 12178 27300 12180
rect 27244 12126 27246 12178
rect 27246 12126 27298 12178
rect 27298 12126 27300 12178
rect 27244 12124 27300 12126
rect 28588 15090 28644 15092
rect 28588 15038 28590 15090
rect 28590 15038 28642 15090
rect 28642 15038 28644 15090
rect 28588 15036 28644 15038
rect 28812 15314 28868 15316
rect 28812 15262 28814 15314
rect 28814 15262 28866 15314
rect 28866 15262 28868 15314
rect 28812 15260 28868 15262
rect 29708 18450 29764 18452
rect 29708 18398 29710 18450
rect 29710 18398 29762 18450
rect 29762 18398 29764 18450
rect 29708 18396 29764 18398
rect 30044 18338 30100 18340
rect 30044 18286 30046 18338
rect 30046 18286 30098 18338
rect 30098 18286 30100 18338
rect 30044 18284 30100 18286
rect 29820 18172 29876 18228
rect 31052 21532 31108 21588
rect 31164 21868 31220 21924
rect 30940 20860 30996 20916
rect 30828 20018 30884 20020
rect 30828 19966 30830 20018
rect 30830 19966 30882 20018
rect 30882 19966 30884 20018
rect 30828 19964 30884 19966
rect 30492 18450 30548 18452
rect 30492 18398 30494 18450
rect 30494 18398 30546 18450
rect 30546 18398 30548 18450
rect 30492 18396 30548 18398
rect 30156 18060 30212 18116
rect 30380 18172 30436 18228
rect 29484 16268 29540 16324
rect 30716 18172 30772 18228
rect 30940 17612 30996 17668
rect 31052 17948 31108 18004
rect 31052 17554 31108 17556
rect 31052 17502 31054 17554
rect 31054 17502 31106 17554
rect 31106 17502 31108 17554
rect 31052 17500 31108 17502
rect 30940 17164 30996 17220
rect 30716 16380 30772 16436
rect 30044 16044 30100 16100
rect 29484 15372 29540 15428
rect 30156 15820 30212 15876
rect 29932 15426 29988 15428
rect 29932 15374 29934 15426
rect 29934 15374 29986 15426
rect 29986 15374 29988 15426
rect 29932 15372 29988 15374
rect 29596 15314 29652 15316
rect 29596 15262 29598 15314
rect 29598 15262 29650 15314
rect 29650 15262 29652 15314
rect 29596 15260 29652 15262
rect 29148 14700 29204 14756
rect 29148 14530 29204 14532
rect 29148 14478 29150 14530
rect 29150 14478 29202 14530
rect 29202 14478 29204 14530
rect 29148 14476 29204 14478
rect 29036 14306 29092 14308
rect 29036 14254 29038 14306
rect 29038 14254 29090 14306
rect 29090 14254 29092 14306
rect 29036 14252 29092 14254
rect 28700 14140 28756 14196
rect 28812 13970 28868 13972
rect 28812 13918 28814 13970
rect 28814 13918 28866 13970
rect 28866 13918 28868 13970
rect 28812 13916 28868 13918
rect 29484 12962 29540 12964
rect 29484 12910 29486 12962
rect 29486 12910 29538 12962
rect 29538 12910 29540 12962
rect 29484 12908 29540 12910
rect 28700 12178 28756 12180
rect 28700 12126 28702 12178
rect 28702 12126 28754 12178
rect 28754 12126 28756 12178
rect 28700 12124 28756 12126
rect 27916 12012 27972 12068
rect 27916 11788 27972 11844
rect 28140 11788 28196 11844
rect 27468 11394 27524 11396
rect 27468 11342 27470 11394
rect 27470 11342 27522 11394
rect 27522 11342 27524 11394
rect 27468 11340 27524 11342
rect 25228 10780 25284 10836
rect 25116 10668 25172 10724
rect 25564 10386 25620 10388
rect 25564 10334 25566 10386
rect 25566 10334 25618 10386
rect 25618 10334 25620 10386
rect 25564 10332 25620 10334
rect 26124 10834 26180 10836
rect 26124 10782 26126 10834
rect 26126 10782 26178 10834
rect 26178 10782 26180 10834
rect 26124 10780 26180 10782
rect 26572 10780 26628 10836
rect 26908 10780 26964 10836
rect 26124 10444 26180 10500
rect 26236 10332 26292 10388
rect 25900 10108 25956 10164
rect 26124 9714 26180 9716
rect 26124 9662 26126 9714
rect 26126 9662 26178 9714
rect 26178 9662 26180 9714
rect 26124 9660 26180 9662
rect 26908 10108 26964 10164
rect 25676 9548 25732 9604
rect 25676 8428 25732 8484
rect 23996 7420 24052 7476
rect 24220 7250 24276 7252
rect 24220 7198 24222 7250
rect 24222 7198 24274 7250
rect 24274 7198 24276 7250
rect 24220 7196 24276 7198
rect 26796 7196 26852 7252
rect 23548 5292 23604 5348
rect 23212 4956 23268 5012
rect 23548 4844 23604 4900
rect 28812 10722 28868 10724
rect 28812 10670 28814 10722
rect 28814 10670 28866 10722
rect 28866 10670 28868 10722
rect 28812 10668 28868 10670
rect 27692 9938 27748 9940
rect 27692 9886 27694 9938
rect 27694 9886 27746 9938
rect 27746 9886 27748 9938
rect 27692 9884 27748 9886
rect 28812 9884 28868 9940
rect 27916 9714 27972 9716
rect 27916 9662 27918 9714
rect 27918 9662 27970 9714
rect 27970 9662 27972 9714
rect 27916 9660 27972 9662
rect 28476 9714 28532 9716
rect 28476 9662 28478 9714
rect 28478 9662 28530 9714
rect 28530 9662 28532 9714
rect 28476 9660 28532 9662
rect 27804 8204 27860 8260
rect 28252 7586 28308 7588
rect 28252 7534 28254 7586
rect 28254 7534 28306 7586
rect 28306 7534 28308 7586
rect 28252 7532 28308 7534
rect 27244 7196 27300 7252
rect 28364 6412 28420 6468
rect 27580 6018 27636 6020
rect 27580 5966 27582 6018
rect 27582 5966 27634 6018
rect 27634 5966 27636 6018
rect 27580 5964 27636 5966
rect 26012 5234 26068 5236
rect 26012 5182 26014 5234
rect 26014 5182 26066 5234
rect 26066 5182 26068 5234
rect 26012 5180 26068 5182
rect 27692 4956 27748 5012
rect 28252 5180 28308 5236
rect 28700 6076 28756 6132
rect 29484 12178 29540 12180
rect 29484 12126 29486 12178
rect 29486 12126 29538 12178
rect 29538 12126 29540 12178
rect 29484 12124 29540 12126
rect 29372 11788 29428 11844
rect 29932 14252 29988 14308
rect 30156 14588 30212 14644
rect 30044 13356 30100 13412
rect 30044 12348 30100 12404
rect 30268 13858 30324 13860
rect 30268 13806 30270 13858
rect 30270 13806 30322 13858
rect 30322 13806 30324 13858
rect 30268 13804 30324 13806
rect 31052 14364 31108 14420
rect 30828 13020 30884 13076
rect 31052 13244 31108 13300
rect 30380 12124 30436 12180
rect 30716 12572 30772 12628
rect 31164 12572 31220 12628
rect 31052 12460 31108 12516
rect 30604 12012 30660 12068
rect 30268 11506 30324 11508
rect 30268 11454 30270 11506
rect 30270 11454 30322 11506
rect 30322 11454 30324 11506
rect 30268 11452 30324 11454
rect 30716 11452 30772 11508
rect 31052 10556 31108 10612
rect 29148 9714 29204 9716
rect 29148 9662 29150 9714
rect 29150 9662 29202 9714
rect 29202 9662 29204 9714
rect 29148 9660 29204 9662
rect 29372 7532 29428 7588
rect 29708 8764 29764 8820
rect 29372 6524 29428 6580
rect 29932 6578 29988 6580
rect 29932 6526 29934 6578
rect 29934 6526 29986 6578
rect 29986 6526 29988 6578
rect 29932 6524 29988 6526
rect 29148 6466 29204 6468
rect 29148 6414 29150 6466
rect 29150 6414 29202 6466
rect 29202 6414 29204 6466
rect 29148 6412 29204 6414
rect 31612 19964 31668 20020
rect 31612 19180 31668 19236
rect 32060 23266 32116 23268
rect 32060 23214 32062 23266
rect 32062 23214 32114 23266
rect 32114 23214 32116 23266
rect 32060 23212 32116 23214
rect 33292 29932 33348 29988
rect 34300 30044 34356 30100
rect 33628 29426 33684 29428
rect 33628 29374 33630 29426
rect 33630 29374 33682 29426
rect 33682 29374 33684 29426
rect 33628 29372 33684 29374
rect 33404 29260 33460 29316
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34748 30434 34804 30436
rect 34748 30382 34750 30434
rect 34750 30382 34802 30434
rect 34802 30382 34804 30434
rect 34748 30380 34804 30382
rect 34636 30268 34692 30324
rect 35420 30156 35476 30212
rect 34860 29986 34916 29988
rect 34860 29934 34862 29986
rect 34862 29934 34914 29986
rect 34914 29934 34916 29986
rect 34860 29932 34916 29934
rect 34972 29820 35028 29876
rect 35084 29932 35140 29988
rect 33852 28364 33908 28420
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35532 28476 35588 28532
rect 35084 28028 35140 28084
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35532 27186 35588 27188
rect 35532 27134 35534 27186
rect 35534 27134 35586 27186
rect 35586 27134 35588 27186
rect 35532 27132 35588 27134
rect 32396 27020 32452 27076
rect 36428 35026 36484 35028
rect 36428 34974 36430 35026
rect 36430 34974 36482 35026
rect 36482 34974 36484 35026
rect 36428 34972 36484 34974
rect 36204 34188 36260 34244
rect 37548 44098 37604 44100
rect 37548 44046 37550 44098
rect 37550 44046 37602 44098
rect 37602 44046 37604 44098
rect 37548 44044 37604 44046
rect 38668 44322 38724 44324
rect 38668 44270 38670 44322
rect 38670 44270 38722 44322
rect 38722 44270 38724 44322
rect 38668 44268 38724 44270
rect 36876 43538 36932 43540
rect 36876 43486 36878 43538
rect 36878 43486 36930 43538
rect 36930 43486 36932 43538
rect 36876 43484 36932 43486
rect 38444 44210 38500 44212
rect 38444 44158 38446 44210
rect 38446 44158 38498 44210
rect 38498 44158 38500 44210
rect 38444 44156 38500 44158
rect 39116 44098 39172 44100
rect 39116 44046 39118 44098
rect 39118 44046 39170 44098
rect 39170 44046 39172 44098
rect 39116 44044 39172 44046
rect 36988 42700 37044 42756
rect 37660 42754 37716 42756
rect 37660 42702 37662 42754
rect 37662 42702 37714 42754
rect 37714 42702 37716 42754
rect 37660 42700 37716 42702
rect 37548 42252 37604 42308
rect 37996 42194 38052 42196
rect 37996 42142 37998 42194
rect 37998 42142 38050 42194
rect 38050 42142 38052 42194
rect 37996 42140 38052 42142
rect 36988 41916 37044 41972
rect 38556 42812 38612 42868
rect 39228 43820 39284 43876
rect 39004 43596 39060 43652
rect 38780 42866 38836 42868
rect 38780 42814 38782 42866
rect 38782 42814 38834 42866
rect 38834 42814 38836 42866
rect 38780 42812 38836 42814
rect 38668 42700 38724 42756
rect 38108 41804 38164 41860
rect 38780 41916 38836 41972
rect 39340 43426 39396 43428
rect 39340 43374 39342 43426
rect 39342 43374 39394 43426
rect 39394 43374 39396 43426
rect 39340 43372 39396 43374
rect 39004 42140 39060 42196
rect 39564 42082 39620 42084
rect 39564 42030 39566 42082
rect 39566 42030 39618 42082
rect 39618 42030 39620 42082
rect 39564 42028 39620 42030
rect 40012 46284 40068 46340
rect 40012 45612 40068 45668
rect 40012 44268 40068 44324
rect 39900 44044 39956 44100
rect 39788 43650 39844 43652
rect 39788 43598 39790 43650
rect 39790 43598 39842 43650
rect 39842 43598 39844 43650
rect 39788 43596 39844 43598
rect 40348 47346 40404 47348
rect 40348 47294 40350 47346
rect 40350 47294 40402 47346
rect 40402 47294 40404 47346
rect 40348 47292 40404 47294
rect 40460 46620 40516 46676
rect 40460 44940 40516 44996
rect 39676 41916 39732 41972
rect 38444 41020 38500 41076
rect 38556 41804 38612 41860
rect 37212 40460 37268 40516
rect 37772 39618 37828 39620
rect 37772 39566 37774 39618
rect 37774 39566 37826 39618
rect 37826 39566 37828 39618
rect 37772 39564 37828 39566
rect 39228 41804 39284 41860
rect 36988 39058 37044 39060
rect 36988 39006 36990 39058
rect 36990 39006 37042 39058
rect 37042 39006 37044 39058
rect 36988 39004 37044 39006
rect 37772 39058 37828 39060
rect 37772 39006 37774 39058
rect 37774 39006 37826 39058
rect 37826 39006 37828 39058
rect 37772 39004 37828 39006
rect 37660 38834 37716 38836
rect 37660 38782 37662 38834
rect 37662 38782 37714 38834
rect 37714 38782 37716 38834
rect 37660 38780 37716 38782
rect 36988 38220 37044 38276
rect 37100 38444 37156 38500
rect 37660 38274 37716 38276
rect 37660 38222 37662 38274
rect 37662 38222 37714 38274
rect 37714 38222 37716 38274
rect 37660 38220 37716 38222
rect 37660 37884 37716 37940
rect 37772 36652 37828 36708
rect 39228 41186 39284 41188
rect 39228 41134 39230 41186
rect 39230 41134 39282 41186
rect 39282 41134 39284 41186
rect 39228 41132 39284 41134
rect 39900 41186 39956 41188
rect 39900 41134 39902 41186
rect 39902 41134 39954 41186
rect 39954 41134 39956 41186
rect 39900 41132 39956 41134
rect 39788 40962 39844 40964
rect 39788 40910 39790 40962
rect 39790 40910 39842 40962
rect 39842 40910 39844 40962
rect 39788 40908 39844 40910
rect 39900 40514 39956 40516
rect 39900 40462 39902 40514
rect 39902 40462 39954 40514
rect 39954 40462 39956 40514
rect 39900 40460 39956 40462
rect 41468 48300 41524 48356
rect 40908 48242 40964 48244
rect 40908 48190 40910 48242
rect 40910 48190 40962 48242
rect 40962 48190 40964 48242
rect 40908 48188 40964 48190
rect 41804 49810 41860 49812
rect 41804 49758 41806 49810
rect 41806 49758 41858 49810
rect 41858 49758 41860 49810
rect 41804 49756 41860 49758
rect 42700 51324 42756 51380
rect 42588 51212 42644 51268
rect 42588 50652 42644 50708
rect 42476 50594 42532 50596
rect 42476 50542 42478 50594
rect 42478 50542 42530 50594
rect 42530 50542 42532 50594
rect 42476 50540 42532 50542
rect 42364 50092 42420 50148
rect 43484 53116 43540 53172
rect 43708 53564 43764 53620
rect 43484 52892 43540 52948
rect 42924 52108 42980 52164
rect 43148 52108 43204 52164
rect 43260 51938 43316 51940
rect 43260 51886 43262 51938
rect 43262 51886 43314 51938
rect 43314 51886 43316 51938
rect 43260 51884 43316 51886
rect 43260 51378 43316 51380
rect 43260 51326 43262 51378
rect 43262 51326 43314 51378
rect 43314 51326 43316 51378
rect 43260 51324 43316 51326
rect 42812 50204 42868 50260
rect 42476 49756 42532 49812
rect 41916 48972 41972 49028
rect 41692 48300 41748 48356
rect 41020 47292 41076 47348
rect 41468 45724 41524 45780
rect 41916 48188 41972 48244
rect 41804 47346 41860 47348
rect 41804 47294 41806 47346
rect 41806 47294 41858 47346
rect 41858 47294 41860 47346
rect 41804 47292 41860 47294
rect 42028 47292 42084 47348
rect 41804 46674 41860 46676
rect 41804 46622 41806 46674
rect 41806 46622 41858 46674
rect 41858 46622 41860 46674
rect 41804 46620 41860 46622
rect 41804 45890 41860 45892
rect 41804 45838 41806 45890
rect 41806 45838 41858 45890
rect 41858 45838 41860 45890
rect 41804 45836 41860 45838
rect 41692 45500 41748 45556
rect 42140 46172 42196 46228
rect 42588 49138 42644 49140
rect 42588 49086 42590 49138
rect 42590 49086 42642 49138
rect 42642 49086 42644 49138
rect 42588 49084 42644 49086
rect 42700 48242 42756 48244
rect 42700 48190 42702 48242
rect 42702 48190 42754 48242
rect 42754 48190 42756 48242
rect 42700 48188 42756 48190
rect 42924 47516 42980 47572
rect 43820 53452 43876 53508
rect 44156 53452 44212 53508
rect 44380 53228 44436 53284
rect 45500 54348 45556 54404
rect 44828 53228 44884 53284
rect 44044 51660 44100 51716
rect 44940 52162 44996 52164
rect 44940 52110 44942 52162
rect 44942 52110 44994 52162
rect 44994 52110 44996 52162
rect 44940 52108 44996 52110
rect 43708 51490 43764 51492
rect 43708 51438 43710 51490
rect 43710 51438 43762 51490
rect 43762 51438 43764 51490
rect 43708 51436 43764 51438
rect 43932 50988 43988 51044
rect 43596 50204 43652 50260
rect 43820 50482 43876 50484
rect 43820 50430 43822 50482
rect 43822 50430 43874 50482
rect 43874 50430 43876 50482
rect 43820 50428 43876 50430
rect 44044 50764 44100 50820
rect 44156 50652 44212 50708
rect 42476 46898 42532 46900
rect 42476 46846 42478 46898
rect 42478 46846 42530 46898
rect 42530 46846 42532 46898
rect 42476 46844 42532 46846
rect 42252 46060 42308 46116
rect 42924 46674 42980 46676
rect 42924 46622 42926 46674
rect 42926 46622 42978 46674
rect 42978 46622 42980 46674
rect 42924 46620 42980 46622
rect 42140 45666 42196 45668
rect 42140 45614 42142 45666
rect 42142 45614 42194 45666
rect 42194 45614 42196 45666
rect 42140 45612 42196 45614
rect 41020 44828 41076 44884
rect 42924 45948 42980 46004
rect 43036 45890 43092 45892
rect 43036 45838 43038 45890
rect 43038 45838 43090 45890
rect 43090 45838 43092 45890
rect 43036 45836 43092 45838
rect 43260 45612 43316 45668
rect 42252 45106 42308 45108
rect 42252 45054 42254 45106
rect 42254 45054 42306 45106
rect 42306 45054 42308 45106
rect 42252 45052 42308 45054
rect 40796 44322 40852 44324
rect 40796 44270 40798 44322
rect 40798 44270 40850 44322
rect 40850 44270 40852 44322
rect 40796 44268 40852 44270
rect 42252 44492 42308 44548
rect 40572 44044 40628 44100
rect 41244 43820 41300 43876
rect 40460 43708 40516 43764
rect 41132 43708 41188 43764
rect 40236 43148 40292 43204
rect 40124 42476 40180 42532
rect 40572 42866 40628 42868
rect 40572 42814 40574 42866
rect 40574 42814 40626 42866
rect 40626 42814 40628 42866
rect 40572 42812 40628 42814
rect 41020 41970 41076 41972
rect 41020 41918 41022 41970
rect 41022 41918 41074 41970
rect 41074 41918 41076 41970
rect 41020 41916 41076 41918
rect 40236 41804 40292 41860
rect 40124 41746 40180 41748
rect 40124 41694 40126 41746
rect 40126 41694 40178 41746
rect 40178 41694 40180 41746
rect 40124 41692 40180 41694
rect 40124 41356 40180 41412
rect 40124 40908 40180 40964
rect 38220 38220 38276 38276
rect 38780 37884 38836 37940
rect 38780 37266 38836 37268
rect 38780 37214 38782 37266
rect 38782 37214 38834 37266
rect 38834 37214 38836 37266
rect 38780 37212 38836 37214
rect 36988 35868 37044 35924
rect 36876 35532 36932 35588
rect 36764 34524 36820 34580
rect 36428 32620 36484 32676
rect 35868 30044 35924 30100
rect 35868 29426 35924 29428
rect 35868 29374 35870 29426
rect 35870 29374 35922 29426
rect 35922 29374 35924 29426
rect 35868 29372 35924 29374
rect 36428 30098 36484 30100
rect 36428 30046 36430 30098
rect 36430 30046 36482 30098
rect 36482 30046 36484 30098
rect 36428 30044 36484 30046
rect 36316 29484 36372 29540
rect 36428 28530 36484 28532
rect 36428 28478 36430 28530
rect 36430 28478 36482 28530
rect 36482 28478 36484 28530
rect 36428 28476 36484 28478
rect 35980 27746 36036 27748
rect 35980 27694 35982 27746
rect 35982 27694 36034 27746
rect 36034 27694 36036 27746
rect 35980 27692 36036 27694
rect 36428 27356 36484 27412
rect 37100 34860 37156 34916
rect 38108 35644 38164 35700
rect 38332 36258 38388 36260
rect 38332 36206 38334 36258
rect 38334 36206 38386 36258
rect 38386 36206 38388 36258
rect 38332 36204 38388 36206
rect 41244 41692 41300 41748
rect 41356 42588 41412 42644
rect 41132 41244 41188 41300
rect 40572 40460 40628 40516
rect 40348 39788 40404 39844
rect 39900 39228 39956 39284
rect 39452 37266 39508 37268
rect 39452 37214 39454 37266
rect 39454 37214 39506 37266
rect 39506 37214 39508 37266
rect 39452 37212 39508 37214
rect 39340 36988 39396 37044
rect 39228 36876 39284 36932
rect 39116 36370 39172 36372
rect 39116 36318 39118 36370
rect 39118 36318 39170 36370
rect 39170 36318 39172 36370
rect 39116 36316 39172 36318
rect 38892 35698 38948 35700
rect 38892 35646 38894 35698
rect 38894 35646 38946 35698
rect 38946 35646 38948 35698
rect 38892 35644 38948 35646
rect 38220 34914 38276 34916
rect 38220 34862 38222 34914
rect 38222 34862 38274 34914
rect 38274 34862 38276 34914
rect 38220 34860 38276 34862
rect 37100 34188 37156 34244
rect 37996 34242 38052 34244
rect 37996 34190 37998 34242
rect 37998 34190 38050 34242
rect 38050 34190 38052 34242
rect 37996 34188 38052 34190
rect 38668 34076 38724 34132
rect 37100 33122 37156 33124
rect 37100 33070 37102 33122
rect 37102 33070 37154 33122
rect 37154 33070 37156 33122
rect 37100 33068 37156 33070
rect 39228 36258 39284 36260
rect 39228 36206 39230 36258
rect 39230 36206 39282 36258
rect 39282 36206 39284 36258
rect 39228 36204 39284 36206
rect 39452 33852 39508 33908
rect 39564 35084 39620 35140
rect 39788 36876 39844 36932
rect 40124 35810 40180 35812
rect 40124 35758 40126 35810
rect 40126 35758 40178 35810
rect 40178 35758 40180 35810
rect 40124 35756 40180 35758
rect 36988 31778 37044 31780
rect 36988 31726 36990 31778
rect 36990 31726 37042 31778
rect 37042 31726 37044 31778
rect 36988 31724 37044 31726
rect 37212 32620 37268 32676
rect 37660 32674 37716 32676
rect 37660 32622 37662 32674
rect 37662 32622 37714 32674
rect 37714 32622 37716 32674
rect 37660 32620 37716 32622
rect 37660 31666 37716 31668
rect 37660 31614 37662 31666
rect 37662 31614 37714 31666
rect 37714 31614 37716 31666
rect 37660 31612 37716 31614
rect 37324 31500 37380 31556
rect 38108 31612 38164 31668
rect 37884 31500 37940 31556
rect 37100 29484 37156 29540
rect 36988 29260 37044 29316
rect 36988 28028 37044 28084
rect 37548 31218 37604 31220
rect 37548 31166 37550 31218
rect 37550 31166 37602 31218
rect 37602 31166 37604 31218
rect 37548 31164 37604 31166
rect 37324 31106 37380 31108
rect 37324 31054 37326 31106
rect 37326 31054 37378 31106
rect 37378 31054 37380 31106
rect 37324 31052 37380 31054
rect 38220 31052 38276 31108
rect 38220 30322 38276 30324
rect 38220 30270 38222 30322
rect 38222 30270 38274 30322
rect 38274 30270 38276 30322
rect 38220 30268 38276 30270
rect 37884 30156 37940 30212
rect 37772 30044 37828 30100
rect 37324 29596 37380 29652
rect 38780 31778 38836 31780
rect 38780 31726 38782 31778
rect 38782 31726 38834 31778
rect 38834 31726 38836 31778
rect 38780 31724 38836 31726
rect 38892 31666 38948 31668
rect 38892 31614 38894 31666
rect 38894 31614 38946 31666
rect 38946 31614 38948 31666
rect 38892 31612 38948 31614
rect 39340 31778 39396 31780
rect 39340 31726 39342 31778
rect 39342 31726 39394 31778
rect 39394 31726 39396 31778
rect 39340 31724 39396 31726
rect 39676 31612 39732 31668
rect 39788 31388 39844 31444
rect 39228 31164 39284 31220
rect 38892 31052 38948 31108
rect 39228 30268 39284 30324
rect 38780 30210 38836 30212
rect 38780 30158 38782 30210
rect 38782 30158 38834 30210
rect 38834 30158 38836 30210
rect 38780 30156 38836 30158
rect 38556 29596 38612 29652
rect 38780 29484 38836 29540
rect 37324 29260 37380 29316
rect 37324 28476 37380 28532
rect 37436 28364 37492 28420
rect 36764 27356 36820 27412
rect 37212 27580 37268 27636
rect 37100 26908 37156 26964
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 32508 24834 32564 24836
rect 32508 24782 32510 24834
rect 32510 24782 32562 24834
rect 32562 24782 32564 24834
rect 32508 24780 32564 24782
rect 32396 23938 32452 23940
rect 32396 23886 32398 23938
rect 32398 23886 32450 23938
rect 32450 23886 32452 23938
rect 32396 23884 32452 23886
rect 33180 23826 33236 23828
rect 33180 23774 33182 23826
rect 33182 23774 33234 23826
rect 33234 23774 33236 23826
rect 33180 23772 33236 23774
rect 32620 23436 32676 23492
rect 33180 23266 33236 23268
rect 33180 23214 33182 23266
rect 33182 23214 33234 23266
rect 33234 23214 33236 23266
rect 33180 23212 33236 23214
rect 33292 22428 33348 22484
rect 33516 22930 33572 22932
rect 33516 22878 33518 22930
rect 33518 22878 33570 22930
rect 33570 22878 33572 22930
rect 33516 22876 33572 22878
rect 32508 22204 32564 22260
rect 33180 22316 33236 22372
rect 32396 21644 32452 21700
rect 32284 21586 32340 21588
rect 32284 21534 32286 21586
rect 32286 21534 32338 21586
rect 32338 21534 32340 21586
rect 32284 21532 32340 21534
rect 32060 20914 32116 20916
rect 32060 20862 32062 20914
rect 32062 20862 32114 20914
rect 32114 20862 32116 20914
rect 32060 20860 32116 20862
rect 33292 22204 33348 22260
rect 32396 20578 32452 20580
rect 32396 20526 32398 20578
rect 32398 20526 32450 20578
rect 32450 20526 32452 20578
rect 32396 20524 32452 20526
rect 31388 16380 31444 16436
rect 31388 15372 31444 15428
rect 32284 19404 32340 19460
rect 32060 18620 32116 18676
rect 32396 18674 32452 18676
rect 32396 18622 32398 18674
rect 32398 18622 32450 18674
rect 32450 18622 32452 18674
rect 32396 18620 32452 18622
rect 32620 19964 32676 20020
rect 36876 26684 36932 26740
rect 37436 27132 37492 27188
rect 38668 29202 38724 29204
rect 38668 29150 38670 29202
rect 38670 29150 38722 29202
rect 38722 29150 38724 29202
rect 38668 29148 38724 29150
rect 38444 28754 38500 28756
rect 38444 28702 38446 28754
rect 38446 28702 38498 28754
rect 38498 28702 38500 28754
rect 38444 28700 38500 28702
rect 39788 30828 39844 30884
rect 40012 30380 40068 30436
rect 39564 29372 39620 29428
rect 39228 28812 39284 28868
rect 39452 28812 39508 28868
rect 39116 28700 39172 28756
rect 39676 28700 39732 28756
rect 40460 39058 40516 39060
rect 40460 39006 40462 39058
rect 40462 39006 40514 39058
rect 40514 39006 40516 39058
rect 40460 39004 40516 39006
rect 40908 41074 40964 41076
rect 40908 41022 40910 41074
rect 40910 41022 40962 41074
rect 40962 41022 40964 41074
rect 40908 41020 40964 41022
rect 40796 40460 40852 40516
rect 41244 41020 41300 41076
rect 41468 42530 41524 42532
rect 41468 42478 41470 42530
rect 41470 42478 41522 42530
rect 41522 42478 41524 42530
rect 41468 42476 41524 42478
rect 41468 42028 41524 42084
rect 41468 41692 41524 41748
rect 41580 41970 41636 41972
rect 41580 41918 41582 41970
rect 41582 41918 41634 41970
rect 41634 41918 41636 41970
rect 41580 41916 41636 41918
rect 41020 40908 41076 40964
rect 41468 39788 41524 39844
rect 41020 39116 41076 39172
rect 40684 38220 40740 38276
rect 41132 38780 41188 38836
rect 41356 39228 41412 39284
rect 43372 45164 43428 45220
rect 42476 44156 42532 44212
rect 43036 44716 43092 44772
rect 43260 44492 43316 44548
rect 42924 43820 42980 43876
rect 43036 44156 43092 44212
rect 42476 43538 42532 43540
rect 42476 43486 42478 43538
rect 42478 43486 42530 43538
rect 42530 43486 42532 43538
rect 42476 43484 42532 43486
rect 42812 43538 42868 43540
rect 42812 43486 42814 43538
rect 42814 43486 42866 43538
rect 42866 43486 42868 43538
rect 42812 43484 42868 43486
rect 43484 43484 43540 43540
rect 42476 42866 42532 42868
rect 42476 42814 42478 42866
rect 42478 42814 42530 42866
rect 42530 42814 42532 42866
rect 42476 42812 42532 42814
rect 42364 42642 42420 42644
rect 42364 42590 42366 42642
rect 42366 42590 42418 42642
rect 42418 42590 42420 42642
rect 42364 42588 42420 42590
rect 42812 42754 42868 42756
rect 42812 42702 42814 42754
rect 42814 42702 42866 42754
rect 42866 42702 42868 42754
rect 42812 42700 42868 42702
rect 42924 42642 42980 42644
rect 42924 42590 42926 42642
rect 42926 42590 42978 42642
rect 42978 42590 42980 42642
rect 42924 42588 42980 42590
rect 43820 49308 43876 49364
rect 43932 49026 43988 49028
rect 43932 48974 43934 49026
rect 43934 48974 43986 49026
rect 43986 48974 43988 49026
rect 43932 48972 43988 48974
rect 43820 48860 43876 48916
rect 43708 47292 43764 47348
rect 43820 46396 43876 46452
rect 43708 45612 43764 45668
rect 43932 45500 43988 45556
rect 43708 44604 43764 44660
rect 43820 45276 43876 45332
rect 45276 51660 45332 51716
rect 45276 51378 45332 51380
rect 45276 51326 45278 51378
rect 45278 51326 45330 51378
rect 45330 51326 45332 51378
rect 45276 51324 45332 51326
rect 46284 54402 46340 54404
rect 46284 54350 46286 54402
rect 46286 54350 46338 54402
rect 46338 54350 46340 54402
rect 46284 54348 46340 54350
rect 46620 53228 46676 53284
rect 45724 51378 45780 51380
rect 45724 51326 45726 51378
rect 45726 51326 45778 51378
rect 45778 51326 45780 51378
rect 45724 51324 45780 51326
rect 44940 49868 44996 49924
rect 44380 48748 44436 48804
rect 44380 48466 44436 48468
rect 44380 48414 44382 48466
rect 44382 48414 44434 48466
rect 44434 48414 44436 48466
rect 44380 48412 44436 48414
rect 44380 47964 44436 48020
rect 44156 47570 44212 47572
rect 44156 47518 44158 47570
rect 44158 47518 44210 47570
rect 44210 47518 44212 47570
rect 44156 47516 44212 47518
rect 44268 47458 44324 47460
rect 44268 47406 44270 47458
rect 44270 47406 44322 47458
rect 44322 47406 44324 47458
rect 44268 47404 44324 47406
rect 44380 46898 44436 46900
rect 44380 46846 44382 46898
rect 44382 46846 44434 46898
rect 44434 46846 44436 46898
rect 44380 46844 44436 46846
rect 44828 49084 44884 49140
rect 45276 48972 45332 49028
rect 44828 48188 44884 48244
rect 45276 48748 45332 48804
rect 46508 51324 46564 51380
rect 46844 52108 46900 52164
rect 46844 50594 46900 50596
rect 46844 50542 46846 50594
rect 46846 50542 46898 50594
rect 46898 50542 46900 50594
rect 46844 50540 46900 50542
rect 46396 50428 46452 50484
rect 47516 53452 47572 53508
rect 47068 53170 47124 53172
rect 47068 53118 47070 53170
rect 47070 53118 47122 53170
rect 47122 53118 47124 53170
rect 47068 53116 47124 53118
rect 48076 53170 48132 53172
rect 48076 53118 48078 53170
rect 48078 53118 48130 53170
rect 48130 53118 48132 53170
rect 48076 53116 48132 53118
rect 47180 51772 47236 51828
rect 47404 51660 47460 51716
rect 47180 50540 47236 50596
rect 45836 49644 45892 49700
rect 45500 49420 45556 49476
rect 45724 49308 45780 49364
rect 45836 49084 45892 49140
rect 45388 48412 45444 48468
rect 45724 48466 45780 48468
rect 45724 48414 45726 48466
rect 45726 48414 45778 48466
rect 45778 48414 45780 48466
rect 45724 48412 45780 48414
rect 46284 49810 46340 49812
rect 46284 49758 46286 49810
rect 46286 49758 46338 49810
rect 46338 49758 46340 49810
rect 46284 49756 46340 49758
rect 46172 49420 46228 49476
rect 46284 49026 46340 49028
rect 46284 48974 46286 49026
rect 46286 48974 46338 49026
rect 46338 48974 46340 49026
rect 46284 48972 46340 48974
rect 46172 48914 46228 48916
rect 46172 48862 46174 48914
rect 46174 48862 46226 48914
rect 46226 48862 46228 48914
rect 46172 48860 46228 48862
rect 46060 48802 46116 48804
rect 46060 48750 46062 48802
rect 46062 48750 46114 48802
rect 46114 48750 46116 48802
rect 46060 48748 46116 48750
rect 46620 50316 46676 50372
rect 48860 53116 48916 53172
rect 49420 53452 49476 53508
rect 48188 52834 48244 52836
rect 48188 52782 48190 52834
rect 48190 52782 48242 52834
rect 48242 52782 48244 52834
rect 48188 52780 48244 52782
rect 48300 52444 48356 52500
rect 48076 52162 48132 52164
rect 48076 52110 48078 52162
rect 48078 52110 48130 52162
rect 48130 52110 48132 52162
rect 48076 52108 48132 52110
rect 47964 51548 48020 51604
rect 47740 51324 47796 51380
rect 47180 50316 47236 50372
rect 46956 49810 47012 49812
rect 46956 49758 46958 49810
rect 46958 49758 47010 49810
rect 47010 49758 47012 49810
rect 46956 49756 47012 49758
rect 46844 49196 46900 49252
rect 46732 49084 46788 49140
rect 47292 49532 47348 49588
rect 48076 49868 48132 49924
rect 47964 49756 48020 49812
rect 45052 48354 45108 48356
rect 45052 48302 45054 48354
rect 45054 48302 45106 48354
rect 45106 48302 45108 48354
rect 45052 48300 45108 48302
rect 45164 48188 45220 48244
rect 45500 47740 45556 47796
rect 44940 47404 44996 47460
rect 44828 47292 44884 47348
rect 44604 46956 44660 47012
rect 44604 46172 44660 46228
rect 44268 45948 44324 46004
rect 44268 45666 44324 45668
rect 44268 45614 44270 45666
rect 44270 45614 44322 45666
rect 44322 45614 44324 45666
rect 44268 45612 44324 45614
rect 44044 45164 44100 45220
rect 44380 44940 44436 44996
rect 43596 42924 43652 42980
rect 43036 41692 43092 41748
rect 41804 41244 41860 41300
rect 41916 41356 41972 41412
rect 41804 41020 41860 41076
rect 42028 40626 42084 40628
rect 42028 40574 42030 40626
rect 42030 40574 42082 40626
rect 42082 40574 42084 40626
rect 42028 40572 42084 40574
rect 42140 39452 42196 39508
rect 41468 38892 41524 38948
rect 41916 39116 41972 39172
rect 41468 38108 41524 38164
rect 43036 40684 43092 40740
rect 42588 39788 42644 39844
rect 42700 40572 42756 40628
rect 42252 39004 42308 39060
rect 42476 38892 42532 38948
rect 41804 38668 41860 38724
rect 41916 38556 41972 38612
rect 41692 37212 41748 37268
rect 41244 36988 41300 37044
rect 40908 36316 40964 36372
rect 41580 35810 41636 35812
rect 41580 35758 41582 35810
rect 41582 35758 41634 35810
rect 41634 35758 41636 35810
rect 41580 35756 41636 35758
rect 41132 35532 41188 35588
rect 40908 35308 40964 35364
rect 40460 35084 40516 35140
rect 40684 34860 40740 34916
rect 40796 34802 40852 34804
rect 40796 34750 40798 34802
rect 40798 34750 40850 34802
rect 40850 34750 40852 34802
rect 40796 34748 40852 34750
rect 41804 34914 41860 34916
rect 41804 34862 41806 34914
rect 41806 34862 41858 34914
rect 41858 34862 41860 34914
rect 41804 34860 41860 34862
rect 41132 33964 41188 34020
rect 42924 40402 42980 40404
rect 42924 40350 42926 40402
rect 42926 40350 42978 40402
rect 42978 40350 42980 40402
rect 42924 40348 42980 40350
rect 42924 39676 42980 39732
rect 42812 39452 42868 39508
rect 42588 38722 42644 38724
rect 42588 38670 42590 38722
rect 42590 38670 42642 38722
rect 42642 38670 42644 38722
rect 42588 38668 42644 38670
rect 42476 37996 42532 38052
rect 42252 37548 42308 37604
rect 42140 36764 42196 36820
rect 42028 35532 42084 35588
rect 41916 33964 41972 34020
rect 42028 34076 42084 34132
rect 40236 33852 40292 33908
rect 42364 37266 42420 37268
rect 42364 37214 42366 37266
rect 42366 37214 42418 37266
rect 42418 37214 42420 37266
rect 42364 37212 42420 37214
rect 42700 38162 42756 38164
rect 42700 38110 42702 38162
rect 42702 38110 42754 38162
rect 42754 38110 42756 38162
rect 42700 38108 42756 38110
rect 42700 37884 42756 37940
rect 43036 36988 43092 37044
rect 42812 35756 42868 35812
rect 42700 34914 42756 34916
rect 42700 34862 42702 34914
rect 42702 34862 42754 34914
rect 42754 34862 42756 34914
rect 42700 34860 42756 34862
rect 43596 41970 43652 41972
rect 43596 41918 43598 41970
rect 43598 41918 43650 41970
rect 43650 41918 43652 41970
rect 43596 41916 43652 41918
rect 43372 40962 43428 40964
rect 43372 40910 43374 40962
rect 43374 40910 43426 40962
rect 43426 40910 43428 40962
rect 43372 40908 43428 40910
rect 43372 40684 43428 40740
rect 43148 36764 43204 36820
rect 43148 36370 43204 36372
rect 43148 36318 43150 36370
rect 43150 36318 43202 36370
rect 43202 36318 43204 36370
rect 43148 36316 43204 36318
rect 43596 40626 43652 40628
rect 43596 40574 43598 40626
rect 43598 40574 43650 40626
rect 43650 40574 43652 40626
rect 43596 40572 43652 40574
rect 43484 40124 43540 40180
rect 43484 39788 43540 39844
rect 43596 38946 43652 38948
rect 43596 38894 43598 38946
rect 43598 38894 43650 38946
rect 43650 38894 43652 38946
rect 43596 38892 43652 38894
rect 43820 41020 43876 41076
rect 43820 40402 43876 40404
rect 43820 40350 43822 40402
rect 43822 40350 43874 40402
rect 43874 40350 43876 40402
rect 43820 40348 43876 40350
rect 44492 44156 44548 44212
rect 44380 43484 44436 43540
rect 44268 42754 44324 42756
rect 44268 42702 44270 42754
rect 44270 42702 44322 42754
rect 44322 42702 44324 42754
rect 44268 42700 44324 42702
rect 44156 41916 44212 41972
rect 44380 40402 44436 40404
rect 44380 40350 44382 40402
rect 44382 40350 44434 40402
rect 44434 40350 44436 40402
rect 44380 40348 44436 40350
rect 43932 39676 43988 39732
rect 44156 39116 44212 39172
rect 43484 38780 43540 38836
rect 43372 37548 43428 37604
rect 44380 39058 44436 39060
rect 44380 39006 44382 39058
rect 44382 39006 44434 39058
rect 44434 39006 44436 39058
rect 44380 39004 44436 39006
rect 44716 45106 44772 45108
rect 44716 45054 44718 45106
rect 44718 45054 44770 45106
rect 44770 45054 44772 45106
rect 44716 45052 44772 45054
rect 44940 45106 44996 45108
rect 44940 45054 44942 45106
rect 44942 45054 44994 45106
rect 44994 45054 44996 45106
rect 44940 45052 44996 45054
rect 46956 48860 47012 48916
rect 46844 48412 46900 48468
rect 46172 47516 46228 47572
rect 45724 47180 45780 47236
rect 45164 46172 45220 46228
rect 45388 45836 45444 45892
rect 45164 45276 45220 45332
rect 45388 45164 45444 45220
rect 45612 46844 45668 46900
rect 45612 46396 45668 46452
rect 45836 45948 45892 46004
rect 46284 46844 46340 46900
rect 46508 46844 46564 46900
rect 46396 46284 46452 46340
rect 45276 44994 45332 44996
rect 45276 44942 45278 44994
rect 45278 44942 45330 44994
rect 45330 44942 45332 44994
rect 45276 44940 45332 44942
rect 45500 44828 45556 44884
rect 45276 44716 45332 44772
rect 45276 43708 45332 43764
rect 45164 43148 45220 43204
rect 44940 42812 44996 42868
rect 45164 42700 45220 42756
rect 45724 44210 45780 44212
rect 45724 44158 45726 44210
rect 45726 44158 45778 44210
rect 45778 44158 45780 44210
rect 45724 44156 45780 44158
rect 46396 46060 46452 46116
rect 46060 45276 46116 45332
rect 45948 44156 46004 44212
rect 46172 43596 46228 43652
rect 45836 43484 45892 43540
rect 44828 41468 44884 41524
rect 44940 40908 44996 40964
rect 45276 41468 45332 41524
rect 44716 40460 44772 40516
rect 44604 39228 44660 39284
rect 45164 39618 45220 39620
rect 45164 39566 45166 39618
rect 45166 39566 45218 39618
rect 45218 39566 45220 39618
rect 45164 39564 45220 39566
rect 44604 38892 44660 38948
rect 44716 38780 44772 38836
rect 43932 38220 43988 38276
rect 43820 37996 43876 38052
rect 45500 40402 45556 40404
rect 45500 40350 45502 40402
rect 45502 40350 45554 40402
rect 45554 40350 45556 40402
rect 45500 40348 45556 40350
rect 45388 39900 45444 39956
rect 45836 42866 45892 42868
rect 45836 42814 45838 42866
rect 45838 42814 45890 42866
rect 45890 42814 45892 42866
rect 45836 42812 45892 42814
rect 46284 41916 46340 41972
rect 45836 41692 45892 41748
rect 45836 39900 45892 39956
rect 46060 39564 46116 39620
rect 46172 40236 46228 40292
rect 45276 38332 45332 38388
rect 44604 37490 44660 37492
rect 44604 37438 44606 37490
rect 44606 37438 44658 37490
rect 44658 37438 44660 37490
rect 44604 37436 44660 37438
rect 43820 37212 43876 37268
rect 43708 37154 43764 37156
rect 43708 37102 43710 37154
rect 43710 37102 43762 37154
rect 43762 37102 43764 37154
rect 43708 37100 43764 37102
rect 43372 36876 43428 36932
rect 43372 36482 43428 36484
rect 43372 36430 43374 36482
rect 43374 36430 43426 36482
rect 43426 36430 43428 36482
rect 43372 36428 43428 36430
rect 43484 36764 43540 36820
rect 44156 36594 44212 36596
rect 44156 36542 44158 36594
rect 44158 36542 44210 36594
rect 44210 36542 44212 36594
rect 44156 36540 44212 36542
rect 43484 35756 43540 35812
rect 43036 35308 43092 35364
rect 43484 34748 43540 34804
rect 43036 34130 43092 34132
rect 43036 34078 43038 34130
rect 43038 34078 43090 34130
rect 43090 34078 43092 34130
rect 43036 34076 43092 34078
rect 42588 33852 42644 33908
rect 44380 36316 44436 36372
rect 44268 35980 44324 36036
rect 44492 35810 44548 35812
rect 44492 35758 44494 35810
rect 44494 35758 44546 35810
rect 44546 35758 44548 35810
rect 44492 35756 44548 35758
rect 45164 37266 45220 37268
rect 45164 37214 45166 37266
rect 45166 37214 45218 37266
rect 45218 37214 45220 37266
rect 45164 37212 45220 37214
rect 45500 36876 45556 36932
rect 45388 35980 45444 36036
rect 45052 34972 45108 35028
rect 45388 34690 45444 34692
rect 45388 34638 45390 34690
rect 45390 34638 45442 34690
rect 45442 34638 45444 34690
rect 45388 34636 45444 34638
rect 43932 34524 43988 34580
rect 43596 33852 43652 33908
rect 44604 33852 44660 33908
rect 40236 31778 40292 31780
rect 40236 31726 40238 31778
rect 40238 31726 40290 31778
rect 40290 31726 40292 31778
rect 40236 31724 40292 31726
rect 40236 31218 40292 31220
rect 40236 31166 40238 31218
rect 40238 31166 40290 31218
rect 40290 31166 40292 31218
rect 40236 31164 40292 31166
rect 40796 31052 40852 31108
rect 40348 30828 40404 30884
rect 41468 32508 41524 32564
rect 41356 31890 41412 31892
rect 41356 31838 41358 31890
rect 41358 31838 41410 31890
rect 41410 31838 41412 31890
rect 41356 31836 41412 31838
rect 41356 31500 41412 31556
rect 41132 31164 41188 31220
rect 41244 31388 41300 31444
rect 40908 30380 40964 30436
rect 40348 30268 40404 30324
rect 41244 30322 41300 30324
rect 41244 30270 41246 30322
rect 41246 30270 41298 30322
rect 41298 30270 41300 30322
rect 41244 30268 41300 30270
rect 42140 32562 42196 32564
rect 42140 32510 42142 32562
rect 42142 32510 42194 32562
rect 42194 32510 42196 32562
rect 42140 32508 42196 32510
rect 41468 30098 41524 30100
rect 41468 30046 41470 30098
rect 41470 30046 41522 30098
rect 41522 30046 41524 30098
rect 41468 30044 41524 30046
rect 41692 31052 41748 31108
rect 45948 38444 46004 38500
rect 46060 38332 46116 38388
rect 46060 37772 46116 37828
rect 45836 36652 45892 36708
rect 45836 36258 45892 36260
rect 45836 36206 45838 36258
rect 45838 36206 45890 36258
rect 45890 36206 45892 36258
rect 45836 36204 45892 36206
rect 45612 33516 45668 33572
rect 45836 34636 45892 34692
rect 46508 43260 46564 43316
rect 46732 42642 46788 42644
rect 46732 42590 46734 42642
rect 46734 42590 46786 42642
rect 46786 42590 46788 42642
rect 46732 42588 46788 42590
rect 46620 41858 46676 41860
rect 46620 41806 46622 41858
rect 46622 41806 46674 41858
rect 46674 41806 46676 41858
rect 46620 41804 46676 41806
rect 47180 48242 47236 48244
rect 47180 48190 47182 48242
rect 47182 48190 47234 48242
rect 47234 48190 47236 48242
rect 47180 48188 47236 48190
rect 48076 48972 48132 49028
rect 48188 47964 48244 48020
rect 48188 47628 48244 47684
rect 47740 47516 47796 47572
rect 47068 47292 47124 47348
rect 48076 47458 48132 47460
rect 48076 47406 48078 47458
rect 48078 47406 48130 47458
rect 48130 47406 48132 47458
rect 48076 47404 48132 47406
rect 47964 47292 48020 47348
rect 46956 41970 47012 41972
rect 46956 41918 46958 41970
rect 46958 41918 47010 41970
rect 47010 41918 47012 41970
rect 46956 41916 47012 41918
rect 47180 46172 47236 46228
rect 47516 45276 47572 45332
rect 47292 43596 47348 43652
rect 47404 43314 47460 43316
rect 47404 43262 47406 43314
rect 47406 43262 47458 43314
rect 47458 43262 47460 43314
rect 47404 43260 47460 43262
rect 47292 42642 47348 42644
rect 47292 42590 47294 42642
rect 47294 42590 47346 42642
rect 47346 42590 47348 42642
rect 47292 42588 47348 42590
rect 47628 43538 47684 43540
rect 47628 43486 47630 43538
rect 47630 43486 47682 43538
rect 47682 43486 47684 43538
rect 47628 43484 47684 43486
rect 47068 41580 47124 41636
rect 46284 37436 46340 37492
rect 46396 37378 46452 37380
rect 46396 37326 46398 37378
rect 46398 37326 46450 37378
rect 46450 37326 46452 37378
rect 46396 37324 46452 37326
rect 46396 36988 46452 37044
rect 47628 42588 47684 42644
rect 47292 42194 47348 42196
rect 47292 42142 47294 42194
rect 47294 42142 47346 42194
rect 47346 42142 47348 42194
rect 47292 42140 47348 42142
rect 47852 42194 47908 42196
rect 47852 42142 47854 42194
rect 47854 42142 47906 42194
rect 47906 42142 47908 42194
rect 47852 42140 47908 42142
rect 47068 40796 47124 40852
rect 46732 39676 46788 39732
rect 46844 39004 46900 39060
rect 46620 37212 46676 37268
rect 46508 36876 46564 36932
rect 46284 36204 46340 36260
rect 47852 41916 47908 41972
rect 47180 36988 47236 37044
rect 48748 53058 48804 53060
rect 48748 53006 48750 53058
rect 48750 53006 48802 53058
rect 48802 53006 48804 53058
rect 48748 53004 48804 53006
rect 48524 52892 48580 52948
rect 48972 52946 49028 52948
rect 48972 52894 48974 52946
rect 48974 52894 49026 52946
rect 49026 52894 49028 52946
rect 48972 52892 49028 52894
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 49756 52892 49812 52948
rect 48860 52834 48916 52836
rect 48860 52782 48862 52834
rect 48862 52782 48914 52834
rect 48914 52782 48916 52834
rect 48860 52780 48916 52782
rect 48748 52444 48804 52500
rect 49308 52162 49364 52164
rect 49308 52110 49310 52162
rect 49310 52110 49362 52162
rect 49362 52110 49364 52162
rect 49308 52108 49364 52110
rect 48748 51602 48804 51604
rect 48748 51550 48750 51602
rect 48750 51550 48802 51602
rect 48802 51550 48804 51602
rect 48748 51548 48804 51550
rect 48860 51436 48916 51492
rect 48412 49644 48468 49700
rect 49084 50540 49140 50596
rect 49532 50482 49588 50484
rect 49532 50430 49534 50482
rect 49534 50430 49586 50482
rect 49586 50430 49588 50482
rect 49532 50428 49588 50430
rect 49084 50370 49140 50372
rect 49084 50318 49086 50370
rect 49086 50318 49138 50370
rect 49138 50318 49140 50370
rect 49084 50316 49140 50318
rect 49308 50092 49364 50148
rect 49420 50316 49476 50372
rect 48636 49644 48692 49700
rect 48748 49196 48804 49252
rect 49084 49586 49140 49588
rect 49084 49534 49086 49586
rect 49086 49534 49138 49586
rect 49138 49534 49140 49586
rect 49084 49532 49140 49534
rect 49084 48636 49140 48692
rect 48860 48466 48916 48468
rect 48860 48414 48862 48466
rect 48862 48414 48914 48466
rect 48914 48414 48916 48466
rect 48860 48412 48916 48414
rect 48636 48300 48692 48356
rect 48972 48300 49028 48356
rect 48748 48076 48804 48132
rect 48748 47516 48804 47572
rect 48972 47458 49028 47460
rect 48972 47406 48974 47458
rect 48974 47406 49026 47458
rect 49026 47406 49028 47458
rect 48972 47404 49028 47406
rect 48860 47234 48916 47236
rect 48860 47182 48862 47234
rect 48862 47182 48914 47234
rect 48914 47182 48916 47234
rect 48860 47180 48916 47182
rect 48636 46002 48692 46004
rect 48636 45950 48638 46002
rect 48638 45950 48690 46002
rect 48690 45950 48692 46002
rect 48636 45948 48692 45950
rect 48524 45164 48580 45220
rect 48748 45388 48804 45444
rect 48188 43538 48244 43540
rect 48188 43486 48190 43538
rect 48190 43486 48242 43538
rect 48242 43486 48244 43538
rect 48188 43484 48244 43486
rect 48300 41804 48356 41860
rect 48300 41468 48356 41524
rect 48524 41804 48580 41860
rect 47964 41244 48020 41300
rect 48524 41132 48580 41188
rect 48076 40348 48132 40404
rect 48412 39394 48468 39396
rect 48412 39342 48414 39394
rect 48414 39342 48466 39394
rect 48466 39342 48468 39394
rect 48412 39340 48468 39342
rect 47404 35980 47460 36036
rect 47516 35868 47572 35924
rect 47628 37100 47684 37156
rect 46732 35420 46788 35476
rect 47068 34914 47124 34916
rect 47068 34862 47070 34914
rect 47070 34862 47122 34914
rect 47122 34862 47124 34914
rect 47068 34860 47124 34862
rect 46284 34636 46340 34692
rect 46172 32956 46228 33012
rect 45388 32562 45444 32564
rect 45388 32510 45390 32562
rect 45390 32510 45442 32562
rect 45442 32510 45444 32562
rect 45388 32508 45444 32510
rect 46732 32562 46788 32564
rect 46732 32510 46734 32562
rect 46734 32510 46786 32562
rect 46786 32510 46788 32562
rect 46732 32508 46788 32510
rect 48412 38556 48468 38612
rect 48412 36988 48468 37044
rect 48188 36876 48244 36932
rect 48188 36540 48244 36596
rect 47852 36204 47908 36260
rect 47740 35922 47796 35924
rect 47740 35870 47742 35922
rect 47742 35870 47794 35922
rect 47794 35870 47796 35922
rect 47740 35868 47796 35870
rect 48300 36258 48356 36260
rect 48300 36206 48302 36258
rect 48302 36206 48354 36258
rect 48354 36206 48356 36258
rect 48300 36204 48356 36206
rect 48748 42028 48804 42084
rect 48972 44210 49028 44212
rect 48972 44158 48974 44210
rect 48974 44158 49026 44210
rect 49026 44158 49028 44210
rect 48972 44156 49028 44158
rect 49308 49810 49364 49812
rect 49308 49758 49310 49810
rect 49310 49758 49362 49810
rect 49362 49758 49364 49810
rect 49308 49756 49364 49758
rect 49308 48466 49364 48468
rect 49308 48414 49310 48466
rect 49310 48414 49362 48466
rect 49362 48414 49364 48466
rect 49308 48412 49364 48414
rect 49868 52050 49924 52052
rect 49868 51998 49870 52050
rect 49870 51998 49922 52050
rect 49922 51998 49924 52050
rect 49868 51996 49924 51998
rect 49868 50482 49924 50484
rect 49868 50430 49870 50482
rect 49870 50430 49922 50482
rect 49922 50430 49924 50482
rect 49868 50428 49924 50430
rect 50092 50428 50148 50484
rect 49980 50370 50036 50372
rect 49980 50318 49982 50370
rect 49982 50318 50034 50370
rect 50034 50318 50036 50370
rect 49980 50316 50036 50318
rect 50764 52780 50820 52836
rect 50876 52332 50932 52388
rect 51548 52444 51604 52500
rect 51436 52050 51492 52052
rect 51436 51998 51438 52050
rect 51438 51998 51490 52050
rect 51490 51998 51492 52050
rect 51436 51996 51492 51998
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 51884 53452 51940 53508
rect 53004 52834 53060 52836
rect 53004 52782 53006 52834
rect 53006 52782 53058 52834
rect 53058 52782 53060 52834
rect 53004 52780 53060 52782
rect 51884 52220 51940 52276
rect 52780 52274 52836 52276
rect 52780 52222 52782 52274
rect 52782 52222 52834 52274
rect 52834 52222 52836 52274
rect 52780 52220 52836 52222
rect 51996 51996 52052 52052
rect 51660 51490 51716 51492
rect 51660 51438 51662 51490
rect 51662 51438 51714 51490
rect 51714 51438 51716 51490
rect 51660 51436 51716 51438
rect 50764 51378 50820 51380
rect 50764 51326 50766 51378
rect 50766 51326 50818 51378
rect 50818 51326 50820 51378
rect 50764 51324 50820 51326
rect 51884 51378 51940 51380
rect 51884 51326 51886 51378
rect 51886 51326 51938 51378
rect 51938 51326 51940 51378
rect 51884 51324 51940 51326
rect 50876 51266 50932 51268
rect 50876 51214 50878 51266
rect 50878 51214 50930 51266
rect 50930 51214 50932 51266
rect 50876 51212 50932 51214
rect 50876 50428 50932 50484
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50204 49922 50260 49924
rect 50204 49870 50206 49922
rect 50206 49870 50258 49922
rect 50258 49870 50260 49922
rect 50204 49868 50260 49870
rect 51772 50482 51828 50484
rect 51772 50430 51774 50482
rect 51774 50430 51826 50482
rect 51826 50430 51828 50482
rect 51772 50428 51828 50430
rect 52780 51212 52836 51268
rect 52780 50594 52836 50596
rect 52780 50542 52782 50594
rect 52782 50542 52834 50594
rect 52834 50542 52836 50594
rect 52780 50540 52836 50542
rect 53340 51266 53396 51268
rect 53340 51214 53342 51266
rect 53342 51214 53394 51266
rect 53394 51214 53396 51266
rect 53340 51212 53396 51214
rect 53004 51100 53060 51156
rect 51100 49868 51156 49924
rect 50764 49756 50820 49812
rect 50092 49698 50148 49700
rect 50092 49646 50094 49698
rect 50094 49646 50146 49698
rect 50146 49646 50148 49698
rect 50092 49644 50148 49646
rect 50204 49532 50260 49588
rect 49868 48748 49924 48804
rect 50092 49196 50148 49252
rect 49980 48018 50036 48020
rect 49980 47966 49982 48018
rect 49982 47966 50034 48018
rect 50034 47966 50036 48018
rect 49980 47964 50036 47966
rect 50092 47852 50148 47908
rect 50764 49196 50820 49252
rect 50540 49026 50596 49028
rect 50540 48974 50542 49026
rect 50542 48974 50594 49026
rect 50594 48974 50596 49026
rect 50540 48972 50596 48974
rect 50428 48860 50484 48916
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50428 47852 50484 47908
rect 50652 47682 50708 47684
rect 50652 47630 50654 47682
rect 50654 47630 50706 47682
rect 50706 47630 50708 47682
rect 50652 47628 50708 47630
rect 49196 44492 49252 44548
rect 49756 47458 49812 47460
rect 49756 47406 49758 47458
rect 49758 47406 49810 47458
rect 49810 47406 49812 47458
rect 49756 47404 49812 47406
rect 49308 47292 49364 47348
rect 49532 47292 49588 47348
rect 49420 46396 49476 46452
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 49196 44156 49252 44212
rect 49084 43484 49140 43540
rect 49196 43596 49252 43652
rect 49420 43538 49476 43540
rect 49420 43486 49422 43538
rect 49422 43486 49474 43538
rect 49474 43486 49476 43538
rect 49420 43484 49476 43486
rect 50204 46674 50260 46676
rect 50204 46622 50206 46674
rect 50206 46622 50258 46674
rect 50258 46622 50260 46674
rect 50204 46620 50260 46622
rect 49868 46562 49924 46564
rect 49868 46510 49870 46562
rect 49870 46510 49922 46562
rect 49922 46510 49924 46562
rect 49868 46508 49924 46510
rect 50316 46508 50372 46564
rect 50092 46396 50148 46452
rect 50764 46562 50820 46564
rect 50764 46510 50766 46562
rect 50766 46510 50818 46562
rect 50818 46510 50820 46562
rect 50764 46508 50820 46510
rect 50540 46284 50596 46340
rect 50540 45836 50596 45892
rect 51324 48242 51380 48244
rect 51324 48190 51326 48242
rect 51326 48190 51378 48242
rect 51378 48190 51380 48242
rect 51324 48188 51380 48190
rect 51884 50316 51940 50372
rect 51548 49084 51604 49140
rect 51660 49308 51716 49364
rect 51996 49138 52052 49140
rect 51996 49086 51998 49138
rect 51998 49086 52050 49138
rect 52050 49086 52052 49138
rect 51996 49084 52052 49086
rect 52108 49026 52164 49028
rect 52108 48974 52110 49026
rect 52110 48974 52162 49026
rect 52162 48974 52164 49026
rect 52108 48972 52164 48974
rect 51548 48300 51604 48356
rect 53900 51100 53956 51156
rect 54460 51100 54516 51156
rect 54460 50540 54516 50596
rect 53340 50370 53396 50372
rect 53340 50318 53342 50370
rect 53342 50318 53394 50370
rect 53394 50318 53396 50370
rect 53340 50316 53396 50318
rect 53116 49810 53172 49812
rect 53116 49758 53118 49810
rect 53118 49758 53170 49810
rect 53170 49758 53172 49810
rect 53116 49756 53172 49758
rect 53788 49810 53844 49812
rect 53788 49758 53790 49810
rect 53790 49758 53842 49810
rect 53842 49758 53844 49810
rect 53788 49756 53844 49758
rect 52780 49698 52836 49700
rect 52780 49646 52782 49698
rect 52782 49646 52834 49698
rect 52834 49646 52836 49698
rect 52780 49644 52836 49646
rect 52668 49308 52724 49364
rect 52780 48972 52836 49028
rect 52332 48860 52388 48916
rect 52668 48188 52724 48244
rect 51996 47570 52052 47572
rect 51996 47518 51998 47570
rect 51998 47518 52050 47570
rect 52050 47518 52052 47570
rect 51996 47516 52052 47518
rect 52668 47516 52724 47572
rect 51100 47068 51156 47124
rect 50764 46284 50820 46340
rect 50876 45890 50932 45892
rect 50876 45838 50878 45890
rect 50878 45838 50930 45890
rect 50930 45838 50932 45890
rect 50876 45836 50932 45838
rect 51324 46284 51380 46340
rect 51436 47180 51492 47236
rect 49756 45388 49812 45444
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50316 45052 50372 45108
rect 50204 44156 50260 44212
rect 50092 44098 50148 44100
rect 50092 44046 50094 44098
rect 50094 44046 50146 44098
rect 50146 44046 50148 44098
rect 50092 44044 50148 44046
rect 49644 43538 49700 43540
rect 49644 43486 49646 43538
rect 49646 43486 49698 43538
rect 49698 43486 49700 43538
rect 49644 43484 49700 43486
rect 48860 41692 48916 41748
rect 49644 42140 49700 42196
rect 49868 43260 49924 43316
rect 49532 42082 49588 42084
rect 49532 42030 49534 42082
rect 49534 42030 49586 42082
rect 49586 42030 49588 42082
rect 49532 42028 49588 42030
rect 49084 41746 49140 41748
rect 49084 41694 49086 41746
rect 49086 41694 49138 41746
rect 49138 41694 49140 41746
rect 49084 41692 49140 41694
rect 49196 41580 49252 41636
rect 48748 40908 48804 40964
rect 48972 41244 49028 41300
rect 49532 41244 49588 41300
rect 49756 40962 49812 40964
rect 49756 40910 49758 40962
rect 49758 40910 49810 40962
rect 49810 40910 49812 40962
rect 49756 40908 49812 40910
rect 49084 40514 49140 40516
rect 49084 40462 49086 40514
rect 49086 40462 49138 40514
rect 49138 40462 49140 40514
rect 49084 40460 49140 40462
rect 49532 40348 49588 40404
rect 48748 39340 48804 39396
rect 48860 39564 48916 39620
rect 48860 38556 48916 38612
rect 49084 39340 49140 39396
rect 51100 45106 51156 45108
rect 51100 45054 51102 45106
rect 51102 45054 51154 45106
rect 51154 45054 51156 45106
rect 51100 45052 51156 45054
rect 50876 44210 50932 44212
rect 50876 44158 50878 44210
rect 50878 44158 50930 44210
rect 50930 44158 50932 44210
rect 50876 44156 50932 44158
rect 51100 44210 51156 44212
rect 51100 44158 51102 44210
rect 51102 44158 51154 44210
rect 51154 44158 51156 44210
rect 51100 44156 51156 44158
rect 50764 44044 50820 44100
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50316 43708 50372 43764
rect 50092 41186 50148 41188
rect 50092 41134 50094 41186
rect 50094 41134 50146 41186
rect 50146 41134 50148 41186
rect 50092 41132 50148 41134
rect 50204 41074 50260 41076
rect 50204 41022 50206 41074
rect 50206 41022 50258 41074
rect 50258 41022 50260 41074
rect 50204 41020 50260 41022
rect 49980 40908 50036 40964
rect 50876 43314 50932 43316
rect 50876 43262 50878 43314
rect 50878 43262 50930 43314
rect 50930 43262 50932 43314
rect 50876 43260 50932 43262
rect 50876 42924 50932 42980
rect 50988 42754 51044 42756
rect 50988 42702 50990 42754
rect 50990 42702 51042 42754
rect 51042 42702 51044 42754
rect 50988 42700 51044 42702
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50540 42028 50596 42084
rect 51100 41858 51156 41860
rect 51100 41806 51102 41858
rect 51102 41806 51154 41858
rect 51154 41806 51156 41858
rect 51100 41804 51156 41806
rect 50652 41692 50708 41748
rect 50540 41580 50596 41636
rect 51436 43708 51492 43764
rect 51324 43426 51380 43428
rect 51324 43374 51326 43426
rect 51326 43374 51378 43426
rect 51378 43374 51380 43426
rect 51324 43372 51380 43374
rect 51324 43036 51380 43092
rect 51436 43260 51492 43316
rect 51884 47404 51940 47460
rect 51884 47068 51940 47124
rect 52108 47068 52164 47124
rect 51660 46786 51716 46788
rect 51660 46734 51662 46786
rect 51662 46734 51714 46786
rect 51714 46734 51716 46786
rect 51660 46732 51716 46734
rect 52220 46674 52276 46676
rect 52220 46622 52222 46674
rect 52222 46622 52274 46674
rect 52274 46622 52276 46674
rect 52220 46620 52276 46622
rect 52780 47292 52836 47348
rect 52556 46956 52612 47012
rect 52332 45724 52388 45780
rect 52444 46620 52500 46676
rect 51548 43148 51604 43204
rect 51772 42924 51828 42980
rect 52444 45276 52500 45332
rect 53452 49196 53508 49252
rect 53004 48972 53060 49028
rect 53340 48914 53396 48916
rect 53340 48862 53342 48914
rect 53342 48862 53394 48914
rect 53394 48862 53396 48914
rect 53340 48860 53396 48862
rect 53564 48242 53620 48244
rect 53564 48190 53566 48242
rect 53566 48190 53618 48242
rect 53618 48190 53620 48242
rect 53564 48188 53620 48190
rect 53004 47458 53060 47460
rect 53004 47406 53006 47458
rect 53006 47406 53058 47458
rect 53058 47406 53060 47458
rect 53004 47404 53060 47406
rect 53788 47516 53844 47572
rect 53116 47292 53172 47348
rect 53788 47346 53844 47348
rect 53788 47294 53790 47346
rect 53790 47294 53842 47346
rect 53842 47294 53844 47346
rect 53788 47292 53844 47294
rect 53452 47234 53508 47236
rect 53452 47182 53454 47234
rect 53454 47182 53506 47234
rect 53506 47182 53508 47234
rect 53452 47180 53508 47182
rect 53452 46956 53508 47012
rect 54124 48076 54180 48132
rect 54012 47964 54068 48020
rect 53900 46956 53956 47012
rect 53228 46732 53284 46788
rect 52668 45836 52724 45892
rect 53452 46674 53508 46676
rect 53452 46622 53454 46674
rect 53454 46622 53506 46674
rect 53506 46622 53508 46674
rect 53452 46620 53508 46622
rect 53228 46396 53284 46452
rect 53564 46508 53620 46564
rect 52108 43148 52164 43204
rect 51324 42476 51380 42532
rect 51212 41580 51268 41636
rect 50988 41186 51044 41188
rect 50988 41134 50990 41186
rect 50990 41134 51042 41186
rect 51042 41134 51044 41186
rect 50988 41132 51044 41134
rect 50540 41020 50596 41076
rect 50876 40908 50932 40964
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 51772 41916 51828 41972
rect 51100 40684 51156 40740
rect 51548 41298 51604 41300
rect 51548 41246 51550 41298
rect 51550 41246 51602 41298
rect 51602 41246 51604 41298
rect 51548 41244 51604 41246
rect 50204 40460 50260 40516
rect 50428 39788 50484 39844
rect 50540 39564 50596 39620
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 51660 41132 51716 41188
rect 51324 41020 51380 41076
rect 50428 38834 50484 38836
rect 50428 38782 50430 38834
rect 50430 38782 50482 38834
rect 50482 38782 50484 38834
rect 50428 38780 50484 38782
rect 50652 38668 50708 38724
rect 48860 36876 48916 36932
rect 48972 37996 49028 38052
rect 48636 36652 48692 36708
rect 47964 35698 48020 35700
rect 47964 35646 47966 35698
rect 47966 35646 48018 35698
rect 48018 35646 48020 35698
rect 47964 35644 48020 35646
rect 47964 35196 48020 35252
rect 47740 34860 47796 34916
rect 47404 33516 47460 33572
rect 47964 33516 48020 33572
rect 46508 32396 46564 32452
rect 45388 31948 45444 32004
rect 43596 31836 43652 31892
rect 45500 31836 45556 31892
rect 47516 32786 47572 32788
rect 47516 32734 47518 32786
rect 47518 32734 47570 32786
rect 47570 32734 47572 32786
rect 47516 32732 47572 32734
rect 47180 32284 47236 32340
rect 48076 34300 48132 34356
rect 47852 33122 47908 33124
rect 47852 33070 47854 33122
rect 47854 33070 47906 33122
rect 47906 33070 47908 33122
rect 47852 33068 47908 33070
rect 48412 34076 48468 34132
rect 48860 32956 48916 33012
rect 49868 38050 49924 38052
rect 49868 37998 49870 38050
rect 49870 37998 49922 38050
rect 49922 37998 49924 38050
rect 49868 37996 49924 37998
rect 49644 36316 49700 36372
rect 50540 37938 50596 37940
rect 50540 37886 50542 37938
rect 50542 37886 50594 37938
rect 50594 37886 50596 37938
rect 50540 37884 50596 37886
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50204 37436 50260 37492
rect 51884 40908 51940 40964
rect 51660 40684 51716 40740
rect 51996 40236 52052 40292
rect 53900 46562 53956 46564
rect 53900 46510 53902 46562
rect 53902 46510 53954 46562
rect 53954 46510 53956 46562
rect 53900 46508 53956 46510
rect 53564 45106 53620 45108
rect 53564 45054 53566 45106
rect 53566 45054 53618 45106
rect 53618 45054 53620 45106
rect 53564 45052 53620 45054
rect 54684 49644 54740 49700
rect 54572 48914 54628 48916
rect 54572 48862 54574 48914
rect 54574 48862 54626 48914
rect 54626 48862 54628 48914
rect 54572 48860 54628 48862
rect 54572 47964 54628 48020
rect 54460 46732 54516 46788
rect 54796 46956 54852 47012
rect 53788 45164 53844 45220
rect 53676 44940 53732 44996
rect 53116 44828 53172 44884
rect 53004 44156 53060 44212
rect 52444 42476 52500 42532
rect 53116 43596 53172 43652
rect 53564 44268 53620 44324
rect 53900 44322 53956 44324
rect 53900 44270 53902 44322
rect 53902 44270 53954 44322
rect 53954 44270 53956 44322
rect 53900 44268 53956 44270
rect 53900 43314 53956 43316
rect 53900 43262 53902 43314
rect 53902 43262 53954 43314
rect 53954 43262 53956 43314
rect 53900 43260 53956 43262
rect 53676 43148 53732 43204
rect 53564 43036 53620 43092
rect 53004 42754 53060 42756
rect 53004 42702 53006 42754
rect 53006 42702 53058 42754
rect 53058 42702 53060 42754
rect 53004 42700 53060 42702
rect 52892 42588 52948 42644
rect 53228 42642 53284 42644
rect 53228 42590 53230 42642
rect 53230 42590 53282 42642
rect 53282 42590 53284 42642
rect 53228 42588 53284 42590
rect 52444 41970 52500 41972
rect 52444 41918 52446 41970
rect 52446 41918 52498 41970
rect 52498 41918 52500 41970
rect 52444 41916 52500 41918
rect 52220 40124 52276 40180
rect 52668 41746 52724 41748
rect 52668 41694 52670 41746
rect 52670 41694 52722 41746
rect 52722 41694 52724 41746
rect 52668 41692 52724 41694
rect 52556 41468 52612 41524
rect 51996 39452 52052 39508
rect 52220 39452 52276 39508
rect 51436 39340 51492 39396
rect 51436 38668 51492 38724
rect 50988 37324 51044 37380
rect 50876 36540 50932 36596
rect 50316 36258 50372 36260
rect 50316 36206 50318 36258
rect 50318 36206 50370 36258
rect 50370 36206 50372 36258
rect 50316 36204 50372 36206
rect 49196 35698 49252 35700
rect 49196 35646 49198 35698
rect 49198 35646 49250 35698
rect 49250 35646 49252 35698
rect 49196 35644 49252 35646
rect 49980 35644 50036 35700
rect 49532 35586 49588 35588
rect 49532 35534 49534 35586
rect 49534 35534 49586 35586
rect 49586 35534 49588 35586
rect 49532 35532 49588 35534
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50764 35532 50820 35588
rect 50988 35420 51044 35476
rect 50428 34914 50484 34916
rect 50428 34862 50430 34914
rect 50430 34862 50482 34914
rect 50482 34862 50484 34914
rect 50428 34860 50484 34862
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50204 34354 50260 34356
rect 50204 34302 50206 34354
rect 50206 34302 50258 34354
rect 50258 34302 50260 34354
rect 50204 34300 50260 34302
rect 50764 34242 50820 34244
rect 50764 34190 50766 34242
rect 50766 34190 50818 34242
rect 50818 34190 50820 34242
rect 50764 34188 50820 34190
rect 49084 33852 49140 33908
rect 48748 32732 48804 32788
rect 48860 32450 48916 32452
rect 48860 32398 48862 32450
rect 48862 32398 48914 32450
rect 48914 32398 48916 32450
rect 48860 32396 48916 32398
rect 47404 32172 47460 32228
rect 48636 32172 48692 32228
rect 48188 31836 48244 31892
rect 44268 31500 44324 31556
rect 42140 31218 42196 31220
rect 42140 31166 42142 31218
rect 42142 31166 42194 31218
rect 42194 31166 42196 31218
rect 42140 31164 42196 31166
rect 40908 29986 40964 29988
rect 40908 29934 40910 29986
rect 40910 29934 40962 29986
rect 40962 29934 40964 29986
rect 40908 29932 40964 29934
rect 41356 29986 41412 29988
rect 41356 29934 41358 29986
rect 41358 29934 41410 29986
rect 41410 29934 41412 29986
rect 41356 29932 41412 29934
rect 40236 29426 40292 29428
rect 40236 29374 40238 29426
rect 40238 29374 40290 29426
rect 40290 29374 40292 29426
rect 40236 29372 40292 29374
rect 40124 29148 40180 29204
rect 41244 28812 41300 28868
rect 40124 28642 40180 28644
rect 40124 28590 40126 28642
rect 40126 28590 40178 28642
rect 40178 28590 40180 28642
rect 40124 28588 40180 28590
rect 39676 28364 39732 28420
rect 38556 28028 38612 28084
rect 37772 26962 37828 26964
rect 37772 26910 37774 26962
rect 37774 26910 37826 26962
rect 37826 26910 37828 26962
rect 37772 26908 37828 26910
rect 38332 27916 38388 27972
rect 39340 27692 39396 27748
rect 37436 26684 37492 26740
rect 39788 28028 39844 28084
rect 40124 27970 40180 27972
rect 40124 27918 40126 27970
rect 40126 27918 40178 27970
rect 40178 27918 40180 27970
rect 40124 27916 40180 27918
rect 39788 27634 39844 27636
rect 39788 27582 39790 27634
rect 39790 27582 39842 27634
rect 39842 27582 39844 27634
rect 39788 27580 39844 27582
rect 42364 31106 42420 31108
rect 42364 31054 42366 31106
rect 42366 31054 42418 31106
rect 42418 31054 42420 31106
rect 42364 31052 42420 31054
rect 43372 29932 43428 29988
rect 42476 29372 42532 29428
rect 44940 31554 44996 31556
rect 44940 31502 44942 31554
rect 44942 31502 44994 31554
rect 44994 31502 44996 31554
rect 44940 31500 44996 31502
rect 45388 31554 45444 31556
rect 45388 31502 45390 31554
rect 45390 31502 45442 31554
rect 45442 31502 45444 31554
rect 45388 31500 45444 31502
rect 45836 31500 45892 31556
rect 48972 31948 49028 32004
rect 49644 33068 49700 33124
rect 50092 34130 50148 34132
rect 50092 34078 50094 34130
rect 50094 34078 50146 34130
rect 50146 34078 50148 34130
rect 50092 34076 50148 34078
rect 50316 33852 50372 33908
rect 52220 38668 52276 38724
rect 51660 37548 51716 37604
rect 51772 37772 51828 37828
rect 51436 36482 51492 36484
rect 51436 36430 51438 36482
rect 51438 36430 51490 36482
rect 51490 36430 51492 36482
rect 51436 36428 51492 36430
rect 51772 35756 51828 35812
rect 51660 35586 51716 35588
rect 51660 35534 51662 35586
rect 51662 35534 51714 35586
rect 51714 35534 51716 35586
rect 51660 35532 51716 35534
rect 51436 34972 51492 35028
rect 51884 36652 51940 36708
rect 51100 34300 51156 34356
rect 50316 33292 50372 33348
rect 49196 31836 49252 31892
rect 49420 32284 49476 32340
rect 50652 33346 50708 33348
rect 50652 33294 50654 33346
rect 50654 33294 50706 33346
rect 50706 33294 50708 33346
rect 50652 33292 50708 33294
rect 51324 33906 51380 33908
rect 51324 33854 51326 33906
rect 51326 33854 51378 33906
rect 51378 33854 51380 33906
rect 51324 33852 51380 33854
rect 50540 33068 50596 33124
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 51436 33068 51492 33124
rect 51548 33852 51604 33908
rect 49980 32172 50036 32228
rect 49980 31778 50036 31780
rect 49980 31726 49982 31778
rect 49982 31726 50034 31778
rect 50034 31726 50036 31778
rect 49980 31724 50036 31726
rect 49644 31612 49700 31668
rect 50540 31500 50596 31556
rect 51660 32732 51716 32788
rect 52444 38610 52500 38612
rect 52444 38558 52446 38610
rect 52446 38558 52498 38610
rect 52498 38558 52500 38610
rect 52444 38556 52500 38558
rect 52332 37548 52388 37604
rect 52220 37378 52276 37380
rect 52220 37326 52222 37378
rect 52222 37326 52274 37378
rect 52274 37326 52276 37378
rect 52220 37324 52276 37326
rect 52220 36876 52276 36932
rect 53564 41580 53620 41636
rect 54124 46284 54180 46340
rect 54460 46172 54516 46228
rect 54908 46284 54964 46340
rect 54908 45948 54964 46004
rect 54460 45724 54516 45780
rect 55244 49810 55300 49812
rect 55244 49758 55246 49810
rect 55246 49758 55298 49810
rect 55298 49758 55300 49810
rect 55244 49756 55300 49758
rect 56140 50428 56196 50484
rect 55468 47068 55524 47124
rect 55356 46674 55412 46676
rect 55356 46622 55358 46674
rect 55358 46622 55410 46674
rect 55410 46622 55412 46674
rect 55356 46620 55412 46622
rect 55692 45778 55748 45780
rect 55692 45726 55694 45778
rect 55694 45726 55746 45778
rect 55746 45726 55748 45778
rect 55692 45724 55748 45726
rect 54124 45106 54180 45108
rect 54124 45054 54126 45106
rect 54126 45054 54178 45106
rect 54178 45054 54180 45106
rect 54124 45052 54180 45054
rect 54348 44882 54404 44884
rect 54348 44830 54350 44882
rect 54350 44830 54402 44882
rect 54402 44830 54404 44882
rect 54348 44828 54404 44830
rect 54348 43596 54404 43652
rect 55692 45500 55748 45556
rect 54684 45052 54740 45108
rect 55580 45218 55636 45220
rect 55580 45166 55582 45218
rect 55582 45166 55634 45218
rect 55634 45166 55636 45218
rect 55580 45164 55636 45166
rect 55132 45052 55188 45108
rect 55020 44994 55076 44996
rect 55020 44942 55022 44994
rect 55022 44942 55074 44994
rect 55074 44942 55076 44994
rect 55020 44940 55076 44942
rect 55020 44210 55076 44212
rect 55020 44158 55022 44210
rect 55022 44158 55074 44210
rect 55074 44158 55076 44210
rect 55020 44156 55076 44158
rect 54908 43372 54964 43428
rect 55356 44044 55412 44100
rect 54460 43148 54516 43204
rect 52668 40348 52724 40404
rect 55804 44156 55860 44212
rect 55468 43538 55524 43540
rect 55468 43486 55470 43538
rect 55470 43486 55522 43538
rect 55522 43486 55524 43538
rect 55468 43484 55524 43486
rect 56028 43650 56084 43652
rect 56028 43598 56030 43650
rect 56030 43598 56082 43650
rect 56082 43598 56084 43650
rect 56028 43596 56084 43598
rect 55692 43260 55748 43316
rect 55356 42700 55412 42756
rect 55580 42924 55636 42980
rect 53900 41692 53956 41748
rect 52892 40236 52948 40292
rect 53116 39564 53172 39620
rect 53004 39506 53060 39508
rect 53004 39454 53006 39506
rect 53006 39454 53058 39506
rect 53058 39454 53060 39506
rect 53004 39452 53060 39454
rect 52668 39394 52724 39396
rect 52668 39342 52670 39394
rect 52670 39342 52722 39394
rect 52722 39342 52724 39394
rect 52668 39340 52724 39342
rect 53228 39340 53284 39396
rect 52892 38834 52948 38836
rect 52892 38782 52894 38834
rect 52894 38782 52946 38834
rect 52946 38782 52948 38834
rect 52892 38780 52948 38782
rect 55580 42140 55636 42196
rect 54124 40460 54180 40516
rect 53788 40348 53844 40404
rect 53676 40290 53732 40292
rect 53676 40238 53678 40290
rect 53678 40238 53730 40290
rect 53730 40238 53732 40290
rect 53676 40236 53732 40238
rect 53900 40124 53956 40180
rect 54348 40402 54404 40404
rect 54348 40350 54350 40402
rect 54350 40350 54402 40402
rect 54402 40350 54404 40402
rect 54348 40348 54404 40350
rect 54124 39730 54180 39732
rect 54124 39678 54126 39730
rect 54126 39678 54178 39730
rect 54178 39678 54180 39730
rect 54124 39676 54180 39678
rect 54348 39506 54404 39508
rect 54348 39454 54350 39506
rect 54350 39454 54402 39506
rect 54402 39454 54404 39506
rect 54348 39452 54404 39454
rect 53788 39394 53844 39396
rect 53788 39342 53790 39394
rect 53790 39342 53842 39394
rect 53842 39342 53844 39394
rect 53788 39340 53844 39342
rect 54124 38722 54180 38724
rect 54124 38670 54126 38722
rect 54126 38670 54178 38722
rect 54178 38670 54180 38722
rect 54124 38668 54180 38670
rect 53116 38556 53172 38612
rect 53116 38050 53172 38052
rect 53116 37998 53118 38050
rect 53118 37998 53170 38050
rect 53170 37998 53172 38050
rect 53116 37996 53172 37998
rect 52892 37938 52948 37940
rect 52892 37886 52894 37938
rect 52894 37886 52946 37938
rect 52946 37886 52948 37938
rect 52892 37884 52948 37886
rect 52668 37436 52724 37492
rect 52892 37660 52948 37716
rect 52556 36652 52612 36708
rect 52668 36540 52724 36596
rect 51996 36316 52052 36372
rect 52444 35474 52500 35476
rect 52444 35422 52446 35474
rect 52446 35422 52498 35474
rect 52498 35422 52500 35474
rect 52444 35420 52500 35422
rect 52108 35084 52164 35140
rect 52108 34188 52164 34244
rect 52220 34860 52276 34916
rect 53340 38556 53396 38612
rect 53564 38050 53620 38052
rect 53564 37998 53566 38050
rect 53566 37998 53618 38050
rect 53618 37998 53620 38050
rect 53564 37996 53620 37998
rect 54908 41692 54964 41748
rect 55020 41244 55076 41300
rect 56028 42028 56084 42084
rect 55692 41858 55748 41860
rect 55692 41806 55694 41858
rect 55694 41806 55746 41858
rect 55746 41806 55748 41858
rect 55692 41804 55748 41806
rect 55692 41580 55748 41636
rect 55244 40460 55300 40516
rect 55692 40460 55748 40516
rect 54684 39676 54740 39732
rect 55020 38892 55076 38948
rect 53676 37884 53732 37940
rect 53228 37324 53284 37380
rect 53004 36482 53060 36484
rect 53004 36430 53006 36482
rect 53006 36430 53058 36482
rect 53058 36430 53060 36482
rect 53004 36428 53060 36430
rect 53452 37548 53508 37604
rect 54124 37378 54180 37380
rect 54124 37326 54126 37378
rect 54126 37326 54178 37378
rect 54178 37326 54180 37378
rect 54124 37324 54180 37326
rect 53788 37266 53844 37268
rect 53788 37214 53790 37266
rect 53790 37214 53842 37266
rect 53842 37214 53844 37266
rect 53788 37212 53844 37214
rect 54236 37266 54292 37268
rect 54236 37214 54238 37266
rect 54238 37214 54290 37266
rect 54290 37214 54292 37266
rect 54236 37212 54292 37214
rect 53452 36876 53508 36932
rect 54348 36876 54404 36932
rect 54236 36652 54292 36708
rect 54012 36258 54068 36260
rect 54012 36206 54014 36258
rect 54014 36206 54066 36258
rect 54066 36206 54068 36258
rect 54012 36204 54068 36206
rect 53788 35868 53844 35924
rect 53228 35810 53284 35812
rect 53228 35758 53230 35810
rect 53230 35758 53282 35810
rect 53282 35758 53284 35810
rect 53228 35756 53284 35758
rect 54348 36482 54404 36484
rect 54348 36430 54350 36482
rect 54350 36430 54402 36482
rect 54402 36430 54404 36482
rect 54348 36428 54404 36430
rect 54236 35756 54292 35812
rect 52892 35420 52948 35476
rect 53004 35532 53060 35588
rect 53004 35308 53060 35364
rect 53564 35698 53620 35700
rect 53564 35646 53566 35698
rect 53566 35646 53618 35698
rect 53618 35646 53620 35698
rect 53564 35644 53620 35646
rect 54124 35532 54180 35588
rect 53788 35474 53844 35476
rect 53788 35422 53790 35474
rect 53790 35422 53842 35474
rect 53842 35422 53844 35474
rect 53788 35420 53844 35422
rect 53676 35084 53732 35140
rect 53340 34972 53396 35028
rect 53228 34914 53284 34916
rect 53228 34862 53230 34914
rect 53230 34862 53282 34914
rect 53282 34862 53284 34914
rect 53228 34860 53284 34862
rect 55356 39452 55412 39508
rect 55356 39004 55412 39060
rect 54684 37938 54740 37940
rect 54684 37886 54686 37938
rect 54686 37886 54738 37938
rect 54738 37886 54740 37938
rect 54684 37884 54740 37886
rect 54908 37378 54964 37380
rect 54908 37326 54910 37378
rect 54910 37326 54962 37378
rect 54962 37326 54964 37378
rect 54908 37324 54964 37326
rect 54684 37266 54740 37268
rect 54684 37214 54686 37266
rect 54686 37214 54738 37266
rect 54738 37214 54740 37266
rect 54684 37212 54740 37214
rect 54572 37100 54628 37156
rect 54908 36988 54964 37044
rect 54908 35980 54964 36036
rect 54684 35868 54740 35924
rect 52220 34130 52276 34132
rect 52220 34078 52222 34130
rect 52222 34078 52274 34130
rect 52274 34078 52276 34130
rect 52220 34076 52276 34078
rect 52780 34130 52836 34132
rect 52780 34078 52782 34130
rect 52782 34078 52834 34130
rect 52834 34078 52836 34130
rect 52780 34076 52836 34078
rect 53228 34130 53284 34132
rect 53228 34078 53230 34130
rect 53230 34078 53282 34130
rect 53282 34078 53284 34130
rect 53228 34076 53284 34078
rect 54572 35756 54628 35812
rect 54012 34076 54068 34132
rect 51884 33404 51940 33460
rect 51660 32562 51716 32564
rect 51660 32510 51662 32562
rect 51662 32510 51714 32562
rect 51714 32510 51716 32562
rect 51660 32508 51716 32510
rect 52780 33458 52836 33460
rect 52780 33406 52782 33458
rect 52782 33406 52834 33458
rect 52834 33406 52836 33458
rect 52780 33404 52836 33406
rect 54796 35586 54852 35588
rect 54796 35534 54798 35586
rect 54798 35534 54850 35586
rect 54850 35534 54852 35586
rect 54796 35532 54852 35534
rect 54684 34860 54740 34916
rect 54684 33964 54740 34020
rect 55244 36876 55300 36932
rect 55804 39730 55860 39732
rect 55804 39678 55806 39730
rect 55806 39678 55858 39730
rect 55858 39678 55860 39730
rect 55804 39676 55860 39678
rect 55916 38946 55972 38948
rect 55916 38894 55918 38946
rect 55918 38894 55970 38946
rect 55970 38894 55972 38946
rect 55916 38892 55972 38894
rect 56476 49810 56532 49812
rect 56476 49758 56478 49810
rect 56478 49758 56530 49810
rect 56530 49758 56532 49810
rect 56476 49756 56532 49758
rect 57484 49138 57540 49140
rect 57484 49086 57486 49138
rect 57486 49086 57538 49138
rect 57538 49086 57540 49138
rect 57484 49084 57540 49086
rect 56588 48130 56644 48132
rect 56588 48078 56590 48130
rect 56590 48078 56642 48130
rect 56642 48078 56644 48130
rect 56588 48076 56644 48078
rect 57148 46172 57204 46228
rect 56588 45218 56644 45220
rect 56588 45166 56590 45218
rect 56590 45166 56642 45218
rect 56642 45166 56644 45218
rect 56588 45164 56644 45166
rect 57820 45500 57876 45556
rect 56364 44322 56420 44324
rect 56364 44270 56366 44322
rect 56366 44270 56418 44322
rect 56418 44270 56420 44322
rect 56364 44268 56420 44270
rect 56588 44210 56644 44212
rect 56588 44158 56590 44210
rect 56590 44158 56642 44210
rect 56642 44158 56644 44210
rect 56588 44156 56644 44158
rect 57148 44210 57204 44212
rect 57148 44158 57150 44210
rect 57150 44158 57202 44210
rect 57202 44158 57204 44210
rect 57148 44156 57204 44158
rect 57596 44044 57652 44100
rect 56252 43596 56308 43652
rect 57036 43650 57092 43652
rect 57036 43598 57038 43650
rect 57038 43598 57090 43650
rect 57090 43598 57092 43650
rect 57036 43596 57092 43598
rect 56588 43538 56644 43540
rect 56588 43486 56590 43538
rect 56590 43486 56642 43538
rect 56642 43486 56644 43538
rect 56588 43484 56644 43486
rect 56812 43372 56868 43428
rect 56700 42140 56756 42196
rect 56588 42028 56644 42084
rect 57036 42028 57092 42084
rect 56700 41074 56756 41076
rect 56700 41022 56702 41074
rect 56702 41022 56754 41074
rect 56754 41022 56756 41074
rect 56700 41020 56756 41022
rect 55468 37660 55524 37716
rect 55804 37660 55860 37716
rect 55692 37490 55748 37492
rect 55692 37438 55694 37490
rect 55694 37438 55746 37490
rect 55746 37438 55748 37490
rect 55692 37436 55748 37438
rect 55580 37378 55636 37380
rect 55580 37326 55582 37378
rect 55582 37326 55634 37378
rect 55634 37326 55636 37378
rect 55580 37324 55636 37326
rect 55804 37100 55860 37156
rect 55356 35756 55412 35812
rect 55580 35698 55636 35700
rect 55580 35646 55582 35698
rect 55582 35646 55634 35698
rect 55634 35646 55636 35698
rect 55580 35644 55636 35646
rect 55132 35420 55188 35476
rect 55468 35308 55524 35364
rect 55132 35026 55188 35028
rect 55132 34974 55134 35026
rect 55134 34974 55186 35026
rect 55186 34974 55188 35026
rect 55132 34972 55188 34974
rect 52108 32732 52164 32788
rect 54236 32562 54292 32564
rect 54236 32510 54238 32562
rect 54238 32510 54290 32562
rect 54290 32510 54292 32562
rect 54236 32508 54292 32510
rect 52108 32450 52164 32452
rect 52108 32398 52110 32450
rect 52110 32398 52162 32450
rect 52162 32398 52164 32450
rect 52108 32396 52164 32398
rect 52780 32396 52836 32452
rect 51324 31836 51380 31892
rect 51996 32172 52052 32228
rect 51212 31778 51268 31780
rect 51212 31726 51214 31778
rect 51214 31726 51266 31778
rect 51266 31726 51268 31778
rect 51212 31724 51268 31726
rect 51772 31778 51828 31780
rect 51772 31726 51774 31778
rect 51774 31726 51826 31778
rect 51826 31726 51828 31778
rect 51772 31724 51828 31726
rect 51548 31666 51604 31668
rect 51548 31614 51550 31666
rect 51550 31614 51602 31666
rect 51602 31614 51604 31666
rect 51548 31612 51604 31614
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 49196 30828 49252 30884
rect 49756 30882 49812 30884
rect 49756 30830 49758 30882
rect 49758 30830 49810 30882
rect 49810 30830 49812 30882
rect 49756 30828 49812 30830
rect 49980 30828 50036 30884
rect 45836 30156 45892 30212
rect 48860 30210 48916 30212
rect 48860 30158 48862 30210
rect 48862 30158 48914 30210
rect 48914 30158 48916 30210
rect 48860 30156 48916 30158
rect 49308 30210 49364 30212
rect 49308 30158 49310 30210
rect 49310 30158 49362 30210
rect 49362 30158 49364 30210
rect 49308 30156 49364 30158
rect 50876 31164 50932 31220
rect 50652 30994 50708 30996
rect 50652 30942 50654 30994
rect 50654 30942 50706 30994
rect 50706 30942 50708 30994
rect 50652 30940 50708 30942
rect 50540 30828 50596 30884
rect 52668 31890 52724 31892
rect 52668 31838 52670 31890
rect 52670 31838 52722 31890
rect 52722 31838 52724 31890
rect 52668 31836 52724 31838
rect 56588 37996 56644 38052
rect 56140 37548 56196 37604
rect 56028 37100 56084 37156
rect 56812 37772 56868 37828
rect 56812 36988 56868 37044
rect 57148 39058 57204 39060
rect 57148 39006 57150 39058
rect 57150 39006 57202 39058
rect 57202 39006 57204 39058
rect 57148 39004 57204 39006
rect 57372 40514 57428 40516
rect 57372 40462 57374 40514
rect 57374 40462 57426 40514
rect 57426 40462 57428 40514
rect 57372 40460 57428 40462
rect 57260 37826 57316 37828
rect 57260 37774 57262 37826
rect 57262 37774 57314 37826
rect 57314 37774 57316 37826
rect 57260 37772 57316 37774
rect 57260 37266 57316 37268
rect 57260 37214 57262 37266
rect 57262 37214 57314 37266
rect 57314 37214 57316 37266
rect 57260 37212 57316 37214
rect 57148 37154 57204 37156
rect 57148 37102 57150 37154
rect 57150 37102 57202 37154
rect 57202 37102 57204 37154
rect 57148 37100 57204 37102
rect 57260 36428 57316 36484
rect 56588 35810 56644 35812
rect 56588 35758 56590 35810
rect 56590 35758 56642 35810
rect 56642 35758 56644 35810
rect 56588 35756 56644 35758
rect 57036 35698 57092 35700
rect 57036 35646 57038 35698
rect 57038 35646 57090 35698
rect 57090 35646 57092 35698
rect 57036 35644 57092 35646
rect 57932 35698 57988 35700
rect 57932 35646 57934 35698
rect 57934 35646 57986 35698
rect 57986 35646 57988 35698
rect 57932 35644 57988 35646
rect 57260 35532 57316 35588
rect 58044 35586 58100 35588
rect 58044 35534 58046 35586
rect 58046 35534 58098 35586
rect 58098 35534 58100 35586
rect 58044 35532 58100 35534
rect 56028 34018 56084 34020
rect 56028 33966 56030 34018
rect 56030 33966 56082 34018
rect 56082 33966 56084 34018
rect 56028 33964 56084 33966
rect 55916 32172 55972 32228
rect 52108 31554 52164 31556
rect 52108 31502 52110 31554
rect 52110 31502 52162 31554
rect 52162 31502 52164 31554
rect 52108 31500 52164 31502
rect 51996 31218 52052 31220
rect 51996 31166 51998 31218
rect 51998 31166 52050 31218
rect 52050 31166 52052 31218
rect 51996 31164 52052 31166
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 42140 28866 42196 28868
rect 42140 28814 42142 28866
rect 42142 28814 42194 28866
rect 42194 28814 42196 28866
rect 42140 28812 42196 28814
rect 42812 28812 42868 28868
rect 41916 28642 41972 28644
rect 41916 28590 41918 28642
rect 41918 28590 41970 28642
rect 41970 28590 41972 28642
rect 41916 28588 41972 28590
rect 42252 28530 42308 28532
rect 42252 28478 42254 28530
rect 42254 28478 42306 28530
rect 42306 28478 42308 28530
rect 42252 28476 42308 28478
rect 41804 27916 41860 27972
rect 40236 27692 40292 27748
rect 40684 27692 40740 27748
rect 40460 27132 40516 27188
rect 39900 26514 39956 26516
rect 39900 26462 39902 26514
rect 39902 26462 39954 26514
rect 39954 26462 39956 26514
rect 39900 26460 39956 26462
rect 40908 27132 40964 27188
rect 40684 26236 40740 26292
rect 39452 25618 39508 25620
rect 39452 25566 39454 25618
rect 39454 25566 39506 25618
rect 39506 25566 39508 25618
rect 39452 25564 39508 25566
rect 41132 27020 41188 27076
rect 41132 26460 41188 26516
rect 41244 26908 41300 26964
rect 42140 27074 42196 27076
rect 42140 27022 42142 27074
rect 42142 27022 42194 27074
rect 42194 27022 42196 27074
rect 42140 27020 42196 27022
rect 40684 25564 40740 25620
rect 42476 26962 42532 26964
rect 42476 26910 42478 26962
rect 42478 26910 42530 26962
rect 42530 26910 42532 26962
rect 42476 26908 42532 26910
rect 41804 26290 41860 26292
rect 41804 26238 41806 26290
rect 41806 26238 41858 26290
rect 41858 26238 41860 26290
rect 41804 26236 41860 26238
rect 44044 28812 44100 28868
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 33852 24834 33908 24836
rect 33852 24782 33854 24834
rect 33854 24782 33906 24834
rect 33906 24782 33908 24834
rect 33852 24780 33908 24782
rect 34860 24556 34916 24612
rect 33852 23884 33908 23940
rect 33740 23436 33796 23492
rect 35980 24610 36036 24612
rect 35980 24558 35982 24610
rect 35982 24558 36034 24610
rect 36034 24558 36036 24610
rect 35980 24556 36036 24558
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34860 23772 34916 23828
rect 33628 22204 33684 22260
rect 33404 21756 33460 21812
rect 32956 20076 33012 20132
rect 32172 16156 32228 16212
rect 32396 15932 32452 15988
rect 32060 15484 32116 15540
rect 33068 20018 33124 20020
rect 33068 19966 33070 20018
rect 33070 19966 33122 20018
rect 33122 19966 33124 20018
rect 33068 19964 33124 19966
rect 33516 21420 33572 21476
rect 36092 23772 36148 23828
rect 33852 22316 33908 22372
rect 33852 21698 33908 21700
rect 33852 21646 33854 21698
rect 33854 21646 33906 21698
rect 33906 21646 33908 21698
rect 33852 21644 33908 21646
rect 33628 21084 33684 21140
rect 33852 20748 33908 20804
rect 33740 19964 33796 20020
rect 33404 19404 33460 19460
rect 32956 19122 33012 19124
rect 32956 19070 32958 19122
rect 32958 19070 33010 19122
rect 33010 19070 33012 19122
rect 32956 19068 33012 19070
rect 33292 18620 33348 18676
rect 33740 18620 33796 18676
rect 33628 18450 33684 18452
rect 33628 18398 33630 18450
rect 33630 18398 33682 18450
rect 33682 18398 33684 18450
rect 33628 18396 33684 18398
rect 33068 18284 33124 18340
rect 32844 18060 32900 18116
rect 33068 17836 33124 17892
rect 33180 17442 33236 17444
rect 33180 17390 33182 17442
rect 33182 17390 33234 17442
rect 33234 17390 33236 17442
rect 33180 17388 33236 17390
rect 33180 17052 33236 17108
rect 33292 16940 33348 16996
rect 33068 16882 33124 16884
rect 33068 16830 33070 16882
rect 33070 16830 33122 16882
rect 33122 16830 33124 16882
rect 33068 16828 33124 16830
rect 35308 22876 35364 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35084 22482 35140 22484
rect 35084 22430 35086 22482
rect 35086 22430 35138 22482
rect 35138 22430 35140 22482
rect 35084 22428 35140 22430
rect 37772 23826 37828 23828
rect 37772 23774 37774 23826
rect 37774 23774 37826 23826
rect 37826 23774 37828 23826
rect 37772 23772 37828 23774
rect 36540 23042 36596 23044
rect 36540 22990 36542 23042
rect 36542 22990 36594 23042
rect 36594 22990 36596 23042
rect 36540 22988 36596 22990
rect 37436 22988 37492 23044
rect 35644 22370 35700 22372
rect 35644 22318 35646 22370
rect 35646 22318 35698 22370
rect 35698 22318 35700 22370
rect 35644 22316 35700 22318
rect 36988 22370 37044 22372
rect 36988 22318 36990 22370
rect 36990 22318 37042 22370
rect 37042 22318 37044 22370
rect 36988 22316 37044 22318
rect 35308 22258 35364 22260
rect 35308 22206 35310 22258
rect 35310 22206 35362 22258
rect 35362 22206 35364 22258
rect 35308 22204 35364 22206
rect 35084 21980 35140 22036
rect 34300 21532 34356 21588
rect 34636 21644 34692 21700
rect 34972 21420 35028 21476
rect 34412 19852 34468 19908
rect 34636 21084 34692 21140
rect 34188 19404 34244 19460
rect 34076 19010 34132 19012
rect 34076 18958 34078 19010
rect 34078 18958 34130 19010
rect 34130 18958 34132 19010
rect 34076 18956 34132 18958
rect 35868 22258 35924 22260
rect 35868 22206 35870 22258
rect 35870 22206 35922 22258
rect 35922 22206 35924 22258
rect 35868 22204 35924 22206
rect 37548 22258 37604 22260
rect 37548 22206 37550 22258
rect 37550 22206 37602 22258
rect 37602 22206 37604 22258
rect 37548 22204 37604 22206
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35308 20018 35364 20020
rect 35308 19966 35310 20018
rect 35310 19966 35362 20018
rect 35362 19966 35364 20018
rect 35308 19964 35364 19966
rect 35420 19740 35476 19796
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35084 19404 35140 19460
rect 34524 18956 34580 19012
rect 32620 14924 32676 14980
rect 31948 14642 32004 14644
rect 31948 14590 31950 14642
rect 31950 14590 32002 14642
rect 32002 14590 32004 14642
rect 31948 14588 32004 14590
rect 32284 14364 32340 14420
rect 31948 14140 32004 14196
rect 31836 12738 31892 12740
rect 31836 12686 31838 12738
rect 31838 12686 31890 12738
rect 31890 12686 31892 12738
rect 31836 12684 31892 12686
rect 31388 11900 31444 11956
rect 31388 8876 31444 8932
rect 31276 8146 31332 8148
rect 31276 8094 31278 8146
rect 31278 8094 31330 8146
rect 31330 8094 31332 8146
rect 31276 8092 31332 8094
rect 32060 13692 32116 13748
rect 32620 14306 32676 14308
rect 32620 14254 32622 14306
rect 32622 14254 32674 14306
rect 32674 14254 32676 14306
rect 32620 14252 32676 14254
rect 32732 14140 32788 14196
rect 33404 15932 33460 15988
rect 32956 14306 33012 14308
rect 32956 14254 32958 14306
rect 32958 14254 33010 14306
rect 33010 14254 33012 14306
rect 32956 14252 33012 14254
rect 32396 13580 32452 13636
rect 32172 13244 32228 13300
rect 32396 12796 32452 12852
rect 32060 12402 32116 12404
rect 32060 12350 32062 12402
rect 32062 12350 32114 12402
rect 32114 12350 32116 12402
rect 32060 12348 32116 12350
rect 32508 10780 32564 10836
rect 32844 12348 32900 12404
rect 31948 8146 32004 8148
rect 31948 8094 31950 8146
rect 31950 8094 32002 8146
rect 32002 8094 32004 8146
rect 31948 8092 32004 8094
rect 31500 7532 31556 7588
rect 33292 13858 33348 13860
rect 33292 13806 33294 13858
rect 33294 13806 33346 13858
rect 33346 13806 33348 13858
rect 33292 13804 33348 13806
rect 34636 18620 34692 18676
rect 33964 17500 34020 17556
rect 33740 16940 33796 16996
rect 33852 17388 33908 17444
rect 36092 22146 36148 22148
rect 36092 22094 36094 22146
rect 36094 22094 36146 22146
rect 36146 22094 36148 22146
rect 36092 22092 36148 22094
rect 36316 22146 36372 22148
rect 36316 22094 36318 22146
rect 36318 22094 36370 22146
rect 36370 22094 36372 22146
rect 36316 22092 36372 22094
rect 37324 21868 37380 21924
rect 36428 21644 36484 21700
rect 35084 18620 35140 18676
rect 35644 21532 35700 21588
rect 38220 22988 38276 23044
rect 38220 22146 38276 22148
rect 38220 22094 38222 22146
rect 38222 22094 38274 22146
rect 38274 22094 38276 22146
rect 38220 22092 38276 22094
rect 38668 23042 38724 23044
rect 38668 22990 38670 23042
rect 38670 22990 38722 23042
rect 38722 22990 38724 23042
rect 38668 22988 38724 22990
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 38556 21980 38612 22036
rect 38108 21868 38164 21924
rect 37996 21532 38052 21588
rect 39228 21756 39284 21812
rect 37772 20860 37828 20916
rect 36428 20802 36484 20804
rect 36428 20750 36430 20802
rect 36430 20750 36482 20802
rect 36482 20750 36484 20802
rect 36428 20748 36484 20750
rect 35980 20636 36036 20692
rect 35644 19852 35700 19908
rect 34412 18284 34468 18340
rect 34524 18396 34580 18452
rect 34524 17948 34580 18004
rect 34412 17052 34468 17108
rect 34636 17500 34692 17556
rect 34524 16716 34580 16772
rect 34524 16156 34580 16212
rect 34300 16098 34356 16100
rect 34300 16046 34302 16098
rect 34302 16046 34354 16098
rect 34354 16046 34356 16098
rect 34300 16044 34356 16046
rect 33516 14924 33572 14980
rect 33852 13804 33908 13860
rect 33292 13634 33348 13636
rect 33292 13582 33294 13634
rect 33294 13582 33346 13634
rect 33346 13582 33348 13634
rect 33292 13580 33348 13582
rect 33180 12850 33236 12852
rect 33180 12798 33182 12850
rect 33182 12798 33234 12850
rect 33234 12798 33236 12850
rect 33180 12796 33236 12798
rect 33180 11452 33236 11508
rect 32396 9826 32452 9828
rect 32396 9774 32398 9826
rect 32398 9774 32450 9826
rect 32450 9774 32452 9826
rect 32396 9772 32452 9774
rect 33404 10834 33460 10836
rect 33404 10782 33406 10834
rect 33406 10782 33458 10834
rect 33458 10782 33460 10834
rect 33404 10780 33460 10782
rect 32844 9602 32900 9604
rect 32844 9550 32846 9602
rect 32846 9550 32898 9602
rect 32898 9550 32900 9602
rect 32844 9548 32900 9550
rect 34300 14252 34356 14308
rect 33964 9996 34020 10052
rect 33404 9826 33460 9828
rect 33404 9774 33406 9826
rect 33406 9774 33458 9826
rect 33458 9774 33460 9826
rect 33404 9772 33460 9774
rect 33628 9548 33684 9604
rect 33628 9324 33684 9380
rect 33404 9212 33460 9268
rect 33180 9154 33236 9156
rect 33180 9102 33182 9154
rect 33182 9102 33234 9154
rect 33234 9102 33236 9154
rect 33180 9100 33236 9102
rect 33852 9212 33908 9268
rect 33628 9100 33684 9156
rect 33068 8764 33124 8820
rect 33068 8540 33124 8596
rect 31500 6636 31556 6692
rect 32844 6748 32900 6804
rect 31276 6578 31332 6580
rect 31276 6526 31278 6578
rect 31278 6526 31330 6578
rect 31330 6526 31332 6578
rect 31276 6524 31332 6526
rect 31052 6076 31108 6132
rect 28924 5794 28980 5796
rect 28924 5742 28926 5794
rect 28926 5742 28978 5794
rect 28978 5742 28980 5794
rect 28924 5740 28980 5742
rect 29260 5180 29316 5236
rect 28476 4956 28532 5012
rect 24332 4562 24388 4564
rect 24332 4510 24334 4562
rect 24334 4510 24386 4562
rect 24386 4510 24388 4562
rect 24332 4508 24388 4510
rect 25564 4562 25620 4564
rect 25564 4510 25566 4562
rect 25566 4510 25618 4562
rect 25618 4510 25620 4562
rect 25564 4508 25620 4510
rect 26012 4508 26068 4564
rect 32060 6578 32116 6580
rect 32060 6526 32062 6578
rect 32062 6526 32114 6578
rect 32114 6526 32116 6578
rect 32060 6524 32116 6526
rect 32844 6076 32900 6132
rect 32956 6412 33012 6468
rect 32172 6018 32228 6020
rect 32172 5966 32174 6018
rect 32174 5966 32226 6018
rect 32226 5966 32228 6018
rect 32172 5964 32228 5966
rect 32396 5964 32452 6020
rect 30156 5628 30212 5684
rect 30828 5180 30884 5236
rect 33404 8540 33460 8596
rect 33516 8764 33572 8820
rect 33964 9100 34020 9156
rect 33740 8988 33796 9044
rect 33404 7980 33460 8036
rect 33740 7980 33796 8036
rect 34412 13746 34468 13748
rect 34412 13694 34414 13746
rect 34414 13694 34466 13746
rect 34466 13694 34468 13746
rect 34412 13692 34468 13694
rect 34300 12290 34356 12292
rect 34300 12238 34302 12290
rect 34302 12238 34354 12290
rect 34354 12238 34356 12290
rect 34300 12236 34356 12238
rect 34188 10780 34244 10836
rect 35084 18450 35140 18452
rect 35084 18398 35086 18450
rect 35086 18398 35138 18450
rect 35138 18398 35140 18450
rect 35084 18396 35140 18398
rect 35420 18674 35476 18676
rect 35420 18622 35422 18674
rect 35422 18622 35474 18674
rect 35474 18622 35476 18674
rect 35420 18620 35476 18622
rect 35308 18284 35364 18340
rect 34860 18060 34916 18116
rect 34972 17724 35028 17780
rect 35084 18172 35140 18228
rect 35532 18172 35588 18228
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 17554 35252 17556
rect 35196 17502 35198 17554
rect 35198 17502 35250 17554
rect 35250 17502 35252 17554
rect 35196 17500 35252 17502
rect 34972 16940 35028 16996
rect 35756 20524 35812 20580
rect 35868 20018 35924 20020
rect 35868 19966 35870 20018
rect 35870 19966 35922 20018
rect 35922 19966 35924 20018
rect 35868 19964 35924 19966
rect 35868 19740 35924 19796
rect 36316 20412 36372 20468
rect 37212 20412 37268 20468
rect 37212 20188 37268 20244
rect 37548 20690 37604 20692
rect 37548 20638 37550 20690
rect 37550 20638 37602 20690
rect 37602 20638 37604 20690
rect 37548 20636 37604 20638
rect 37996 20914 38052 20916
rect 37996 20862 37998 20914
rect 37998 20862 38050 20914
rect 38050 20862 38052 20914
rect 37996 20860 38052 20862
rect 38668 20860 38724 20916
rect 38444 20748 38500 20804
rect 37772 20636 37828 20692
rect 38332 20690 38388 20692
rect 38332 20638 38334 20690
rect 38334 20638 38386 20690
rect 38386 20638 38388 20690
rect 38332 20636 38388 20638
rect 36316 18284 36372 18340
rect 37212 19906 37268 19908
rect 37212 19854 37214 19906
rect 37214 19854 37266 19906
rect 37266 19854 37268 19906
rect 37212 19852 37268 19854
rect 36652 19292 36708 19348
rect 37660 20188 37716 20244
rect 39004 20802 39060 20804
rect 39004 20750 39006 20802
rect 39006 20750 39058 20802
rect 39058 20750 39060 20802
rect 39004 20748 39060 20750
rect 38892 20636 38948 20692
rect 38892 20300 38948 20356
rect 36540 18284 36596 18340
rect 36316 17836 36372 17892
rect 35980 17724 36036 17780
rect 36204 17778 36260 17780
rect 36204 17726 36206 17778
rect 36206 17726 36258 17778
rect 36258 17726 36260 17778
rect 36204 17724 36260 17726
rect 36428 17948 36484 18004
rect 35532 16828 35588 16884
rect 36204 16828 36260 16884
rect 35980 16770 36036 16772
rect 35980 16718 35982 16770
rect 35982 16718 36034 16770
rect 36034 16718 36036 16770
rect 35980 16716 36036 16718
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 37100 17948 37156 18004
rect 36876 17666 36932 17668
rect 36876 17614 36878 17666
rect 36878 17614 36930 17666
rect 36930 17614 36932 17666
rect 36876 17612 36932 17614
rect 37100 17612 37156 17668
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35084 14418 35140 14420
rect 35084 14366 35086 14418
rect 35086 14366 35138 14418
rect 35138 14366 35140 14418
rect 35084 14364 35140 14366
rect 34860 13692 34916 13748
rect 34972 13132 35028 13188
rect 35420 13468 35476 13524
rect 35644 13522 35700 13524
rect 35644 13470 35646 13522
rect 35646 13470 35698 13522
rect 35698 13470 35700 13522
rect 35644 13468 35700 13470
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35868 13858 35924 13860
rect 35868 13806 35870 13858
rect 35870 13806 35922 13858
rect 35922 13806 35924 13858
rect 35868 13804 35924 13806
rect 35308 13132 35364 13188
rect 34972 12962 35028 12964
rect 34972 12910 34974 12962
rect 34974 12910 35026 12962
rect 35026 12910 35028 12962
rect 34972 12908 35028 12910
rect 34748 12796 34804 12852
rect 34636 12178 34692 12180
rect 34636 12126 34638 12178
rect 34638 12126 34690 12178
rect 34690 12126 34692 12178
rect 34636 12124 34692 12126
rect 34972 11900 35028 11956
rect 34524 10668 34580 10724
rect 34300 9996 34356 10052
rect 34972 10722 35028 10724
rect 34972 10670 34974 10722
rect 34974 10670 35026 10722
rect 35026 10670 35028 10722
rect 34972 10668 35028 10670
rect 34524 9996 34580 10052
rect 34300 9266 34356 9268
rect 34300 9214 34302 9266
rect 34302 9214 34354 9266
rect 34354 9214 34356 9266
rect 34300 9212 34356 9214
rect 34748 9100 34804 9156
rect 35532 13074 35588 13076
rect 35532 13022 35534 13074
rect 35534 13022 35586 13074
rect 35586 13022 35588 13074
rect 35532 13020 35588 13022
rect 35420 12850 35476 12852
rect 35420 12798 35422 12850
rect 35422 12798 35474 12850
rect 35474 12798 35476 12850
rect 35420 12796 35476 12798
rect 35532 12572 35588 12628
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 9996 35252 10052
rect 35756 12962 35812 12964
rect 35756 12910 35758 12962
rect 35758 12910 35810 12962
rect 35810 12910 35812 12962
rect 35756 12908 35812 12910
rect 36092 13746 36148 13748
rect 36092 13694 36094 13746
rect 36094 13694 36146 13746
rect 36146 13694 36148 13746
rect 36092 13692 36148 13694
rect 36988 15484 37044 15540
rect 36540 15314 36596 15316
rect 36540 15262 36542 15314
rect 36542 15262 36594 15314
rect 36594 15262 36596 15314
rect 36540 15260 36596 15262
rect 36428 14418 36484 14420
rect 36428 14366 36430 14418
rect 36430 14366 36482 14418
rect 36482 14366 36484 14418
rect 36428 14364 36484 14366
rect 36876 15148 36932 15204
rect 37548 18284 37604 18340
rect 37436 17724 37492 17780
rect 37436 15820 37492 15876
rect 38892 19964 38948 20020
rect 37772 19346 37828 19348
rect 37772 19294 37774 19346
rect 37774 19294 37826 19346
rect 37826 19294 37828 19346
rect 37772 19292 37828 19294
rect 38108 19292 38164 19348
rect 38444 18732 38500 18788
rect 37996 18338 38052 18340
rect 37996 18286 37998 18338
rect 37998 18286 38050 18338
rect 38050 18286 38052 18338
rect 37996 18284 38052 18286
rect 38220 16716 38276 16772
rect 38108 15874 38164 15876
rect 38108 15822 38110 15874
rect 38110 15822 38162 15874
rect 38162 15822 38164 15874
rect 38108 15820 38164 15822
rect 39116 20076 39172 20132
rect 39676 21644 39732 21700
rect 40124 21756 40180 21812
rect 39340 21532 39396 21588
rect 42812 21756 42868 21812
rect 40908 21644 40964 21700
rect 39788 20690 39844 20692
rect 39788 20638 39790 20690
rect 39790 20638 39842 20690
rect 39842 20638 39844 20690
rect 39788 20636 39844 20638
rect 40796 20860 40852 20916
rect 40236 20636 40292 20692
rect 40460 20636 40516 20692
rect 39340 20188 39396 20244
rect 39676 20300 39732 20356
rect 40236 20242 40292 20244
rect 40236 20190 40238 20242
rect 40238 20190 40290 20242
rect 40290 20190 40292 20242
rect 40236 20188 40292 20190
rect 40012 20130 40068 20132
rect 40012 20078 40014 20130
rect 40014 20078 40066 20130
rect 40066 20078 40068 20130
rect 40012 20076 40068 20078
rect 39900 19346 39956 19348
rect 39900 19294 39902 19346
rect 39902 19294 39954 19346
rect 39954 19294 39956 19346
rect 39900 19292 39956 19294
rect 39228 18060 39284 18116
rect 39900 18338 39956 18340
rect 39900 18286 39902 18338
rect 39902 18286 39954 18338
rect 39954 18286 39956 18338
rect 39900 18284 39956 18286
rect 39340 17948 39396 18004
rect 39004 17778 39060 17780
rect 39004 17726 39006 17778
rect 39006 17726 39058 17778
rect 39058 17726 39060 17778
rect 39004 17724 39060 17726
rect 40684 20524 40740 20580
rect 40460 18396 40516 18452
rect 41692 20860 41748 20916
rect 42364 21420 42420 21476
rect 42252 20690 42308 20692
rect 42252 20638 42254 20690
rect 42254 20638 42306 20690
rect 42306 20638 42308 20690
rect 42252 20636 42308 20638
rect 40908 19852 40964 19908
rect 41132 20018 41188 20020
rect 41132 19966 41134 20018
rect 41134 19966 41186 20018
rect 41186 19966 41188 20018
rect 41132 19964 41188 19966
rect 42252 19906 42308 19908
rect 42252 19854 42254 19906
rect 42254 19854 42306 19906
rect 42306 19854 42308 19906
rect 42252 19852 42308 19854
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 43820 21474 43876 21476
rect 43820 21422 43822 21474
rect 43822 21422 43874 21474
rect 43874 21422 43876 21474
rect 43820 21420 43876 21422
rect 43372 19852 43428 19908
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 44268 19852 44324 19908
rect 41244 19292 41300 19348
rect 42812 19346 42868 19348
rect 42812 19294 42814 19346
rect 42814 19294 42866 19346
rect 42866 19294 42868 19346
rect 42812 19292 42868 19294
rect 41692 18338 41748 18340
rect 41692 18286 41694 18338
rect 41694 18286 41746 18338
rect 41746 18286 41748 18338
rect 41692 18284 41748 18286
rect 40012 18172 40068 18228
rect 40572 17778 40628 17780
rect 40572 17726 40574 17778
rect 40574 17726 40626 17778
rect 40626 17726 40628 17778
rect 40572 17724 40628 17726
rect 39900 17666 39956 17668
rect 39900 17614 39902 17666
rect 39902 17614 39954 17666
rect 39954 17614 39956 17666
rect 39900 17612 39956 17614
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 43372 18172 43428 18228
rect 42812 17612 42868 17668
rect 39116 16828 39172 16884
rect 41916 16882 41972 16884
rect 41916 16830 41918 16882
rect 41918 16830 41970 16882
rect 41970 16830 41972 16882
rect 41916 16828 41972 16830
rect 39228 16770 39284 16772
rect 39228 16718 39230 16770
rect 39230 16718 39282 16770
rect 39282 16718 39284 16770
rect 39228 16716 39284 16718
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 43148 16156 43204 16212
rect 43820 16156 43876 16212
rect 38668 15372 38724 15428
rect 37884 14642 37940 14644
rect 37884 14590 37886 14642
rect 37886 14590 37938 14642
rect 37938 14590 37940 14642
rect 37884 14588 37940 14590
rect 37660 14476 37716 14532
rect 36428 13468 36484 13524
rect 36540 12236 36596 12292
rect 36428 12178 36484 12180
rect 36428 12126 36430 12178
rect 36430 12126 36482 12178
rect 36482 12126 36484 12178
rect 36428 12124 36484 12126
rect 38668 15202 38724 15204
rect 38668 15150 38670 15202
rect 38670 15150 38722 15202
rect 38722 15150 38724 15202
rect 38668 15148 38724 15150
rect 37996 12796 38052 12852
rect 38220 12402 38276 12404
rect 38220 12350 38222 12402
rect 38222 12350 38274 12402
rect 38274 12350 38276 12402
rect 38220 12348 38276 12350
rect 37100 11788 37156 11844
rect 36316 11452 36372 11508
rect 36204 10668 36260 10724
rect 36428 10556 36484 10612
rect 36876 9996 36932 10052
rect 35196 9436 35252 9492
rect 34524 8876 34580 8932
rect 34524 8204 34580 8260
rect 34636 8764 34692 8820
rect 33180 5964 33236 6020
rect 33852 6018 33908 6020
rect 33852 5966 33854 6018
rect 33854 5966 33906 6018
rect 33906 5966 33908 6018
rect 33852 5964 33908 5966
rect 33068 5740 33124 5796
rect 33180 5682 33236 5684
rect 33180 5630 33182 5682
rect 33182 5630 33234 5682
rect 33234 5630 33236 5682
rect 33180 5628 33236 5630
rect 32508 5180 32564 5236
rect 34300 5740 34356 5796
rect 35756 9602 35812 9604
rect 35756 9550 35758 9602
rect 35758 9550 35810 9602
rect 35810 9550 35812 9602
rect 35756 9548 35812 9550
rect 36204 9436 36260 9492
rect 35756 9212 35812 9268
rect 35308 9154 35364 9156
rect 35308 9102 35310 9154
rect 35310 9102 35362 9154
rect 35362 9102 35364 9154
rect 35308 9100 35364 9102
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35868 8316 35924 8372
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35420 6748 35476 6804
rect 36092 8258 36148 8260
rect 36092 8206 36094 8258
rect 36094 8206 36146 8258
rect 36146 8206 36148 8258
rect 36092 8204 36148 8206
rect 35532 5740 35588 5796
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34076 5234 34132 5236
rect 34076 5182 34078 5234
rect 34078 5182 34130 5234
rect 34130 5182 34132 5234
rect 34076 5180 34132 5182
rect 36428 9324 36484 9380
rect 36988 9324 37044 9380
rect 36540 9212 36596 9268
rect 37548 11954 37604 11956
rect 37548 11902 37550 11954
rect 37550 11902 37602 11954
rect 37602 11902 37604 11954
rect 37548 11900 37604 11902
rect 37212 10556 37268 10612
rect 37884 11452 37940 11508
rect 37324 9324 37380 9380
rect 37660 10556 37716 10612
rect 37436 9042 37492 9044
rect 37436 8990 37438 9042
rect 37438 8990 37490 9042
rect 37490 8990 37492 9042
rect 37436 8988 37492 8990
rect 37436 8370 37492 8372
rect 37436 8318 37438 8370
rect 37438 8318 37490 8370
rect 37490 8318 37492 8370
rect 37436 8316 37492 8318
rect 39004 14588 39060 14644
rect 38444 13858 38500 13860
rect 38444 13806 38446 13858
rect 38446 13806 38498 13858
rect 38498 13806 38500 13858
rect 38444 13804 38500 13806
rect 42700 15372 42756 15428
rect 42476 15148 42532 15204
rect 42140 14418 42196 14420
rect 42140 14366 42142 14418
rect 42142 14366 42194 14418
rect 42194 14366 42196 14418
rect 42140 14364 42196 14366
rect 39004 13468 39060 13524
rect 39788 13468 39844 13524
rect 39116 12850 39172 12852
rect 39116 12798 39118 12850
rect 39118 12798 39170 12850
rect 39170 12798 39172 12850
rect 39116 12796 39172 12798
rect 39340 12962 39396 12964
rect 39340 12910 39342 12962
rect 39342 12910 39394 12962
rect 39394 12910 39396 12962
rect 39340 12908 39396 12910
rect 39676 12850 39732 12852
rect 39676 12798 39678 12850
rect 39678 12798 39730 12850
rect 39730 12798 39732 12850
rect 39676 12796 39732 12798
rect 39228 12348 39284 12404
rect 39676 12290 39732 12292
rect 39676 12238 39678 12290
rect 39678 12238 39730 12290
rect 39730 12238 39732 12290
rect 39676 12236 39732 12238
rect 38892 11954 38948 11956
rect 38892 11902 38894 11954
rect 38894 11902 38946 11954
rect 38946 11902 38948 11954
rect 38892 11900 38948 11902
rect 37996 9266 38052 9268
rect 37996 9214 37998 9266
rect 37998 9214 38050 9266
rect 38050 9214 38052 9266
rect 37996 9212 38052 9214
rect 38444 9212 38500 9268
rect 38892 10780 38948 10836
rect 39452 9996 39508 10052
rect 38556 8988 38612 9044
rect 42140 13692 42196 13748
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 44268 15314 44324 15316
rect 44268 15262 44270 15314
rect 44270 15262 44322 15314
rect 44322 15262 44324 15314
rect 44268 15260 44324 15262
rect 45276 15260 45332 15316
rect 43820 15202 43876 15204
rect 43820 15150 43822 15202
rect 43822 15150 43874 15202
rect 43874 15150 43876 15202
rect 43820 15148 43876 15150
rect 42588 13858 42644 13860
rect 42588 13806 42590 13858
rect 42590 13806 42642 13858
rect 42642 13806 42644 13858
rect 42588 13804 42644 13806
rect 39788 10780 39844 10836
rect 39788 9996 39844 10052
rect 40012 9884 40068 9940
rect 42812 13858 42868 13860
rect 42812 13806 42814 13858
rect 42814 13806 42866 13858
rect 42866 13806 42868 13858
rect 42812 13804 42868 13806
rect 42812 13468 42868 13524
rect 43596 13858 43652 13860
rect 43596 13806 43598 13858
rect 43598 13806 43650 13858
rect 43650 13806 43652 13858
rect 43596 13804 43652 13806
rect 43260 13468 43316 13524
rect 44380 13746 44436 13748
rect 44380 13694 44382 13746
rect 44382 13694 44434 13746
rect 44434 13694 44436 13746
rect 44380 13692 44436 13694
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 47068 13692 47124 13748
rect 44604 13020 44660 13076
rect 43820 12908 43876 12964
rect 43148 12290 43204 12292
rect 43148 12238 43150 12290
rect 43150 12238 43202 12290
rect 43202 12238 43204 12290
rect 43148 12236 43204 12238
rect 44268 12850 44324 12852
rect 44268 12798 44270 12850
rect 44270 12798 44322 12850
rect 44322 12798 44324 12850
rect 44268 12796 44324 12798
rect 44044 12348 44100 12404
rect 43932 12290 43988 12292
rect 43932 12238 43934 12290
rect 43934 12238 43986 12290
rect 43986 12238 43988 12290
rect 43932 12236 43988 12238
rect 43260 11900 43316 11956
rect 44604 11900 44660 11956
rect 47740 13074 47796 13076
rect 47740 13022 47742 13074
rect 47742 13022 47794 13074
rect 47794 13022 47796 13074
rect 47740 13020 47796 13022
rect 42476 11564 42532 11620
rect 44268 11564 44324 11620
rect 45612 12850 45668 12852
rect 45612 12798 45614 12850
rect 45614 12798 45666 12850
rect 45666 12798 45668 12850
rect 45612 12796 45668 12798
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 44940 12402 44996 12404
rect 44940 12350 44942 12402
rect 44942 12350 44994 12402
rect 44994 12350 44996 12402
rect 44940 12348 44996 12350
rect 41356 9996 41412 10052
rect 42252 9996 42308 10052
rect 41580 9938 41636 9940
rect 41580 9886 41582 9938
rect 41582 9886 41634 9938
rect 41634 9886 41636 9938
rect 41580 9884 41636 9886
rect 42812 9996 42868 10052
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 44828 9772 44884 9828
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 37996 8204 38052 8260
rect 38220 8204 38276 8260
rect 39340 8258 39396 8260
rect 39340 8206 39342 8258
rect 39342 8206 39394 8258
rect 39394 8206 39396 8258
rect 39340 8204 39396 8206
rect 38444 7586 38500 7588
rect 38444 7534 38446 7586
rect 38446 7534 38498 7586
rect 38498 7534 38500 7586
rect 38444 7532 38500 7534
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 39788 6524 39844 6580
rect 40348 6578 40404 6580
rect 40348 6526 40350 6578
rect 40350 6526 40402 6578
rect 40402 6526 40404 6578
rect 40348 6524 40404 6526
rect 36316 5180 36372 5236
rect 36652 4508 36708 4564
rect 36988 5234 37044 5236
rect 36988 5182 36990 5234
rect 36990 5182 37042 5234
rect 37042 5182 37044 5234
rect 36988 5180 37044 5182
rect 39900 5180 39956 5236
rect 37324 5068 37380 5124
rect 39116 5122 39172 5124
rect 39116 5070 39118 5122
rect 39118 5070 39170 5122
rect 39170 5070 39172 5122
rect 39116 5068 39172 5070
rect 40348 5234 40404 5236
rect 40348 5182 40350 5234
rect 40350 5182 40402 5234
rect 40402 5182 40404 5234
rect 40348 5180 40404 5182
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 41132 5180 41188 5236
rect 37772 4562 37828 4564
rect 37772 4510 37774 4562
rect 37774 4510 37826 4562
rect 37826 4510 37828 4562
rect 37772 4508 37828 4510
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 39900 4508 39956 4564
rect 34748 4172 34804 4228
rect 35868 4226 35924 4228
rect 35868 4174 35870 4226
rect 35870 4174 35922 4226
rect 35922 4174 35924 4226
rect 35868 4172 35924 4174
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 33170 57036 33180 57092
rect 33236 57036 34636 57092
rect 34692 57036 34702 57092
rect 36754 57036 36764 57092
rect 36820 57036 37996 57092
rect 38052 57036 38062 57092
rect 38098 56924 38108 56980
rect 38164 56924 40572 56980
rect 40628 56924 40638 56980
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4610 56252 4620 56308
rect 4676 56252 5516 56308
rect 5572 56252 5582 56308
rect 14354 56252 14364 56308
rect 14420 56252 16604 56308
rect 16660 56252 16670 56308
rect 30034 56252 30044 56308
rect 30100 56252 31052 56308
rect 31108 56252 31118 56308
rect 31378 56252 31388 56308
rect 31444 56252 32620 56308
rect 32676 56252 32686 56308
rect 33618 56252 33628 56308
rect 33684 56252 35308 56308
rect 35364 56252 35374 56308
rect 36306 56252 36316 56308
rect 36372 56252 39116 56308
rect 39172 56252 39182 56308
rect 39890 56252 39900 56308
rect 39956 56252 41132 56308
rect 41188 56252 41580 56308
rect 41636 56252 41646 56308
rect 5842 56140 5852 56196
rect 5908 56140 9100 56196
rect 9156 56140 9166 56196
rect 15026 56140 15036 56196
rect 15092 56140 15372 56196
rect 15428 56140 15438 56196
rect 37426 56140 37436 56196
rect 37492 56140 41356 56196
rect 41412 56140 41422 56196
rect 15922 56028 15932 56084
rect 15988 56028 16772 56084
rect 27458 56028 27468 56084
rect 27524 56028 28700 56084
rect 28756 56028 28766 56084
rect 38546 56028 38556 56084
rect 38612 56028 39788 56084
rect 39844 56028 39854 56084
rect 41234 56028 41244 56084
rect 41300 56028 41580 56084
rect 41636 56028 42028 56084
rect 42084 56028 42094 56084
rect 16716 55972 16772 56028
rect 13906 55916 13916 55972
rect 13972 55916 16156 55972
rect 16212 55916 16222 55972
rect 16706 55916 16716 55972
rect 16772 55916 19068 55972
rect 19124 55916 19852 55972
rect 19908 55916 19918 55972
rect 40338 55916 40348 55972
rect 40404 55916 42700 55972
rect 42756 55916 42766 55972
rect 28578 55692 28588 55748
rect 28644 55692 30268 55748
rect 30324 55692 30334 55748
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 16482 55580 16492 55636
rect 16548 55580 18060 55636
rect 18116 55580 18126 55636
rect 34066 55580 34076 55636
rect 34132 55580 34972 55636
rect 35028 55580 35038 55636
rect 15362 55468 15372 55524
rect 15428 55468 16380 55524
rect 16436 55468 16446 55524
rect 16818 55468 16828 55524
rect 16884 55468 17220 55524
rect 17164 55412 17220 55468
rect 14802 55356 14812 55412
rect 14868 55356 16940 55412
rect 16996 55356 17006 55412
rect 17164 55356 18844 55412
rect 18900 55356 19292 55412
rect 19348 55356 19358 55412
rect 19954 55356 19964 55412
rect 20020 55356 20524 55412
rect 20580 55356 21084 55412
rect 21140 55356 21150 55412
rect 27346 55356 27356 55412
rect 27412 55356 29596 55412
rect 29652 55356 29662 55412
rect 39442 55356 39452 55412
rect 39508 55356 40684 55412
rect 40740 55356 40750 55412
rect 15922 55244 15932 55300
rect 15988 55244 17500 55300
rect 17556 55244 17836 55300
rect 17892 55244 17902 55300
rect 18386 55244 18396 55300
rect 18452 55244 19628 55300
rect 19684 55244 19694 55300
rect 24658 55244 24668 55300
rect 24724 55244 25676 55300
rect 25732 55244 25742 55300
rect 18834 55132 18844 55188
rect 18900 55132 19180 55188
rect 19236 55132 19246 55188
rect 26450 55132 26460 55188
rect 26516 55132 27804 55188
rect 27860 55132 27870 55188
rect 34850 55132 34860 55188
rect 34916 55132 36204 55188
rect 36260 55132 36270 55188
rect 17602 55020 17612 55076
rect 17668 55020 18060 55076
rect 18116 55020 18956 55076
rect 19012 55020 23548 55076
rect 23604 55020 23614 55076
rect 30370 55020 30380 55076
rect 30436 55020 30828 55076
rect 30884 55020 30894 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 15586 54684 15596 54740
rect 15652 54684 16604 54740
rect 16660 54684 16670 54740
rect 21410 54684 21420 54740
rect 21476 54684 21980 54740
rect 22036 54684 22652 54740
rect 22708 54684 24668 54740
rect 24724 54684 24734 54740
rect 37650 54684 37660 54740
rect 37716 54684 38892 54740
rect 38948 54684 38958 54740
rect 16604 54628 16660 54684
rect 9986 54572 9996 54628
rect 10052 54572 10668 54628
rect 10724 54572 11452 54628
rect 11508 54572 11518 54628
rect 16604 54572 19404 54628
rect 19460 54572 20748 54628
rect 20804 54572 20814 54628
rect 16370 54460 16380 54516
rect 16436 54460 18732 54516
rect 18788 54460 18798 54516
rect 19282 54460 19292 54516
rect 19348 54460 20300 54516
rect 20356 54460 20366 54516
rect 31266 54460 31276 54516
rect 31332 54460 32396 54516
rect 32452 54460 32462 54516
rect 35746 54460 35756 54516
rect 35812 54460 37100 54516
rect 37156 54460 38780 54516
rect 38836 54460 40908 54516
rect 40964 54460 40974 54516
rect 19366 54348 19404 54404
rect 19460 54348 19470 54404
rect 28914 54348 28924 54404
rect 28980 54348 32284 54404
rect 32340 54348 32350 54404
rect 45490 54348 45500 54404
rect 45556 54348 46284 54404
rect 46340 54348 46350 54404
rect 3490 54236 3500 54292
rect 3556 54236 5516 54292
rect 5572 54236 5582 54292
rect 6962 54236 6972 54292
rect 7028 54236 8876 54292
rect 8932 54236 9884 54292
rect 9940 54236 9950 54292
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 34178 53900 34188 53956
rect 34244 53900 37436 53956
rect 37492 53900 37502 53956
rect 1586 53788 1596 53844
rect 1652 53788 4060 53844
rect 4116 53788 4126 53844
rect 18162 53788 18172 53844
rect 18228 53788 18844 53844
rect 18900 53788 19852 53844
rect 19908 53788 19918 53844
rect 23314 53788 23324 53844
rect 23380 53788 23660 53844
rect 23716 53788 23726 53844
rect 35196 53788 35756 53844
rect 35812 53788 35822 53844
rect 35970 53788 35980 53844
rect 36036 53788 37100 53844
rect 37156 53788 37772 53844
rect 37828 53788 37838 53844
rect 41570 53788 41580 53844
rect 41636 53788 42476 53844
rect 42532 53788 42542 53844
rect 35196 53732 35252 53788
rect 3826 53676 3836 53732
rect 3892 53676 4844 53732
rect 4900 53676 4910 53732
rect 22866 53676 22876 53732
rect 22932 53676 24332 53732
rect 24388 53676 24398 53732
rect 25554 53676 25564 53732
rect 25620 53676 29372 53732
rect 29428 53676 29438 53732
rect 31938 53676 31948 53732
rect 32004 53676 33180 53732
rect 33236 53676 35252 53732
rect 42354 53676 42364 53732
rect 42420 53676 43484 53732
rect 43540 53676 43550 53732
rect 12786 53564 12796 53620
rect 12852 53564 13580 53620
rect 13636 53564 15148 53620
rect 15204 53564 15820 53620
rect 15876 53564 15886 53620
rect 43026 53564 43036 53620
rect 43092 53564 43708 53620
rect 43764 53564 44212 53620
rect 44156 53508 44212 53564
rect 2370 53452 2380 53508
rect 2436 53452 3164 53508
rect 3220 53452 3230 53508
rect 16370 53452 16380 53508
rect 16436 53452 17052 53508
rect 17108 53452 23436 53508
rect 23492 53452 23502 53508
rect 42578 53452 42588 53508
rect 42644 53452 43820 53508
rect 43876 53452 43886 53508
rect 44146 53452 44156 53508
rect 44212 53452 47516 53508
rect 47572 53452 49420 53508
rect 49476 53452 51884 53508
rect 51940 53452 51950 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 44370 53228 44380 53284
rect 44436 53228 44828 53284
rect 44884 53228 46620 53284
rect 46676 53228 46686 53284
rect 14242 53116 14252 53172
rect 14308 53116 16044 53172
rect 16100 53116 16110 53172
rect 43474 53116 43484 53172
rect 43540 53116 47068 53172
rect 47124 53116 47134 53172
rect 48066 53116 48076 53172
rect 48132 53116 48860 53172
rect 48916 53116 48926 53172
rect 47068 53060 47124 53116
rect 6066 53004 6076 53060
rect 6132 53004 6972 53060
rect 7028 53004 7420 53060
rect 7476 53004 7486 53060
rect 28354 53004 28364 53060
rect 28420 53004 29596 53060
rect 29652 53004 29662 53060
rect 29922 53004 29932 53060
rect 29988 53004 30716 53060
rect 30772 53004 30940 53060
rect 30996 53004 31006 53060
rect 36418 53004 36428 53060
rect 36484 53004 37548 53060
rect 37604 53004 37614 53060
rect 47068 53004 48748 53060
rect 48804 53004 48814 53060
rect 6290 52892 6300 52948
rect 6356 52892 7308 52948
rect 7364 52892 7374 52948
rect 16594 52892 16604 52948
rect 16660 52892 19628 52948
rect 19684 52892 19694 52948
rect 28018 52892 28028 52948
rect 28084 52892 29148 52948
rect 29204 52892 29214 52948
rect 40786 52892 40796 52948
rect 40852 52892 41692 52948
rect 41748 52892 42140 52948
rect 42196 52892 43484 52948
rect 43540 52892 43550 52948
rect 48514 52892 48524 52948
rect 48580 52892 48972 52948
rect 49028 52892 49756 52948
rect 49812 52892 49822 52948
rect 5170 52780 5180 52836
rect 5236 52780 6188 52836
rect 6244 52780 6860 52836
rect 6916 52780 6926 52836
rect 18722 52780 18732 52836
rect 18788 52780 19404 52836
rect 19460 52780 19470 52836
rect 28802 52780 28812 52836
rect 28868 52780 30268 52836
rect 30324 52780 30334 52836
rect 39442 52780 39452 52836
rect 39508 52780 42364 52836
rect 42420 52780 42430 52836
rect 48178 52780 48188 52836
rect 48244 52780 48860 52836
rect 48916 52780 48926 52836
rect 50754 52780 50764 52836
rect 50820 52780 53004 52836
rect 53060 52780 53070 52836
rect 2482 52668 2492 52724
rect 2548 52668 5516 52724
rect 5572 52668 5582 52724
rect 23426 52668 23436 52724
rect 23492 52668 24220 52724
rect 24276 52668 24286 52724
rect 24546 52668 24556 52724
rect 24612 52668 26908 52724
rect 26964 52668 26974 52724
rect 27906 52668 27916 52724
rect 27972 52668 29820 52724
rect 29876 52668 31276 52724
rect 31332 52668 31342 52724
rect 21858 52556 21868 52612
rect 21924 52556 23884 52612
rect 23940 52556 24892 52612
rect 24948 52556 34300 52612
rect 34356 52556 34366 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 27458 52444 27468 52500
rect 27524 52444 28924 52500
rect 28980 52444 28990 52500
rect 48290 52444 48300 52500
rect 48356 52444 48748 52500
rect 48804 52444 51548 52500
rect 51604 52444 51614 52500
rect 3714 52332 3724 52388
rect 3780 52332 5180 52388
rect 5236 52332 5740 52388
rect 5796 52332 5806 52388
rect 11666 52332 11676 52388
rect 11732 52332 11742 52388
rect 15810 52332 15820 52388
rect 15876 52332 16268 52388
rect 16324 52332 16334 52388
rect 17490 52332 17500 52388
rect 17556 52332 18284 52388
rect 18340 52332 18350 52388
rect 28130 52332 28140 52388
rect 28196 52332 30044 52388
rect 30100 52332 30110 52388
rect 50866 52332 50876 52388
rect 50932 52332 50942 52388
rect 4834 52220 4844 52276
rect 4900 52220 5628 52276
rect 5684 52220 5694 52276
rect 4610 52108 4620 52164
rect 4676 52108 5852 52164
rect 5908 52108 7868 52164
rect 7924 52108 7934 52164
rect 11676 52052 11732 52332
rect 18498 52220 18508 52276
rect 18564 52220 21980 52276
rect 22036 52220 22046 52276
rect 27458 52220 27468 52276
rect 27524 52220 28588 52276
rect 28644 52220 28654 52276
rect 28914 52220 28924 52276
rect 28980 52220 33292 52276
rect 33348 52220 34076 52276
rect 34132 52220 34142 52276
rect 34962 52220 34972 52276
rect 35028 52220 35644 52276
rect 35700 52220 35710 52276
rect 38882 52220 38892 52276
rect 38948 52220 40796 52276
rect 40852 52220 40862 52276
rect 17042 52108 17052 52164
rect 17108 52108 17612 52164
rect 17668 52108 17678 52164
rect 19730 52108 19740 52164
rect 19796 52108 21532 52164
rect 21588 52108 21598 52164
rect 23202 52108 23212 52164
rect 23268 52108 24444 52164
rect 24500 52108 24510 52164
rect 26114 52108 26124 52164
rect 26180 52108 27132 52164
rect 27188 52108 27198 52164
rect 27794 52108 27804 52164
rect 27860 52108 29148 52164
rect 29204 52108 29214 52164
rect 33394 52108 33404 52164
rect 33460 52108 33852 52164
rect 33908 52108 33918 52164
rect 37874 52108 37884 52164
rect 37940 52108 42140 52164
rect 42196 52108 42206 52164
rect 42354 52108 42364 52164
rect 42420 52108 42924 52164
rect 42980 52108 42990 52164
rect 43138 52108 43148 52164
rect 43204 52108 44940 52164
rect 44996 52108 45006 52164
rect 46834 52108 46844 52164
rect 46900 52108 48076 52164
rect 48132 52108 49308 52164
rect 49364 52108 49374 52164
rect 50876 52052 50932 52332
rect 51874 52220 51884 52276
rect 51940 52220 52780 52276
rect 52836 52220 52846 52276
rect 11442 51996 11452 52052
rect 11508 51996 11900 52052
rect 11956 51996 11966 52052
rect 15474 51996 15484 52052
rect 15540 51996 16604 52052
rect 16660 51996 17948 52052
rect 18004 51996 18014 52052
rect 23650 51996 23660 52052
rect 23716 51996 24668 52052
rect 24724 51996 24734 52052
rect 39666 51996 39676 52052
rect 39732 51996 40348 52052
rect 40404 51996 41076 52052
rect 49746 51996 49756 52052
rect 49812 51996 49868 52052
rect 49924 51996 51436 52052
rect 51492 51996 51996 52052
rect 52052 51996 52062 52052
rect 41020 51940 41076 51996
rect 16930 51884 16940 51940
rect 16996 51884 18396 51940
rect 18452 51884 18462 51940
rect 23314 51884 23324 51940
rect 23380 51884 23772 51940
rect 23828 51884 23838 51940
rect 32274 51884 32284 51940
rect 32340 51884 33180 51940
rect 33236 51884 33246 51940
rect 41010 51884 41020 51940
rect 41076 51884 41086 51940
rect 42130 51884 42140 51940
rect 42196 51884 43260 51940
rect 43316 51884 43326 51940
rect 26338 51772 26348 51828
rect 26404 51772 26908 51828
rect 38098 51772 38108 51828
rect 38164 51772 39116 51828
rect 39172 51772 41580 51828
rect 41636 51772 47180 51828
rect 47236 51772 47246 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 26450 51660 26460 51716
rect 26516 51660 26526 51716
rect 9650 51548 9660 51604
rect 9716 51548 11004 51604
rect 11060 51548 11070 51604
rect 11330 51548 11340 51604
rect 11396 51548 12348 51604
rect 12404 51548 12414 51604
rect 18274 51548 18284 51604
rect 18340 51548 19292 51604
rect 19348 51548 21756 51604
rect 21812 51548 22540 51604
rect 22596 51548 22606 51604
rect 16156 51436 16716 51492
rect 16772 51436 18060 51492
rect 18116 51436 23884 51492
rect 23940 51436 23950 51492
rect 16156 51380 16212 51436
rect 26460 51380 26516 51660
rect 26852 51492 26908 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 37090 51660 37100 51716
rect 37156 51660 38668 51716
rect 38724 51660 41860 51716
rect 44034 51660 44044 51716
rect 44100 51660 45276 51716
rect 45332 51660 47404 51716
rect 47460 51660 47470 51716
rect 41804 51604 41860 51660
rect 28914 51548 28924 51604
rect 28980 51548 29708 51604
rect 29764 51548 30604 51604
rect 30660 51548 33852 51604
rect 33908 51548 33918 51604
rect 40114 51548 40124 51604
rect 40180 51548 40908 51604
rect 40964 51548 40974 51604
rect 41794 51548 41804 51604
rect 41860 51548 45780 51604
rect 47954 51548 47964 51604
rect 48020 51548 48748 51604
rect 48804 51548 48814 51604
rect 26852 51436 28700 51492
rect 28756 51436 28766 51492
rect 38098 51436 38108 51492
rect 38164 51436 43708 51492
rect 43764 51436 43774 51492
rect 45724 51380 45780 51548
rect 48850 51436 48860 51492
rect 48916 51436 51660 51492
rect 51716 51436 51726 51492
rect 5394 51324 5404 51380
rect 5460 51324 6076 51380
rect 6132 51324 8876 51380
rect 8932 51324 9772 51380
rect 9828 51324 9838 51380
rect 10210 51324 10220 51380
rect 10276 51324 11340 51380
rect 11396 51324 11406 51380
rect 13122 51324 13132 51380
rect 13188 51324 15148 51380
rect 15204 51324 15932 51380
rect 15988 51324 15998 51380
rect 16146 51324 16156 51380
rect 16212 51324 16222 51380
rect 22642 51324 22652 51380
rect 22708 51324 25564 51380
rect 25620 51324 25630 51380
rect 26460 51324 27132 51380
rect 27188 51324 27916 51380
rect 27972 51324 27982 51380
rect 35074 51324 35084 51380
rect 35140 51324 35868 51380
rect 35924 51324 37436 51380
rect 37492 51324 37502 51380
rect 40226 51324 40236 51380
rect 40292 51324 40460 51380
rect 40516 51324 40526 51380
rect 42130 51324 42140 51380
rect 42196 51324 42700 51380
rect 42756 51324 43260 51380
rect 43316 51324 45276 51380
rect 45332 51324 45342 51380
rect 45714 51324 45724 51380
rect 45780 51324 46508 51380
rect 46564 51324 46574 51380
rect 47730 51324 47740 51380
rect 47796 51324 50428 51380
rect 50754 51324 50764 51380
rect 50820 51324 51884 51380
rect 51940 51324 51950 51380
rect 50372 51268 50428 51324
rect 19170 51212 19180 51268
rect 19236 51212 19964 51268
rect 20020 51212 20030 51268
rect 22978 51212 22988 51268
rect 23044 51212 23772 51268
rect 23828 51212 23838 51268
rect 29586 51212 29596 51268
rect 29652 51212 30268 51268
rect 30324 51212 30334 51268
rect 41794 51212 41804 51268
rect 41860 51212 42588 51268
rect 42644 51212 42654 51268
rect 50372 51212 50876 51268
rect 50932 51212 52780 51268
rect 52836 51212 53340 51268
rect 53396 51212 53406 51268
rect 6962 51100 6972 51156
rect 7028 51100 8428 51156
rect 8484 51100 8494 51156
rect 25554 51100 25564 51156
rect 25620 51100 27468 51156
rect 27524 51100 27534 51156
rect 36530 51100 36540 51156
rect 36596 51100 37660 51156
rect 37716 51100 37726 51156
rect 38546 51100 38556 51156
rect 38612 51100 53004 51156
rect 53060 51100 53900 51156
rect 53956 51100 54460 51156
rect 54516 51100 54526 51156
rect 41906 50988 41916 51044
rect 41972 50988 43932 51044
rect 43988 50988 43998 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 19954 50876 19964 50932
rect 20020 50876 22092 50932
rect 22148 50876 23324 50932
rect 23380 50876 23390 50932
rect 10434 50764 10444 50820
rect 10500 50764 11340 50820
rect 11396 50764 11406 50820
rect 27458 50764 27468 50820
rect 27524 50764 28140 50820
rect 28196 50764 28206 50820
rect 30258 50764 30268 50820
rect 30324 50764 31948 50820
rect 32004 50764 33404 50820
rect 33460 50764 33470 50820
rect 40012 50764 41020 50820
rect 41076 50764 44044 50820
rect 44100 50764 44110 50820
rect 40012 50708 40068 50764
rect 9874 50652 9884 50708
rect 9940 50652 11228 50708
rect 11284 50652 12572 50708
rect 12628 50652 12638 50708
rect 15922 50652 15932 50708
rect 15988 50652 18172 50708
rect 18228 50652 18238 50708
rect 21522 50652 21532 50708
rect 21588 50652 24668 50708
rect 24724 50652 24734 50708
rect 28466 50652 28476 50708
rect 28532 50652 29932 50708
rect 29988 50652 31276 50708
rect 31332 50652 31342 50708
rect 31826 50652 31836 50708
rect 31892 50652 33068 50708
rect 33124 50652 33134 50708
rect 40002 50652 40012 50708
rect 40068 50652 40078 50708
rect 40348 50652 41692 50708
rect 41748 50652 41758 50708
rect 42578 50652 42588 50708
rect 42644 50652 44156 50708
rect 44212 50652 44222 50708
rect 40348 50596 40404 50652
rect 10882 50540 10892 50596
rect 10948 50540 11900 50596
rect 11956 50540 11966 50596
rect 18946 50540 18956 50596
rect 19012 50540 22652 50596
rect 22708 50540 22718 50596
rect 23650 50540 23660 50596
rect 23716 50540 24108 50596
rect 24164 50540 24174 50596
rect 24332 50540 24444 50596
rect 24500 50540 24510 50596
rect 26786 50540 26796 50596
rect 26852 50540 27692 50596
rect 27748 50540 28252 50596
rect 28308 50540 28318 50596
rect 28802 50540 28812 50596
rect 28868 50540 32172 50596
rect 32228 50540 32238 50596
rect 40114 50540 40124 50596
rect 40180 50540 40404 50596
rect 41234 50540 41244 50596
rect 41300 50540 42476 50596
rect 42532 50540 42542 50596
rect 46834 50540 46844 50596
rect 46900 50540 47180 50596
rect 47236 50540 47246 50596
rect 49046 50540 49084 50596
rect 49140 50540 49150 50596
rect 52770 50540 52780 50596
rect 52836 50540 54460 50596
rect 54516 50540 54526 50596
rect 24332 50484 24388 50540
rect 5730 50428 5740 50484
rect 5796 50428 6860 50484
rect 6916 50428 6926 50484
rect 10098 50428 10108 50484
rect 10164 50428 10780 50484
rect 10836 50428 10846 50484
rect 11442 50428 11452 50484
rect 11508 50428 12460 50484
rect 12516 50428 12526 50484
rect 16706 50428 16716 50484
rect 16772 50428 17388 50484
rect 17444 50428 17454 50484
rect 18834 50428 18844 50484
rect 18900 50428 19516 50484
rect 19572 50428 19582 50484
rect 22418 50428 22428 50484
rect 22484 50428 23772 50484
rect 23828 50428 24388 50484
rect 24546 50428 24556 50484
rect 24612 50428 26236 50484
rect 26292 50428 27132 50484
rect 27188 50428 27198 50484
rect 29810 50428 29820 50484
rect 29876 50428 30492 50484
rect 30548 50428 30558 50484
rect 33282 50428 33292 50484
rect 33348 50428 34300 50484
rect 34356 50428 34366 50484
rect 36306 50428 36316 50484
rect 36372 50428 37548 50484
rect 37604 50428 38444 50484
rect 38500 50428 38510 50484
rect 40338 50428 40348 50484
rect 40404 50428 40796 50484
rect 40852 50428 40862 50484
rect 41346 50428 41356 50484
rect 41412 50428 42420 50484
rect 42364 50372 42420 50428
rect 42812 50428 43820 50484
rect 43876 50428 43886 50484
rect 46386 50428 46396 50484
rect 46452 50428 49532 50484
rect 49588 50428 49868 50484
rect 49924 50428 49934 50484
rect 50082 50428 50092 50484
rect 50148 50428 50186 50484
rect 50866 50428 50876 50484
rect 50932 50428 51772 50484
rect 51828 50428 56140 50484
rect 56196 50428 56206 50484
rect 42812 50372 42868 50428
rect 13906 50316 13916 50372
rect 13972 50316 16380 50372
rect 16436 50316 16446 50372
rect 19618 50316 19628 50372
rect 19684 50316 20412 50372
rect 20468 50316 20478 50372
rect 27346 50316 27356 50372
rect 27412 50316 28364 50372
rect 28420 50316 28430 50372
rect 31826 50316 31836 50372
rect 31892 50316 32508 50372
rect 32564 50316 32574 50372
rect 33170 50316 33180 50372
rect 33236 50316 33246 50372
rect 42364 50316 42868 50372
rect 46610 50316 46620 50372
rect 46676 50316 47180 50372
rect 47236 50316 49084 50372
rect 49140 50316 49150 50372
rect 49410 50316 49420 50372
rect 49476 50316 49980 50372
rect 50036 50316 50046 50372
rect 51874 50316 51884 50372
rect 51940 50316 53340 50372
rect 53396 50316 53406 50372
rect 33180 50260 33236 50316
rect 32274 50204 32284 50260
rect 32340 50204 33236 50260
rect 37874 50204 37884 50260
rect 37940 50204 40012 50260
rect 40068 50204 42812 50260
rect 42868 50204 43596 50260
rect 43652 50204 43662 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 5842 50092 5852 50148
rect 5908 50092 7644 50148
rect 7700 50092 7710 50148
rect 31378 50092 31388 50148
rect 31444 50092 32396 50148
rect 32452 50092 32462 50148
rect 41682 50092 41692 50148
rect 41748 50092 42364 50148
rect 42420 50092 42430 50148
rect 49270 50092 49308 50148
rect 49364 50092 49374 50148
rect 2034 49980 2044 50036
rect 2100 49980 2716 50036
rect 2772 49980 2782 50036
rect 6290 49980 6300 50036
rect 6356 49980 9548 50036
rect 9604 49980 9614 50036
rect 29362 49980 29372 50036
rect 29428 49980 29932 50036
rect 29988 49980 29998 50036
rect 25442 49868 25452 49924
rect 25508 49868 26684 49924
rect 26740 49868 27580 49924
rect 27636 49868 27646 49924
rect 28018 49868 28028 49924
rect 28084 49868 31164 49924
rect 31220 49868 31612 49924
rect 31668 49868 32284 49924
rect 32340 49868 32350 49924
rect 44930 49868 44940 49924
rect 44996 49868 48076 49924
rect 48132 49868 49588 49924
rect 50194 49868 50204 49924
rect 50260 49868 51100 49924
rect 51156 49868 51166 49924
rect 49532 49812 49588 49868
rect 3490 49756 3500 49812
rect 3556 49756 4620 49812
rect 4676 49756 5964 49812
rect 6020 49756 6412 49812
rect 6468 49756 6972 49812
rect 7028 49756 7038 49812
rect 7186 49756 7196 49812
rect 7252 49756 8204 49812
rect 8260 49756 8270 49812
rect 10658 49756 10668 49812
rect 10724 49756 11564 49812
rect 11620 49756 11630 49812
rect 11890 49756 11900 49812
rect 11956 49756 12460 49812
rect 12516 49756 12526 49812
rect 16818 49756 16828 49812
rect 16884 49756 17724 49812
rect 17780 49756 18956 49812
rect 19012 49756 20636 49812
rect 20692 49756 20702 49812
rect 26786 49756 26796 49812
rect 26852 49756 28140 49812
rect 28196 49756 28924 49812
rect 28980 49756 28990 49812
rect 29362 49756 29372 49812
rect 29428 49756 29438 49812
rect 30342 49756 30380 49812
rect 30436 49756 30446 49812
rect 30706 49756 30716 49812
rect 30772 49756 31836 49812
rect 31892 49756 31902 49812
rect 7196 49700 7252 49756
rect 6178 49644 6188 49700
rect 6244 49644 7252 49700
rect 12338 49644 12348 49700
rect 12404 49644 12684 49700
rect 12740 49644 12750 49700
rect 29372 49588 29428 49756
rect 38612 49700 38668 49812
rect 38724 49756 38734 49812
rect 40114 49756 40124 49812
rect 40180 49756 41804 49812
rect 41860 49756 42476 49812
rect 42532 49756 42542 49812
rect 46274 49756 46284 49812
rect 46340 49756 46956 49812
rect 47012 49756 47022 49812
rect 47954 49756 47964 49812
rect 48020 49756 49308 49812
rect 49364 49756 49374 49812
rect 49532 49756 50764 49812
rect 50820 49756 50830 49812
rect 53106 49756 53116 49812
rect 53172 49756 53788 49812
rect 53844 49756 53854 49812
rect 55234 49756 55244 49812
rect 55300 49756 56476 49812
rect 56532 49756 56542 49812
rect 30034 49644 30044 49700
rect 30100 49644 31052 49700
rect 31108 49644 32172 49700
rect 32228 49644 32238 49700
rect 32722 49644 32732 49700
rect 32788 49644 34188 49700
rect 34244 49644 34254 49700
rect 36642 49644 36652 49700
rect 36708 49644 38668 49700
rect 45826 49644 45836 49700
rect 45892 49644 48412 49700
rect 48468 49644 48478 49700
rect 48626 49644 48636 49700
rect 48692 49644 49084 49700
rect 49140 49644 50092 49700
rect 50148 49644 50158 49700
rect 52770 49644 52780 49700
rect 52836 49644 54684 49700
rect 54740 49644 54750 49700
rect 11218 49532 11228 49588
rect 11284 49532 11788 49588
rect 11844 49532 11854 49588
rect 17042 49532 17052 49588
rect 17108 49532 18620 49588
rect 18676 49532 18732 49588
rect 18788 49532 18798 49588
rect 19058 49532 19068 49588
rect 19124 49532 19964 49588
rect 20020 49532 20030 49588
rect 25330 49532 25340 49588
rect 25396 49532 27356 49588
rect 27412 49532 27422 49588
rect 27794 49532 27804 49588
rect 27860 49532 31164 49588
rect 31220 49532 31230 49588
rect 36306 49532 36316 49588
rect 36372 49532 36764 49588
rect 36820 49532 36830 49588
rect 47282 49532 47292 49588
rect 47348 49532 49084 49588
rect 49140 49532 50204 49588
rect 50260 49532 50270 49588
rect 16594 49420 16604 49476
rect 16660 49420 17164 49476
rect 17220 49420 17948 49476
rect 18004 49420 23660 49476
rect 23716 49420 23726 49476
rect 26562 49420 26572 49476
rect 26628 49420 28812 49476
rect 28868 49420 28878 49476
rect 29586 49420 29596 49476
rect 29652 49420 31052 49476
rect 31108 49420 31724 49476
rect 31780 49420 32060 49476
rect 32116 49420 32126 49476
rect 45490 49420 45500 49476
rect 45556 49420 46172 49476
rect 46228 49420 46238 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 12002 49308 12012 49364
rect 12068 49308 12796 49364
rect 12852 49308 12862 49364
rect 18694 49308 18732 49364
rect 18788 49308 18798 49364
rect 19142 49308 19180 49364
rect 19236 49308 19246 49364
rect 20066 49308 20076 49364
rect 20132 49308 20524 49364
rect 20580 49308 20590 49364
rect 21298 49308 21308 49364
rect 21364 49308 21868 49364
rect 21924 49308 21934 49364
rect 27346 49308 27356 49364
rect 27412 49308 28700 49364
rect 28756 49308 28766 49364
rect 29026 49308 29036 49364
rect 29092 49308 31276 49364
rect 31332 49308 31612 49364
rect 31668 49308 31678 49364
rect 43810 49308 43820 49364
rect 43876 49308 45724 49364
rect 45780 49308 51660 49364
rect 51716 49308 52668 49364
rect 52724 49308 52734 49364
rect 2706 49196 2716 49252
rect 2772 49196 3500 49252
rect 3556 49196 3566 49252
rect 11666 49196 11676 49252
rect 11732 49196 11742 49252
rect 20178 49196 20188 49252
rect 20244 49196 20254 49252
rect 21634 49196 21644 49252
rect 21700 49196 22092 49252
rect 22148 49196 22158 49252
rect 26562 49196 26572 49252
rect 26628 49196 27132 49252
rect 27188 49196 27198 49252
rect 28354 49196 28364 49252
rect 28420 49196 29260 49252
rect 29316 49196 29326 49252
rect 30258 49196 30268 49252
rect 30324 49196 30940 49252
rect 30996 49196 31006 49252
rect 44828 49196 46844 49252
rect 46900 49196 48748 49252
rect 48804 49196 50092 49252
rect 50148 49196 50158 49252
rect 50754 49196 50764 49252
rect 50820 49196 53452 49252
rect 53508 49196 53518 49252
rect 11676 49140 11732 49196
rect 20188 49140 20244 49196
rect 44828 49140 44884 49196
rect 10098 49084 10108 49140
rect 10164 49084 10332 49140
rect 10388 49084 11732 49140
rect 19058 49084 19068 49140
rect 19124 49084 20244 49140
rect 26852 49084 27524 49140
rect 28578 49084 28588 49140
rect 28644 49084 29148 49140
rect 29204 49084 30660 49140
rect 30818 49084 30828 49140
rect 30884 49084 30940 49140
rect 30996 49084 31006 49140
rect 42578 49084 42588 49140
rect 42644 49084 44828 49140
rect 44884 49084 44894 49140
rect 45826 49084 45836 49140
rect 45892 49084 46732 49140
rect 46788 49084 46798 49140
rect 51538 49084 51548 49140
rect 51604 49084 51996 49140
rect 52052 49084 57484 49140
rect 57540 49084 57550 49140
rect 26852 49028 26908 49084
rect 27468 49028 27524 49084
rect 4722 48972 4732 49028
rect 4788 48972 7084 49028
rect 7140 48972 7150 49028
rect 8978 48972 8988 49028
rect 9044 48972 9996 49028
rect 10052 48972 11228 49028
rect 11284 48972 11294 49028
rect 18582 48972 18620 49028
rect 18676 48972 18686 49028
rect 19618 48972 19628 49028
rect 19684 48972 20860 49028
rect 20916 48972 21420 49028
rect 21476 48972 21868 49028
rect 21924 48972 21934 49028
rect 26226 48972 26236 49028
rect 26292 48972 26908 49028
rect 27458 48972 27468 49028
rect 27524 48972 27534 49028
rect 28242 48972 28252 49028
rect 28308 48972 29372 49028
rect 29428 48972 29438 49028
rect 28252 48916 28308 48972
rect 2930 48860 2940 48916
rect 2996 48860 3388 48916
rect 3444 48860 4396 48916
rect 4452 48860 5628 48916
rect 5684 48860 5694 48916
rect 11106 48860 11116 48916
rect 11172 48860 11900 48916
rect 11956 48860 12796 48916
rect 12852 48860 12862 48916
rect 17266 48860 17276 48916
rect 17332 48860 18508 48916
rect 18564 48860 18574 48916
rect 20514 48860 20524 48916
rect 20580 48860 21532 48916
rect 21588 48860 21598 48916
rect 23986 48860 23996 48916
rect 24052 48860 26124 48916
rect 26180 48860 26190 48916
rect 26898 48860 26908 48916
rect 26964 48860 28308 48916
rect 28802 48860 28812 48916
rect 28868 48860 29540 48916
rect 29484 48804 29540 48860
rect 30604 48804 30660 49084
rect 31602 48972 31612 49028
rect 31668 48972 32732 49028
rect 32788 48972 32798 49028
rect 39666 48972 39676 49028
rect 39732 48972 40012 49028
rect 40068 48972 41916 49028
rect 41972 48972 41982 49028
rect 43922 48972 43932 49028
rect 43988 48972 45276 49028
rect 45332 48972 46284 49028
rect 46340 48972 46676 49028
rect 48066 48972 48076 49028
rect 48132 48972 50540 49028
rect 50596 48972 50606 49028
rect 52098 48972 52108 49028
rect 52164 48972 52780 49028
rect 52836 48972 53004 49028
rect 53060 48972 53070 49028
rect 46620 48916 46676 48972
rect 36306 48860 36316 48916
rect 36372 48860 37324 48916
rect 37380 48860 37390 48916
rect 43810 48860 43820 48916
rect 43876 48860 46172 48916
rect 46228 48860 46238 48916
rect 46620 48860 46956 48916
rect 47012 48860 50428 48916
rect 50484 48860 50494 48916
rect 50764 48860 52332 48916
rect 52388 48860 52398 48916
rect 53330 48860 53340 48916
rect 53396 48860 54572 48916
rect 54628 48860 54638 48916
rect 50764 48804 50820 48860
rect 17826 48748 17836 48804
rect 17892 48748 20412 48804
rect 20468 48748 21084 48804
rect 21140 48748 21150 48804
rect 27234 48748 27244 48804
rect 27300 48748 28476 48804
rect 28532 48748 29260 48804
rect 29316 48748 29326 48804
rect 29484 48748 29708 48804
rect 29764 48748 29774 48804
rect 30594 48748 30604 48804
rect 30660 48748 30670 48804
rect 44370 48748 44380 48804
rect 44436 48748 45276 48804
rect 45332 48748 46060 48804
rect 46116 48748 46126 48804
rect 49858 48748 49868 48804
rect 49924 48748 50820 48804
rect 20738 48636 20748 48692
rect 20804 48636 21756 48692
rect 21812 48636 21822 48692
rect 30146 48636 30156 48692
rect 30212 48636 30828 48692
rect 30884 48636 30894 48692
rect 49074 48636 49084 48692
rect 49140 48636 49308 48692
rect 49364 48636 49374 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 20748 48468 20804 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 49308 48524 50204 48580
rect 50260 48524 50270 48580
rect 49308 48468 49364 48524
rect 3826 48412 3836 48468
rect 3892 48412 6972 48468
rect 7028 48412 7038 48468
rect 19730 48412 19740 48468
rect 19796 48412 20804 48468
rect 20962 48412 20972 48468
rect 21028 48412 22540 48468
rect 22596 48412 22606 48468
rect 27682 48412 27692 48468
rect 27748 48412 31052 48468
rect 31108 48412 31118 48468
rect 44370 48412 44380 48468
rect 44436 48412 45388 48468
rect 45444 48412 45454 48468
rect 45714 48412 45724 48468
rect 45780 48412 46844 48468
rect 46900 48412 48860 48468
rect 48916 48412 49308 48468
rect 49364 48412 49374 48468
rect 11554 48300 11564 48356
rect 11620 48300 13580 48356
rect 13636 48300 13646 48356
rect 15026 48300 15036 48356
rect 15092 48300 16044 48356
rect 16100 48300 16110 48356
rect 27010 48300 27020 48356
rect 27076 48300 27468 48356
rect 27524 48300 28252 48356
rect 28308 48300 28318 48356
rect 28578 48300 28588 48356
rect 28644 48300 30380 48356
rect 30436 48300 31948 48356
rect 32004 48300 32014 48356
rect 41458 48300 41468 48356
rect 41524 48300 41692 48356
rect 41748 48300 45052 48356
rect 45108 48300 48636 48356
rect 48692 48300 48702 48356
rect 48962 48300 48972 48356
rect 49028 48300 51548 48356
rect 51604 48300 51614 48356
rect 16146 48188 16156 48244
rect 16212 48188 17500 48244
rect 17556 48188 17566 48244
rect 29810 48188 29820 48244
rect 29876 48188 31612 48244
rect 31668 48188 31678 48244
rect 38546 48188 38556 48244
rect 38612 48188 39116 48244
rect 39172 48188 40908 48244
rect 40964 48188 40974 48244
rect 41906 48188 41916 48244
rect 41972 48188 42700 48244
rect 42756 48188 42766 48244
rect 44818 48188 44828 48244
rect 44884 48188 45164 48244
rect 45220 48188 45230 48244
rect 47170 48188 47180 48244
rect 47236 48188 51324 48244
rect 51380 48188 51390 48244
rect 52658 48188 52668 48244
rect 52724 48188 53564 48244
rect 53620 48188 53630 48244
rect 8866 48076 8876 48132
rect 8932 48076 9884 48132
rect 9940 48076 9950 48132
rect 32946 48076 32956 48132
rect 33012 48076 35644 48132
rect 35700 48076 37996 48132
rect 38052 48076 38062 48132
rect 48738 48076 48748 48132
rect 48804 48076 54124 48132
rect 54180 48076 56588 48132
rect 56644 48076 56654 48132
rect 37996 48020 38052 48076
rect 7746 47964 7756 48020
rect 7812 47964 9548 48020
rect 9604 47964 9614 48020
rect 37996 47964 38892 48020
rect 38948 47964 44380 48020
rect 44436 47964 44446 48020
rect 48178 47964 48188 48020
rect 48244 47964 49980 48020
rect 50036 47964 50046 48020
rect 50194 47964 50204 48020
rect 50260 47964 54012 48020
rect 54068 47964 54572 48020
rect 54628 47964 54638 48020
rect 6962 47852 6972 47908
rect 7028 47852 9660 47908
rect 9716 47852 10108 47908
rect 10164 47852 10174 47908
rect 50082 47852 50092 47908
rect 50148 47852 50428 47908
rect 50484 47852 50494 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 45490 47740 45500 47796
rect 45556 47740 50092 47796
rect 50148 47740 50158 47796
rect 20514 47628 20524 47684
rect 20580 47628 21420 47684
rect 21476 47628 22540 47684
rect 22596 47628 22606 47684
rect 48178 47628 48188 47684
rect 48244 47628 50652 47684
rect 50708 47628 50718 47684
rect 5730 47516 5740 47572
rect 5796 47516 6636 47572
rect 6692 47516 11228 47572
rect 11284 47516 11294 47572
rect 14802 47516 14812 47572
rect 14868 47516 15260 47572
rect 15316 47516 16604 47572
rect 16660 47516 19852 47572
rect 19908 47516 19918 47572
rect 42914 47516 42924 47572
rect 42980 47516 44156 47572
rect 44212 47516 44222 47572
rect 46162 47516 46172 47572
rect 46228 47516 47740 47572
rect 47796 47516 48748 47572
rect 48804 47516 48814 47572
rect 51986 47516 51996 47572
rect 52052 47516 52668 47572
rect 52724 47516 52734 47572
rect 53778 47516 53788 47572
rect 53844 47516 53854 47572
rect 53788 47460 53844 47516
rect 4946 47404 4956 47460
rect 5012 47404 5964 47460
rect 6020 47404 6030 47460
rect 8978 47404 8988 47460
rect 9044 47404 11004 47460
rect 11060 47404 12572 47460
rect 12628 47404 12638 47460
rect 16258 47404 16268 47460
rect 16324 47404 18620 47460
rect 18676 47404 21420 47460
rect 21476 47404 21486 47460
rect 36754 47404 36764 47460
rect 36820 47404 37100 47460
rect 37156 47404 37166 47460
rect 44258 47404 44268 47460
rect 44324 47404 44940 47460
rect 44996 47404 45006 47460
rect 48066 47404 48076 47460
rect 48132 47404 48972 47460
rect 49028 47404 49038 47460
rect 49718 47404 49756 47460
rect 49812 47404 49822 47460
rect 51874 47404 51884 47460
rect 51940 47404 53004 47460
rect 53060 47404 53844 47460
rect 3332 47292 5628 47348
rect 5684 47292 5694 47348
rect 19366 47292 19404 47348
rect 19460 47292 19470 47348
rect 20738 47292 20748 47348
rect 20804 47292 22316 47348
rect 22372 47292 25228 47348
rect 25284 47292 25294 47348
rect 40338 47292 40348 47348
rect 40404 47292 41020 47348
rect 41076 47292 41086 47348
rect 41794 47292 41804 47348
rect 41860 47292 42028 47348
rect 42084 47292 43708 47348
rect 43764 47292 44828 47348
rect 44884 47292 47068 47348
rect 47124 47292 47134 47348
rect 47954 47292 47964 47348
rect 48020 47292 49308 47348
rect 49364 47292 49374 47348
rect 49522 47292 49532 47348
rect 49588 47292 50092 47348
rect 50148 47292 50158 47348
rect 52770 47292 52780 47348
rect 52836 47292 53116 47348
rect 53172 47292 53788 47348
rect 53844 47292 53854 47348
rect 3332 47124 3388 47292
rect 11218 47180 11228 47236
rect 11284 47180 11788 47236
rect 11844 47180 11854 47236
rect 22978 47180 22988 47236
rect 23044 47180 32956 47236
rect 33012 47180 33022 47236
rect 45714 47180 45724 47236
rect 45780 47180 48860 47236
rect 48916 47180 48926 47236
rect 51426 47180 51436 47236
rect 51492 47180 53452 47236
rect 53508 47180 53518 47236
rect 2930 47068 2940 47124
rect 2996 47068 3388 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 22988 47012 23044 47180
rect 51090 47068 51100 47124
rect 51156 47068 51884 47124
rect 51940 47068 51950 47124
rect 52098 47068 52108 47124
rect 52164 47068 55468 47124
rect 55524 47068 55534 47124
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 8754 46956 8764 47012
rect 8820 46956 9884 47012
rect 9940 46956 9950 47012
rect 20402 46956 20412 47012
rect 20468 46956 23044 47012
rect 34178 46956 34188 47012
rect 34244 46956 37548 47012
rect 37604 46956 37614 47012
rect 37986 46956 37996 47012
rect 38052 46956 38892 47012
rect 38948 46956 38958 47012
rect 39788 46956 44604 47012
rect 44660 46956 44670 47012
rect 52546 46956 52556 47012
rect 52612 46956 53452 47012
rect 53508 46956 53518 47012
rect 53890 46956 53900 47012
rect 53956 46956 54796 47012
rect 54852 46956 54862 47012
rect 39788 46900 39844 46956
rect 10546 46844 10556 46900
rect 10612 46844 11900 46900
rect 11956 46844 12796 46900
rect 12852 46844 12862 46900
rect 33506 46844 33516 46900
rect 33572 46844 35532 46900
rect 35588 46844 36204 46900
rect 36260 46844 36270 46900
rect 36418 46844 36428 46900
rect 36484 46844 37100 46900
rect 37156 46844 37166 46900
rect 38322 46844 38332 46900
rect 38388 46844 39844 46900
rect 40002 46844 40012 46900
rect 40068 46844 42476 46900
rect 42532 46844 42542 46900
rect 44370 46844 44380 46900
rect 44436 46844 45612 46900
rect 45668 46844 46284 46900
rect 46340 46844 46350 46900
rect 46498 46844 46508 46900
rect 46564 46844 50428 46900
rect 5954 46732 5964 46788
rect 6020 46732 6860 46788
rect 6916 46732 8652 46788
rect 8708 46732 10668 46788
rect 10724 46732 10734 46788
rect 11666 46732 11676 46788
rect 11732 46732 14028 46788
rect 14084 46732 14094 46788
rect 21746 46732 21756 46788
rect 21812 46732 23660 46788
rect 23716 46732 23726 46788
rect 40012 46676 40068 46844
rect 50372 46788 50428 46844
rect 50372 46732 51660 46788
rect 51716 46732 51726 46788
rect 53218 46732 53228 46788
rect 53284 46732 54460 46788
rect 54516 46732 54526 46788
rect 4834 46620 4844 46676
rect 4900 46620 6300 46676
rect 6356 46620 7196 46676
rect 7252 46620 7644 46676
rect 7700 46620 7710 46676
rect 8418 46620 8428 46676
rect 8484 46620 10220 46676
rect 10276 46620 10286 46676
rect 17938 46620 17948 46676
rect 18004 46620 20412 46676
rect 20468 46620 20478 46676
rect 30146 46620 30156 46676
rect 30212 46620 30828 46676
rect 30884 46620 31388 46676
rect 31444 46620 31454 46676
rect 36194 46620 36204 46676
rect 36260 46620 36876 46676
rect 36932 46620 40068 46676
rect 40450 46620 40460 46676
rect 40516 46620 41804 46676
rect 41860 46620 41870 46676
rect 42354 46620 42364 46676
rect 42420 46620 42924 46676
rect 42980 46620 42990 46676
rect 50194 46620 50204 46676
rect 50260 46620 52220 46676
rect 52276 46620 52286 46676
rect 52434 46620 52444 46676
rect 52500 46620 53452 46676
rect 53508 46620 55356 46676
rect 55412 46620 55422 46676
rect 21298 46508 21308 46564
rect 21364 46508 24332 46564
rect 24388 46508 24398 46564
rect 25778 46508 25788 46564
rect 25844 46508 27356 46564
rect 27412 46508 27422 46564
rect 31042 46508 31052 46564
rect 31108 46508 32060 46564
rect 32116 46508 32126 46564
rect 37874 46508 37884 46564
rect 37940 46508 38780 46564
rect 38836 46508 38846 46564
rect 49858 46508 49868 46564
rect 49924 46508 50316 46564
rect 50372 46508 50764 46564
rect 50820 46508 50830 46564
rect 53554 46508 53564 46564
rect 53620 46508 53900 46564
rect 53956 46508 53966 46564
rect 4946 46396 4956 46452
rect 5012 46396 5740 46452
rect 5796 46396 5806 46452
rect 32386 46396 32396 46452
rect 32452 46396 37212 46452
rect 37268 46396 37278 46452
rect 37538 46396 37548 46452
rect 37604 46396 43820 46452
rect 43876 46396 43886 46452
rect 45602 46396 45612 46452
rect 45668 46396 49420 46452
rect 49476 46396 49486 46452
rect 50082 46396 50092 46452
rect 50148 46396 53228 46452
rect 53284 46396 53294 46452
rect 36418 46284 36428 46340
rect 36484 46284 37996 46340
rect 38052 46284 38062 46340
rect 40002 46284 40012 46340
rect 40068 46284 46396 46340
rect 46452 46284 46462 46340
rect 50530 46284 50540 46340
rect 50596 46284 50764 46340
rect 50820 46284 51324 46340
rect 51380 46284 51390 46340
rect 54114 46284 54124 46340
rect 54180 46284 54908 46340
rect 54964 46284 54974 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 36754 46172 36764 46228
rect 36820 46172 42140 46228
rect 42196 46172 42206 46228
rect 44594 46172 44604 46228
rect 44660 46172 45164 46228
rect 45220 46172 45230 46228
rect 47170 46172 47180 46228
rect 47236 46172 54460 46228
rect 54516 46172 57148 46228
rect 57204 46172 57214 46228
rect 5058 46060 5068 46116
rect 5124 46060 6076 46116
rect 6132 46060 6412 46116
rect 6468 46060 6478 46116
rect 11330 46060 11340 46116
rect 11396 46060 13356 46116
rect 13412 46060 13422 46116
rect 31714 46060 31724 46116
rect 31780 46060 36540 46116
rect 36596 46060 37548 46116
rect 37604 46060 37614 46116
rect 42242 46060 42252 46116
rect 42308 46060 46396 46116
rect 46452 46060 46462 46116
rect 2258 45948 2268 46004
rect 2324 45948 4396 46004
rect 4452 45948 6972 46004
rect 7028 45948 7038 46004
rect 16930 45948 16940 46004
rect 16996 45948 17612 46004
rect 17668 45948 17678 46004
rect 17826 45948 17836 46004
rect 17892 45948 27916 46004
rect 27972 45948 29820 46004
rect 29876 45948 29886 46004
rect 34738 45948 34748 46004
rect 34804 45948 35868 46004
rect 35924 45948 37324 46004
rect 37380 45948 37390 46004
rect 42914 45948 42924 46004
rect 42980 45948 43316 46004
rect 44258 45948 44268 46004
rect 44324 45948 45836 46004
rect 45892 45948 45902 46004
rect 48626 45948 48636 46004
rect 48692 45948 54908 46004
rect 54964 45948 54974 46004
rect 43260 45892 43316 45948
rect 31938 45836 31948 45892
rect 32004 45836 33180 45892
rect 33236 45836 33246 45892
rect 41794 45836 41804 45892
rect 41860 45836 43036 45892
rect 43092 45836 43102 45892
rect 43260 45836 45388 45892
rect 45444 45836 45454 45892
rect 47012 45836 50540 45892
rect 50596 45836 50606 45892
rect 50866 45836 50876 45892
rect 50932 45836 52668 45892
rect 52724 45836 52734 45892
rect 47012 45780 47068 45836
rect 8978 45724 8988 45780
rect 9044 45724 9660 45780
rect 9716 45724 9726 45780
rect 14802 45724 14812 45780
rect 14868 45724 15372 45780
rect 15428 45724 15438 45780
rect 19180 45724 20076 45780
rect 20132 45724 20142 45780
rect 37538 45724 37548 45780
rect 37604 45724 38108 45780
rect 38164 45724 39004 45780
rect 39060 45724 39070 45780
rect 41458 45724 41468 45780
rect 41524 45724 47068 45780
rect 52322 45724 52332 45780
rect 52388 45724 52398 45780
rect 54450 45724 54460 45780
rect 54516 45724 55692 45780
rect 55748 45724 55758 45780
rect 19180 45668 19236 45724
rect 52332 45668 52388 45724
rect 9090 45612 9100 45668
rect 9156 45612 13244 45668
rect 13300 45612 13310 45668
rect 19170 45612 19180 45668
rect 19236 45612 19246 45668
rect 19618 45612 19628 45668
rect 19684 45612 21196 45668
rect 21252 45612 21262 45668
rect 25778 45612 25788 45668
rect 25844 45612 26236 45668
rect 26292 45612 26684 45668
rect 26740 45612 28924 45668
rect 28980 45612 31052 45668
rect 31108 45612 31118 45668
rect 37090 45612 37100 45668
rect 37156 45612 37660 45668
rect 37716 45612 40012 45668
rect 40068 45612 40078 45668
rect 42130 45612 42140 45668
rect 42196 45612 43260 45668
rect 43316 45612 43326 45668
rect 43698 45612 43708 45668
rect 43764 45612 44268 45668
rect 44324 45612 44334 45668
rect 50372 45612 52388 45668
rect 41682 45500 41692 45556
rect 41748 45500 43932 45556
rect 43988 45500 43998 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50372 45444 50428 45612
rect 55682 45500 55692 45556
rect 55748 45500 57820 45556
rect 57876 45500 57886 45556
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 6962 45388 6972 45444
rect 7028 45388 8092 45444
rect 8148 45388 8764 45444
rect 8820 45388 9660 45444
rect 9716 45388 17948 45444
rect 18004 45388 18014 45444
rect 25330 45388 25340 45444
rect 25396 45388 26348 45444
rect 26404 45388 26414 45444
rect 39218 45388 39228 45444
rect 39284 45388 48748 45444
rect 48804 45388 49756 45444
rect 49812 45388 50428 45444
rect 7634 45276 7644 45332
rect 7700 45276 10556 45332
rect 10612 45276 10622 45332
rect 12786 45276 12796 45332
rect 12852 45276 32788 45332
rect 37986 45276 37996 45332
rect 38052 45276 38780 45332
rect 38836 45276 38846 45332
rect 43810 45276 43820 45332
rect 43876 45276 45164 45332
rect 45220 45276 46060 45332
rect 46116 45276 46126 45332
rect 47506 45276 47516 45332
rect 47572 45276 52444 45332
rect 52500 45276 52510 45332
rect 12796 45220 12852 45276
rect 8082 45164 8092 45220
rect 8148 45164 10220 45220
rect 10276 45164 12852 45220
rect 16258 45164 16268 45220
rect 16324 45164 17836 45220
rect 17892 45164 17902 45220
rect 19506 45164 19516 45220
rect 19572 45164 20860 45220
rect 20916 45164 20926 45220
rect 21746 45164 21756 45220
rect 21812 45164 23100 45220
rect 23156 45164 23166 45220
rect 14130 45052 14140 45108
rect 14196 45052 14588 45108
rect 14644 45052 16716 45108
rect 16772 45052 16782 45108
rect 29250 44940 29260 44996
rect 29316 44940 31388 44996
rect 31444 44940 31454 44996
rect 32732 44884 32788 45276
rect 38612 45164 39508 45220
rect 43362 45164 43372 45220
rect 43428 45164 44044 45220
rect 44100 45164 44996 45220
rect 45378 45164 45388 45220
rect 45444 45164 48524 45220
rect 48580 45164 48590 45220
rect 53778 45164 53788 45220
rect 53844 45164 55580 45220
rect 55636 45164 56588 45220
rect 56644 45164 56654 45220
rect 38612 45108 38668 45164
rect 34514 45052 34524 45108
rect 34580 45052 35308 45108
rect 35364 45052 35374 45108
rect 38434 45052 38444 45108
rect 38500 45052 38668 45108
rect 39452 44996 39508 45164
rect 44940 45108 44996 45164
rect 42242 45052 42252 45108
rect 42308 45052 44716 45108
rect 44772 45052 44782 45108
rect 44930 45052 44940 45108
rect 44996 45052 45006 45108
rect 50306 45052 50316 45108
rect 50372 45052 51100 45108
rect 51156 45052 51166 45108
rect 53554 45052 53564 45108
rect 53620 45052 54124 45108
rect 54180 45052 54190 45108
rect 54674 45052 54684 45108
rect 54740 45052 55132 45108
rect 55188 45052 55198 45108
rect 39442 44940 39452 44996
rect 39508 44940 40460 44996
rect 40516 44940 40526 44996
rect 44370 44940 44380 44996
rect 44436 44940 45276 44996
rect 45332 44940 45342 44996
rect 53666 44940 53676 44996
rect 53732 44940 55020 44996
rect 55076 44940 55086 44996
rect 20066 44828 20076 44884
rect 20132 44828 25676 44884
rect 25732 44828 25742 44884
rect 26002 44828 26012 44884
rect 26068 44828 27580 44884
rect 27636 44828 27646 44884
rect 32732 44828 38668 44884
rect 38994 44828 39004 44884
rect 39060 44828 41020 44884
rect 41076 44828 45500 44884
rect 45556 44828 45566 44884
rect 53106 44828 53116 44884
rect 53172 44828 54348 44884
rect 54404 44828 54414 44884
rect 38612 44772 38668 44828
rect 38612 44716 43036 44772
rect 43092 44716 45276 44772
rect 45332 44716 45342 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 36866 44604 36876 44660
rect 36932 44604 43708 44660
rect 43764 44604 43774 44660
rect 42242 44492 42252 44548
rect 42308 44492 43260 44548
rect 43316 44492 43326 44548
rect 49158 44492 49196 44548
rect 49252 44492 49262 44548
rect 7410 44380 7420 44436
rect 7476 44380 7980 44436
rect 8036 44380 12124 44436
rect 12180 44380 12190 44436
rect 13234 44380 13244 44436
rect 13300 44380 14812 44436
rect 14868 44380 15148 44436
rect 15204 44380 15214 44436
rect 18946 44380 18956 44436
rect 19012 44380 19516 44436
rect 19572 44380 19582 44436
rect 30370 44380 30380 44436
rect 30436 44380 38220 44436
rect 38276 44380 38286 44436
rect 7298 44268 7308 44324
rect 7364 44268 9548 44324
rect 9604 44268 9614 44324
rect 20402 44268 20412 44324
rect 20468 44268 24444 44324
rect 24500 44268 25452 44324
rect 25508 44268 25518 44324
rect 31378 44268 31388 44324
rect 31444 44268 32172 44324
rect 32228 44268 32238 44324
rect 32498 44268 32508 44324
rect 32564 44268 33292 44324
rect 33348 44268 33358 44324
rect 33954 44268 33964 44324
rect 34020 44268 35980 44324
rect 36036 44268 36046 44324
rect 37650 44268 37660 44324
rect 37716 44268 38668 44324
rect 38724 44268 38734 44324
rect 40002 44268 40012 44324
rect 40068 44268 40796 44324
rect 40852 44268 40862 44324
rect 53554 44268 53564 44324
rect 53620 44268 53900 44324
rect 53956 44268 56364 44324
rect 56420 44268 56430 44324
rect 7186 44156 7196 44212
rect 7252 44156 9772 44212
rect 9828 44156 9838 44212
rect 18162 44156 18172 44212
rect 18228 44156 19852 44212
rect 19908 44156 19918 44212
rect 21298 44156 21308 44212
rect 21364 44156 22092 44212
rect 22148 44156 22158 44212
rect 31042 44156 31052 44212
rect 31108 44156 34188 44212
rect 34244 44156 34254 44212
rect 35298 44156 35308 44212
rect 35364 44156 35644 44212
rect 35700 44156 35710 44212
rect 38434 44156 38444 44212
rect 38500 44156 38668 44212
rect 42466 44156 42476 44212
rect 42532 44156 43036 44212
rect 43092 44156 43102 44212
rect 44482 44156 44492 44212
rect 44548 44156 45724 44212
rect 45780 44156 45790 44212
rect 45938 44156 45948 44212
rect 46004 44156 48972 44212
rect 49028 44156 49038 44212
rect 49186 44156 49196 44212
rect 49252 44156 50204 44212
rect 50260 44156 50876 44212
rect 50932 44156 50942 44212
rect 51090 44156 51100 44212
rect 51156 44156 53004 44212
rect 53060 44156 53070 44212
rect 55010 44156 55020 44212
rect 55076 44156 55804 44212
rect 55860 44156 56588 44212
rect 56644 44156 57148 44212
rect 57204 44156 57214 44212
rect 38612 44100 38668 44156
rect 11666 44044 11676 44100
rect 11732 44044 12348 44100
rect 12404 44044 15484 44100
rect 15540 44044 15550 44100
rect 28690 44044 28700 44100
rect 28756 44044 29260 44100
rect 29316 44044 29326 44100
rect 33506 44044 33516 44100
rect 33572 44044 34636 44100
rect 34692 44044 36652 44100
rect 36708 44044 37548 44100
rect 37604 44044 37614 44100
rect 38612 44044 39116 44100
rect 39172 44044 39900 44100
rect 39956 44044 39966 44100
rect 40562 44044 40572 44100
rect 40628 44044 40638 44100
rect 50082 44044 50092 44100
rect 50148 44044 50764 44100
rect 50820 44044 50830 44100
rect 55346 44044 55356 44100
rect 55412 44044 57596 44100
rect 57652 44044 57662 44100
rect 7858 43932 7868 43988
rect 7924 43932 9436 43988
rect 9492 43932 10556 43988
rect 10612 43932 10622 43988
rect 16706 43932 16716 43988
rect 16772 43932 18060 43988
rect 18116 43932 19628 43988
rect 19684 43932 19694 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 40572 43876 40628 44044
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 39218 43820 39228 43876
rect 39284 43820 41244 43876
rect 41300 43820 41310 43876
rect 42914 43820 42924 43876
rect 42980 43820 42990 43876
rect 7634 43708 7644 43764
rect 7700 43708 10108 43764
rect 10164 43708 10174 43764
rect 21522 43708 21532 43764
rect 21588 43708 22988 43764
rect 23044 43708 23054 43764
rect 40450 43708 40460 43764
rect 40516 43708 41132 43764
rect 41188 43708 41198 43764
rect 42924 43652 42980 43820
rect 45266 43708 45276 43764
rect 45332 43708 50316 43764
rect 50372 43708 51436 43764
rect 51492 43708 51502 43764
rect 11442 43596 11452 43652
rect 11508 43596 17052 43652
rect 17108 43596 17118 43652
rect 17826 43596 17836 43652
rect 17892 43596 18396 43652
rect 18452 43596 18462 43652
rect 21186 43596 21196 43652
rect 21252 43596 24108 43652
rect 24164 43596 24174 43652
rect 26852 43596 27244 43652
rect 27300 43596 28700 43652
rect 28756 43596 28766 43652
rect 30482 43596 30492 43652
rect 30548 43596 31948 43652
rect 32004 43596 32014 43652
rect 34738 43596 34748 43652
rect 34804 43596 35644 43652
rect 35700 43596 35710 43652
rect 38994 43596 39004 43652
rect 39060 43596 39788 43652
rect 39844 43596 39854 43652
rect 42476 43596 42980 43652
rect 46162 43596 46172 43652
rect 46228 43596 47292 43652
rect 47348 43596 47358 43652
rect 49158 43596 49196 43652
rect 49252 43596 53116 43652
rect 53172 43596 54348 43652
rect 54404 43596 54414 43652
rect 56018 43596 56028 43652
rect 56084 43596 56252 43652
rect 56308 43596 57036 43652
rect 57092 43596 57102 43652
rect 26852 43540 26908 43596
rect 42476 43540 42532 43596
rect 22418 43484 22428 43540
rect 22484 43484 23324 43540
rect 23380 43484 26908 43540
rect 27122 43484 27132 43540
rect 27188 43484 28588 43540
rect 28644 43484 28654 43540
rect 32834 43484 32844 43540
rect 32900 43484 33628 43540
rect 33684 43484 34412 43540
rect 34468 43484 34478 43540
rect 34850 43484 34860 43540
rect 34916 43484 36092 43540
rect 36148 43484 36158 43540
rect 36866 43484 36876 43540
rect 36932 43484 42476 43540
rect 42532 43484 42542 43540
rect 42802 43484 42812 43540
rect 42868 43484 43484 43540
rect 43540 43484 43550 43540
rect 44370 43484 44380 43540
rect 44436 43484 45836 43540
rect 45892 43484 47628 43540
rect 47684 43484 47694 43540
rect 48178 43484 48188 43540
rect 48244 43484 49084 43540
rect 49140 43484 49150 43540
rect 49410 43484 49420 43540
rect 49476 43484 49486 43540
rect 49634 43484 49644 43540
rect 49700 43484 55468 43540
rect 55524 43484 56588 43540
rect 56644 43484 56654 43540
rect 49420 43428 49476 43484
rect 22642 43372 22652 43428
rect 22708 43372 23884 43428
rect 23940 43372 23950 43428
rect 35298 43372 35308 43428
rect 35364 43372 39340 43428
rect 39396 43372 39406 43428
rect 49420 43372 51324 43428
rect 51380 43372 51390 43428
rect 54898 43372 54908 43428
rect 54964 43372 56812 43428
rect 56868 43372 56878 43428
rect 20402 43260 20412 43316
rect 20468 43260 24780 43316
rect 24836 43260 24846 43316
rect 35410 43260 35420 43316
rect 35476 43260 36204 43316
rect 36260 43260 36270 43316
rect 46498 43260 46508 43316
rect 46564 43260 47404 43316
rect 47460 43260 49868 43316
rect 49924 43260 49934 43316
rect 50866 43260 50876 43316
rect 50932 43260 51436 43316
rect 51492 43260 51502 43316
rect 53890 43260 53900 43316
rect 53956 43260 55692 43316
rect 55748 43260 55758 43316
rect 40198 43148 40236 43204
rect 40292 43148 40302 43204
rect 45154 43148 45164 43204
rect 45220 43148 51548 43204
rect 51604 43148 52108 43204
rect 52164 43148 52174 43204
rect 53666 43148 53676 43204
rect 53732 43148 54460 43204
rect 54516 43148 54526 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 51314 43036 51324 43092
rect 51380 43036 53564 43092
rect 53620 43036 53630 43092
rect 16706 42924 16716 42980
rect 16772 42924 18060 42980
rect 18116 42924 18126 42980
rect 34626 42924 34636 42980
rect 34692 42924 36540 42980
rect 36596 42924 36606 42980
rect 43558 42924 43596 42980
rect 43652 42924 43662 42980
rect 50866 42924 50876 42980
rect 50932 42924 51772 42980
rect 51828 42924 55580 42980
rect 55636 42924 55646 42980
rect 17042 42812 17052 42868
rect 17108 42812 17164 42868
rect 17220 42812 17836 42868
rect 17892 42812 17902 42868
rect 23090 42812 23100 42868
rect 23156 42812 24332 42868
rect 24388 42812 24398 42868
rect 33730 42812 33740 42868
rect 33796 42812 35868 42868
rect 35924 42812 35934 42868
rect 36306 42812 36316 42868
rect 36372 42812 38556 42868
rect 38612 42812 38780 42868
rect 38836 42812 40572 42868
rect 40628 42812 40638 42868
rect 42466 42812 42476 42868
rect 42532 42812 44940 42868
rect 44996 42812 45836 42868
rect 45892 42812 45902 42868
rect 6738 42700 6748 42756
rect 6804 42700 7532 42756
rect 7588 42700 7598 42756
rect 17266 42700 17276 42756
rect 17332 42700 20188 42756
rect 20244 42700 20254 42756
rect 23538 42700 23548 42756
rect 23604 42700 24556 42756
rect 24612 42700 25340 42756
rect 25396 42700 25406 42756
rect 30706 42700 30716 42756
rect 30772 42700 30828 42756
rect 30884 42700 30894 42756
rect 36194 42700 36204 42756
rect 36260 42700 36988 42756
rect 37044 42700 37054 42756
rect 37650 42700 37660 42756
rect 37716 42700 38668 42756
rect 38724 42700 38734 42756
rect 42242 42700 42252 42756
rect 42308 42700 42812 42756
rect 42868 42700 42878 42756
rect 44258 42700 44268 42756
rect 44324 42700 45164 42756
rect 45220 42700 45230 42756
rect 50978 42700 50988 42756
rect 51044 42700 53004 42756
rect 53060 42700 55356 42756
rect 55412 42700 55422 42756
rect 17948 42588 21308 42644
rect 21364 42588 21374 42644
rect 41346 42588 41356 42644
rect 41412 42588 42364 42644
rect 42420 42588 42430 42644
rect 42690 42588 42700 42644
rect 42756 42588 42924 42644
rect 42980 42588 42990 42644
rect 46722 42588 46732 42644
rect 46788 42588 47292 42644
rect 47348 42588 47358 42644
rect 47618 42588 47628 42644
rect 47684 42588 52892 42644
rect 52948 42588 53228 42644
rect 53284 42588 53294 42644
rect 9986 42476 9996 42532
rect 10052 42476 10780 42532
rect 10836 42476 11116 42532
rect 11172 42476 11788 42532
rect 11844 42476 12236 42532
rect 12292 42476 12302 42532
rect 17948 42420 18004 42588
rect 47628 42532 47684 42588
rect 18806 42476 18844 42532
rect 18900 42476 19516 42532
rect 19572 42476 19582 42532
rect 21186 42476 21196 42532
rect 21252 42476 21868 42532
rect 21924 42476 21934 42532
rect 31266 42476 31276 42532
rect 31332 42476 35308 42532
rect 40114 42476 40124 42532
rect 40180 42476 41468 42532
rect 41524 42476 47684 42532
rect 51314 42476 51324 42532
rect 51380 42476 52444 42532
rect 52500 42476 52510 42532
rect 17938 42364 17948 42420
rect 18004 42364 18014 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 35252 42308 35308 42476
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 18610 42252 18620 42308
rect 18676 42252 19628 42308
rect 19684 42252 19694 42308
rect 21522 42252 21532 42308
rect 21588 42252 26460 42308
rect 26516 42252 26526 42308
rect 35252 42252 37548 42308
rect 37604 42252 39620 42308
rect 19628 42196 19684 42252
rect 19628 42140 22092 42196
rect 22148 42140 23212 42196
rect 23268 42140 23278 42196
rect 32498 42140 32508 42196
rect 32564 42140 32574 42196
rect 37986 42140 37996 42196
rect 38052 42140 39004 42196
rect 39060 42140 39070 42196
rect 32508 42084 32564 42140
rect 39564 42084 39620 42252
rect 47282 42140 47292 42196
rect 47348 42140 47852 42196
rect 47908 42140 49644 42196
rect 49700 42140 49710 42196
rect 55570 42140 55580 42196
rect 55636 42140 56700 42196
rect 56756 42140 56766 42196
rect 19842 42028 19852 42084
rect 19908 42028 20860 42084
rect 20916 42028 20926 42084
rect 32508 42028 39284 42084
rect 39554 42028 39564 42084
rect 39620 42028 41468 42084
rect 41524 42028 41534 42084
rect 47852 42028 48748 42084
rect 48804 42028 48814 42084
rect 49522 42028 49532 42084
rect 49588 42028 50540 42084
rect 50596 42028 51156 42084
rect 56018 42028 56028 42084
rect 56084 42028 56588 42084
rect 56644 42028 57036 42084
rect 57092 42028 57102 42084
rect 39228 41972 39284 42028
rect 47852 41972 47908 42028
rect 8978 41916 8988 41972
rect 9044 41916 10108 41972
rect 10164 41916 10556 41972
rect 10612 41916 10622 41972
rect 14354 41916 14364 41972
rect 14420 41916 16044 41972
rect 16100 41916 16110 41972
rect 17714 41916 17724 41972
rect 17780 41916 17790 41972
rect 18834 41916 18844 41972
rect 18900 41916 20972 41972
rect 21028 41916 21038 41972
rect 21522 41916 21532 41972
rect 21588 41916 21756 41972
rect 21812 41916 21822 41972
rect 29138 41916 29148 41972
rect 29204 41916 30828 41972
rect 30884 41916 31164 41972
rect 31220 41916 31230 41972
rect 36978 41916 36988 41972
rect 37044 41916 38780 41972
rect 38836 41916 38846 41972
rect 39228 41916 39676 41972
rect 39732 41916 39742 41972
rect 41010 41916 41020 41972
rect 41076 41916 41580 41972
rect 41636 41916 41646 41972
rect 43586 41916 43596 41972
rect 43652 41916 44156 41972
rect 44212 41916 44222 41972
rect 46274 41916 46284 41972
rect 46340 41916 46956 41972
rect 47012 41916 47022 41972
rect 47842 41916 47852 41972
rect 47908 41916 47918 41972
rect 17724 41860 17780 41916
rect 21532 41860 21588 41916
rect 39228 41860 39284 41916
rect 51100 41860 51156 42028
rect 51762 41916 51772 41972
rect 51828 41916 52444 41972
rect 52500 41916 52510 41972
rect 6850 41804 6860 41860
rect 6916 41804 8876 41860
rect 8932 41804 8942 41860
rect 14252 41804 17780 41860
rect 18386 41804 18396 41860
rect 18452 41804 19292 41860
rect 19348 41804 19358 41860
rect 19954 41804 19964 41860
rect 20020 41804 21588 41860
rect 27906 41804 27916 41860
rect 27972 41804 28812 41860
rect 28868 41804 28878 41860
rect 38098 41804 38108 41860
rect 38164 41804 38556 41860
rect 38612 41804 38622 41860
rect 39218 41804 39228 41860
rect 39284 41804 39294 41860
rect 40226 41804 40236 41860
rect 40292 41804 46620 41860
rect 46676 41804 48300 41860
rect 48356 41804 48366 41860
rect 48514 41804 48524 41860
rect 48580 41804 50932 41860
rect 51090 41804 51100 41860
rect 51156 41804 55692 41860
rect 55748 41804 55758 41860
rect 14252 41748 14308 41804
rect 50876 41748 50932 41804
rect 14242 41692 14252 41748
rect 14308 41692 14318 41748
rect 17378 41692 17388 41748
rect 17444 41692 17948 41748
rect 18004 41692 18014 41748
rect 18162 41692 18172 41748
rect 18228 41692 19068 41748
rect 19124 41692 19134 41748
rect 33730 41692 33740 41748
rect 33796 41692 40124 41748
rect 40180 41692 40190 41748
rect 41234 41692 41244 41748
rect 41300 41692 41310 41748
rect 41458 41692 41468 41748
rect 41524 41692 43036 41748
rect 43092 41692 43102 41748
rect 45826 41692 45836 41748
rect 45892 41692 48860 41748
rect 48916 41692 48926 41748
rect 49074 41692 49084 41748
rect 49140 41692 50652 41748
rect 50708 41692 50718 41748
rect 50876 41692 52668 41748
rect 52724 41692 53900 41748
rect 53956 41692 54908 41748
rect 54964 41692 54974 41748
rect 41244 41636 41300 41692
rect 18050 41580 18060 41636
rect 18116 41580 19964 41636
rect 20020 41580 20030 41636
rect 41244 41580 47068 41636
rect 47124 41580 49196 41636
rect 49252 41580 49262 41636
rect 50530 41580 50540 41636
rect 50596 41580 51212 41636
rect 51268 41580 51278 41636
rect 53554 41580 53564 41636
rect 53620 41580 55692 41636
rect 55748 41580 55758 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 41916 41468 44828 41524
rect 44884 41468 45276 41524
rect 45332 41468 45342 41524
rect 48290 41468 48300 41524
rect 48356 41468 52556 41524
rect 52612 41468 52622 41524
rect 41916 41412 41972 41468
rect 17266 41356 17276 41412
rect 17332 41356 18732 41412
rect 18788 41356 18798 41412
rect 40114 41356 40124 41412
rect 40180 41356 41916 41412
rect 41972 41356 41982 41412
rect 18386 41244 18396 41300
rect 18452 41244 22092 41300
rect 22148 41244 22158 41300
rect 22418 41244 22428 41300
rect 22484 41244 23212 41300
rect 23268 41244 23278 41300
rect 41122 41244 41132 41300
rect 41188 41244 41804 41300
rect 41860 41244 41870 41300
rect 47954 41244 47964 41300
rect 48020 41244 48972 41300
rect 49028 41244 49532 41300
rect 49588 41244 49598 41300
rect 51538 41244 51548 41300
rect 51604 41244 55020 41300
rect 55076 41244 55086 41300
rect 15250 41132 15260 41188
rect 15316 41132 15820 41188
rect 15876 41132 15886 41188
rect 16258 41132 16268 41188
rect 16324 41132 19292 41188
rect 19348 41132 19358 41188
rect 19730 41132 19740 41188
rect 19796 41132 21980 41188
rect 22036 41132 22046 41188
rect 28578 41132 28588 41188
rect 28644 41132 29260 41188
rect 29316 41132 31724 41188
rect 31780 41132 31790 41188
rect 39218 41132 39228 41188
rect 39284 41132 39900 41188
rect 39956 41132 48524 41188
rect 48580 41132 48590 41188
rect 50082 41132 50092 41188
rect 50148 41132 50988 41188
rect 51044 41132 51660 41188
rect 51716 41132 51726 41188
rect 14802 41020 14812 41076
rect 14868 41020 16044 41076
rect 16100 41020 16110 41076
rect 16370 41020 16380 41076
rect 16436 41020 17612 41076
rect 17668 41020 17678 41076
rect 19506 41020 19516 41076
rect 19572 41020 20636 41076
rect 20692 41020 20702 41076
rect 32498 41020 32508 41076
rect 32564 41020 33516 41076
rect 33572 41020 33582 41076
rect 38434 41020 38444 41076
rect 38500 41020 40908 41076
rect 40964 41020 40974 41076
rect 41234 41020 41244 41076
rect 41300 41020 41804 41076
rect 41860 41020 43820 41076
rect 43876 41020 43886 41076
rect 50194 41020 50204 41076
rect 50260 41020 50540 41076
rect 50596 41020 50606 41076
rect 51314 41020 51324 41076
rect 51380 41020 56700 41076
rect 56756 41020 56766 41076
rect 5058 40908 5068 40964
rect 5124 40908 6076 40964
rect 6132 40908 8092 40964
rect 8148 40908 9212 40964
rect 9268 40908 9996 40964
rect 10052 40908 10062 40964
rect 14242 40908 14252 40964
rect 14308 40908 15260 40964
rect 15316 40908 15326 40964
rect 17826 40908 17836 40964
rect 17892 40908 19068 40964
rect 19124 40908 20300 40964
rect 20356 40908 20366 40964
rect 33394 40908 33404 40964
rect 33460 40908 34860 40964
rect 34916 40908 34926 40964
rect 35186 40908 35196 40964
rect 35252 40908 36092 40964
rect 36148 40908 36158 40964
rect 36530 40908 36540 40964
rect 36596 40908 39788 40964
rect 39844 40908 39854 40964
rect 40114 40908 40124 40964
rect 40180 40908 40236 40964
rect 40292 40908 41020 40964
rect 41076 40908 41086 40964
rect 43362 40908 43372 40964
rect 43428 40908 44940 40964
rect 44996 40908 48748 40964
rect 48804 40908 49756 40964
rect 49812 40908 49822 40964
rect 49970 40908 49980 40964
rect 50036 40908 50876 40964
rect 50932 40908 51884 40964
rect 51940 40908 51950 40964
rect 41020 40852 41076 40908
rect 7858 40796 7868 40852
rect 7924 40796 14980 40852
rect 15138 40796 15148 40852
rect 15204 40796 16156 40852
rect 16212 40796 16222 40852
rect 41020 40796 47068 40852
rect 47124 40796 47134 40852
rect 14924 40740 14980 40796
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 12450 40684 12460 40740
rect 12516 40684 14868 40740
rect 14924 40684 18508 40740
rect 18564 40684 18574 40740
rect 22306 40684 22316 40740
rect 22372 40684 23324 40740
rect 23380 40684 23390 40740
rect 43026 40684 43036 40740
rect 43092 40684 43372 40740
rect 43428 40684 43438 40740
rect 51090 40684 51100 40740
rect 51156 40684 51660 40740
rect 51716 40684 51726 40740
rect 14812 40628 14868 40684
rect 10630 40572 10668 40628
rect 10724 40572 10734 40628
rect 11442 40572 11452 40628
rect 11508 40572 13468 40628
rect 13524 40572 13534 40628
rect 14802 40572 14812 40628
rect 14868 40572 16940 40628
rect 16996 40572 17006 40628
rect 19282 40572 19292 40628
rect 19348 40572 20636 40628
rect 20692 40572 21756 40628
rect 21812 40572 21822 40628
rect 23202 40572 23212 40628
rect 23268 40572 24556 40628
rect 24612 40572 24622 40628
rect 42018 40572 42028 40628
rect 42084 40572 42700 40628
rect 42756 40572 43596 40628
rect 43652 40572 43662 40628
rect 9772 40460 10108 40516
rect 10164 40460 11564 40516
rect 11620 40460 11630 40516
rect 12898 40460 12908 40516
rect 12964 40460 14588 40516
rect 14644 40460 14654 40516
rect 16006 40460 16044 40516
rect 16100 40460 16110 40516
rect 21634 40460 21644 40516
rect 21700 40460 25676 40516
rect 25732 40460 25742 40516
rect 25900 40460 30492 40516
rect 30548 40460 30558 40516
rect 35634 40460 35644 40516
rect 35700 40460 37212 40516
rect 37268 40460 37278 40516
rect 39890 40460 39900 40516
rect 39956 40460 40572 40516
rect 40628 40460 40638 40516
rect 40786 40460 40796 40516
rect 40852 40460 44716 40516
rect 44772 40460 44782 40516
rect 49074 40460 49084 40516
rect 49140 40460 50204 40516
rect 50260 40460 50270 40516
rect 54114 40460 54124 40516
rect 54180 40460 55244 40516
rect 55300 40460 55310 40516
rect 55682 40460 55692 40516
rect 55748 40460 57372 40516
rect 57428 40460 57438 40516
rect 1810 40348 1820 40404
rect 1876 40348 4060 40404
rect 4116 40348 5068 40404
rect 5124 40348 5134 40404
rect 7410 40348 7420 40404
rect 7476 40348 8316 40404
rect 8372 40348 8382 40404
rect 9772 40292 9828 40460
rect 25900 40404 25956 40460
rect 10210 40348 10220 40404
rect 10276 40348 10892 40404
rect 10948 40348 10958 40404
rect 13570 40348 13580 40404
rect 13636 40348 14476 40404
rect 14532 40348 14542 40404
rect 16818 40348 16828 40404
rect 16884 40348 17836 40404
rect 17892 40348 18284 40404
rect 18340 40348 18350 40404
rect 18834 40348 18844 40404
rect 18900 40348 19068 40404
rect 19124 40348 22540 40404
rect 22596 40348 22606 40404
rect 22764 40348 25956 40404
rect 26450 40348 26460 40404
rect 26516 40348 27804 40404
rect 27860 40348 27870 40404
rect 31042 40348 31052 40404
rect 31108 40348 32060 40404
rect 32116 40348 33516 40404
rect 33572 40348 33582 40404
rect 36082 40348 36092 40404
rect 36148 40348 38668 40404
rect 42914 40348 42924 40404
rect 42980 40348 43820 40404
rect 43876 40348 44380 40404
rect 44436 40348 45500 40404
rect 45556 40348 45566 40404
rect 48066 40348 48076 40404
rect 48132 40348 49532 40404
rect 49588 40348 52668 40404
rect 52724 40348 52734 40404
rect 53778 40348 53788 40404
rect 53844 40348 54348 40404
rect 54404 40348 54414 40404
rect 22764 40292 22820 40348
rect 38612 40292 38668 40348
rect 3266 40236 3276 40292
rect 3332 40236 9604 40292
rect 9762 40236 9772 40292
rect 9828 40236 9838 40292
rect 10108 40236 12012 40292
rect 12068 40236 12078 40292
rect 15138 40236 15148 40292
rect 15204 40236 15820 40292
rect 15876 40236 15886 40292
rect 17042 40236 17052 40292
rect 17108 40236 22820 40292
rect 26562 40236 26572 40292
rect 26628 40236 27580 40292
rect 27636 40236 27646 40292
rect 31154 40236 31164 40292
rect 31220 40236 32508 40292
rect 32564 40236 33068 40292
rect 33124 40236 33134 40292
rect 38612 40236 46172 40292
rect 46228 40236 46238 40292
rect 51986 40236 51996 40292
rect 52052 40236 52892 40292
rect 52948 40236 53676 40292
rect 53732 40236 53742 40292
rect 9548 40180 9604 40236
rect 10108 40180 10164 40236
rect 3042 40124 3052 40180
rect 3108 40124 3948 40180
rect 4004 40124 4014 40180
rect 9548 40124 10164 40180
rect 10322 40124 10332 40180
rect 10388 40124 10398 40180
rect 13458 40124 13468 40180
rect 13524 40124 23436 40180
rect 23492 40124 23502 40180
rect 43474 40124 43484 40180
rect 43540 40124 43596 40180
rect 43652 40124 43662 40180
rect 52210 40124 52220 40180
rect 52276 40124 53900 40180
rect 53956 40124 53966 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 10332 39844 10388 40124
rect 15362 40012 15372 40068
rect 15428 40012 16268 40068
rect 16324 40012 16334 40068
rect 17154 40012 17164 40068
rect 17220 40012 34300 40068
rect 34356 40012 34366 40068
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 16818 39900 16828 39956
rect 16884 39900 18284 39956
rect 18340 39900 19292 39956
rect 19348 39900 19628 39956
rect 19684 39900 19694 39956
rect 26338 39900 26348 39956
rect 26404 39900 26572 39956
rect 26628 39900 26638 39956
rect 41468 39900 45388 39956
rect 45444 39900 45836 39956
rect 45892 39900 45902 39956
rect 41468 39844 41524 39900
rect 7970 39788 7980 39844
rect 8036 39788 10108 39844
rect 10164 39788 10174 39844
rect 10332 39788 11116 39844
rect 11172 39788 13468 39844
rect 13524 39788 13534 39844
rect 21046 39788 21084 39844
rect 21140 39788 21150 39844
rect 21746 39788 21756 39844
rect 21812 39788 22988 39844
rect 23044 39788 28028 39844
rect 28084 39788 28094 39844
rect 40338 39788 40348 39844
rect 40404 39788 41468 39844
rect 41524 39788 41534 39844
rect 42578 39788 42588 39844
rect 42644 39788 42654 39844
rect 43474 39788 43484 39844
rect 43540 39788 50428 39844
rect 50484 39788 50494 39844
rect 42588 39732 42644 39788
rect 4834 39676 4844 39732
rect 4900 39676 5740 39732
rect 5796 39676 5806 39732
rect 7074 39676 7084 39732
rect 7140 39676 8764 39732
rect 8820 39676 8830 39732
rect 12338 39676 12348 39732
rect 12404 39676 13580 39732
rect 13636 39676 13646 39732
rect 16594 39676 16604 39732
rect 16660 39676 17500 39732
rect 17556 39676 17566 39732
rect 17714 39676 17724 39732
rect 17780 39676 18844 39732
rect 18900 39676 18910 39732
rect 19404 39676 30268 39732
rect 30324 39676 31164 39732
rect 31220 39676 31230 39732
rect 34290 39676 34300 39732
rect 34356 39676 42924 39732
rect 42980 39676 42990 39732
rect 43922 39676 43932 39732
rect 43988 39676 46732 39732
rect 46788 39676 54124 39732
rect 54180 39676 54190 39732
rect 54674 39676 54684 39732
rect 54740 39676 55804 39732
rect 55860 39676 55870 39732
rect 17724 39620 17780 39676
rect 6066 39564 6076 39620
rect 6132 39564 7196 39620
rect 7252 39564 7262 39620
rect 8306 39564 8316 39620
rect 8372 39564 9660 39620
rect 9716 39564 11004 39620
rect 11060 39564 11070 39620
rect 12786 39564 12796 39620
rect 12852 39564 13468 39620
rect 13524 39564 13534 39620
rect 15810 39564 15820 39620
rect 15876 39564 17780 39620
rect 18498 39564 18508 39620
rect 18564 39564 19180 39620
rect 19236 39564 19246 39620
rect 7196 39508 7252 39564
rect 12796 39508 12852 39564
rect 19404 39508 19460 39676
rect 22082 39564 22092 39620
rect 22148 39564 28028 39620
rect 28084 39564 28094 39620
rect 30706 39564 30716 39620
rect 30772 39564 33964 39620
rect 34020 39564 34030 39620
rect 34402 39564 34412 39620
rect 34468 39564 36092 39620
rect 36148 39564 36158 39620
rect 36642 39564 36652 39620
rect 36708 39564 37772 39620
rect 37828 39564 37838 39620
rect 45154 39564 45164 39620
rect 45220 39564 46060 39620
rect 46116 39564 46126 39620
rect 48850 39564 48860 39620
rect 48916 39564 50540 39620
rect 50596 39564 53116 39620
rect 53172 39564 53182 39620
rect 4050 39452 4060 39508
rect 4116 39452 5628 39508
rect 5684 39452 5694 39508
rect 7196 39452 12852 39508
rect 14914 39452 14924 39508
rect 14980 39452 15932 39508
rect 15988 39452 19460 39508
rect 20066 39452 20076 39508
rect 20132 39452 20636 39508
rect 20692 39452 21532 39508
rect 21588 39452 21598 39508
rect 21858 39452 21868 39508
rect 21924 39452 24220 39508
rect 24276 39452 25228 39508
rect 25284 39452 25294 39508
rect 42130 39452 42140 39508
rect 42196 39452 42812 39508
rect 42868 39452 42878 39508
rect 50372 39452 51996 39508
rect 52052 39452 52062 39508
rect 52210 39452 52220 39508
rect 52276 39452 53004 39508
rect 53060 39452 53070 39508
rect 54338 39452 54348 39508
rect 54404 39452 55356 39508
rect 55412 39452 55422 39508
rect 50372 39396 50428 39452
rect 9202 39340 9212 39396
rect 9268 39340 9884 39396
rect 9940 39340 9950 39396
rect 10546 39340 10556 39396
rect 10612 39340 11900 39396
rect 11956 39340 13132 39396
rect 13188 39340 30828 39396
rect 30884 39340 31052 39396
rect 31108 39340 31612 39396
rect 31668 39340 31678 39396
rect 48374 39340 48412 39396
rect 48468 39340 48748 39396
rect 48804 39340 48814 39396
rect 49074 39340 49084 39396
rect 49140 39340 50428 39396
rect 51426 39340 51436 39396
rect 51492 39340 52668 39396
rect 52724 39340 52734 39396
rect 53218 39340 53228 39396
rect 53284 39340 53788 39396
rect 53844 39340 53854 39396
rect 3602 39228 3612 39284
rect 3668 39228 6412 39284
rect 6468 39228 10780 39284
rect 10836 39228 10846 39284
rect 24556 39228 26236 39284
rect 26292 39228 26796 39284
rect 26852 39228 26862 39284
rect 35970 39228 35980 39284
rect 36036 39228 39900 39284
rect 39956 39228 39966 39284
rect 41346 39228 41356 39284
rect 41412 39228 44604 39284
rect 44660 39228 44670 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 11330 39116 11340 39172
rect 11396 39116 12684 39172
rect 12740 39116 12750 39172
rect 13356 39116 18844 39172
rect 18900 39116 18910 39172
rect 13356 39060 13412 39116
rect 18844 39060 18900 39116
rect 24556 39060 24612 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 25218 39116 25228 39172
rect 25284 39116 27692 39172
rect 27748 39116 28028 39172
rect 28084 39116 28094 39172
rect 31602 39116 31612 39172
rect 31668 39116 31836 39172
rect 31892 39116 41020 39172
rect 41076 39116 41916 39172
rect 41972 39116 44156 39172
rect 44212 39116 44222 39172
rect 9874 39004 9884 39060
rect 9940 39004 11396 39060
rect 11554 39004 11564 39060
rect 11620 39004 13412 39060
rect 14690 39004 14700 39060
rect 14756 39004 16828 39060
rect 16884 39004 16894 39060
rect 18844 39004 21084 39060
rect 21140 39004 21150 39060
rect 22092 39004 24556 39060
rect 24612 39004 24622 39060
rect 26674 39004 26684 39060
rect 26740 39004 26852 39060
rect 30034 39004 30044 39060
rect 30100 39004 30940 39060
rect 30996 39004 31006 39060
rect 34290 39004 34300 39060
rect 34356 39004 34636 39060
rect 34692 39004 34702 39060
rect 36978 39004 36988 39060
rect 37044 39004 37772 39060
rect 37828 39004 37838 39060
rect 40450 39004 40460 39060
rect 40516 39004 42252 39060
rect 42308 39004 42318 39060
rect 44370 39004 44380 39060
rect 44436 39004 46844 39060
rect 46900 39004 46910 39060
rect 55346 39004 55356 39060
rect 55412 39004 57148 39060
rect 57204 39004 57214 39060
rect 2930 38892 2940 38948
rect 2996 38892 3836 38948
rect 3892 38892 4284 38948
rect 4340 38892 5180 38948
rect 5236 38892 5246 38948
rect 10182 38892 10220 38948
rect 10276 38892 10286 38948
rect 3042 38780 3052 38836
rect 3108 38780 3388 38836
rect 3444 38780 3724 38836
rect 3780 38780 3790 38836
rect 4722 38780 4732 38836
rect 4788 38780 5460 38836
rect 8754 38780 8764 38836
rect 8820 38780 9996 38836
rect 10052 38780 10062 38836
rect 5404 38724 5460 38780
rect 5404 38668 7644 38724
rect 7700 38668 7710 38724
rect 11340 38668 11396 39004
rect 22092 38948 22148 39004
rect 12002 38892 12012 38948
rect 12068 38892 12796 38948
rect 12852 38892 12862 38948
rect 13570 38892 13580 38948
rect 13636 38892 14364 38948
rect 14420 38892 14430 38948
rect 19170 38892 19180 38948
rect 19236 38892 22092 38948
rect 22148 38892 22158 38948
rect 23538 38892 23548 38948
rect 23604 38892 24108 38948
rect 24164 38892 26572 38948
rect 26628 38892 26638 38948
rect 26796 38836 26852 39004
rect 27122 38892 27132 38948
rect 27188 38892 28924 38948
rect 28980 38892 28990 38948
rect 29698 38892 29708 38948
rect 29764 38892 32284 38948
rect 32340 38892 32350 38948
rect 36530 38892 36540 38948
rect 36596 38892 41468 38948
rect 41524 38892 42476 38948
rect 42532 38892 42542 38948
rect 43586 38892 43596 38948
rect 43652 38892 44604 38948
rect 44660 38892 44670 38948
rect 55010 38892 55020 38948
rect 55076 38892 55916 38948
rect 55972 38892 55982 38948
rect 12450 38780 12460 38836
rect 12516 38780 14252 38836
rect 14308 38780 14318 38836
rect 16818 38780 16828 38836
rect 16884 38780 17052 38836
rect 17108 38780 17118 38836
rect 17826 38780 17836 38836
rect 17892 38780 18284 38836
rect 18340 38780 18350 38836
rect 20290 38780 20300 38836
rect 20356 38780 20748 38836
rect 20804 38780 23212 38836
rect 23268 38780 23278 38836
rect 24322 38780 24332 38836
rect 24388 38780 25340 38836
rect 25396 38780 26348 38836
rect 26404 38780 26414 38836
rect 26684 38780 26852 38836
rect 27458 38780 27468 38836
rect 27524 38780 27534 38836
rect 35186 38780 35196 38836
rect 35252 38780 35980 38836
rect 36036 38780 36046 38836
rect 36306 38780 36316 38836
rect 36372 38780 37660 38836
rect 37716 38780 37726 38836
rect 41122 38780 41132 38836
rect 41188 38780 43484 38836
rect 43540 38780 44716 38836
rect 44772 38780 44782 38836
rect 50418 38780 50428 38836
rect 50484 38780 52892 38836
rect 52948 38780 52958 38836
rect 26684 38724 26740 38780
rect 27468 38724 27524 38780
rect 11788 38668 12628 38724
rect 13010 38668 13020 38724
rect 13076 38668 13356 38724
rect 13412 38668 13422 38724
rect 13580 38668 15148 38724
rect 15204 38668 15214 38724
rect 17490 38668 17500 38724
rect 17556 38668 18172 38724
rect 18228 38668 18238 38724
rect 19394 38668 19404 38724
rect 19460 38668 20076 38724
rect 20132 38668 21532 38724
rect 21588 38668 21598 38724
rect 25218 38668 25228 38724
rect 25284 38668 26236 38724
rect 26292 38668 27524 38724
rect 41794 38668 41804 38724
rect 41860 38668 42588 38724
rect 42644 38668 42654 38724
rect 50642 38668 50652 38724
rect 50708 38668 51436 38724
rect 51492 38668 52220 38724
rect 52276 38668 52286 38724
rect 53340 38668 54124 38724
rect 54180 38668 54190 38724
rect 5404 38612 5460 38668
rect 11340 38612 11844 38668
rect 12572 38612 12628 38668
rect 13580 38612 13636 38668
rect 53340 38612 53396 38668
rect 4610 38556 4620 38612
rect 4676 38556 4900 38612
rect 5394 38556 5404 38612
rect 5460 38556 5470 38612
rect 5730 38556 5740 38612
rect 5796 38556 6300 38612
rect 6356 38556 6366 38612
rect 6850 38556 6860 38612
rect 6916 38556 7532 38612
rect 7588 38556 7598 38612
rect 10210 38556 10220 38612
rect 10276 38556 10500 38612
rect 12562 38556 12572 38612
rect 12628 38556 12638 38612
rect 12796 38556 13636 38612
rect 20626 38556 20636 38612
rect 20692 38556 21308 38612
rect 21364 38556 21374 38612
rect 23650 38556 23660 38612
rect 23716 38556 24332 38612
rect 24388 38556 24398 38612
rect 27570 38556 27580 38612
rect 27636 38556 28364 38612
rect 28420 38556 28430 38612
rect 30370 38556 30380 38612
rect 30436 38556 41916 38612
rect 41972 38556 41982 38612
rect 48402 38556 48412 38612
rect 48468 38556 48860 38612
rect 48916 38556 48926 38612
rect 52434 38556 52444 38612
rect 52500 38556 53116 38612
rect 53172 38556 53182 38612
rect 53302 38556 53340 38612
rect 53396 38556 53406 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 4844 38388 4900 38556
rect 10444 38500 10500 38556
rect 12796 38500 12852 38556
rect 10434 38444 10444 38500
rect 10500 38444 10510 38500
rect 11554 38444 11564 38500
rect 11620 38444 12852 38500
rect 13458 38444 13468 38500
rect 13524 38444 14476 38500
rect 14532 38444 14542 38500
rect 20150 38444 20188 38500
rect 20244 38444 20254 38500
rect 20374 38444 20412 38500
rect 20468 38444 20478 38500
rect 21186 38444 21196 38500
rect 21252 38444 21532 38500
rect 21588 38444 21598 38500
rect 4834 38332 4844 38388
rect 4900 38332 4910 38388
rect 8306 38332 8316 38388
rect 8372 38332 10332 38388
rect 10388 38332 10668 38388
rect 10724 38332 10734 38388
rect 15474 38332 15484 38388
rect 15540 38332 20524 38388
rect 20580 38332 20590 38388
rect 9762 38220 9772 38276
rect 9828 38220 10220 38276
rect 10276 38220 10286 38276
rect 12786 38220 12796 38276
rect 12852 38220 15036 38276
rect 15092 38220 20636 38276
rect 20692 38220 24220 38276
rect 24276 38220 24892 38276
rect 24948 38220 24958 38276
rect 30380 38164 30436 38556
rect 53340 38500 53396 38556
rect 36642 38444 36652 38500
rect 36708 38444 37100 38500
rect 37156 38444 37166 38500
rect 40450 38444 40460 38500
rect 40516 38444 45948 38500
rect 46004 38444 53396 38500
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 36988 38332 38668 38388
rect 45266 38332 45276 38388
rect 45332 38332 46060 38388
rect 46116 38332 46126 38388
rect 36988 38276 37044 38332
rect 38612 38276 38668 38332
rect 36978 38220 36988 38276
rect 37044 38220 37054 38276
rect 37650 38220 37660 38276
rect 37716 38220 38220 38276
rect 38276 38220 38286 38276
rect 38612 38220 40684 38276
rect 40740 38220 43932 38276
rect 43988 38220 43998 38276
rect 9650 38108 9660 38164
rect 9716 38108 10668 38164
rect 10724 38108 12908 38164
rect 12964 38108 15708 38164
rect 15764 38108 15774 38164
rect 16594 38108 16604 38164
rect 16660 38108 17164 38164
rect 17220 38108 17230 38164
rect 18498 38108 18508 38164
rect 18564 38108 19628 38164
rect 19684 38108 19694 38164
rect 26852 38108 30436 38164
rect 41458 38108 41468 38164
rect 41524 38108 42700 38164
rect 42756 38108 42766 38164
rect 26852 38052 26908 38108
rect 7522 37996 7532 38052
rect 7588 37996 13804 38052
rect 13860 37996 13870 38052
rect 15092 37996 26908 38052
rect 28578 37996 28588 38052
rect 28644 37996 30044 38052
rect 30100 37996 30110 38052
rect 30930 37996 30940 38052
rect 30996 37996 31612 38052
rect 31668 37996 31678 38052
rect 34738 37996 34748 38052
rect 34804 37996 35420 38052
rect 35476 37996 35756 38052
rect 35812 37996 35822 38052
rect 42466 37996 42476 38052
rect 42532 37996 43820 38052
rect 43876 37996 43886 38052
rect 48962 37996 48972 38052
rect 49028 37996 49868 38052
rect 49924 37996 53116 38052
rect 53172 37996 53182 38052
rect 53554 37996 53564 38052
rect 53620 37996 56588 38052
rect 56644 37996 56654 38052
rect 2706 37884 2716 37940
rect 2772 37884 3948 37940
rect 4004 37884 4014 37940
rect 10434 37884 10444 37940
rect 10500 37884 13468 37940
rect 13524 37884 13534 37940
rect 15092 37828 15148 37996
rect 17126 37884 17164 37940
rect 17220 37884 17230 37940
rect 20626 37884 20636 37940
rect 20692 37884 22204 37940
rect 22260 37884 22270 37940
rect 22530 37884 22540 37940
rect 22596 37884 23436 37940
rect 23492 37884 23772 37940
rect 23828 37884 23838 37940
rect 27794 37884 27804 37940
rect 27860 37884 28364 37940
rect 28420 37884 29260 37940
rect 29316 37884 29326 37940
rect 37650 37884 37660 37940
rect 37716 37884 38780 37940
rect 38836 37884 38846 37940
rect 42662 37884 42700 37940
rect 42756 37884 42766 37940
rect 50530 37884 50540 37940
rect 50596 37884 52892 37940
rect 52948 37884 52958 37940
rect 53666 37884 53676 37940
rect 53732 37884 54684 37940
rect 54740 37884 54750 37940
rect 3714 37772 3724 37828
rect 3780 37772 5068 37828
rect 5124 37772 5134 37828
rect 8418 37772 8428 37828
rect 8484 37772 9212 37828
rect 9268 37772 15148 37828
rect 17378 37772 17388 37828
rect 17444 37772 20188 37828
rect 20244 37772 20254 37828
rect 21270 37772 21308 37828
rect 21364 37772 21374 37828
rect 21634 37772 21644 37828
rect 21700 37772 22316 37828
rect 22372 37772 22382 37828
rect 26674 37772 26684 37828
rect 26740 37772 26908 37828
rect 34402 37772 34412 37828
rect 34468 37772 35084 37828
rect 35140 37772 36316 37828
rect 36372 37772 36382 37828
rect 46050 37772 46060 37828
rect 46116 37772 51772 37828
rect 51828 37772 51838 37828
rect 56802 37772 56812 37828
rect 56868 37772 57260 37828
rect 57316 37772 57326 37828
rect 20188 37716 20244 37772
rect 10546 37660 10556 37716
rect 10612 37660 10668 37716
rect 10724 37660 11116 37716
rect 11172 37660 11182 37716
rect 20188 37660 22764 37716
rect 22820 37660 23996 37716
rect 24052 37660 24062 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 17154 37548 17164 37604
rect 17220 37548 17836 37604
rect 17892 37548 17902 37604
rect 20178 37548 20188 37604
rect 20244 37548 20524 37604
rect 20580 37548 25676 37604
rect 25732 37548 26348 37604
rect 26404 37548 26414 37604
rect 2370 37436 2380 37492
rect 2436 37436 3500 37492
rect 3556 37436 3566 37492
rect 15922 37436 15932 37492
rect 15988 37436 17388 37492
rect 17444 37436 17454 37492
rect 17938 37436 17948 37492
rect 18004 37436 18956 37492
rect 19012 37436 19022 37492
rect 19170 37436 19180 37492
rect 19236 37436 19852 37492
rect 19908 37436 19918 37492
rect 20710 37436 20748 37492
rect 20804 37436 20814 37492
rect 26852 37380 26908 37772
rect 52882 37660 52892 37716
rect 52948 37660 55468 37716
rect 55524 37660 55804 37716
rect 55860 37660 55870 37716
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 42242 37548 42252 37604
rect 42308 37548 43372 37604
rect 43428 37548 43438 37604
rect 51650 37548 51660 37604
rect 51716 37548 52332 37604
rect 52388 37548 53452 37604
rect 53508 37548 56140 37604
rect 56196 37548 56206 37604
rect 51660 37492 51716 37548
rect 28242 37436 28252 37492
rect 28308 37436 29148 37492
rect 29204 37436 29214 37492
rect 31266 37436 31276 37492
rect 31332 37436 31836 37492
rect 31892 37436 31902 37492
rect 36306 37436 36316 37492
rect 36372 37436 44604 37492
rect 44660 37436 46284 37492
rect 46340 37436 46350 37492
rect 50194 37436 50204 37492
rect 50260 37436 51716 37492
rect 52658 37436 52668 37492
rect 52724 37436 55692 37492
rect 55748 37436 55758 37492
rect 6178 37324 6188 37380
rect 6244 37324 7756 37380
rect 7812 37324 7822 37380
rect 13010 37324 13020 37380
rect 13076 37324 22540 37380
rect 22596 37324 22606 37380
rect 26852 37324 27580 37380
rect 27636 37324 27804 37380
rect 27860 37324 27870 37380
rect 33506 37324 33516 37380
rect 33572 37324 46396 37380
rect 46452 37324 46462 37380
rect 50978 37324 50988 37380
rect 51044 37324 52220 37380
rect 52276 37324 52286 37380
rect 53218 37324 53228 37380
rect 53284 37324 54124 37380
rect 54180 37324 54908 37380
rect 54964 37324 55580 37380
rect 55636 37324 55646 37380
rect 3714 37212 3724 37268
rect 3780 37212 4620 37268
rect 4676 37212 4686 37268
rect 5170 37212 5180 37268
rect 5236 37212 5852 37268
rect 5908 37212 5918 37268
rect 14130 37212 14140 37268
rect 14196 37212 14812 37268
rect 14868 37212 20300 37268
rect 20356 37212 20366 37268
rect 21298 37212 21308 37268
rect 21364 37212 21980 37268
rect 22036 37212 22046 37268
rect 31938 37212 31948 37268
rect 32004 37212 35532 37268
rect 35588 37212 35598 37268
rect 38770 37212 38780 37268
rect 38836 37212 39452 37268
rect 39508 37212 39518 37268
rect 41682 37212 41692 37268
rect 41748 37212 42364 37268
rect 42420 37212 43820 37268
rect 43876 37212 43886 37268
rect 45154 37212 45164 37268
rect 45220 37212 46620 37268
rect 46676 37212 53788 37268
rect 53844 37212 53854 37268
rect 54226 37212 54236 37268
rect 54292 37212 54684 37268
rect 54740 37212 54750 37268
rect 55804 37212 57260 37268
rect 57316 37212 57326 37268
rect 21308 37156 21364 37212
rect 53788 37156 53844 37212
rect 55804 37156 55860 37212
rect 3042 37100 3052 37156
rect 3108 37100 6076 37156
rect 6132 37100 6142 37156
rect 6290 37100 6300 37156
rect 6356 37100 9884 37156
rect 9940 37100 11788 37156
rect 11844 37100 11854 37156
rect 16818 37100 16828 37156
rect 16884 37100 17612 37156
rect 17668 37100 21364 37156
rect 24210 37100 24220 37156
rect 24276 37100 27244 37156
rect 27300 37100 27310 37156
rect 43698 37100 43708 37156
rect 43764 37100 47628 37156
rect 47684 37100 47694 37156
rect 53788 37100 54572 37156
rect 54628 37100 54638 37156
rect 55794 37100 55804 37156
rect 55860 37100 55870 37156
rect 56018 37100 56028 37156
rect 56084 37100 57148 37156
rect 57204 37100 57214 37156
rect 2482 36988 2492 37044
rect 2548 36988 3948 37044
rect 4004 36988 4014 37044
rect 5058 36988 5068 37044
rect 5124 36988 6188 37044
rect 6244 36988 6254 37044
rect 11330 36988 11340 37044
rect 11396 36988 14700 37044
rect 14756 36988 14766 37044
rect 15586 36988 15596 37044
rect 15652 36988 16940 37044
rect 16996 36988 17006 37044
rect 20402 36988 20412 37044
rect 20468 36988 20860 37044
rect 20916 36988 20926 37044
rect 39330 36988 39340 37044
rect 39396 36988 41076 37044
rect 41234 36988 41244 37044
rect 41300 36988 43036 37044
rect 43092 36988 43102 37044
rect 46386 36988 46396 37044
rect 46452 36988 47180 37044
rect 47236 36988 48412 37044
rect 48468 36988 48478 37044
rect 54898 36988 54908 37044
rect 54964 36988 56812 37044
rect 56868 36988 56878 37044
rect 41020 36932 41076 36988
rect 15362 36876 15372 36932
rect 15428 36876 19628 36932
rect 19684 36876 19694 36932
rect 39218 36876 39228 36932
rect 39284 36876 39788 36932
rect 39844 36876 39854 36932
rect 41020 36876 43372 36932
rect 43428 36876 43438 36932
rect 45490 36876 45500 36932
rect 45556 36876 46508 36932
rect 46564 36876 46574 36932
rect 48178 36876 48188 36932
rect 48244 36876 48860 36932
rect 48916 36876 48926 36932
rect 52210 36876 52220 36932
rect 52276 36876 53452 36932
rect 53508 36876 54348 36932
rect 54404 36876 55244 36932
rect 55300 36876 55310 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 9090 36764 9100 36820
rect 9156 36764 9660 36820
rect 9716 36764 14476 36820
rect 14532 36764 14542 36820
rect 19954 36764 19964 36820
rect 20020 36764 22988 36820
rect 23044 36764 23054 36820
rect 26226 36764 26236 36820
rect 26292 36764 26908 36820
rect 26964 36764 26974 36820
rect 42130 36764 42140 36820
rect 42196 36764 43148 36820
rect 43204 36764 43484 36820
rect 43540 36764 43550 36820
rect 5282 36652 5292 36708
rect 5348 36652 6412 36708
rect 6468 36652 6478 36708
rect 8306 36652 8316 36708
rect 8372 36652 10108 36708
rect 10164 36652 10174 36708
rect 11554 36652 11564 36708
rect 11620 36652 15036 36708
rect 15092 36652 21532 36708
rect 21588 36652 21598 36708
rect 26786 36652 26796 36708
rect 26852 36652 29260 36708
rect 29316 36652 29326 36708
rect 34514 36652 34524 36708
rect 34580 36652 35308 36708
rect 35364 36652 37772 36708
rect 37828 36652 37838 36708
rect 45826 36652 45836 36708
rect 45892 36652 48636 36708
rect 48692 36652 51884 36708
rect 51940 36652 51950 36708
rect 52546 36652 52556 36708
rect 52612 36652 54236 36708
rect 54292 36652 54302 36708
rect 8194 36540 8204 36596
rect 8260 36540 12124 36596
rect 12180 36540 12190 36596
rect 13458 36540 13468 36596
rect 13524 36540 14588 36596
rect 14644 36540 15148 36596
rect 21410 36540 21420 36596
rect 21476 36540 22764 36596
rect 22820 36540 22830 36596
rect 22988 36540 34076 36596
rect 34132 36540 34142 36596
rect 44146 36540 44156 36596
rect 44212 36540 48188 36596
rect 48244 36540 48254 36596
rect 50866 36540 50876 36596
rect 50932 36540 52668 36596
rect 52724 36540 52734 36596
rect 15092 36484 15148 36540
rect 22988 36484 23044 36540
rect 44156 36484 44212 36540
rect 5730 36428 5740 36484
rect 5796 36428 6076 36484
rect 6132 36428 8876 36484
rect 8932 36428 9436 36484
rect 9492 36428 9502 36484
rect 10098 36428 10108 36484
rect 10164 36428 10780 36484
rect 10836 36428 10846 36484
rect 11666 36428 11676 36484
rect 11732 36428 14028 36484
rect 14084 36428 14094 36484
rect 14802 36428 14812 36484
rect 14868 36428 14878 36484
rect 15092 36428 18732 36484
rect 18788 36428 18798 36484
rect 21532 36428 23044 36484
rect 23426 36428 23436 36484
rect 23492 36428 24108 36484
rect 24164 36428 24174 36484
rect 26450 36428 26460 36484
rect 26516 36428 27580 36484
rect 27636 36428 27646 36484
rect 28578 36428 28588 36484
rect 28644 36428 29596 36484
rect 29652 36428 29662 36484
rect 30034 36428 30044 36484
rect 30100 36428 34188 36484
rect 34244 36428 34860 36484
rect 34916 36428 34926 36484
rect 35074 36428 35084 36484
rect 35140 36428 35420 36484
rect 35476 36428 35980 36484
rect 36036 36428 36046 36484
rect 43362 36428 43372 36484
rect 43428 36428 44212 36484
rect 51426 36428 51436 36484
rect 51492 36428 53004 36484
rect 53060 36428 53070 36484
rect 54338 36428 54348 36484
rect 54404 36428 57260 36484
rect 57316 36428 57326 36484
rect 14812 36372 14868 36428
rect 4610 36316 4620 36372
rect 4676 36316 4956 36372
rect 5012 36316 5022 36372
rect 7298 36316 7308 36372
rect 7364 36316 7532 36372
rect 7588 36316 10668 36372
rect 10724 36316 10734 36372
rect 12786 36316 12796 36372
rect 12852 36316 14364 36372
rect 14420 36316 14868 36372
rect 15138 36316 15148 36372
rect 15204 36316 16156 36372
rect 16212 36316 16222 36372
rect 17938 36316 17948 36372
rect 18004 36316 18844 36372
rect 18900 36316 18910 36372
rect 20598 36316 20636 36372
rect 20692 36316 20702 36372
rect 14812 36260 14868 36316
rect 5954 36204 5964 36260
rect 6020 36204 8204 36260
rect 8260 36204 8270 36260
rect 12114 36204 12124 36260
rect 12180 36204 13916 36260
rect 13972 36204 13982 36260
rect 14130 36204 14140 36260
rect 14196 36204 14234 36260
rect 14550 36204 14588 36260
rect 14644 36204 14654 36260
rect 14812 36204 16044 36260
rect 16100 36204 16110 36260
rect 16258 36204 16268 36260
rect 16324 36204 16362 36260
rect 19628 36204 21308 36260
rect 21364 36204 21374 36260
rect 19628 36148 19684 36204
rect 21532 36148 21588 36428
rect 22754 36316 22764 36372
rect 22820 36316 24556 36372
rect 24612 36316 24622 36372
rect 25666 36316 25676 36372
rect 25732 36316 26796 36372
rect 26852 36316 26862 36372
rect 39106 36316 39116 36372
rect 39172 36316 40908 36372
rect 40964 36316 40974 36372
rect 43138 36316 43148 36372
rect 43204 36316 44380 36372
rect 44436 36316 44446 36372
rect 49634 36316 49644 36372
rect 49700 36316 51996 36372
rect 52052 36316 52062 36372
rect 24434 36204 24444 36260
rect 24500 36204 27804 36260
rect 27860 36204 27870 36260
rect 30258 36204 30268 36260
rect 30324 36204 31388 36260
rect 31444 36204 33628 36260
rect 33684 36204 34188 36260
rect 34244 36204 34860 36260
rect 34916 36204 34926 36260
rect 38322 36204 38332 36260
rect 38388 36204 39228 36260
rect 39284 36204 39294 36260
rect 45826 36204 45836 36260
rect 45892 36204 46284 36260
rect 46340 36204 46350 36260
rect 47842 36204 47852 36260
rect 47908 36204 48300 36260
rect 48356 36204 48366 36260
rect 50306 36204 50316 36260
rect 50372 36204 54012 36260
rect 54068 36204 54078 36260
rect 11218 36092 11228 36148
rect 11284 36092 19684 36148
rect 21084 36092 21588 36148
rect 26674 36092 26684 36148
rect 26740 36092 27020 36148
rect 27076 36092 31052 36148
rect 31108 36092 31118 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 2146 35980 2156 36036
rect 2212 35980 3052 36036
rect 3108 35980 5292 36036
rect 5348 35980 5358 36036
rect 12674 35980 12684 36036
rect 12740 35980 14924 36036
rect 14980 35980 14990 36036
rect 15082 35980 15092 36036
rect 15148 35980 19628 36036
rect 19684 35980 19694 36036
rect 21084 35924 21140 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 10882 35868 10892 35924
rect 10948 35868 11564 35924
rect 11620 35868 11630 35924
rect 14690 35868 14700 35924
rect 14756 35868 15372 35924
rect 15428 35868 15438 35924
rect 16818 35868 16828 35924
rect 16884 35868 19516 35924
rect 19572 35868 21140 35924
rect 21196 35980 26908 36036
rect 27794 35980 27804 36036
rect 27860 35980 29148 36036
rect 29204 35980 29214 36036
rect 35074 35980 35084 36036
rect 35140 35980 43708 36036
rect 44258 35980 44268 36036
rect 44324 35980 45388 36036
rect 45444 35980 45454 36036
rect 47394 35980 47404 36036
rect 47460 35980 48020 36036
rect 21196 35812 21252 35980
rect 26852 35924 26908 35980
rect 43652 35924 43708 35980
rect 47964 35924 48020 35980
rect 53564 35980 54908 36036
rect 54964 35980 54974 36036
rect 53564 35924 53620 35980
rect 14802 35756 14812 35812
rect 14868 35756 15148 35812
rect 15922 35756 15932 35812
rect 15988 35756 21252 35812
rect 21644 35868 22540 35924
rect 22596 35868 22606 35924
rect 23314 35868 23324 35924
rect 23380 35868 23996 35924
rect 24052 35868 26236 35924
rect 26292 35868 26302 35924
rect 26852 35868 31500 35924
rect 31556 35868 36988 35924
rect 37044 35868 37054 35924
rect 43652 35868 47516 35924
rect 47572 35868 47740 35924
rect 47796 35868 47806 35924
rect 47964 35868 53620 35924
rect 53778 35868 53788 35924
rect 53844 35868 54684 35924
rect 54740 35868 54750 35924
rect 6738 35644 6748 35700
rect 6804 35644 13468 35700
rect 13524 35644 13804 35700
rect 13860 35644 13870 35700
rect 15092 35588 15148 35756
rect 15586 35644 15596 35700
rect 15652 35644 16492 35700
rect 16548 35644 16558 35700
rect 20626 35644 20636 35700
rect 20692 35644 21084 35700
rect 21140 35644 21150 35700
rect 21644 35588 21700 35868
rect 22418 35756 22428 35812
rect 22484 35756 26796 35812
rect 26852 35756 26862 35812
rect 33842 35756 33852 35812
rect 33908 35756 34412 35812
rect 34468 35756 35308 35812
rect 35364 35756 35374 35812
rect 40114 35756 40124 35812
rect 40180 35756 41580 35812
rect 41636 35756 42812 35812
rect 42868 35756 42878 35812
rect 43474 35756 43484 35812
rect 43540 35756 44492 35812
rect 44548 35756 44558 35812
rect 51762 35756 51772 35812
rect 51828 35756 53228 35812
rect 53284 35756 53294 35812
rect 54226 35756 54236 35812
rect 54292 35756 54572 35812
rect 54628 35756 54638 35812
rect 55346 35756 55356 35812
rect 55412 35756 56588 35812
rect 56644 35756 56654 35812
rect 22642 35644 22652 35700
rect 22708 35644 23548 35700
rect 23604 35644 23614 35700
rect 23762 35644 23772 35700
rect 23828 35644 23838 35700
rect 24882 35644 24892 35700
rect 24948 35644 28588 35700
rect 28644 35644 28654 35700
rect 29250 35644 29260 35700
rect 29316 35644 29820 35700
rect 29876 35644 29886 35700
rect 32722 35644 32732 35700
rect 32788 35644 36932 35700
rect 38098 35644 38108 35700
rect 38164 35644 38892 35700
rect 38948 35644 38958 35700
rect 47954 35644 47964 35700
rect 48020 35644 49196 35700
rect 49252 35644 49980 35700
rect 50036 35644 50046 35700
rect 53554 35644 53564 35700
rect 53620 35644 55580 35700
rect 55636 35644 57036 35700
rect 57092 35644 57932 35700
rect 57988 35644 57998 35700
rect 23772 35588 23828 35644
rect 36876 35588 36932 35644
rect 3938 35532 3948 35588
rect 4004 35532 4284 35588
rect 4340 35532 8652 35588
rect 8708 35532 9324 35588
rect 9380 35532 9390 35588
rect 13906 35532 13916 35588
rect 13972 35532 14924 35588
rect 14980 35532 14990 35588
rect 15092 35532 16716 35588
rect 16772 35532 17388 35588
rect 17444 35532 17454 35588
rect 20850 35532 20860 35588
rect 20916 35532 21196 35588
rect 21252 35532 21644 35588
rect 21700 35532 21710 35588
rect 22194 35532 22204 35588
rect 22260 35532 22540 35588
rect 22596 35532 23828 35588
rect 27794 35532 27804 35588
rect 27860 35532 29932 35588
rect 29988 35532 29998 35588
rect 32834 35532 32844 35588
rect 32900 35532 33740 35588
rect 33796 35532 33806 35588
rect 34066 35532 34076 35588
rect 34132 35532 34636 35588
rect 34692 35532 35084 35588
rect 35140 35532 35150 35588
rect 36866 35532 36876 35588
rect 36932 35532 41132 35588
rect 41188 35532 42028 35588
rect 42084 35532 42094 35588
rect 49522 35532 49532 35588
rect 49588 35532 50764 35588
rect 50820 35532 50830 35588
rect 51650 35532 51660 35588
rect 51716 35532 53004 35588
rect 53060 35532 53070 35588
rect 54114 35532 54124 35588
rect 54180 35532 54796 35588
rect 54852 35532 54862 35588
rect 57250 35532 57260 35588
rect 57316 35532 58044 35588
rect 58100 35532 58110 35588
rect 5394 35420 5404 35476
rect 5460 35420 7420 35476
rect 7476 35420 7486 35476
rect 16006 35420 16044 35476
rect 16100 35420 16110 35476
rect 17714 35420 17724 35476
rect 17780 35420 18284 35476
rect 18340 35420 18350 35476
rect 21644 35364 21700 35532
rect 32498 35420 32508 35476
rect 32564 35420 34972 35476
rect 35028 35420 35038 35476
rect 46722 35420 46732 35476
rect 46788 35420 48412 35476
rect 48468 35420 50988 35476
rect 51044 35420 52444 35476
rect 52500 35420 52510 35476
rect 52780 35420 52892 35476
rect 52948 35420 52958 35476
rect 53778 35420 53788 35476
rect 53844 35420 55132 35476
rect 55188 35420 55198 35476
rect 4844 35308 6076 35364
rect 6132 35308 6142 35364
rect 15894 35308 15932 35364
rect 15988 35308 15998 35364
rect 16380 35308 16884 35364
rect 19282 35308 19292 35364
rect 19348 35308 20748 35364
rect 20804 35308 20814 35364
rect 21644 35308 22428 35364
rect 22484 35308 22494 35364
rect 24882 35308 24892 35364
rect 24948 35308 28252 35364
rect 28308 35308 28318 35364
rect 28914 35308 28924 35364
rect 28980 35308 32172 35364
rect 32228 35308 32238 35364
rect 40898 35308 40908 35364
rect 40964 35308 43036 35364
rect 43092 35308 43102 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 4844 35140 4900 35308
rect 16380 35252 16436 35308
rect 8642 35196 8652 35252
rect 8708 35196 9660 35252
rect 9716 35196 11452 35252
rect 11508 35196 13804 35252
rect 13860 35196 13870 35252
rect 14242 35196 14252 35252
rect 14308 35196 16436 35252
rect 16828 35140 16884 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 52780 35252 52836 35420
rect 52994 35308 53004 35364
rect 53060 35308 55468 35364
rect 55524 35308 55534 35364
rect 22642 35196 22652 35252
rect 22708 35196 22988 35252
rect 23044 35196 23054 35252
rect 23426 35196 23436 35252
rect 23492 35196 29708 35252
rect 29764 35196 30268 35252
rect 30324 35196 30334 35252
rect 47954 35196 47964 35252
rect 48020 35196 52836 35252
rect 4610 35084 4620 35140
rect 4676 35084 4900 35140
rect 10322 35084 10332 35140
rect 10388 35084 11116 35140
rect 11172 35084 11182 35140
rect 15250 35084 15260 35140
rect 15316 35084 15326 35140
rect 16828 35084 24332 35140
rect 24388 35084 24398 35140
rect 24658 35084 24668 35140
rect 24724 35084 25676 35140
rect 25732 35084 25742 35140
rect 25890 35084 25900 35140
rect 25956 35084 25994 35140
rect 28578 35084 28588 35140
rect 28644 35084 29484 35140
rect 29540 35084 31276 35140
rect 31332 35084 31342 35140
rect 39554 35084 39564 35140
rect 39620 35084 40460 35140
rect 40516 35084 40526 35140
rect 52098 35084 52108 35140
rect 52164 35084 53676 35140
rect 53732 35084 53742 35140
rect 1810 34972 1820 35028
rect 1876 34972 3276 35028
rect 3332 34972 4844 35028
rect 4900 34972 4910 35028
rect 6748 34972 9884 35028
rect 9940 34972 9950 35028
rect 6748 34916 6804 34972
rect 15260 34916 15316 35084
rect 15446 34972 15484 35028
rect 15540 34972 15550 35028
rect 18844 34972 20188 35028
rect 20244 34972 32284 35028
rect 32340 34972 32350 35028
rect 33954 34972 33964 35028
rect 34020 34972 34412 35028
rect 34468 34972 34860 35028
rect 34916 34972 35644 35028
rect 35700 34972 35710 35028
rect 36418 34972 36428 35028
rect 36484 34972 45052 35028
rect 45108 34972 45118 35028
rect 51426 34972 51436 35028
rect 51492 34972 52500 35028
rect 53330 34972 53340 35028
rect 53396 34972 55132 35028
rect 55188 34972 55198 35028
rect 18844 34916 18900 34972
rect 52444 34916 52500 34972
rect 6066 34860 6076 34916
rect 6132 34860 6748 34916
rect 6804 34860 6814 34916
rect 7186 34860 7196 34916
rect 7252 34860 7756 34916
rect 7812 34860 8428 34916
rect 8484 34860 8494 34916
rect 9548 34860 11844 34916
rect 15260 34860 15372 34916
rect 15428 34860 15438 34916
rect 16230 34860 16268 34916
rect 16324 34860 16334 34916
rect 17490 34860 17500 34916
rect 17556 34860 18900 34916
rect 19506 34860 19516 34916
rect 19572 34860 19964 34916
rect 20020 34860 24332 34916
rect 24388 34860 24398 34916
rect 25666 34860 25676 34916
rect 25732 34860 26012 34916
rect 26068 34860 26078 34916
rect 26450 34860 26460 34916
rect 26516 34860 26796 34916
rect 26852 34860 27132 34916
rect 27188 34860 27198 34916
rect 28802 34860 28812 34916
rect 28868 34860 29148 34916
rect 29204 34860 29214 34916
rect 29362 34860 29372 34916
rect 29428 34860 30828 34916
rect 30884 34860 30894 34916
rect 37090 34860 37100 34916
rect 37156 34860 38220 34916
rect 38276 34860 40684 34916
rect 40740 34860 40750 34916
rect 41794 34860 41804 34916
rect 41860 34860 42700 34916
rect 42756 34860 42766 34916
rect 47058 34860 47068 34916
rect 47124 34860 47740 34916
rect 47796 34860 50428 34916
rect 50484 34860 52220 34916
rect 52276 34860 52286 34916
rect 52444 34860 53228 34916
rect 53284 34860 54684 34916
rect 54740 34860 54750 34916
rect 9548 34804 9604 34860
rect 11788 34804 11844 34860
rect 6962 34748 6972 34804
rect 7028 34748 7868 34804
rect 7924 34748 8204 34804
rect 8260 34748 9604 34804
rect 9986 34748 9996 34804
rect 10052 34748 10892 34804
rect 10948 34748 11564 34804
rect 11620 34748 11630 34804
rect 11788 34748 21084 34804
rect 21140 34748 21420 34804
rect 21476 34748 21486 34804
rect 21644 34692 21700 34860
rect 23874 34748 23884 34804
rect 23940 34748 24892 34804
rect 24948 34748 24958 34804
rect 31826 34748 31836 34804
rect 31892 34748 32620 34804
rect 32676 34748 33068 34804
rect 33124 34748 33134 34804
rect 40786 34748 40796 34804
rect 40852 34748 43484 34804
rect 43540 34748 43550 34804
rect 5282 34636 5292 34692
rect 5348 34636 7420 34692
rect 7476 34636 7486 34692
rect 10994 34636 11004 34692
rect 11060 34636 11788 34692
rect 11844 34636 14028 34692
rect 14084 34636 14094 34692
rect 14252 34636 18396 34692
rect 18452 34636 18462 34692
rect 20178 34636 20188 34692
rect 20244 34636 20412 34692
rect 20468 34636 20478 34692
rect 20626 34636 20636 34692
rect 20692 34636 21700 34692
rect 24098 34636 24108 34692
rect 24164 34636 25340 34692
rect 25396 34636 25406 34692
rect 26002 34636 26012 34692
rect 26068 34636 26908 34692
rect 26964 34636 27804 34692
rect 27860 34636 31052 34692
rect 31108 34636 31118 34692
rect 45378 34636 45388 34692
rect 45444 34636 45836 34692
rect 45892 34636 46284 34692
rect 46340 34636 46350 34692
rect 5058 34524 5068 34580
rect 5124 34524 13468 34580
rect 13524 34524 13534 34580
rect 14252 34468 14308 34636
rect 15586 34524 15596 34580
rect 15652 34524 16380 34580
rect 16436 34524 16446 34580
rect 21634 34524 21644 34580
rect 21700 34524 21980 34580
rect 22036 34524 22046 34580
rect 36754 34524 36764 34580
rect 36820 34524 43932 34580
rect 43988 34524 43998 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 10434 34412 10444 34468
rect 10500 34412 11564 34468
rect 11620 34412 11630 34468
rect 13570 34412 13580 34468
rect 13636 34412 14252 34468
rect 14308 34412 14318 34468
rect 14578 34412 14588 34468
rect 14644 34412 17612 34468
rect 17668 34412 17678 34468
rect 24210 34412 24220 34468
rect 24276 34412 30044 34468
rect 30100 34412 30110 34468
rect 13458 34300 13468 34356
rect 13524 34300 20188 34356
rect 20244 34300 20254 34356
rect 21634 34300 21644 34356
rect 21700 34300 22204 34356
rect 22260 34300 22270 34356
rect 48066 34300 48076 34356
rect 48132 34300 50204 34356
rect 50260 34300 51100 34356
rect 51156 34300 51166 34356
rect 16258 34188 16268 34244
rect 16324 34188 23884 34244
rect 23940 34188 23950 34244
rect 25666 34188 25676 34244
rect 25732 34188 26908 34244
rect 26964 34188 26974 34244
rect 31714 34188 31724 34244
rect 31780 34188 36204 34244
rect 36260 34188 37100 34244
rect 37156 34188 37166 34244
rect 37986 34188 37996 34244
rect 38052 34188 38062 34244
rect 50754 34188 50764 34244
rect 50820 34188 52108 34244
rect 52164 34188 52174 34244
rect 5954 34076 5964 34132
rect 6020 34076 7196 34132
rect 7252 34076 7262 34132
rect 10434 34076 10444 34132
rect 10500 34076 11004 34132
rect 11060 34076 11070 34132
rect 12786 34076 12796 34132
rect 12852 34076 13244 34132
rect 13300 34076 13310 34132
rect 14690 34076 14700 34132
rect 14756 34076 15148 34132
rect 15204 34076 16492 34132
rect 16548 34076 17500 34132
rect 17556 34076 17566 34132
rect 18386 34076 18396 34132
rect 18452 34076 22652 34132
rect 22708 34076 22718 34132
rect 30930 34076 30940 34132
rect 30996 34076 31948 34132
rect 32004 34076 32014 34132
rect 12796 34020 12852 34076
rect 37996 34020 38052 34188
rect 38658 34076 38668 34132
rect 38724 34076 42028 34132
rect 42084 34076 43036 34132
rect 43092 34076 43102 34132
rect 48402 34076 48412 34132
rect 48468 34076 50092 34132
rect 50148 34076 50158 34132
rect 50764 34020 50820 34188
rect 9874 33964 9884 34020
rect 9940 33964 12852 34020
rect 15474 33964 15484 34020
rect 15540 33964 18284 34020
rect 18340 33964 18350 34020
rect 20738 33964 20748 34020
rect 20804 33964 28588 34020
rect 28644 33964 30604 34020
rect 30660 33964 30670 34020
rect 33170 33964 33180 34020
rect 33236 33964 34300 34020
rect 34356 33964 34366 34020
rect 37996 33964 41132 34020
rect 41188 33964 41198 34020
rect 41906 33964 41916 34020
rect 41972 33964 50820 34020
rect 51548 33908 51604 34188
rect 52210 34076 52220 34132
rect 52276 34076 52780 34132
rect 52836 34076 53228 34132
rect 53284 34076 54012 34132
rect 54068 34076 54078 34132
rect 54674 33964 54684 34020
rect 54740 33964 56028 34020
rect 56084 33964 56094 34020
rect 2930 33852 2940 33908
rect 2996 33852 5068 33908
rect 5124 33852 5134 33908
rect 14802 33852 14812 33908
rect 14868 33852 16604 33908
rect 16660 33852 16670 33908
rect 17602 33852 17612 33908
rect 17668 33852 19740 33908
rect 19796 33852 20300 33908
rect 20356 33852 20366 33908
rect 24210 33852 24220 33908
rect 24276 33852 26012 33908
rect 26068 33852 26078 33908
rect 27010 33852 27020 33908
rect 27076 33852 27580 33908
rect 27636 33852 28364 33908
rect 28420 33852 28430 33908
rect 30930 33852 30940 33908
rect 30996 33852 32172 33908
rect 32228 33852 32238 33908
rect 39442 33852 39452 33908
rect 39508 33852 40236 33908
rect 40292 33852 42588 33908
rect 42644 33852 42654 33908
rect 43586 33852 43596 33908
rect 43652 33852 44604 33908
rect 44660 33852 44670 33908
rect 49074 33852 49084 33908
rect 49140 33852 50316 33908
rect 50372 33852 51324 33908
rect 51380 33852 51390 33908
rect 51538 33852 51548 33908
rect 51604 33852 51614 33908
rect 22642 33740 22652 33796
rect 22708 33740 26796 33796
rect 26852 33740 26862 33796
rect 30706 33740 30716 33796
rect 30772 33740 31500 33796
rect 31556 33740 31566 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 23986 33628 23996 33684
rect 24052 33628 26908 33684
rect 26964 33628 28476 33684
rect 28532 33628 28542 33684
rect 9314 33516 9324 33572
rect 9380 33516 20748 33572
rect 20804 33516 20814 33572
rect 21186 33516 21196 33572
rect 21252 33516 22092 33572
rect 22148 33516 22158 33572
rect 27794 33516 27804 33572
rect 27860 33516 28812 33572
rect 28868 33516 28878 33572
rect 45602 33516 45612 33572
rect 45668 33516 47404 33572
rect 47460 33516 47964 33572
rect 48020 33516 48030 33572
rect 19282 33404 19292 33460
rect 19348 33404 19964 33460
rect 20020 33404 20030 33460
rect 20290 33404 20300 33460
rect 20356 33404 27692 33460
rect 27748 33404 27758 33460
rect 28018 33404 28028 33460
rect 28084 33404 32508 33460
rect 32564 33404 32574 33460
rect 51874 33404 51884 33460
rect 51940 33404 52780 33460
rect 52836 33404 52846 33460
rect 14130 33292 14140 33348
rect 14196 33292 15036 33348
rect 15092 33292 15102 33348
rect 21634 33292 21644 33348
rect 21700 33292 25116 33348
rect 25172 33292 25182 33348
rect 27458 33292 27468 33348
rect 27524 33292 30604 33348
rect 30660 33292 30670 33348
rect 50306 33292 50316 33348
rect 50372 33292 50652 33348
rect 50708 33292 50718 33348
rect 18610 33180 18620 33236
rect 18676 33180 19068 33236
rect 19124 33180 19134 33236
rect 21746 33180 21756 33236
rect 21812 33180 23100 33236
rect 23156 33180 25900 33236
rect 25956 33180 26236 33236
rect 26292 33180 26302 33236
rect 26852 33180 27356 33236
rect 27412 33180 27422 33236
rect 27682 33180 27692 33236
rect 27748 33180 28252 33236
rect 28308 33180 29148 33236
rect 29204 33180 29214 33236
rect 32722 33180 32732 33236
rect 32788 33180 34300 33236
rect 34356 33180 34366 33236
rect 8530 33068 8540 33124
rect 8596 33068 13916 33124
rect 13972 33068 13982 33124
rect 15250 33068 15260 33124
rect 15316 33068 15596 33124
rect 15652 33068 15662 33124
rect 17154 33068 17164 33124
rect 17220 33068 17948 33124
rect 18004 33068 19180 33124
rect 19236 33068 19246 33124
rect 20738 33068 20748 33124
rect 20804 33068 21420 33124
rect 21476 33068 21486 33124
rect 22082 33068 22092 33124
rect 22148 33068 25452 33124
rect 25508 33068 25676 33124
rect 25732 33068 25742 33124
rect 26852 33012 26908 33180
rect 33618 33068 33628 33124
rect 33684 33068 34524 33124
rect 34580 33068 37100 33124
rect 37156 33068 37166 33124
rect 47842 33068 47852 33124
rect 47908 33068 49644 33124
rect 49700 33068 49710 33124
rect 50530 33068 50540 33124
rect 50596 33068 51436 33124
rect 51492 33068 51502 33124
rect 14662 32956 14700 33012
rect 14756 32956 14766 33012
rect 18274 32956 18284 33012
rect 18340 32956 19292 33012
rect 19348 32956 19358 33012
rect 24546 32956 24556 33012
rect 24612 32956 26908 33012
rect 33170 32956 33180 33012
rect 33236 32956 33740 33012
rect 33796 32956 34636 33012
rect 34692 32956 34702 33012
rect 46162 32956 46172 33012
rect 46228 32956 48860 33012
rect 48916 32956 48926 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 24658 32844 24668 32900
rect 24724 32844 25228 32900
rect 25284 32844 25294 32900
rect 4834 32732 4844 32788
rect 4900 32732 6524 32788
rect 6580 32732 6590 32788
rect 9090 32732 9100 32788
rect 9156 32732 13916 32788
rect 13972 32732 15820 32788
rect 15876 32732 17052 32788
rect 17108 32732 17388 32788
rect 17444 32732 17454 32788
rect 19506 32732 19516 32788
rect 19572 32732 20132 32788
rect 24210 32732 24220 32788
rect 24276 32732 24780 32788
rect 24836 32732 27020 32788
rect 27076 32732 27804 32788
rect 27860 32732 27870 32788
rect 29362 32732 29372 32788
rect 29428 32732 29438 32788
rect 32050 32732 32060 32788
rect 32116 32732 35196 32788
rect 35252 32732 35262 32788
rect 47506 32732 47516 32788
rect 47572 32732 48748 32788
rect 48804 32732 48814 32788
rect 51650 32732 51660 32788
rect 51716 32732 52108 32788
rect 52164 32732 52174 32788
rect 20076 32676 20132 32732
rect 29372 32676 29428 32732
rect 15586 32620 15596 32676
rect 15652 32620 16156 32676
rect 16212 32620 16940 32676
rect 16996 32620 17006 32676
rect 18162 32620 18172 32676
rect 18228 32620 18620 32676
rect 18676 32620 18686 32676
rect 19058 32620 19068 32676
rect 19124 32620 19134 32676
rect 20076 32620 24388 32676
rect 25442 32620 25452 32676
rect 25508 32620 27692 32676
rect 27748 32620 29428 32676
rect 36418 32620 36428 32676
rect 36484 32620 37212 32676
rect 37268 32620 37660 32676
rect 37716 32620 37726 32676
rect 19068 32452 19124 32620
rect 24332 32564 24388 32620
rect 20962 32508 20972 32564
rect 21028 32508 22204 32564
rect 22260 32508 22270 32564
rect 24322 32508 24332 32564
rect 24388 32508 24780 32564
rect 24836 32508 24846 32564
rect 25106 32508 25116 32564
rect 25172 32508 25788 32564
rect 25844 32508 25854 32564
rect 26114 32508 26124 32564
rect 26180 32508 28588 32564
rect 28644 32508 28654 32564
rect 29250 32508 29260 32564
rect 29316 32508 30828 32564
rect 30884 32508 30894 32564
rect 31826 32508 31836 32564
rect 31892 32508 33068 32564
rect 33124 32508 33134 32564
rect 41458 32508 41468 32564
rect 41524 32508 42140 32564
rect 42196 32508 42206 32564
rect 45378 32508 45388 32564
rect 45444 32508 46732 32564
rect 46788 32508 46798 32564
rect 51650 32508 51660 32564
rect 51716 32508 54236 32564
rect 54292 32508 54302 32564
rect 6738 32396 6748 32452
rect 6804 32396 15372 32452
rect 15428 32396 15438 32452
rect 15810 32396 15820 32452
rect 15876 32396 17948 32452
rect 18004 32396 18014 32452
rect 18610 32396 18620 32452
rect 18676 32396 19124 32452
rect 21298 32396 21308 32452
rect 21364 32396 21980 32452
rect 22036 32396 22046 32452
rect 24994 32396 25004 32452
rect 25060 32396 29820 32452
rect 29876 32396 29886 32452
rect 31602 32396 31612 32452
rect 31668 32396 31948 32452
rect 32004 32396 32396 32452
rect 32452 32396 32462 32452
rect 46498 32396 46508 32452
rect 46564 32396 48860 32452
rect 48916 32396 48926 32452
rect 52098 32396 52108 32452
rect 52164 32396 52780 32452
rect 52836 32396 52846 32452
rect 18834 32284 18844 32340
rect 18900 32284 20748 32340
rect 20804 32284 20814 32340
rect 31378 32284 31388 32340
rect 31444 32284 33628 32340
rect 33684 32284 43708 32340
rect 47170 32284 47180 32340
rect 47236 32284 49420 32340
rect 49476 32284 49486 32340
rect 29810 32172 29820 32228
rect 29876 32172 30716 32228
rect 30772 32172 31164 32228
rect 31220 32172 31230 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 15334 32060 15372 32116
rect 15428 32060 21644 32116
rect 21700 32060 21710 32116
rect 21970 32060 21980 32116
rect 22036 32060 23772 32116
rect 23828 32060 23838 32116
rect 43652 32004 43708 32284
rect 47394 32172 47404 32228
rect 47460 32172 48636 32228
rect 48692 32172 49980 32228
rect 50036 32172 50046 32228
rect 50372 32172 51996 32228
rect 52052 32172 55916 32228
rect 55972 32172 55982 32228
rect 50372 32004 50428 32172
rect 8316 31948 8764 32004
rect 8820 31948 9660 32004
rect 9716 31948 10892 32004
rect 10948 31948 11228 32004
rect 11284 31948 11294 32004
rect 12002 31948 12012 32004
rect 12068 31948 18620 32004
rect 18676 31948 18686 32004
rect 24546 31948 24556 32004
rect 24612 31948 25900 32004
rect 25956 31948 25966 32004
rect 30594 31948 30604 32004
rect 30660 31948 32060 32004
rect 32116 31948 32126 32004
rect 43652 31948 45388 32004
rect 45444 31948 45454 32004
rect 48962 31948 48972 32004
rect 49028 31948 50428 32004
rect 8316 31892 8372 31948
rect 6514 31836 6524 31892
rect 6580 31836 7756 31892
rect 7812 31836 8204 31892
rect 8260 31836 8372 31892
rect 10546 31836 10556 31892
rect 10612 31836 11452 31892
rect 11508 31836 11518 31892
rect 21186 31836 21196 31892
rect 21252 31836 21868 31892
rect 21924 31836 21934 31892
rect 22418 31836 22428 31892
rect 22484 31836 23548 31892
rect 23604 31836 23614 31892
rect 41346 31836 41356 31892
rect 41412 31836 43596 31892
rect 43652 31836 43662 31892
rect 45490 31836 45500 31892
rect 45556 31836 48188 31892
rect 48244 31836 49196 31892
rect 49252 31836 49262 31892
rect 51314 31836 51324 31892
rect 51380 31836 52668 31892
rect 52724 31836 52734 31892
rect 12226 31724 12236 31780
rect 12292 31724 13020 31780
rect 13076 31724 13468 31780
rect 13524 31724 13534 31780
rect 14812 31724 15036 31780
rect 15092 31724 15102 31780
rect 16034 31724 16044 31780
rect 16100 31724 16604 31780
rect 16660 31724 16670 31780
rect 18386 31724 18396 31780
rect 18452 31724 20412 31780
rect 20468 31724 20478 31780
rect 20738 31724 20748 31780
rect 20804 31724 22540 31780
rect 22596 31724 22606 31780
rect 23202 31724 23212 31780
rect 23268 31724 25340 31780
rect 25396 31724 25406 31780
rect 25890 31724 25900 31780
rect 25956 31724 27020 31780
rect 27076 31724 27356 31780
rect 27412 31724 27422 31780
rect 27906 31724 27916 31780
rect 27972 31724 28252 31780
rect 28308 31724 29260 31780
rect 29316 31724 29326 31780
rect 30034 31724 30044 31780
rect 30100 31724 30492 31780
rect 30548 31724 33068 31780
rect 33124 31724 34188 31780
rect 34244 31724 34254 31780
rect 36978 31724 36988 31780
rect 37044 31724 38780 31780
rect 38836 31724 38846 31780
rect 39330 31724 39340 31780
rect 39396 31724 40236 31780
rect 40292 31724 40302 31780
rect 49970 31724 49980 31780
rect 50036 31724 51212 31780
rect 51268 31724 51772 31780
rect 51828 31724 51838 31780
rect 14812 31668 14868 31724
rect 14018 31612 14028 31668
rect 14084 31612 14812 31668
rect 14868 31612 14878 31668
rect 15092 31612 19628 31668
rect 19684 31612 19694 31668
rect 21074 31612 21084 31668
rect 21140 31612 22652 31668
rect 22708 31612 22718 31668
rect 22866 31612 22876 31668
rect 22932 31612 26236 31668
rect 26292 31612 26302 31668
rect 26852 31612 29148 31668
rect 29204 31612 29214 31668
rect 34402 31612 34412 31668
rect 34468 31612 37660 31668
rect 37716 31612 38108 31668
rect 38164 31612 38174 31668
rect 38882 31612 38892 31668
rect 38948 31612 39676 31668
rect 39732 31612 39742 31668
rect 49634 31612 49644 31668
rect 49700 31612 51548 31668
rect 51604 31612 51614 31668
rect 15092 31556 15148 31612
rect 26852 31556 26908 31612
rect 13906 31500 13916 31556
rect 13972 31500 15148 31556
rect 15250 31500 15260 31556
rect 15316 31500 16268 31556
rect 16324 31500 16334 31556
rect 17378 31500 17388 31556
rect 17444 31500 20188 31556
rect 20244 31500 20254 31556
rect 26562 31500 26572 31556
rect 26628 31500 26908 31556
rect 29474 31500 29484 31556
rect 29540 31500 33292 31556
rect 33348 31500 33358 31556
rect 37314 31500 37324 31556
rect 37380 31500 37884 31556
rect 37940 31500 41356 31556
rect 41412 31500 41422 31556
rect 44258 31500 44268 31556
rect 44324 31500 44940 31556
rect 44996 31500 45388 31556
rect 45444 31500 45836 31556
rect 45892 31500 45902 31556
rect 50530 31500 50540 31556
rect 50596 31500 52108 31556
rect 52164 31500 52174 31556
rect 10546 31388 10556 31444
rect 10612 31388 11116 31444
rect 11172 31388 18284 31444
rect 18340 31388 18350 31444
rect 24546 31388 24556 31444
rect 24612 31388 25004 31444
rect 25060 31388 25788 31444
rect 25844 31388 27468 31444
rect 27524 31388 28028 31444
rect 28084 31388 28094 31444
rect 39778 31388 39788 31444
rect 39844 31388 41244 31444
rect 41300 31388 41310 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 7858 31276 7868 31332
rect 7924 31276 11340 31332
rect 11396 31276 16044 31332
rect 16100 31276 16110 31332
rect 23314 31276 23324 31332
rect 23380 31276 24444 31332
rect 24500 31276 27132 31332
rect 27188 31276 27198 31332
rect 10322 31164 10332 31220
rect 10388 31164 12460 31220
rect 12516 31164 17388 31220
rect 17444 31164 17454 31220
rect 18050 31164 18060 31220
rect 18116 31164 21084 31220
rect 21140 31164 21150 31220
rect 21298 31164 21308 31220
rect 21364 31164 24892 31220
rect 24948 31164 24958 31220
rect 25330 31164 25340 31220
rect 25396 31164 26460 31220
rect 26516 31164 26526 31220
rect 37538 31164 37548 31220
rect 37604 31164 39228 31220
rect 39284 31164 40236 31220
rect 40292 31164 40302 31220
rect 41122 31164 41132 31220
rect 41188 31164 42140 31220
rect 42196 31164 42206 31220
rect 50866 31164 50876 31220
rect 50932 31164 51996 31220
rect 52052 31164 52062 31220
rect 15138 31052 15148 31108
rect 15204 31052 15708 31108
rect 15764 31052 16604 31108
rect 16660 31052 17612 31108
rect 17668 31052 17678 31108
rect 21186 31052 21196 31108
rect 21252 31052 22764 31108
rect 22820 31052 22830 31108
rect 32386 31052 32396 31108
rect 32452 31052 33964 31108
rect 34020 31052 34030 31108
rect 37314 31052 37324 31108
rect 37380 31052 38220 31108
rect 38276 31052 38892 31108
rect 38948 31052 38958 31108
rect 40786 31052 40796 31108
rect 40852 31052 41692 31108
rect 41748 31052 42364 31108
rect 42420 31052 42430 31108
rect 11106 30940 11116 30996
rect 11172 30940 12012 30996
rect 12068 30940 12078 30996
rect 12562 30940 12572 30996
rect 12628 30940 13916 30996
rect 13972 30940 13982 30996
rect 16258 30940 16268 30996
rect 16324 30940 18396 30996
rect 18452 30940 18462 30996
rect 19618 30940 19628 30996
rect 19684 30940 20972 30996
rect 21028 30940 23996 30996
rect 24052 30940 24062 30996
rect 29474 30940 29484 30996
rect 29540 30940 30940 30996
rect 30996 30940 31006 30996
rect 49756 30940 50652 30996
rect 50708 30940 50718 30996
rect 49756 30884 49812 30940
rect 8978 30828 8988 30884
rect 9044 30828 14028 30884
rect 14084 30828 14094 30884
rect 19394 30828 19404 30884
rect 19460 30828 29820 30884
rect 29876 30828 29886 30884
rect 39778 30828 39788 30884
rect 39844 30828 40348 30884
rect 40404 30828 40414 30884
rect 49186 30828 49196 30884
rect 49252 30828 49756 30884
rect 49812 30828 49822 30884
rect 49970 30828 49980 30884
rect 50036 30828 50540 30884
rect 50596 30828 50606 30884
rect 7298 30716 7308 30772
rect 7364 30716 10220 30772
rect 10276 30716 10286 30772
rect 12338 30716 12348 30772
rect 12404 30716 17164 30772
rect 17220 30716 17230 30772
rect 20514 30716 20524 30772
rect 20580 30716 21868 30772
rect 21924 30716 23100 30772
rect 23156 30716 23166 30772
rect 23314 30716 23324 30772
rect 23380 30716 24332 30772
rect 24388 30716 24892 30772
rect 24948 30716 24958 30772
rect 12786 30604 12796 30660
rect 12852 30604 13804 30660
rect 13860 30604 13870 30660
rect 15026 30604 15036 30660
rect 15092 30604 20188 30660
rect 20244 30604 20254 30660
rect 24210 30604 24220 30660
rect 24276 30604 24286 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 24220 30548 24276 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 13122 30492 13132 30548
rect 13188 30492 13692 30548
rect 13748 30492 15596 30548
rect 15652 30492 15662 30548
rect 18386 30492 18396 30548
rect 18452 30492 24276 30548
rect 14242 30380 14252 30436
rect 14308 30380 14924 30436
rect 14980 30380 14990 30436
rect 33394 30380 33404 30436
rect 33460 30380 34748 30436
rect 34804 30380 34814 30436
rect 40002 30380 40012 30436
rect 40068 30380 40908 30436
rect 40964 30380 40974 30436
rect 9202 30268 9212 30324
rect 9268 30268 11452 30324
rect 11508 30268 12852 30324
rect 15026 30268 15036 30324
rect 15092 30268 15260 30324
rect 15316 30268 15326 30324
rect 15484 30268 15708 30324
rect 15764 30268 15774 30324
rect 18498 30268 18508 30324
rect 18564 30268 18956 30324
rect 19012 30268 21196 30324
rect 21252 30268 21262 30324
rect 24882 30268 24892 30324
rect 24948 30268 26684 30324
rect 26740 30268 26750 30324
rect 30930 30268 30940 30324
rect 30996 30268 33180 30324
rect 33236 30268 34636 30324
rect 34692 30268 35476 30324
rect 38210 30268 38220 30324
rect 38276 30268 39228 30324
rect 39284 30268 39294 30324
rect 40338 30268 40348 30324
rect 40404 30268 41244 30324
rect 41300 30268 41310 30324
rect 12796 30212 12852 30268
rect 12786 30156 12796 30212
rect 12852 30156 12862 30212
rect 14130 30156 14140 30212
rect 14196 30156 14206 30212
rect 14140 30100 14196 30156
rect 15484 30100 15540 30268
rect 35420 30212 35476 30268
rect 17490 30156 17500 30212
rect 17556 30156 18172 30212
rect 18228 30156 18238 30212
rect 18610 30156 18620 30212
rect 18676 30156 19068 30212
rect 19124 30156 19134 30212
rect 21522 30156 21532 30212
rect 21588 30156 23548 30212
rect 23604 30156 23614 30212
rect 25218 30156 25228 30212
rect 25284 30156 26348 30212
rect 26404 30156 26414 30212
rect 30370 30156 30380 30212
rect 30436 30156 33068 30212
rect 33124 30156 33134 30212
rect 35410 30156 35420 30212
rect 35476 30156 35486 30212
rect 37874 30156 37884 30212
rect 37940 30156 38780 30212
rect 38836 30156 38846 30212
rect 45826 30156 45836 30212
rect 45892 30156 48860 30212
rect 48916 30156 49308 30212
rect 49364 30156 49374 30212
rect 25228 30100 25284 30156
rect 11554 30044 11564 30100
rect 11620 30044 13468 30100
rect 13524 30044 14196 30100
rect 14690 30044 14700 30100
rect 14756 30044 15540 30100
rect 19842 30044 19852 30100
rect 19908 30044 22428 30100
rect 22484 30044 22494 30100
rect 22642 30044 22652 30100
rect 22708 30044 25284 30100
rect 34290 30044 34300 30100
rect 34356 30044 35868 30100
rect 35924 30044 35934 30100
rect 36418 30044 36428 30100
rect 36484 30044 37772 30100
rect 37828 30044 37838 30100
rect 40908 30044 41468 30100
rect 41524 30044 41534 30100
rect 40908 29988 40964 30044
rect 1586 29932 1596 29988
rect 1652 29932 28700 29988
rect 28756 29932 28766 29988
rect 33282 29932 33292 29988
rect 33348 29932 34860 29988
rect 34916 29932 34926 29988
rect 35074 29932 35084 29988
rect 35140 29932 40908 29988
rect 40964 29932 40974 29988
rect 41346 29932 41356 29988
rect 41412 29932 43372 29988
rect 43428 29932 43438 29988
rect 14466 29820 14476 29876
rect 14532 29820 17836 29876
rect 17892 29820 19292 29876
rect 19348 29820 19358 29876
rect 32610 29820 32620 29876
rect 32676 29820 34972 29876
rect 35028 29820 35038 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 14802 29708 14812 29764
rect 14868 29708 15932 29764
rect 15988 29708 15998 29764
rect 12002 29596 12012 29652
rect 12068 29596 13356 29652
rect 13412 29596 13422 29652
rect 15138 29596 15148 29652
rect 15204 29596 17948 29652
rect 18004 29596 18014 29652
rect 18274 29596 18284 29652
rect 18340 29596 18620 29652
rect 18676 29596 18956 29652
rect 19012 29596 21308 29652
rect 21364 29596 21374 29652
rect 27234 29596 27244 29652
rect 27300 29596 31948 29652
rect 32004 29596 32014 29652
rect 37314 29596 37324 29652
rect 37380 29596 38556 29652
rect 38612 29596 40292 29652
rect 15026 29484 15036 29540
rect 15092 29484 16156 29540
rect 16212 29484 16222 29540
rect 19954 29484 19964 29540
rect 20020 29484 20188 29540
rect 20244 29484 20254 29540
rect 20514 29484 20524 29540
rect 20580 29484 20860 29540
rect 20916 29484 20926 29540
rect 23650 29484 23660 29540
rect 23716 29484 25340 29540
rect 25396 29484 25406 29540
rect 28690 29484 28700 29540
rect 28756 29484 29596 29540
rect 29652 29484 29662 29540
rect 32274 29484 32284 29540
rect 32340 29484 36316 29540
rect 36372 29484 37100 29540
rect 37156 29484 38780 29540
rect 38836 29484 38846 29540
rect 40236 29428 40292 29596
rect 12786 29372 12796 29428
rect 12852 29372 13804 29428
rect 13860 29372 13870 29428
rect 15810 29372 15820 29428
rect 15876 29372 16716 29428
rect 16772 29372 17500 29428
rect 17556 29372 17566 29428
rect 26898 29372 26908 29428
rect 26964 29372 27804 29428
rect 27860 29372 27870 29428
rect 32498 29372 32508 29428
rect 32564 29372 32844 29428
rect 32900 29372 33628 29428
rect 33684 29372 33694 29428
rect 35858 29372 35868 29428
rect 35924 29372 39564 29428
rect 39620 29372 39630 29428
rect 40226 29372 40236 29428
rect 40292 29372 42476 29428
rect 42532 29372 42542 29428
rect 5170 29260 5180 29316
rect 5236 29260 6188 29316
rect 6244 29260 6748 29316
rect 6804 29260 8204 29316
rect 8260 29260 9772 29316
rect 9828 29260 9838 29316
rect 14242 29260 14252 29316
rect 14308 29260 20300 29316
rect 20356 29260 22540 29316
rect 22596 29260 22606 29316
rect 25218 29260 25228 29316
rect 25284 29260 25452 29316
rect 25508 29260 25900 29316
rect 25956 29260 26460 29316
rect 26516 29260 26526 29316
rect 33394 29260 33404 29316
rect 33460 29260 36988 29316
rect 37044 29260 37324 29316
rect 37380 29260 37390 29316
rect 12450 29148 12460 29204
rect 12516 29148 15708 29204
rect 15764 29148 15774 29204
rect 24434 29148 24444 29204
rect 24500 29148 30828 29204
rect 30884 29148 30894 29204
rect 38658 29148 38668 29204
rect 38724 29148 40124 29204
rect 40180 29148 40190 29204
rect 6514 29036 6524 29092
rect 6580 29036 6972 29092
rect 7028 29036 28364 29092
rect 28420 29036 28430 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 13458 28924 13468 28980
rect 13524 28924 13804 28980
rect 13860 28924 14756 28980
rect 14700 28868 14756 28924
rect 13346 28812 13356 28868
rect 13412 28812 14476 28868
rect 14532 28812 14542 28868
rect 14690 28812 14700 28868
rect 14756 28812 26908 28868
rect 39218 28812 39228 28868
rect 39284 28812 39452 28868
rect 39508 28812 41244 28868
rect 41300 28812 42140 28868
rect 42196 28812 42206 28868
rect 42802 28812 42812 28868
rect 42868 28812 44044 28868
rect 44100 28812 44110 28868
rect 26852 28756 26908 28812
rect 17948 28700 18732 28756
rect 18788 28700 19516 28756
rect 19572 28700 20636 28756
rect 20692 28700 21532 28756
rect 21588 28700 21598 28756
rect 26852 28700 27468 28756
rect 27524 28700 27534 28756
rect 29922 28700 29932 28756
rect 29988 28700 29998 28756
rect 38434 28700 38444 28756
rect 38500 28700 39116 28756
rect 39172 28700 39676 28756
rect 39732 28700 39742 28756
rect 13234 28588 13244 28644
rect 13300 28588 13468 28644
rect 13524 28588 13534 28644
rect 17042 28588 17052 28644
rect 17108 28588 17724 28644
rect 17780 28588 17790 28644
rect 14354 28476 14364 28532
rect 14420 28476 16044 28532
rect 16100 28476 16110 28532
rect 16268 28476 17276 28532
rect 17332 28476 17342 28532
rect 16268 28420 16324 28476
rect 17948 28420 18004 28700
rect 29932 28644 29988 28700
rect 18162 28588 18172 28644
rect 18228 28588 19068 28644
rect 19124 28588 19134 28644
rect 19394 28588 19404 28644
rect 19460 28588 19964 28644
rect 20020 28588 20030 28644
rect 29932 28588 30604 28644
rect 30660 28588 32620 28644
rect 32676 28588 32686 28644
rect 40114 28588 40124 28644
rect 40180 28588 41916 28644
rect 41972 28588 41982 28644
rect 40124 28532 40180 28588
rect 18610 28476 18620 28532
rect 18676 28476 20188 28532
rect 20244 28476 20254 28532
rect 21410 28476 21420 28532
rect 21476 28476 22428 28532
rect 22484 28476 23324 28532
rect 23380 28476 23390 28532
rect 35522 28476 35532 28532
rect 35588 28476 36428 28532
rect 36484 28476 36494 28532
rect 37314 28476 37324 28532
rect 37380 28476 40180 28532
rect 42214 28476 42252 28532
rect 42308 28476 42318 28532
rect 14018 28364 14028 28420
rect 14084 28364 16324 28420
rect 16482 28364 16492 28420
rect 16548 28364 17724 28420
rect 17780 28364 17790 28420
rect 17938 28364 17948 28420
rect 18004 28364 18014 28420
rect 18172 28364 21868 28420
rect 21924 28364 24444 28420
rect 24500 28364 24510 28420
rect 32498 28364 32508 28420
rect 32564 28364 33852 28420
rect 33908 28364 33918 28420
rect 37426 28364 37436 28420
rect 37492 28364 39676 28420
rect 39732 28364 39742 28420
rect 18172 28308 18228 28364
rect 16034 28252 16044 28308
rect 16100 28252 18228 28308
rect 22530 28252 22540 28308
rect 22596 28252 23324 28308
rect 23380 28252 23390 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 16146 28140 16156 28196
rect 16212 28140 19628 28196
rect 19684 28140 19694 28196
rect 12898 28028 12908 28084
rect 12964 28028 15148 28084
rect 17938 28028 17948 28084
rect 18004 28028 24780 28084
rect 24836 28028 25452 28084
rect 25508 28028 35084 28084
rect 35140 28028 35150 28084
rect 36978 28028 36988 28084
rect 37044 28028 38556 28084
rect 38612 28028 39788 28084
rect 39844 28028 39854 28084
rect 9650 27916 9660 27972
rect 9716 27916 10220 27972
rect 10276 27916 10286 27972
rect 7746 27804 7756 27860
rect 7812 27804 8428 27860
rect 8484 27804 9884 27860
rect 9940 27804 9950 27860
rect 10546 27804 10556 27860
rect 10612 27804 13580 27860
rect 13636 27804 14700 27860
rect 14756 27804 14766 27860
rect 15092 27748 15148 28028
rect 30146 27916 30156 27972
rect 30212 27916 30716 27972
rect 30772 27916 32060 27972
rect 32116 27916 32126 27972
rect 38322 27916 38332 27972
rect 38388 27916 40124 27972
rect 40180 27916 41804 27972
rect 41860 27916 41870 27972
rect 22866 27804 22876 27860
rect 22932 27804 23436 27860
rect 23492 27804 24108 27860
rect 24164 27804 24668 27860
rect 24724 27804 24734 27860
rect 32274 27804 32284 27860
rect 32340 27804 32844 27860
rect 32900 27804 32910 27860
rect 15092 27692 15596 27748
rect 15652 27692 16380 27748
rect 16436 27692 16446 27748
rect 35970 27692 35980 27748
rect 36036 27692 39340 27748
rect 39396 27692 40236 27748
rect 40292 27692 40684 27748
rect 40740 27692 40750 27748
rect 7970 27580 7980 27636
rect 8036 27580 13020 27636
rect 13076 27580 14364 27636
rect 14420 27580 14430 27636
rect 37202 27580 37212 27636
rect 37268 27580 39788 27636
rect 39844 27580 39854 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 6514 27356 6524 27412
rect 6580 27356 9548 27412
rect 9604 27356 24332 27412
rect 24388 27356 25228 27412
rect 25284 27356 25294 27412
rect 36418 27356 36428 27412
rect 36484 27356 36764 27412
rect 36820 27356 38668 27412
rect 38612 27188 38668 27356
rect 15474 27132 15484 27188
rect 15540 27132 15820 27188
rect 15876 27132 15886 27188
rect 35522 27132 35532 27188
rect 35588 27132 37436 27188
rect 37492 27132 37502 27188
rect 38612 27132 40460 27188
rect 40516 27132 40908 27188
rect 40964 27132 40974 27188
rect 11116 27020 12236 27076
rect 12292 27020 13132 27076
rect 13188 27020 13198 27076
rect 14242 27020 14252 27076
rect 14308 27020 15036 27076
rect 15092 27020 15102 27076
rect 17826 27020 17836 27076
rect 17892 27020 17902 27076
rect 29250 27020 29260 27076
rect 29316 27020 32396 27076
rect 32452 27020 32462 27076
rect 41122 27020 41132 27076
rect 41188 27020 42140 27076
rect 42196 27020 42206 27076
rect 11116 26964 11172 27020
rect 17836 26964 17892 27020
rect 7634 26908 7644 26964
rect 7700 26908 8540 26964
rect 8596 26908 9996 26964
rect 10052 26908 10062 26964
rect 11106 26908 11116 26964
rect 11172 26908 11182 26964
rect 17836 26908 18060 26964
rect 18116 26908 18126 26964
rect 21868 26908 22428 26964
rect 22484 26908 22494 26964
rect 37090 26908 37100 26964
rect 37156 26908 37772 26964
rect 37828 26908 37838 26964
rect 41234 26908 41244 26964
rect 41300 26908 42476 26964
rect 42532 26908 42542 26964
rect 21868 26852 21924 26908
rect 17826 26796 17836 26852
rect 17892 26796 20524 26852
rect 20580 26796 21924 26852
rect 36866 26684 36876 26740
rect 36932 26684 37436 26740
rect 37492 26684 37502 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 15810 26460 15820 26516
rect 15876 26460 22092 26516
rect 22148 26460 22158 26516
rect 39890 26460 39900 26516
rect 39956 26460 41132 26516
rect 41188 26460 41198 26516
rect 11330 26348 11340 26404
rect 11396 26348 12236 26404
rect 12292 26348 12302 26404
rect 15138 26348 15148 26404
rect 15204 26348 19180 26404
rect 19236 26348 19852 26404
rect 19908 26348 19918 26404
rect 3490 26236 3500 26292
rect 3556 26236 4956 26292
rect 5012 26236 5022 26292
rect 7298 26236 7308 26292
rect 7364 26236 7756 26292
rect 7812 26236 7822 26292
rect 8754 26236 8764 26292
rect 8820 26236 9436 26292
rect 9492 26236 10108 26292
rect 10164 26236 10174 26292
rect 14130 26236 14140 26292
rect 14196 26236 14476 26292
rect 14532 26236 15260 26292
rect 15316 26236 15326 26292
rect 16706 26236 16716 26292
rect 16772 26236 17388 26292
rect 17444 26236 17454 26292
rect 18274 26236 18284 26292
rect 18340 26236 18844 26292
rect 18900 26236 18910 26292
rect 40674 26236 40684 26292
rect 40740 26236 41804 26292
rect 41860 26236 41870 26292
rect 4162 26124 4172 26180
rect 4228 26124 5628 26180
rect 5684 26124 5694 26180
rect 5954 26124 5964 26180
rect 6020 26124 9660 26180
rect 9716 26124 9726 26180
rect 16594 26124 16604 26180
rect 16660 26124 30716 26180
rect 30772 26124 31612 26180
rect 31668 26124 31678 26180
rect 6962 26012 6972 26068
rect 7028 26012 9548 26068
rect 9604 26012 9614 26068
rect 14914 26012 14924 26068
rect 14980 26012 15484 26068
rect 15540 26012 15550 26068
rect 18274 26012 18284 26068
rect 18340 26012 19068 26068
rect 19124 26012 19134 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 7634 25564 7644 25620
rect 7700 25564 10332 25620
rect 10388 25564 10398 25620
rect 39442 25564 39452 25620
rect 39508 25564 40684 25620
rect 40740 25564 40750 25620
rect 6290 25452 6300 25508
rect 6356 25452 7308 25508
rect 7364 25452 9324 25508
rect 9380 25452 9390 25508
rect 14130 25452 14140 25508
rect 14196 25452 14700 25508
rect 14756 25452 14766 25508
rect 7410 25340 7420 25396
rect 7476 25340 7980 25396
rect 8036 25340 8764 25396
rect 8820 25340 8830 25396
rect 17042 25340 17052 25396
rect 17108 25340 17500 25396
rect 17556 25340 20300 25396
rect 20356 25340 20366 25396
rect 13682 25228 13692 25284
rect 13748 25228 14588 25284
rect 14644 25228 14654 25284
rect 16034 25228 16044 25284
rect 16100 25228 16268 25284
rect 16324 25228 16334 25284
rect 24658 25228 24668 25284
rect 24724 25228 25340 25284
rect 25396 25228 25788 25284
rect 25844 25228 25854 25284
rect 11890 25116 11900 25172
rect 11956 25116 13356 25172
rect 13412 25116 13422 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 7634 25004 7644 25060
rect 7700 25004 9548 25060
rect 9604 25004 11452 25060
rect 11508 25004 13804 25060
rect 13860 25004 13870 25060
rect 8418 24892 8428 24948
rect 8484 24892 9212 24948
rect 9268 24892 10780 24948
rect 10836 24892 10846 24948
rect 10322 24780 10332 24836
rect 10388 24780 10668 24836
rect 10724 24780 10734 24836
rect 13010 24780 13020 24836
rect 13076 24780 14588 24836
rect 14644 24780 14654 24836
rect 16818 24780 16828 24836
rect 16884 24780 19348 24836
rect 32498 24780 32508 24836
rect 32564 24780 33852 24836
rect 33908 24780 33918 24836
rect 19292 24724 19348 24780
rect 16034 24668 16044 24724
rect 16100 24668 17612 24724
rect 17668 24668 19068 24724
rect 19124 24668 19134 24724
rect 19282 24668 19292 24724
rect 19348 24668 19628 24724
rect 19684 24668 20748 24724
rect 20804 24668 20814 24724
rect 14802 24556 14812 24612
rect 14868 24556 18284 24612
rect 18340 24556 18350 24612
rect 34850 24556 34860 24612
rect 34916 24556 35980 24612
rect 36036 24556 36046 24612
rect 8642 24444 8652 24500
rect 8708 24444 12348 24500
rect 12404 24444 12414 24500
rect 17826 24444 17836 24500
rect 17892 24444 18732 24500
rect 18788 24444 18798 24500
rect 12226 24332 12236 24388
rect 12292 24332 12908 24388
rect 12964 24332 12974 24388
rect 16146 24332 16156 24388
rect 16212 24332 16492 24388
rect 16548 24332 16558 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 18498 24220 18508 24276
rect 18564 24220 20076 24276
rect 20132 24220 20860 24276
rect 20916 24220 20926 24276
rect 8530 24108 8540 24164
rect 8596 24108 9324 24164
rect 9380 24108 9390 24164
rect 16230 24108 16268 24164
rect 16324 24108 16334 24164
rect 14018 23996 14028 24052
rect 14084 23996 16044 24052
rect 16100 23996 16110 24052
rect 26450 23996 26460 24052
rect 26516 23996 27804 24052
rect 27860 23996 27870 24052
rect 15810 23884 15820 23940
rect 15876 23884 18060 23940
rect 18116 23884 18126 23940
rect 18722 23884 18732 23940
rect 18788 23884 20412 23940
rect 20468 23884 20478 23940
rect 32386 23884 32396 23940
rect 32452 23884 33852 23940
rect 33908 23884 33918 23940
rect 7074 23772 7084 23828
rect 7140 23772 8428 23828
rect 8484 23772 9212 23828
rect 9268 23772 9278 23828
rect 10770 23772 10780 23828
rect 10836 23772 14476 23828
rect 14532 23772 14542 23828
rect 15922 23772 15932 23828
rect 15988 23772 20188 23828
rect 20244 23772 20972 23828
rect 21028 23772 21308 23828
rect 21364 23772 21374 23828
rect 21746 23772 21756 23828
rect 21812 23772 23548 23828
rect 23604 23772 23614 23828
rect 27122 23772 27132 23828
rect 27188 23772 27692 23828
rect 27748 23772 28812 23828
rect 28868 23772 28878 23828
rect 33170 23772 33180 23828
rect 33236 23772 34860 23828
rect 34916 23772 34926 23828
rect 36082 23772 36092 23828
rect 36148 23772 37772 23828
rect 37828 23772 37838 23828
rect 3938 23660 3948 23716
rect 4004 23660 5852 23716
rect 5908 23660 5918 23716
rect 12338 23660 12348 23716
rect 12404 23660 13468 23716
rect 13524 23660 13534 23716
rect 23202 23660 23212 23716
rect 23268 23660 23996 23716
rect 24052 23660 24668 23716
rect 24724 23660 24734 23716
rect 7298 23548 7308 23604
rect 7364 23548 7374 23604
rect 20402 23548 20412 23604
rect 20468 23548 20748 23604
rect 20804 23548 21532 23604
rect 21588 23548 21598 23604
rect 7308 23492 7364 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 6514 23436 6524 23492
rect 6580 23436 7364 23492
rect 7858 23436 7868 23492
rect 7924 23436 10332 23492
rect 10388 23436 10398 23492
rect 21410 23436 21420 23492
rect 21476 23436 32620 23492
rect 32676 23436 33740 23492
rect 33796 23436 33806 23492
rect 5954 23324 5964 23380
rect 6020 23324 7532 23380
rect 7588 23324 7598 23380
rect 7970 23324 7980 23380
rect 8036 23324 8046 23380
rect 10882 23324 10892 23380
rect 10948 23324 14140 23380
rect 14196 23324 14206 23380
rect 20626 23324 20636 23380
rect 20692 23324 21644 23380
rect 21700 23324 21710 23380
rect 24770 23324 24780 23380
rect 24836 23324 25564 23380
rect 25620 23324 25630 23380
rect 7980 23268 8036 23324
rect 7410 23212 7420 23268
rect 7476 23212 8036 23268
rect 32050 23212 32060 23268
rect 32116 23212 33180 23268
rect 33236 23212 33246 23268
rect 3266 23100 3276 23156
rect 3332 23100 5740 23156
rect 5796 23100 5806 23156
rect 20962 23100 20972 23156
rect 21028 23100 22204 23156
rect 22260 23100 22270 23156
rect 26450 23100 26460 23156
rect 26516 23100 27244 23156
rect 27300 23100 27310 23156
rect 6066 22988 6076 23044
rect 6132 22988 7420 23044
rect 7476 22988 7486 23044
rect 19730 22988 19740 23044
rect 19796 22988 22764 23044
rect 22820 22988 22830 23044
rect 24210 22988 24220 23044
rect 24276 22988 26236 23044
rect 26292 22988 26302 23044
rect 28466 22988 28476 23044
rect 28532 22988 29260 23044
rect 29316 22988 29326 23044
rect 36530 22988 36540 23044
rect 36596 22988 37436 23044
rect 37492 22988 37502 23044
rect 38210 22988 38220 23044
rect 38276 22988 38668 23044
rect 38724 22988 38734 23044
rect 19058 22876 19068 22932
rect 19124 22876 21980 22932
rect 22036 22876 22046 22932
rect 27010 22876 27020 22932
rect 27076 22876 28028 22932
rect 28084 22876 29036 22932
rect 29092 22876 29102 22932
rect 33506 22876 33516 22932
rect 33572 22876 35308 22932
rect 35364 22876 35374 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14242 22540 14252 22596
rect 14308 22540 15148 22596
rect 15204 22540 17388 22596
rect 17444 22540 17454 22596
rect 18946 22540 18956 22596
rect 19012 22540 20412 22596
rect 20468 22540 20478 22596
rect 23650 22540 23660 22596
rect 23716 22540 24780 22596
rect 24836 22540 25900 22596
rect 25956 22540 25966 22596
rect 5730 22428 5740 22484
rect 5796 22428 6748 22484
rect 6804 22428 7980 22484
rect 8036 22428 8988 22484
rect 9044 22428 10220 22484
rect 10276 22428 11004 22484
rect 11060 22428 12908 22484
rect 12964 22428 13804 22484
rect 13860 22428 13870 22484
rect 25442 22428 25452 22484
rect 25508 22428 27356 22484
rect 27412 22428 27422 22484
rect 29148 22428 29484 22484
rect 29540 22428 29550 22484
rect 33282 22428 33292 22484
rect 33348 22428 35084 22484
rect 35140 22428 35150 22484
rect 29148 22372 29204 22428
rect 14130 22316 14140 22372
rect 14196 22316 15708 22372
rect 15764 22316 15774 22372
rect 24098 22316 24108 22372
rect 24164 22316 25116 22372
rect 25172 22316 29204 22372
rect 29362 22316 29372 22372
rect 29428 22316 30940 22372
rect 30996 22316 31006 22372
rect 33170 22316 33180 22372
rect 33236 22316 33852 22372
rect 33908 22316 33918 22372
rect 35634 22316 35644 22372
rect 35700 22316 36988 22372
rect 37044 22316 37054 22372
rect 16818 22204 16828 22260
rect 16884 22204 17388 22260
rect 17444 22204 17454 22260
rect 32498 22204 32508 22260
rect 32564 22204 33292 22260
rect 33348 22204 33628 22260
rect 33684 22204 33694 22260
rect 35298 22204 35308 22260
rect 35364 22204 35868 22260
rect 35924 22204 37548 22260
rect 37604 22204 37614 22260
rect 15474 22092 15484 22148
rect 15540 22092 16604 22148
rect 16660 22092 16670 22148
rect 21410 22092 21420 22148
rect 21476 22092 22652 22148
rect 22708 22092 22718 22148
rect 24658 22092 24668 22148
rect 24724 22092 25564 22148
rect 25620 22092 25630 22148
rect 30258 22092 30268 22148
rect 30324 22092 36092 22148
rect 36148 22092 36158 22148
rect 36306 22092 36316 22148
rect 36372 22092 38220 22148
rect 38276 22092 38286 22148
rect 36092 22036 36148 22092
rect 21970 21980 21980 22036
rect 22036 21980 27020 22036
rect 27076 21980 27086 22036
rect 29474 21980 29484 22036
rect 29540 21980 35084 22036
rect 35140 21980 35150 22036
rect 36092 21980 38556 22036
rect 38612 21980 38622 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 11666 21868 11676 21924
rect 11732 21868 14028 21924
rect 14084 21868 14094 21924
rect 16156 21868 18172 21924
rect 18228 21868 18238 21924
rect 24658 21868 24668 21924
rect 24724 21868 26908 21924
rect 31154 21868 31164 21924
rect 31220 21868 37324 21924
rect 37380 21868 38108 21924
rect 38164 21868 38174 21924
rect 16156 21812 16212 21868
rect 11330 21756 11340 21812
rect 11396 21756 12124 21812
rect 12180 21756 16212 21812
rect 26852 21700 26908 21868
rect 28018 21756 28028 21812
rect 28084 21756 28588 21812
rect 28644 21756 33404 21812
rect 33460 21756 33470 21812
rect 39218 21756 39228 21812
rect 39284 21756 40124 21812
rect 40180 21756 42812 21812
rect 42868 21756 42878 21812
rect 16258 21644 16268 21700
rect 16324 21644 17500 21700
rect 17556 21644 17566 21700
rect 18162 21644 18172 21700
rect 18228 21644 19180 21700
rect 19236 21644 19246 21700
rect 26852 21644 27244 21700
rect 27300 21644 32396 21700
rect 32452 21644 32462 21700
rect 33842 21644 33852 21700
rect 33908 21644 34636 21700
rect 34692 21644 36428 21700
rect 36484 21644 36494 21700
rect 39666 21644 39676 21700
rect 39732 21644 40908 21700
rect 40964 21644 40974 21700
rect 12012 21532 14812 21588
rect 14868 21532 15148 21588
rect 15810 21532 15820 21588
rect 15876 21532 16716 21588
rect 16772 21532 18396 21588
rect 18452 21532 18462 21588
rect 19618 21532 19628 21588
rect 19684 21532 21980 21588
rect 22036 21532 22988 21588
rect 23044 21532 23054 21588
rect 29250 21532 29260 21588
rect 29316 21532 31052 21588
rect 31108 21532 32284 21588
rect 32340 21532 34300 21588
rect 34356 21532 35644 21588
rect 35700 21532 35710 21588
rect 37986 21532 37996 21588
rect 38052 21532 39340 21588
rect 39396 21532 39406 21588
rect 12012 21476 12068 21532
rect 15092 21476 15148 21532
rect 37996 21476 38052 21532
rect 12002 21420 12012 21476
rect 12068 21420 12078 21476
rect 13010 21420 13020 21476
rect 13076 21420 14252 21476
rect 14308 21420 14318 21476
rect 15092 21420 16380 21476
rect 16436 21420 16446 21476
rect 22642 21420 22652 21476
rect 22708 21420 33516 21476
rect 33572 21420 33582 21476
rect 34962 21420 34972 21476
rect 35028 21420 38052 21476
rect 42354 21420 42364 21476
rect 42420 21420 43820 21476
rect 43876 21420 43886 21476
rect 13458 21308 13468 21364
rect 13524 21308 14588 21364
rect 14644 21308 16716 21364
rect 16772 21308 16782 21364
rect 15138 21196 15148 21252
rect 15204 21196 16268 21252
rect 16324 21196 16334 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 15092 21084 16604 21140
rect 16660 21084 16670 21140
rect 29474 21084 29484 21140
rect 29540 21084 30044 21140
rect 30100 21084 33628 21140
rect 33684 21084 34636 21140
rect 34692 21084 34702 21140
rect 15092 20916 15148 21084
rect 12450 20860 12460 20916
rect 12516 20860 13468 20916
rect 13524 20860 13534 20916
rect 14914 20860 14924 20916
rect 14980 20860 15148 20916
rect 19058 20860 19068 20916
rect 19124 20860 20524 20916
rect 20580 20860 20590 20916
rect 20860 20860 22876 20916
rect 22932 20860 22942 20916
rect 30930 20860 30940 20916
rect 30996 20860 32060 20916
rect 32116 20860 32126 20916
rect 35084 20860 37772 20916
rect 37828 20860 37838 20916
rect 37986 20860 37996 20916
rect 38052 20860 38668 20916
rect 38724 20860 38734 20916
rect 40786 20860 40796 20916
rect 40852 20860 41692 20916
rect 41748 20860 41758 20916
rect 14018 20748 14028 20804
rect 14084 20748 16492 20804
rect 16548 20748 20412 20804
rect 20468 20748 20478 20804
rect 20860 20692 20916 20860
rect 35084 20804 35140 20860
rect 21074 20748 21084 20804
rect 21140 20748 33852 20804
rect 33908 20748 35140 20804
rect 36418 20748 36428 20804
rect 36484 20748 38444 20804
rect 38500 20748 38510 20804
rect 38612 20748 39004 20804
rect 39060 20748 39070 20804
rect 38612 20692 38668 20748
rect 16706 20636 16716 20692
rect 16772 20636 18508 20692
rect 18564 20636 20916 20692
rect 21970 20636 21980 20692
rect 22036 20636 22988 20692
rect 23044 20636 23054 20692
rect 35970 20636 35980 20692
rect 36036 20636 37548 20692
rect 37604 20636 37614 20692
rect 37762 20636 37772 20692
rect 37828 20636 38332 20692
rect 38388 20636 38668 20692
rect 38882 20636 38892 20692
rect 38948 20636 39788 20692
rect 39844 20636 40236 20692
rect 40292 20636 40302 20692
rect 40450 20636 40460 20692
rect 40516 20636 42252 20692
rect 42308 20636 42318 20692
rect 40236 20580 40292 20636
rect 8082 20524 8092 20580
rect 8148 20524 11340 20580
rect 11396 20524 11406 20580
rect 16818 20524 16828 20580
rect 16884 20524 19068 20580
rect 19124 20524 21756 20580
rect 21812 20524 21822 20580
rect 22194 20524 22204 20580
rect 22260 20524 23660 20580
rect 23716 20524 23996 20580
rect 24052 20524 24062 20580
rect 32386 20524 32396 20580
rect 32452 20524 35756 20580
rect 35812 20524 35822 20580
rect 40236 20524 40684 20580
rect 40740 20524 40750 20580
rect 11218 20412 11228 20468
rect 11284 20412 12012 20468
rect 12068 20412 12078 20468
rect 13570 20412 13580 20468
rect 13636 20412 15372 20468
rect 15428 20412 19180 20468
rect 19236 20412 19246 20468
rect 20402 20412 20412 20468
rect 20468 20412 21532 20468
rect 21588 20412 22428 20468
rect 22484 20412 22494 20468
rect 26852 20412 36316 20468
rect 36372 20412 37212 20468
rect 37268 20412 37278 20468
rect 13580 20244 13636 20412
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 26852 20356 26908 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 22316 20300 26908 20356
rect 33628 20300 38892 20356
rect 38948 20300 39676 20356
rect 39732 20300 39742 20356
rect 22316 20244 22372 20300
rect 33628 20244 33684 20300
rect 12348 20188 13636 20244
rect 19730 20188 19740 20244
rect 19796 20188 22372 20244
rect 22530 20188 22540 20244
rect 22596 20188 23772 20244
rect 23828 20188 23838 20244
rect 33516 20188 33684 20244
rect 37202 20188 37212 20244
rect 37268 20188 37660 20244
rect 37716 20188 37726 20244
rect 39330 20188 39340 20244
rect 39396 20188 40236 20244
rect 40292 20188 40302 20244
rect 12348 20020 12404 20188
rect 33516 20132 33572 20188
rect 13346 20076 13356 20132
rect 13412 20076 14924 20132
rect 14980 20076 14990 20132
rect 23090 20076 23100 20132
rect 23156 20076 24220 20132
rect 24276 20076 24286 20132
rect 26450 20076 26460 20132
rect 26516 20076 27692 20132
rect 27748 20076 27758 20132
rect 27906 20076 27916 20132
rect 27972 20076 29372 20132
rect 29428 20076 29438 20132
rect 32946 20076 32956 20132
rect 33012 20076 33572 20132
rect 39106 20076 39116 20132
rect 39172 20076 40012 20132
rect 40068 20076 40078 20132
rect 12338 19964 12348 20020
rect 12404 19964 12414 20020
rect 16706 19964 16716 20020
rect 16772 19964 17388 20020
rect 17444 19964 17454 20020
rect 24434 19964 24444 20020
rect 24500 19964 25452 20020
rect 25508 19964 25518 20020
rect 29586 19964 29596 20020
rect 29652 19964 29932 20020
rect 29988 19964 30828 20020
rect 30884 19964 30894 20020
rect 31602 19964 31612 20020
rect 31668 19964 32620 20020
rect 32676 19964 33068 20020
rect 33124 19964 33740 20020
rect 33796 19964 33806 20020
rect 35298 19964 35308 20020
rect 35364 19964 35868 20020
rect 35924 19964 35934 20020
rect 38882 19964 38892 20020
rect 38948 19964 41132 20020
rect 41188 19964 41198 20020
rect 21074 19852 21084 19908
rect 21140 19852 22092 19908
rect 22148 19852 22158 19908
rect 23090 19852 23100 19908
rect 23156 19852 26348 19908
rect 26404 19852 26908 19908
rect 26964 19852 34412 19908
rect 34468 19852 34478 19908
rect 35634 19852 35644 19908
rect 35700 19852 37212 19908
rect 37268 19852 37278 19908
rect 40898 19852 40908 19908
rect 40964 19852 42252 19908
rect 42308 19852 43372 19908
rect 43428 19852 44268 19908
rect 44324 19852 44334 19908
rect 22306 19740 22316 19796
rect 22372 19740 23548 19796
rect 23604 19740 23614 19796
rect 27794 19740 27804 19796
rect 27860 19740 28364 19796
rect 28420 19740 28430 19796
rect 35410 19740 35420 19796
rect 35476 19740 35868 19796
rect 35924 19740 35934 19796
rect 27122 19628 27132 19684
rect 27188 19628 28028 19684
rect 28084 19628 28094 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 15138 19516 15148 19572
rect 15204 19516 17724 19572
rect 17780 19516 17790 19572
rect 8642 19404 8652 19460
rect 8708 19404 12124 19460
rect 12180 19404 12190 19460
rect 27010 19404 27020 19460
rect 27076 19404 32284 19460
rect 32340 19404 33404 19460
rect 33460 19404 34188 19460
rect 34244 19404 35084 19460
rect 35140 19404 35150 19460
rect 16146 19292 16156 19348
rect 16212 19292 18844 19348
rect 18900 19292 20412 19348
rect 20468 19292 20478 19348
rect 22418 19292 22428 19348
rect 22484 19292 23996 19348
rect 24052 19292 25116 19348
rect 25172 19292 25182 19348
rect 36642 19292 36652 19348
rect 36708 19292 37772 19348
rect 37828 19292 37838 19348
rect 38098 19292 38108 19348
rect 38164 19292 39900 19348
rect 39956 19292 39966 19348
rect 41234 19292 41244 19348
rect 41300 19292 42812 19348
rect 42868 19292 42878 19348
rect 21634 19180 21644 19236
rect 21700 19180 31612 19236
rect 31668 19180 31678 19236
rect 23874 19068 23884 19124
rect 23940 19068 24444 19124
rect 24500 19068 32956 19124
rect 33012 19068 33022 19124
rect 12114 18956 12124 19012
rect 12180 18956 14476 19012
rect 14532 18956 20188 19012
rect 20244 18956 21308 19012
rect 21364 18956 21374 19012
rect 23426 18956 23436 19012
rect 23492 18956 23502 19012
rect 26086 18956 26124 19012
rect 26180 18956 26684 19012
rect 26740 18956 26750 19012
rect 27010 18956 27020 19012
rect 27076 18956 27356 19012
rect 27412 18956 27422 19012
rect 28130 18956 28140 19012
rect 28196 18956 29596 19012
rect 29652 18956 29662 19012
rect 34066 18956 34076 19012
rect 34132 18956 34524 19012
rect 34580 18956 34590 19012
rect 23436 18900 23492 18956
rect 23436 18844 30156 18900
rect 30212 18844 30222 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 20514 18732 20524 18788
rect 20580 18732 27020 18788
rect 27076 18732 27086 18788
rect 27570 18732 27580 18788
rect 27636 18732 28140 18788
rect 28196 18732 28206 18788
rect 28812 18732 38444 18788
rect 38500 18732 38510 18788
rect 28812 18676 28868 18732
rect 19618 18620 19628 18676
rect 19684 18620 23548 18676
rect 27458 18620 27468 18676
rect 27524 18620 28868 18676
rect 29026 18620 29036 18676
rect 29092 18620 29820 18676
rect 29876 18620 32060 18676
rect 32116 18620 32396 18676
rect 32452 18620 33292 18676
rect 33348 18620 33358 18676
rect 33730 18620 33740 18676
rect 33796 18620 34636 18676
rect 34692 18620 34702 18676
rect 35074 18620 35084 18676
rect 35140 18620 35420 18676
rect 35476 18620 35486 18676
rect 23492 18452 23548 18620
rect 24658 18508 24668 18564
rect 24724 18508 27244 18564
rect 27300 18508 29484 18564
rect 29540 18508 29550 18564
rect 6066 18396 6076 18452
rect 6132 18396 7420 18452
rect 7476 18396 8428 18452
rect 8484 18396 8494 18452
rect 9650 18396 9660 18452
rect 9716 18396 10668 18452
rect 10724 18396 12012 18452
rect 12068 18396 12348 18452
rect 12404 18396 12414 18452
rect 23492 18396 27132 18452
rect 27188 18396 27198 18452
rect 27346 18396 27356 18452
rect 27412 18396 28028 18452
rect 28084 18396 28094 18452
rect 28354 18396 28364 18452
rect 28420 18396 28812 18452
rect 28868 18396 29708 18452
rect 29764 18396 30492 18452
rect 30548 18396 30558 18452
rect 33618 18396 33628 18452
rect 33684 18396 34524 18452
rect 34580 18396 34590 18452
rect 35074 18396 35084 18452
rect 35140 18396 40460 18452
rect 40516 18396 40526 18452
rect 18498 18284 18508 18340
rect 18564 18284 19628 18340
rect 19684 18284 19694 18340
rect 27010 18284 27020 18340
rect 27076 18284 30044 18340
rect 30100 18284 30110 18340
rect 33058 18284 33068 18340
rect 33124 18284 34412 18340
rect 34468 18284 34478 18340
rect 35298 18284 35308 18340
rect 35364 18284 36316 18340
rect 36372 18284 36382 18340
rect 36530 18284 36540 18340
rect 36596 18284 37548 18340
rect 37604 18284 37996 18340
rect 38052 18284 38062 18340
rect 39890 18284 39900 18340
rect 39956 18284 41692 18340
rect 41748 18284 41758 18340
rect 34412 18228 34468 18284
rect 7858 18172 7868 18228
rect 7924 18172 10780 18228
rect 10836 18172 10846 18228
rect 18946 18172 18956 18228
rect 19012 18172 20972 18228
rect 21028 18172 21038 18228
rect 24770 18172 24780 18228
rect 24836 18172 25676 18228
rect 25732 18172 25742 18228
rect 26338 18172 26348 18228
rect 26404 18172 27356 18228
rect 27412 18172 27422 18228
rect 28018 18172 28028 18228
rect 28084 18172 29820 18228
rect 29876 18172 30380 18228
rect 30436 18172 30716 18228
rect 30772 18172 30782 18228
rect 34412 18172 35084 18228
rect 35140 18172 35150 18228
rect 35522 18172 35532 18228
rect 35588 18172 40012 18228
rect 40068 18172 43372 18228
rect 43428 18172 43438 18228
rect 8866 18060 8876 18116
rect 8932 18060 23996 18116
rect 24052 18060 24332 18116
rect 24388 18060 24398 18116
rect 26002 18060 26012 18116
rect 26068 18060 26852 18116
rect 26908 18060 26918 18116
rect 30146 18060 30156 18116
rect 30212 18060 32844 18116
rect 32900 18060 34860 18116
rect 34916 18060 34926 18116
rect 36092 18060 39228 18116
rect 39284 18060 39294 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 18274 17948 18284 18004
rect 18340 17948 19292 18004
rect 19348 17948 19358 18004
rect 22418 17948 22428 18004
rect 22484 17948 22988 18004
rect 23044 17948 23054 18004
rect 25554 17948 25564 18004
rect 25620 17948 31052 18004
rect 31108 17948 31118 18004
rect 34514 17948 34524 18004
rect 34580 17948 34590 18004
rect 34524 17892 34580 17948
rect 36092 17892 36148 18060
rect 36418 17948 36428 18004
rect 36484 17948 37100 18004
rect 37156 17948 37166 18004
rect 38612 17948 39340 18004
rect 39396 17948 39406 18004
rect 38612 17892 38668 17948
rect 11106 17836 11116 17892
rect 11172 17836 14476 17892
rect 14532 17836 14542 17892
rect 18386 17836 18396 17892
rect 18452 17836 26180 17892
rect 27010 17836 27020 17892
rect 27076 17836 33068 17892
rect 33124 17836 33134 17892
rect 34524 17836 36148 17892
rect 36306 17836 36316 17892
rect 36372 17836 38668 17892
rect 12450 17724 12460 17780
rect 12516 17724 15148 17780
rect 17826 17724 17836 17780
rect 17892 17724 18844 17780
rect 18900 17724 20524 17780
rect 20580 17724 20590 17780
rect 15092 17668 15148 17724
rect 26124 17668 26180 17836
rect 34962 17724 34972 17780
rect 35028 17724 35980 17780
rect 36036 17724 36046 17780
rect 36194 17724 36204 17780
rect 36260 17724 37436 17780
rect 37492 17724 37502 17780
rect 38994 17724 39004 17780
rect 39060 17724 40572 17780
rect 40628 17724 40638 17780
rect 35980 17668 36036 17724
rect 15092 17612 15484 17668
rect 15540 17612 15550 17668
rect 19618 17612 19628 17668
rect 19684 17612 21756 17668
rect 21812 17612 25900 17668
rect 25956 17612 25966 17668
rect 26124 17612 27020 17668
rect 27076 17612 27086 17668
rect 27570 17612 27580 17668
rect 27636 17612 30940 17668
rect 30996 17612 31006 17668
rect 35980 17612 36876 17668
rect 36932 17612 36942 17668
rect 37090 17612 37100 17668
rect 37156 17612 39900 17668
rect 39956 17612 42812 17668
rect 42868 17612 42878 17668
rect 18610 17500 18620 17556
rect 18676 17500 19852 17556
rect 19908 17500 19918 17556
rect 23314 17500 23324 17556
rect 23380 17500 23772 17556
rect 23828 17500 26348 17556
rect 26404 17500 27468 17556
rect 27524 17500 27534 17556
rect 31042 17500 31052 17556
rect 31108 17500 33964 17556
rect 34020 17500 34636 17556
rect 34692 17500 35196 17556
rect 35252 17500 35262 17556
rect 14578 17388 14588 17444
rect 14644 17388 18284 17444
rect 18340 17388 18350 17444
rect 19618 17388 19628 17444
rect 19684 17388 20300 17444
rect 20356 17388 22092 17444
rect 22148 17388 22158 17444
rect 25778 17388 25788 17444
rect 25844 17388 27916 17444
rect 27972 17388 27982 17444
rect 33170 17388 33180 17444
rect 33236 17388 33852 17444
rect 33908 17388 33918 17444
rect 15026 17276 15036 17332
rect 15092 17276 17500 17332
rect 17556 17276 18396 17332
rect 18452 17276 18462 17332
rect 24546 17276 24556 17332
rect 24612 17276 25396 17332
rect 25554 17276 25564 17332
rect 25620 17276 26124 17332
rect 26180 17276 26572 17332
rect 26628 17276 26638 17332
rect 27122 17276 27132 17332
rect 27188 17276 27468 17332
rect 27524 17276 27534 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 25340 17220 25396 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 11890 17164 11900 17220
rect 11956 17164 19180 17220
rect 19236 17164 19246 17220
rect 20962 17164 20972 17220
rect 21028 17164 22428 17220
rect 22484 17164 22494 17220
rect 25340 17164 30940 17220
rect 30996 17164 31006 17220
rect 11554 17052 11564 17108
rect 11620 17052 24444 17108
rect 24500 17052 24510 17108
rect 27122 17052 27132 17108
rect 27188 17052 28028 17108
rect 28084 17052 28094 17108
rect 30156 17052 33180 17108
rect 33236 17052 34412 17108
rect 34468 17052 34478 17108
rect 16818 16940 16828 16996
rect 16884 16940 17500 16996
rect 17556 16940 17566 16996
rect 20178 16940 20188 16996
rect 20244 16940 23660 16996
rect 23716 16940 23726 16996
rect 26562 16940 26572 16996
rect 26628 16940 28252 16996
rect 28308 16940 28318 16996
rect 13122 16828 13132 16884
rect 13188 16828 16044 16884
rect 16100 16828 16716 16884
rect 16772 16828 23884 16884
rect 23940 16828 23950 16884
rect 25442 16828 25452 16884
rect 25508 16828 26124 16884
rect 26180 16828 27132 16884
rect 27188 16828 27198 16884
rect 30156 16772 30212 17052
rect 33282 16940 33292 16996
rect 33348 16940 33740 16996
rect 33796 16940 33806 16996
rect 34962 16940 34972 16996
rect 35028 16940 38668 16996
rect 38612 16884 38668 16940
rect 33058 16828 33068 16884
rect 33124 16828 35532 16884
rect 35588 16828 36204 16884
rect 36260 16828 36270 16884
rect 38612 16828 39116 16884
rect 39172 16828 41916 16884
rect 41972 16828 41982 16884
rect 12786 16716 12796 16772
rect 12852 16716 14924 16772
rect 14980 16716 15820 16772
rect 15876 16716 15886 16772
rect 18274 16716 18284 16772
rect 18340 16716 22988 16772
rect 23044 16716 23054 16772
rect 24994 16716 25004 16772
rect 25060 16716 30212 16772
rect 34514 16716 34524 16772
rect 34580 16716 35980 16772
rect 36036 16716 36046 16772
rect 38210 16716 38220 16772
rect 38276 16716 39228 16772
rect 39284 16716 39294 16772
rect 23314 16604 23324 16660
rect 23380 16604 23996 16660
rect 24052 16604 24062 16660
rect 20290 16492 20300 16548
rect 20356 16492 26684 16548
rect 26740 16492 26750 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 22866 16380 22876 16436
rect 22932 16380 24668 16436
rect 24724 16380 24734 16436
rect 30706 16380 30716 16436
rect 30772 16380 31388 16436
rect 31444 16380 31454 16436
rect 9874 16268 9884 16324
rect 9940 16268 11228 16324
rect 11284 16268 11294 16324
rect 11778 16268 11788 16324
rect 11844 16268 14700 16324
rect 14756 16268 15036 16324
rect 15092 16268 15102 16324
rect 16258 16268 16268 16324
rect 16324 16268 20188 16324
rect 20244 16268 20254 16324
rect 24434 16268 24444 16324
rect 24500 16268 29484 16324
rect 29540 16268 29550 16324
rect 20066 16156 20076 16212
rect 20132 16156 22764 16212
rect 22820 16156 23324 16212
rect 23380 16156 23390 16212
rect 24770 16156 24780 16212
rect 24836 16156 28364 16212
rect 28420 16156 32172 16212
rect 32228 16156 34524 16212
rect 34580 16156 34590 16212
rect 43138 16156 43148 16212
rect 43204 16156 43820 16212
rect 43876 16156 43886 16212
rect 24210 16044 24220 16100
rect 24276 16044 24444 16100
rect 24500 16044 30044 16100
rect 30100 16044 34300 16100
rect 34356 16044 34366 16100
rect 13794 15932 13804 15988
rect 13860 15932 14812 15988
rect 14868 15932 15932 15988
rect 15988 15932 15998 15988
rect 32386 15932 32396 15988
rect 32452 15932 33404 15988
rect 33460 15932 33470 15988
rect 30146 15820 30156 15876
rect 30212 15820 37436 15876
rect 37492 15820 38108 15876
rect 38164 15820 38174 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 8866 15484 8876 15540
rect 8932 15484 19908 15540
rect 26674 15484 26684 15540
rect 26740 15484 27916 15540
rect 27972 15484 27982 15540
rect 29932 15484 32060 15540
rect 32116 15484 36988 15540
rect 37044 15484 37054 15540
rect 19852 15428 19908 15484
rect 29932 15428 29988 15484
rect 16930 15372 16940 15428
rect 16996 15372 19292 15428
rect 19348 15372 19358 15428
rect 19852 15372 25900 15428
rect 25956 15372 26124 15428
rect 26180 15372 26190 15428
rect 26786 15372 26796 15428
rect 26852 15372 28028 15428
rect 28084 15372 28094 15428
rect 29474 15372 29484 15428
rect 29540 15372 29932 15428
rect 29988 15372 29998 15428
rect 31378 15372 31388 15428
rect 31444 15372 38668 15428
rect 38724 15372 42700 15428
rect 42756 15372 42766 15428
rect 19618 15260 19628 15316
rect 19684 15260 21308 15316
rect 21364 15260 21374 15316
rect 24210 15260 24220 15316
rect 24276 15260 25788 15316
rect 25844 15260 25854 15316
rect 28802 15260 28812 15316
rect 28868 15260 29596 15316
rect 29652 15260 36540 15316
rect 36596 15260 36606 15316
rect 44258 15260 44268 15316
rect 44324 15260 45276 15316
rect 45332 15260 45342 15316
rect 6066 15148 6076 15204
rect 6132 15148 7980 15204
rect 8036 15148 8540 15204
rect 8596 15148 9660 15204
rect 9716 15148 10444 15204
rect 10500 15148 11900 15204
rect 11956 15148 12796 15204
rect 12852 15148 12862 15204
rect 15586 15148 15596 15204
rect 15652 15148 17388 15204
rect 17444 15148 17454 15204
rect 21746 15148 21756 15204
rect 21812 15148 22876 15204
rect 22932 15148 26908 15204
rect 26964 15148 26974 15204
rect 36866 15148 36876 15204
rect 36932 15148 38668 15204
rect 38724 15148 38734 15204
rect 42466 15148 42476 15204
rect 42532 15148 43820 15204
rect 43876 15148 43886 15204
rect 17714 15036 17724 15092
rect 17780 15036 28588 15092
rect 28644 15036 28654 15092
rect 32610 14924 32620 14980
rect 32676 14924 33516 14980
rect 33572 14924 33582 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 17378 14700 17388 14756
rect 17444 14700 20076 14756
rect 20132 14700 20748 14756
rect 20804 14700 20814 14756
rect 27682 14700 27692 14756
rect 27748 14700 29148 14756
rect 29204 14700 29214 14756
rect 26114 14588 26124 14644
rect 26180 14588 29988 14644
rect 30146 14588 30156 14644
rect 30212 14588 31948 14644
rect 32004 14588 32014 14644
rect 37874 14588 37884 14644
rect 37940 14588 39004 14644
rect 39060 14588 39070 14644
rect 29932 14532 29988 14588
rect 19170 14476 19180 14532
rect 19236 14476 20636 14532
rect 20692 14476 20702 14532
rect 26786 14476 26796 14532
rect 26852 14476 29148 14532
rect 29204 14476 29214 14532
rect 29932 14476 37660 14532
rect 37716 14476 37726 14532
rect 11890 14364 11900 14420
rect 11956 14364 12236 14420
rect 12292 14364 16380 14420
rect 16436 14364 16446 14420
rect 20850 14364 20860 14420
rect 20916 14364 21980 14420
rect 22036 14364 22204 14420
rect 22260 14364 22270 14420
rect 23874 14364 23884 14420
rect 23940 14364 24332 14420
rect 24388 14364 24398 14420
rect 25666 14364 25676 14420
rect 25732 14364 26908 14420
rect 26964 14364 31052 14420
rect 31108 14364 31118 14420
rect 32274 14364 32284 14420
rect 32340 14364 35084 14420
rect 35140 14364 35150 14420
rect 36418 14364 36428 14420
rect 36484 14364 42140 14420
rect 42196 14364 42206 14420
rect 25778 14252 25788 14308
rect 25844 14252 27468 14308
rect 27524 14252 27534 14308
rect 28354 14252 28364 14308
rect 28420 14252 29036 14308
rect 29092 14252 29102 14308
rect 29922 14252 29932 14308
rect 29988 14252 32620 14308
rect 32676 14252 32686 14308
rect 32946 14252 32956 14308
rect 33012 14252 34300 14308
rect 34356 14252 34366 14308
rect 28690 14140 28700 14196
rect 28756 14140 31948 14196
rect 32004 14140 32732 14196
rect 32788 14140 32798 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 25778 14028 25788 14084
rect 25844 14028 26124 14084
rect 26180 14028 26190 14084
rect 23314 13916 23324 13972
rect 23380 13916 25340 13972
rect 25396 13916 25406 13972
rect 28242 13916 28252 13972
rect 28308 13916 28812 13972
rect 28868 13916 28878 13972
rect 11442 13804 11452 13860
rect 11508 13804 13692 13860
rect 13748 13804 13758 13860
rect 15092 13804 17612 13860
rect 17668 13804 17678 13860
rect 21746 13804 21756 13860
rect 21812 13804 25116 13860
rect 25172 13804 25182 13860
rect 27906 13804 27916 13860
rect 27972 13804 30268 13860
rect 30324 13804 30334 13860
rect 32060 13804 33292 13860
rect 33348 13804 33358 13860
rect 33842 13804 33852 13860
rect 33908 13804 35868 13860
rect 35924 13804 35934 13860
rect 38434 13804 38444 13860
rect 38500 13804 42588 13860
rect 42644 13804 42654 13860
rect 42802 13804 42812 13860
rect 42868 13804 43596 13860
rect 43652 13804 43662 13860
rect 9874 13692 9884 13748
rect 9940 13692 11116 13748
rect 11172 13692 11182 13748
rect 15092 13636 15148 13804
rect 32060 13748 32116 13804
rect 33292 13748 33348 13804
rect 18610 13692 18620 13748
rect 18676 13692 22540 13748
rect 22596 13692 22606 13748
rect 23314 13692 23324 13748
rect 23380 13692 24444 13748
rect 24500 13692 24510 13748
rect 25666 13692 25676 13748
rect 25732 13692 26572 13748
rect 26628 13692 26638 13748
rect 32050 13692 32060 13748
rect 32116 13692 32126 13748
rect 33292 13692 34412 13748
rect 34468 13692 34860 13748
rect 34916 13692 34926 13748
rect 36082 13692 36092 13748
rect 36148 13692 42140 13748
rect 42196 13692 42206 13748
rect 44370 13692 44380 13748
rect 44436 13692 47068 13748
rect 47124 13692 47134 13748
rect 11330 13580 11340 13636
rect 11396 13580 15148 13636
rect 16482 13580 16492 13636
rect 16548 13580 19180 13636
rect 19236 13580 19246 13636
rect 23874 13580 23884 13636
rect 23940 13580 25228 13636
rect 25284 13580 25294 13636
rect 32386 13580 32396 13636
rect 32452 13580 33292 13636
rect 33348 13580 33358 13636
rect 44380 13524 44436 13692
rect 8978 13468 8988 13524
rect 9044 13468 10220 13524
rect 10276 13468 10286 13524
rect 14690 13468 14700 13524
rect 14756 13468 21812 13524
rect 24210 13468 24220 13524
rect 24276 13468 24556 13524
rect 24612 13468 24622 13524
rect 25666 13468 25676 13524
rect 25732 13468 26460 13524
rect 26516 13468 26526 13524
rect 34972 13468 35420 13524
rect 35476 13468 35486 13524
rect 35634 13468 35644 13524
rect 35700 13468 36428 13524
rect 36484 13468 36494 13524
rect 38994 13468 39004 13524
rect 39060 13468 39788 13524
rect 39844 13468 42812 13524
rect 42868 13468 42878 13524
rect 43250 13468 43260 13524
rect 43316 13468 44436 13524
rect 21756 13412 21812 13468
rect 34972 13412 35028 13468
rect 21756 13356 23996 13412
rect 24052 13356 24062 13412
rect 25330 13356 25340 13412
rect 25396 13356 26012 13412
rect 26068 13356 26078 13412
rect 30034 13356 30044 13412
rect 30100 13356 35028 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 17266 13244 17276 13300
rect 17332 13244 18060 13300
rect 18116 13244 18126 13300
rect 24098 13244 24108 13300
rect 24164 13244 26348 13300
rect 26404 13244 26414 13300
rect 31042 13244 31052 13300
rect 31108 13244 32172 13300
rect 32228 13244 32238 13300
rect 15362 13132 15372 13188
rect 15428 13132 16716 13188
rect 16772 13132 18508 13188
rect 18564 13132 18574 13188
rect 24546 13132 24556 13188
rect 24612 13132 25452 13188
rect 25508 13132 25518 13188
rect 34962 13132 34972 13188
rect 35028 13132 35308 13188
rect 35364 13132 35374 13188
rect 10994 13020 11004 13076
rect 11060 13020 11564 13076
rect 11620 13020 14028 13076
rect 14084 13020 14364 13076
rect 14420 13020 17500 13076
rect 17556 13020 17566 13076
rect 25554 13020 25564 13076
rect 25620 13020 25630 13076
rect 30818 13020 30828 13076
rect 30884 13020 35532 13076
rect 35588 13020 35598 13076
rect 44594 13020 44604 13076
rect 44660 13020 47740 13076
rect 47796 13020 47806 13076
rect 25564 12964 25620 13020
rect 15810 12908 15820 12964
rect 15876 12908 17724 12964
rect 17780 12908 17790 12964
rect 25564 12908 25900 12964
rect 25956 12908 26572 12964
rect 26628 12908 29484 12964
rect 29540 12908 29550 12964
rect 34962 12908 34972 12964
rect 35028 12908 35756 12964
rect 35812 12908 35822 12964
rect 39330 12908 39340 12964
rect 39396 12908 43820 12964
rect 43876 12908 43886 12964
rect 24770 12796 24780 12852
rect 24836 12796 25564 12852
rect 25620 12796 25630 12852
rect 27570 12796 27580 12852
rect 27636 12796 28252 12852
rect 28308 12796 28318 12852
rect 32386 12796 32396 12852
rect 32452 12796 33180 12852
rect 33236 12796 33246 12852
rect 34738 12796 34748 12852
rect 34804 12796 35420 12852
rect 35476 12796 35486 12852
rect 37986 12796 37996 12852
rect 38052 12796 39116 12852
rect 39172 12796 39676 12852
rect 39732 12796 39742 12852
rect 44258 12796 44268 12852
rect 44324 12796 45612 12852
rect 45668 12796 45678 12852
rect 8530 12684 8540 12740
rect 8596 12684 22988 12740
rect 23044 12684 23548 12740
rect 23604 12684 25228 12740
rect 25284 12684 25900 12740
rect 25956 12684 25966 12740
rect 30716 12684 31836 12740
rect 31892 12684 31902 12740
rect 30716 12628 30772 12684
rect 30706 12572 30716 12628
rect 30772 12572 30782 12628
rect 31154 12572 31164 12628
rect 31220 12572 35532 12628
rect 35588 12572 35598 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 22950 12460 22988 12516
rect 23044 12460 23054 12516
rect 27458 12460 27468 12516
rect 27524 12460 31052 12516
rect 31108 12460 31118 12516
rect 22754 12348 22764 12404
rect 22820 12348 23212 12404
rect 23268 12348 24220 12404
rect 24276 12348 24286 12404
rect 25890 12348 25900 12404
rect 25956 12348 27244 12404
rect 27300 12348 27580 12404
rect 27636 12348 27646 12404
rect 28354 12348 28364 12404
rect 28420 12348 30044 12404
rect 30100 12348 30110 12404
rect 32050 12348 32060 12404
rect 32116 12348 32844 12404
rect 32900 12348 32910 12404
rect 38210 12348 38220 12404
rect 38276 12348 39228 12404
rect 39284 12348 39294 12404
rect 44034 12348 44044 12404
rect 44100 12348 44940 12404
rect 44996 12348 45006 12404
rect 26852 12236 34300 12292
rect 34356 12236 36540 12292
rect 36596 12236 36606 12292
rect 39666 12236 39676 12292
rect 39732 12236 43148 12292
rect 43204 12236 43932 12292
rect 43988 12236 43998 12292
rect 26852 12180 26908 12236
rect 17154 12124 17164 12180
rect 17220 12124 19852 12180
rect 19908 12124 19918 12180
rect 24434 12124 24444 12180
rect 24500 12124 24780 12180
rect 24836 12124 25340 12180
rect 25396 12124 26908 12180
rect 27234 12124 27244 12180
rect 27300 12124 27310 12180
rect 28690 12124 28700 12180
rect 28756 12124 29484 12180
rect 29540 12124 30380 12180
rect 30436 12124 34636 12180
rect 34692 12124 36428 12180
rect 36484 12124 36494 12180
rect 27244 12068 27300 12124
rect 21746 12012 21756 12068
rect 21812 12012 22764 12068
rect 22820 12012 27300 12068
rect 27906 12012 27916 12068
rect 27972 12012 30604 12068
rect 30660 12012 30670 12068
rect 12450 11900 12460 11956
rect 12516 11900 14252 11956
rect 14308 11900 14318 11956
rect 23426 11900 23436 11956
rect 23492 11900 24164 11956
rect 25218 11900 25228 11956
rect 25284 11900 31388 11956
rect 31444 11900 31454 11956
rect 34962 11900 34972 11956
rect 35028 11900 37156 11956
rect 37538 11900 37548 11956
rect 37604 11900 38892 11956
rect 38948 11900 38958 11956
rect 43250 11900 43260 11956
rect 43316 11900 44604 11956
rect 44660 11900 44670 11956
rect 24108 11844 24164 11900
rect 37100 11844 37156 11900
rect 15138 11788 15148 11844
rect 15204 11788 23884 11844
rect 23940 11788 23950 11844
rect 24108 11788 27916 11844
rect 27972 11788 27982 11844
rect 28130 11788 28140 11844
rect 28196 11788 29372 11844
rect 29428 11788 29438 11844
rect 37090 11788 37100 11844
rect 37156 11788 37166 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 16034 11676 16044 11732
rect 16100 11676 17500 11732
rect 17556 11676 17566 11732
rect 19842 11676 19852 11732
rect 19908 11676 20636 11732
rect 20692 11676 22540 11732
rect 22596 11676 22606 11732
rect 42466 11564 42476 11620
rect 42532 11564 44268 11620
rect 44324 11564 44334 11620
rect 20178 11452 20188 11508
rect 20244 11452 21644 11508
rect 21700 11452 21710 11508
rect 23874 11452 23884 11508
rect 23940 11452 30268 11508
rect 30324 11452 30716 11508
rect 30772 11452 30782 11508
rect 33170 11452 33180 11508
rect 33236 11452 36316 11508
rect 36372 11452 37884 11508
rect 37940 11452 37950 11508
rect 21970 11340 21980 11396
rect 22036 11340 23100 11396
rect 23156 11340 23166 11396
rect 24322 11340 24332 11396
rect 24388 11340 27468 11396
rect 27524 11340 27534 11396
rect 16706 11228 16716 11284
rect 16772 11228 24220 11284
rect 24276 11228 24286 11284
rect 16258 11116 16268 11172
rect 16324 11116 23212 11172
rect 23268 11116 23278 11172
rect 18498 11004 18508 11060
rect 18564 11004 19180 11060
rect 19236 11004 19246 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 17602 10780 17612 10836
rect 17668 10780 23548 10836
rect 23604 10780 25228 10836
rect 25284 10780 25294 10836
rect 26086 10780 26124 10836
rect 26180 10780 26572 10836
rect 26628 10780 26638 10836
rect 26898 10780 26908 10836
rect 26964 10780 32508 10836
rect 32564 10780 33404 10836
rect 33460 10780 34188 10836
rect 34244 10780 34254 10836
rect 38882 10780 38892 10836
rect 38948 10780 39788 10836
rect 39844 10780 39854 10836
rect 13458 10668 13468 10724
rect 13524 10668 14476 10724
rect 14532 10668 15708 10724
rect 15764 10668 15774 10724
rect 22054 10668 22092 10724
rect 22148 10668 22158 10724
rect 22306 10668 22316 10724
rect 22372 10668 22764 10724
rect 22820 10668 22830 10724
rect 25106 10668 25116 10724
rect 25172 10668 25182 10724
rect 28802 10668 28812 10724
rect 28868 10668 34524 10724
rect 34580 10668 34590 10724
rect 34962 10668 34972 10724
rect 35028 10668 36204 10724
rect 36260 10668 36270 10724
rect 25116 10612 25172 10668
rect 17826 10556 17836 10612
rect 17892 10556 18620 10612
rect 18676 10556 18686 10612
rect 18946 10556 18956 10612
rect 19012 10556 19628 10612
rect 19684 10556 19694 10612
rect 20738 10556 20748 10612
rect 20804 10556 21980 10612
rect 22036 10556 22046 10612
rect 23202 10556 23212 10612
rect 23268 10556 24332 10612
rect 24388 10556 25172 10612
rect 31042 10556 31052 10612
rect 31108 10556 36428 10612
rect 36484 10556 37212 10612
rect 37268 10556 37660 10612
rect 37716 10556 37726 10612
rect 13234 10444 13244 10500
rect 13300 10444 14364 10500
rect 14420 10444 14700 10500
rect 14756 10444 14766 10500
rect 17378 10444 17388 10500
rect 17444 10444 18284 10500
rect 18340 10444 26124 10500
rect 26180 10444 26190 10500
rect 25554 10332 25564 10388
rect 25620 10332 26236 10388
rect 26292 10332 26302 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 22082 10108 22092 10164
rect 22148 10108 22428 10164
rect 22484 10108 22494 10164
rect 25890 10108 25900 10164
rect 25956 10108 26908 10164
rect 26964 10108 26974 10164
rect 15250 9996 15260 10052
rect 15316 9996 19628 10052
rect 19684 9996 20524 10052
rect 20580 9996 21196 10052
rect 21252 9996 21262 10052
rect 22642 9996 22652 10052
rect 22708 9996 22718 10052
rect 33954 9996 33964 10052
rect 34020 9996 34300 10052
rect 34356 9996 34366 10052
rect 34514 9996 34524 10052
rect 34580 9996 35196 10052
rect 35252 9996 35262 10052
rect 36866 9996 36876 10052
rect 36932 9996 39452 10052
rect 39508 9996 39788 10052
rect 39844 9996 39854 10052
rect 41346 9996 41356 10052
rect 41412 9996 42252 10052
rect 42308 9996 42812 10052
rect 42868 9996 43708 10052
rect 22652 9940 22708 9996
rect 17490 9884 17500 9940
rect 17556 9884 18060 9940
rect 18116 9884 22708 9940
rect 27682 9884 27692 9940
rect 27748 9884 28812 9940
rect 28868 9884 28878 9940
rect 40002 9884 40012 9940
rect 40068 9884 41580 9940
rect 41636 9884 41646 9940
rect 43652 9828 43708 9996
rect 18722 9772 18732 9828
rect 18788 9772 22092 9828
rect 22148 9772 22540 9828
rect 22596 9772 22606 9828
rect 22764 9772 32396 9828
rect 32452 9772 33404 9828
rect 33460 9772 33470 9828
rect 43652 9772 44828 9828
rect 44884 9772 44894 9828
rect 22764 9716 22820 9772
rect 11666 9660 11676 9716
rect 11732 9660 14028 9716
rect 14084 9660 14094 9716
rect 14802 9660 14812 9716
rect 14868 9660 15148 9716
rect 16930 9660 16940 9716
rect 16996 9660 17948 9716
rect 18004 9660 19180 9716
rect 19236 9660 19246 9716
rect 19506 9660 19516 9716
rect 19572 9660 19740 9716
rect 19796 9660 22820 9716
rect 22978 9660 22988 9716
rect 23044 9660 26124 9716
rect 26180 9660 27916 9716
rect 27972 9660 27982 9716
rect 28466 9660 28476 9716
rect 28532 9660 29148 9716
rect 29204 9660 29214 9716
rect 15092 9604 15148 9660
rect 15092 9548 15932 9604
rect 15988 9548 17164 9604
rect 17220 9548 17230 9604
rect 19282 9548 19292 9604
rect 19348 9548 20188 9604
rect 20244 9548 25676 9604
rect 25732 9548 25742 9604
rect 32834 9548 32844 9604
rect 32900 9548 33628 9604
rect 33684 9548 35756 9604
rect 35812 9548 35822 9604
rect 18610 9436 18620 9492
rect 18676 9436 19516 9492
rect 19572 9436 19582 9492
rect 35186 9436 35196 9492
rect 35252 9436 36204 9492
rect 36260 9436 36270 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 33618 9324 33628 9380
rect 33684 9324 36428 9380
rect 36484 9324 36988 9380
rect 37044 9324 37324 9380
rect 37380 9324 37390 9380
rect 22754 9212 22764 9268
rect 22820 9212 23660 9268
rect 23716 9212 23726 9268
rect 33394 9212 33404 9268
rect 33460 9212 33852 9268
rect 33908 9212 34300 9268
rect 34356 9212 34366 9268
rect 35746 9212 35756 9268
rect 35812 9212 36540 9268
rect 36596 9212 37996 9268
rect 38052 9212 38444 9268
rect 38500 9212 38510 9268
rect 14914 9100 14924 9156
rect 14980 9100 21868 9156
rect 21924 9100 21934 9156
rect 22978 9100 22988 9156
rect 23044 9100 33180 9156
rect 33236 9100 33628 9156
rect 33684 9100 33694 9156
rect 33954 9100 33964 9156
rect 34020 9100 34748 9156
rect 34804 9100 35308 9156
rect 35364 9100 35374 9156
rect 15026 8988 15036 9044
rect 15092 8988 16156 9044
rect 16212 8988 17724 9044
rect 17780 8988 17790 9044
rect 33730 8988 33740 9044
rect 33796 8988 37436 9044
rect 37492 8988 38556 9044
rect 38612 8988 38622 9044
rect 21522 8876 21532 8932
rect 21588 8876 22204 8932
rect 22260 8876 23212 8932
rect 23268 8876 31388 8932
rect 31444 8876 34524 8932
rect 34580 8876 34590 8932
rect 11890 8764 11900 8820
rect 11956 8764 13916 8820
rect 13972 8764 13982 8820
rect 19954 8764 19964 8820
rect 20020 8764 20524 8820
rect 20580 8764 20590 8820
rect 29698 8764 29708 8820
rect 29764 8764 33068 8820
rect 33124 8764 33516 8820
rect 33572 8764 34636 8820
rect 34692 8764 34702 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 33058 8540 33068 8596
rect 33124 8540 33404 8596
rect 33460 8540 33470 8596
rect 23772 8428 25676 8484
rect 25732 8428 25742 8484
rect 23772 8372 23828 8428
rect 15138 8316 15148 8372
rect 15204 8316 16380 8372
rect 16436 8316 16446 8372
rect 16706 8316 16716 8372
rect 16772 8316 17836 8372
rect 17892 8316 19404 8372
rect 19460 8316 20636 8372
rect 20692 8316 22540 8372
rect 22596 8316 23548 8372
rect 23604 8316 23772 8372
rect 23828 8316 23838 8372
rect 35858 8316 35868 8372
rect 35924 8316 37436 8372
rect 37492 8316 37502 8372
rect 18162 8204 18172 8260
rect 18228 8204 19516 8260
rect 19572 8204 27804 8260
rect 27860 8204 27870 8260
rect 34514 8204 34524 8260
rect 34580 8204 36092 8260
rect 36148 8204 37996 8260
rect 38052 8204 38062 8260
rect 38210 8204 38220 8260
rect 38276 8204 39340 8260
rect 39396 8204 39406 8260
rect 21970 8092 21980 8148
rect 22036 8092 23212 8148
rect 23268 8092 26908 8148
rect 31266 8092 31276 8148
rect 31332 8092 31948 8148
rect 32004 8092 32014 8148
rect 26852 8036 26908 8092
rect 26852 7980 33404 8036
rect 33460 7980 33740 8036
rect 33796 7980 33806 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 18834 7532 18844 7588
rect 18900 7532 22316 7588
rect 22372 7532 22382 7588
rect 26852 7532 28252 7588
rect 28308 7532 29372 7588
rect 29428 7532 29438 7588
rect 31490 7532 31500 7588
rect 31556 7532 38444 7588
rect 38500 7532 38510 7588
rect 26852 7476 26908 7532
rect 12226 7420 12236 7476
rect 12292 7420 13580 7476
rect 13636 7420 13646 7476
rect 23426 7420 23436 7476
rect 23492 7420 23996 7476
rect 24052 7420 26908 7476
rect 20402 7308 20412 7364
rect 20468 7308 22316 7364
rect 22372 7308 23548 7364
rect 23604 7308 23614 7364
rect 24210 7196 24220 7252
rect 24276 7196 26796 7252
rect 26852 7196 27244 7252
rect 27300 7196 27310 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 15474 6860 15484 6916
rect 15540 6860 15932 6916
rect 15988 6860 15998 6916
rect 32834 6748 32844 6804
rect 32900 6748 35420 6804
rect 35476 6748 35486 6804
rect 21746 6636 21756 6692
rect 21812 6636 22652 6692
rect 22708 6636 22718 6692
rect 29932 6636 31500 6692
rect 31556 6636 31566 6692
rect 29932 6580 29988 6636
rect 23202 6524 23212 6580
rect 23268 6524 29372 6580
rect 29428 6524 29932 6580
rect 29988 6524 29998 6580
rect 31266 6524 31276 6580
rect 31332 6524 32060 6580
rect 32116 6524 32126 6580
rect 39778 6524 39788 6580
rect 39844 6524 40348 6580
rect 40404 6524 40414 6580
rect 28354 6412 28364 6468
rect 28420 6412 29148 6468
rect 29204 6412 32956 6468
rect 33012 6412 33022 6468
rect 22530 6300 22540 6356
rect 22596 6300 23212 6356
rect 23268 6300 23278 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 28690 6076 28700 6132
rect 28756 6076 31052 6132
rect 31108 6076 31118 6132
rect 32172 6076 32844 6132
rect 32900 6076 32910 6132
rect 32172 6020 32228 6076
rect 16034 5964 16044 6020
rect 16100 5964 18396 6020
rect 18452 5964 21756 6020
rect 21812 5964 21822 6020
rect 27570 5964 27580 6020
rect 27636 5964 32172 6020
rect 32228 5964 32238 6020
rect 32386 5964 32396 6020
rect 32452 5964 33180 6020
rect 33236 5964 33852 6020
rect 33908 5964 33918 6020
rect 16930 5740 16940 5796
rect 16996 5740 17836 5796
rect 17892 5740 28924 5796
rect 28980 5740 28990 5796
rect 33058 5740 33068 5796
rect 33124 5740 34300 5796
rect 34356 5740 35532 5796
rect 35588 5740 35598 5796
rect 21410 5628 21420 5684
rect 21476 5628 22988 5684
rect 23044 5628 23054 5684
rect 30146 5628 30156 5684
rect 30212 5628 33180 5684
rect 33236 5628 33246 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19282 5292 19292 5348
rect 19348 5292 20636 5348
rect 20692 5292 23548 5348
rect 23604 5292 23614 5348
rect 22306 5180 22316 5236
rect 22372 5180 26012 5236
rect 26068 5180 28252 5236
rect 28308 5180 28318 5236
rect 29250 5180 29260 5236
rect 29316 5180 30828 5236
rect 30884 5180 32508 5236
rect 32564 5180 34076 5236
rect 34132 5180 34142 5236
rect 36306 5180 36316 5236
rect 36372 5180 36988 5236
rect 37044 5180 37054 5236
rect 39890 5180 39900 5236
rect 39956 5180 40348 5236
rect 40404 5180 41132 5236
rect 41188 5180 41198 5236
rect 14466 5068 14476 5124
rect 14532 5068 15148 5124
rect 15204 5068 15214 5124
rect 15474 5068 15484 5124
rect 15540 5068 15550 5124
rect 37314 5068 37324 5124
rect 37380 5068 39116 5124
rect 39172 5068 39182 5124
rect 15484 5012 15540 5068
rect 13458 4956 13468 5012
rect 13524 4956 14028 5012
rect 14084 4956 16828 5012
rect 16884 4956 17164 5012
rect 17220 4956 17230 5012
rect 20402 4956 20412 5012
rect 20468 4956 20972 5012
rect 21028 4956 22876 5012
rect 22932 4956 23212 5012
rect 23268 4956 23278 5012
rect 27682 4956 27692 5012
rect 27748 4956 28476 5012
rect 28532 4956 28542 5012
rect 22642 4844 22652 4900
rect 22708 4844 23548 4900
rect 23604 4844 23614 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 24322 4508 24332 4564
rect 24388 4508 25564 4564
rect 25620 4508 26012 4564
rect 26068 4508 26078 4564
rect 36642 4508 36652 4564
rect 36708 4508 37772 4564
rect 37828 4508 39900 4564
rect 39956 4508 39966 4564
rect 14690 4396 14700 4452
rect 14756 4396 17388 4452
rect 17444 4396 17454 4452
rect 18722 4396 18732 4452
rect 18788 4396 21868 4452
rect 21924 4396 21934 4452
rect 34738 4172 34748 4228
rect 34804 4172 35868 4228
rect 35924 4172 35934 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19180 55132 19236 55188
rect 30828 55020 30884 55076
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 18732 54460 18788 54516
rect 19404 54348 19460 54404
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 30940 53004 30996 53060
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 49756 51996 49812 52052
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 40460 51324 40516 51380
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 49084 50540 49140 50596
rect 50092 50428 50148 50484
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 49308 50092 49364 50148
rect 30380 49756 30436 49812
rect 49084 49644 49140 49700
rect 18620 49532 18676 49588
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 18732 49308 18788 49364
rect 19180 49308 19236 49364
rect 30940 49084 30996 49140
rect 18620 48972 18676 49028
rect 49308 48636 49364 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 50204 48524 50260 48580
rect 30380 48300 30436 48356
rect 50204 47964 50260 48020
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 50092 47740 50148 47796
rect 49756 47404 49812 47460
rect 19404 47292 19460 47348
rect 50092 47292 50148 47348
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 42364 46620 42420 46676
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 49196 44492 49252 44548
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 49196 43596 49252 43652
rect 40236 43148 40292 43204
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 43596 42924 43652 42980
rect 17164 42812 17220 42868
rect 30828 42700 30884 42756
rect 42252 42700 42308 42756
rect 42364 42588 42420 42644
rect 42700 42588 42756 42644
rect 18844 42476 18900 42532
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 40236 40908 40292 40964
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 10668 40572 10724 40628
rect 16044 40460 16100 40516
rect 17052 40236 17108 40292
rect 43596 40124 43652 40180
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 21084 39788 21140 39844
rect 20636 39452 20692 39508
rect 48412 39340 48468 39396
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 14700 39004 14756 39060
rect 10220 38892 10276 38948
rect 17052 38780 17108 38836
rect 20748 38780 20804 38836
rect 10220 38556 10276 38612
rect 21308 38556 21364 38612
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 20188 38444 20244 38500
rect 20412 38444 20468 38500
rect 40460 38444 40516 38500
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 17164 37884 17220 37940
rect 42700 37884 42756 37940
rect 21308 37772 21364 37828
rect 10668 37660 10724 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 20188 37548 20244 37604
rect 20748 37436 20804 37492
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 14140 37212 14196 37268
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 14588 36540 14644 36596
rect 18844 36316 18900 36372
rect 20636 36316 20692 36372
rect 14140 36204 14196 36260
rect 14588 36204 14644 36260
rect 16268 36204 16324 36260
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 15092 35980 15148 36036
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 15932 35756 15988 35812
rect 21084 35644 21140 35700
rect 14924 35532 14980 35588
rect 16044 35420 16100 35476
rect 48412 35420 48468 35476
rect 15932 35308 15988 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 25900 35084 25956 35140
rect 15484 34972 15540 35028
rect 20188 34972 20244 35028
rect 15372 34860 15428 34916
rect 16268 34860 16324 34916
rect 20412 34636 20468 34692
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 25900 33180 25956 33236
rect 14700 32956 14756 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 17948 32396 18004 32452
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 15372 32060 15428 32116
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 20188 29484 20244 29540
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 42252 28476 42308 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 17948 28028 18004 28084
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 15484 27132 15540 27188
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 17052 25340 17108 25396
rect 16268 25228 16324 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 16268 24108 16324 24164
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 22988 21532 23044 21588
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 26124 18956 26180 19012
rect 27020 18956 27076 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 27468 18620 27524 18676
rect 27132 18396 27188 18452
rect 26852 18060 26908 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 27020 17836 27076 17892
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 26124 14588 26180 14644
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 22988 12460 23044 12516
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 26124 10780 26180 10836
rect 22092 10668 22148 10724
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 22092 10108 22148 10164
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19180 55188 19236 55198
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 18732 54516 18788 54526
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 18620 49588 18676 49598
rect 18620 49028 18676 49532
rect 18732 49364 18788 54460
rect 18732 49298 18788 49308
rect 19180 49364 19236 55132
rect 19808 54908 20128 56420
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19180 49298 19236 49308
rect 19404 54404 19460 54414
rect 18620 48962 18676 48972
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 19404 47348 19460 54348
rect 19404 47282 19460 47292
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 30828 55076 30884 55086
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 19808 47068 20128 48580
rect 30380 49812 30436 49822
rect 30380 48356 30436 49756
rect 30380 48290 30436 48300
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 17164 42868 17220 42878
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 10668 40628 10724 40638
rect 10220 38948 10276 38958
rect 10220 38612 10276 38892
rect 10220 38546 10276 38556
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 10668 37716 10724 40572
rect 16044 40516 16100 40526
rect 10668 37650 10724 37660
rect 14700 39060 14756 39070
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 14140 37268 14196 37278
rect 14140 36260 14196 37212
rect 14140 36194 14196 36204
rect 14588 36596 14644 36606
rect 14588 36260 14644 36540
rect 14588 36194 14644 36204
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 14700 33012 14756 39004
rect 15092 36036 15148 36046
rect 15092 35938 15148 35980
rect 15036 35882 15148 35938
rect 15036 35758 15092 35882
rect 14924 35702 15092 35758
rect 15932 35812 15988 35822
rect 14924 35588 14980 35702
rect 14924 35522 14980 35532
rect 15932 35364 15988 35756
rect 16044 35476 16100 40460
rect 17052 40292 17108 40302
rect 17052 38836 17108 40236
rect 16044 35410 16100 35420
rect 16268 36260 16324 36270
rect 15932 35298 15988 35308
rect 15484 35028 15540 35038
rect 14700 32946 14756 32956
rect 15372 34916 15428 34926
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 15372 32116 15428 34860
rect 15372 32050 15428 32060
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 15484 27188 15540 34972
rect 16268 34916 16324 36204
rect 16268 34850 16324 34860
rect 15484 27122 15540 27132
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 17052 25396 17108 38780
rect 17164 37940 17220 42812
rect 17164 37874 17220 37884
rect 18844 42532 18900 42542
rect 18844 36372 18900 42476
rect 18844 36306 18900 36316
rect 19808 42364 20128 43876
rect 30828 42756 30884 55020
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 30940 53060 30996 53070
rect 30940 49140 30996 53004
rect 30940 49074 30996 49084
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 49756 52052 49812 52062
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 30828 42690 30884 42700
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 40460 51380 40516 51390
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 40236 43204 40292 43214
rect 40236 40964 40292 43148
rect 40236 40898 40292 40908
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 21084 39844 21140 39854
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 20636 39508 20692 39518
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 20188 38500 20244 38510
rect 20188 37604 20244 38444
rect 20188 37538 20244 37548
rect 20412 38500 20468 38510
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 17948 32452 18004 32462
rect 17948 28084 18004 32396
rect 17948 28018 18004 28028
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 20188 35028 20244 35038
rect 20188 29540 20244 34972
rect 20412 34692 20468 38444
rect 20636 36372 20692 39452
rect 20748 38836 20804 38846
rect 20748 37492 20804 38780
rect 20748 37426 20804 37436
rect 20636 36306 20692 36316
rect 21084 35700 21140 39788
rect 21308 38612 21364 38622
rect 21308 37828 21364 38556
rect 21308 37762 21364 37772
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 40460 38500 40516 51324
rect 49084 50596 49140 50606
rect 49084 49700 49140 50540
rect 49084 49634 49140 49644
rect 49308 50148 49364 50158
rect 49308 48692 49364 50092
rect 49308 48626 49364 48636
rect 49756 47460 49812 51996
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 49756 47394 49812 47404
rect 50092 50484 50148 50494
rect 50092 47796 50148 50428
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50204 48580 50260 48590
rect 50204 48020 50260 48524
rect 50204 47954 50260 47964
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50092 47348 50148 47740
rect 50092 47282 50148 47292
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 42364 46676 42420 46686
rect 40460 38434 40516 38444
rect 42252 42756 42308 42766
rect 21084 35634 21140 35644
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 20412 34626 20468 34636
rect 25900 35140 25956 35150
rect 25900 33236 25956 35084
rect 25900 33170 25956 33180
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 20188 29474 20244 29484
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 17052 25330 17108 25340
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 16268 25284 16324 25294
rect 16268 24164 16324 25228
rect 16268 24098 16324 24108
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 42252 28532 42308 42700
rect 42364 42644 42420 46620
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 49196 44548 49252 44558
rect 49196 43652 49252 44492
rect 49196 43586 49252 43596
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 43596 42980 43652 42990
rect 42364 42578 42420 42588
rect 42700 42644 42756 42654
rect 42700 37940 42756 42588
rect 43596 40180 43652 42924
rect 43596 40114 43652 40124
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 42700 37874 42756 37884
rect 48412 39396 48468 39406
rect 48412 35476 48468 39340
rect 48412 35410 48468 35420
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 42252 28466 42308 28476
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 22988 21588 23044 21598
rect 22988 12516 23044 21532
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 22988 12450 23044 12460
rect 26124 19012 26180 19022
rect 26124 14644 26180 18956
rect 27020 19012 27076 19022
rect 26852 18118 26908 18126
rect 27020 18118 27076 18956
rect 27468 18676 27524 18686
rect 27132 18452 27188 18462
rect 27468 18452 27524 18620
rect 27188 18396 27524 18452
rect 27132 18386 27188 18396
rect 26852 18116 27076 18118
rect 26908 18062 27076 18116
rect 26852 18050 26908 18060
rect 27020 17892 27076 18062
rect 27020 17826 27076 17836
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 26124 10836 26180 14588
rect 26124 10770 26180 10780
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 22092 10724 22148 10734
rect 22092 10164 22148 10668
rect 22092 10098 22148 10108
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1341_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15232 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1342_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17136 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1343_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17920 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1344_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1345_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1346_
timestamp 1698431365
transform -1 0 18928 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1347_
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1348_
timestamp 1698431365
transform 1 0 25872 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1349_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24080 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1350_
timestamp 1698431365
transform 1 0 24976 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1351_
timestamp 1698431365
transform -1 0 31584 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1352_
timestamp 1698431365
transform 1 0 30912 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1353_
timestamp 1698431365
transform 1 0 31584 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1354_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1355_
timestamp 1698431365
transform 1 0 24192 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1356_
timestamp 1698431365
transform 1 0 29344 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1357_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29456 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1358_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27104 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1359_
timestamp 1698431365
transform -1 0 24192 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1360_
timestamp 1698431365
transform -1 0 23744 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1361_
timestamp 1698431365
transform 1 0 22960 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1362_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1363_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1364_
timestamp 1698431365
transform 1 0 24080 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1365_
timestamp 1698431365
transform -1 0 30912 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1366_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30464 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1367_
timestamp 1698431365
transform -1 0 29568 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1368_
timestamp 1698431365
transform 1 0 31584 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1369_
timestamp 1698431365
transform -1 0 38416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1370_
timestamp 1698431365
transform -1 0 24640 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1371_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1372_
timestamp 1698431365
transform 1 0 29456 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1373_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30352 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1374_
timestamp 1698431365
transform 1 0 27440 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1375_
timestamp 1698431365
transform 1 0 29120 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1376_
timestamp 1698431365
transform 1 0 27440 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1377_
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1378_
timestamp 1698431365
transform 1 0 25088 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1379_
timestamp 1698431365
transform 1 0 30800 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1380_
timestamp 1698431365
transform -1 0 30912 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1381_
timestamp 1698431365
transform -1 0 38416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1382_
timestamp 1698431365
transform -1 0 31248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1383_
timestamp 1698431365
transform 1 0 26768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1384_
timestamp 1698431365
transform -1 0 31136 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1385_
timestamp 1698431365
transform -1 0 30128 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1386_
timestamp 1698431365
transform 1 0 22848 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1387_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26880 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1388_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1389_
timestamp 1698431365
transform 1 0 25984 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1390_
timestamp 1698431365
transform -1 0 18928 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1391_
timestamp 1698431365
transform 1 0 31696 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1392_
timestamp 1698431365
transform -1 0 23856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1393_
timestamp 1698431365
transform -1 0 16464 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1394_
timestamp 1698431365
transform 1 0 14336 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1395_
timestamp 1698431365
transform 1 0 29568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1396_
timestamp 1698431365
transform 1 0 22400 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1397_
timestamp 1698431365
transform -1 0 23856 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1398_
timestamp 1698431365
transform 1 0 22400 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1399_
timestamp 1698431365
transform 1 0 25200 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1400_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26320 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1401_
timestamp 1698431365
transform 1 0 31584 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1402_
timestamp 1698431365
transform -1 0 42224 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1403_
timestamp 1698431365
transform -1 0 35056 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1404_
timestamp 1698431365
transform -1 0 35280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1405_
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1406_
timestamp 1698431365
transform -1 0 35056 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1407_
timestamp 1698431365
transform 1 0 31696 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1408_
timestamp 1698431365
transform 1 0 41888 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1409_
timestamp 1698431365
transform -1 0 38304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1410_
timestamp 1698431365
transform -1 0 39200 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1411_
timestamp 1698431365
transform -1 0 37520 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1412_
timestamp 1698431365
transform -1 0 36624 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1413_
timestamp 1698431365
transform 1 0 35280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1414_
timestamp 1698431365
transform -1 0 31584 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1415_
timestamp 1698431365
transform -1 0 42560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1416_
timestamp 1698431365
transform -1 0 27888 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1417_
timestamp 1698431365
transform -1 0 35168 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1418_
timestamp 1698431365
transform 1 0 34048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1419_
timestamp 1698431365
transform -1 0 35056 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1420_
timestamp 1698431365
transform -1 0 34272 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1421_
timestamp 1698431365
transform 1 0 32480 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1422_
timestamp 1698431365
transform -1 0 33376 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1423_
timestamp 1698431365
transform -1 0 29120 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1424_
timestamp 1698431365
transform -1 0 27104 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1425_
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1426_
timestamp 1698431365
transform 1 0 27888 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1427_
timestamp 1698431365
transform -1 0 29120 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1428_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1429_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28784 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1430_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1431_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1432_
timestamp 1698431365
transform -1 0 29120 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1433_
timestamp 1698431365
transform 1 0 27664 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1434_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1435_
timestamp 1698431365
transform -1 0 15344 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1436_
timestamp 1698431365
transform 1 0 23744 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1437_
timestamp 1698431365
transform -1 0 24192 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1438_
timestamp 1698431365
transform -1 0 34720 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1439_
timestamp 1698431365
transform -1 0 25760 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1440_
timestamp 1698431365
transform -1 0 25200 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1441_
timestamp 1698431365
transform 1 0 23520 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1442_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1443_
timestamp 1698431365
transform -1 0 38864 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1444_
timestamp 1698431365
transform -1 0 30352 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1445_
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1446_
timestamp 1698431365
transform -1 0 28784 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1447_
timestamp 1698431365
transform -1 0 27664 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1448_
timestamp 1698431365
transform 1 0 25760 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1449_
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1450_
timestamp 1698431365
transform -1 0 15008 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1451_
timestamp 1698431365
transform -1 0 25760 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1452_
timestamp 1698431365
transform 1 0 24304 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1453_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1454_
timestamp 1698431365
transform 1 0 23856 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1455_
timestamp 1698431365
transform 1 0 25424 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1456_
timestamp 1698431365
transform -1 0 26320 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1457_
timestamp 1698431365
transform -1 0 43680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1458_
timestamp 1698431365
transform -1 0 35728 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1459_
timestamp 1698431365
transform -1 0 35504 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1460_
timestamp 1698431365
transform 1 0 35616 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1461_
timestamp 1698431365
transform 1 0 35952 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1462_
timestamp 1698431365
transform 1 0 41888 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1463_
timestamp 1698431365
transform -1 0 38192 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1464_
timestamp 1698431365
transform -1 0 37744 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1465_
timestamp 1698431365
transform -1 0 37408 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1466_
timestamp 1698431365
transform -1 0 36288 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1467_
timestamp 1698431365
transform -1 0 35952 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1468_
timestamp 1698431365
transform -1 0 43120 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1469_
timestamp 1698431365
transform -1 0 33824 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1470_
timestamp 1698431365
transform 1 0 31808 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1471_
timestamp 1698431365
transform -1 0 33376 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1472_
timestamp 1698431365
transform -1 0 32704 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1473_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1474_
timestamp 1698431365
transform -1 0 32592 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1475_
timestamp 1698431365
transform -1 0 24864 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1476_
timestamp 1698431365
transform 1 0 23408 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1477_
timestamp 1698431365
transform 1 0 15792 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1478_
timestamp 1698431365
transform -1 0 24640 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1479_
timestamp 1698431365
transform 1 0 23744 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1480_
timestamp 1698431365
transform 1 0 26208 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1481_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1482_
timestamp 1698431365
transform -1 0 28784 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1483_
timestamp 1698431365
transform 1 0 25872 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1484_
timestamp 1698431365
transform 1 0 27216 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1485_
timestamp 1698431365
transform 1 0 14560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1486_
timestamp 1698431365
transform 1 0 4816 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1487_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5824 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1488_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9744 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1489_
timestamp 1698431365
transform 1 0 14224 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1490_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14672 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1491_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10752 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1492_
timestamp 1698431365
transform 1 0 7392 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1493_
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1494_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14448 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1495_
timestamp 1698431365
transform -1 0 12208 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1496_
timestamp 1698431365
transform 1 0 14784 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1497_
timestamp 1698431365
transform 1 0 15120 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1498_
timestamp 1698431365
transform 1 0 15008 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1499_
timestamp 1698431365
transform 1 0 15792 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1500_
timestamp 1698431365
transform 1 0 29680 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1501_
timestamp 1698431365
transform -1 0 30240 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1502_
timestamp 1698431365
transform 1 0 15792 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1503_
timestamp 1698431365
transform -1 0 11984 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1504_
timestamp 1698431365
transform -1 0 8736 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1505_
timestamp 1698431365
transform 1 0 10864 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1506_
timestamp 1698431365
transform 1 0 11760 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1507_
timestamp 1698431365
transform -1 0 6384 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1508_
timestamp 1698431365
transform 1 0 7168 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1509_
timestamp 1698431365
transform 1 0 4592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1510_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5040 0 -1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1511_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12320 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1512_
timestamp 1698431365
transform -1 0 10304 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1513_
timestamp 1698431365
transform -1 0 11088 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1514_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10416 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1515_
timestamp 1698431365
transform -1 0 10752 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1516_
timestamp 1698431365
transform -1 0 7504 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1517_
timestamp 1698431365
transform 1 0 30016 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1518_
timestamp 1698431365
transform 1 0 31136 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1519_
timestamp 1698431365
transform 1 0 22400 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1520_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11424 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1521_
timestamp 1698431365
transform 1 0 19712 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1522_
timestamp 1698431365
transform 1 0 16128 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1523_
timestamp 1698431365
transform 1 0 11872 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1524_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1525_
timestamp 1698431365
transform -1 0 20496 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1526_
timestamp 1698431365
transform 1 0 16352 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1527_
timestamp 1698431365
transform 1 0 16464 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1528_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1529_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19376 0 1 54880
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1530_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17360 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1531_
timestamp 1698431365
transform 1 0 20720 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1532_
timestamp 1698431365
transform -1 0 22288 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1533_
timestamp 1698431365
transform -1 0 17248 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1534_
timestamp 1698431365
transform 1 0 10416 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1535_
timestamp 1698431365
transform -1 0 4592 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1536_
timestamp 1698431365
transform 1 0 4592 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1537_
timestamp 1698431365
transform 1 0 5040 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1538_
timestamp 1698431365
transform 1 0 7840 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1539_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8512 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1540_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11648 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1541_
timestamp 1698431365
transform 1 0 14560 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1542_
timestamp 1698431365
transform 1 0 9072 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1543_
timestamp 1698431365
transform -1 0 9744 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1544_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1545_
timestamp 1698431365
transform 1 0 10528 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1546_
timestamp 1698431365
transform -1 0 14448 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1547_
timestamp 1698431365
transform -1 0 7504 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1548_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6496 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1549_
timestamp 1698431365
transform 1 0 10080 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1550_
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1551_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7056 0 -1 25088
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1552_
timestamp 1698431365
transform 1 0 13664 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1553_
timestamp 1698431365
transform -1 0 15792 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1554_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1555_
timestamp 1698431365
transform -1 0 9072 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1556_
timestamp 1698431365
transform 1 0 9632 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1557_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15008 0 -1 23520
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1558_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1559_
timestamp 1698431365
transform 1 0 9968 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1560_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14224 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1561_
timestamp 1698431365
transform -1 0 11984 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1562_
timestamp 1698431365
transform 1 0 10640 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1563_
timestamp 1698431365
transform 1 0 11984 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1564_
timestamp 1698431365
transform -1 0 24752 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1565_
timestamp 1698431365
transform -1 0 16352 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1566_
timestamp 1698431365
transform -1 0 15120 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1567_
timestamp 1698431365
transform 1 0 9744 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1568_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13216 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1569_
timestamp 1698431365
transform 1 0 10416 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1570_
timestamp 1698431365
transform -1 0 22064 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1571_
timestamp 1698431365
transform 1 0 21280 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1572_
timestamp 1698431365
transform -1 0 23408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1573_
timestamp 1698431365
transform -1 0 13888 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1574_
timestamp 1698431365
transform 1 0 13664 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1575_
timestamp 1698431365
transform 1 0 11312 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1576_
timestamp 1698431365
transform 1 0 15456 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1577_
timestamp 1698431365
transform 1 0 14672 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1578_
timestamp 1698431365
transform -1 0 14896 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1579_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1580_
timestamp 1698431365
transform 1 0 13776 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1581_
timestamp 1698431365
transform 1 0 24192 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1582_
timestamp 1698431365
transform -1 0 34384 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1583_
timestamp 1698431365
transform -1 0 33824 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1584_
timestamp 1698431365
transform 1 0 33824 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1585_
timestamp 1698431365
transform 1 0 35504 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1586_
timestamp 1698431365
transform -1 0 37296 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1587_
timestamp 1698431365
transform 1 0 29456 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1588_
timestamp 1698431365
transform 1 0 22624 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1589_
timestamp 1698431365
transform 1 0 23632 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1590_
timestamp 1698431365
transform 1 0 22736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1591_
timestamp 1698431365
transform 1 0 23072 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1592_
timestamp 1698431365
transform -1 0 24864 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1593_
timestamp 1698431365
transform 1 0 18704 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1594_
timestamp 1698431365
transform -1 0 23072 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1595_
timestamp 1698431365
transform -1 0 23072 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1596_
timestamp 1698431365
transform 1 0 25536 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1597_
timestamp 1698431365
transform 1 0 26880 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1598_
timestamp 1698431365
transform -1 0 24304 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1599_
timestamp 1698431365
transform 1 0 26096 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1600_
timestamp 1698431365
transform 1 0 23296 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1601_
timestamp 1698431365
transform 1 0 23744 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1602_
timestamp 1698431365
transform 1 0 25760 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1603_
timestamp 1698431365
transform 1 0 27888 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1604_
timestamp 1698431365
transform -1 0 34720 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1605_
timestamp 1698431365
transform 1 0 32480 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1606_
timestamp 1698431365
transform 1 0 23632 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1607_
timestamp 1698431365
transform 1 0 26096 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1608_
timestamp 1698431365
transform -1 0 24864 0 -1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1609_
timestamp 1698431365
transform 1 0 27104 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1610_
timestamp 1698431365
transform 1 0 31024 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1611_
timestamp 1698431365
transform 1 0 31584 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1612_
timestamp 1698431365
transform 1 0 26432 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1613_
timestamp 1698431365
transform 1 0 27888 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1614_
timestamp 1698431365
transform 1 0 27104 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1615_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1616_
timestamp 1698431365
transform 1 0 27776 0 -1 48608
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1617_
timestamp 1698431365
transform -1 0 32704 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1618_
timestamp 1698431365
transform 1 0 30464 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1619_
timestamp 1698431365
transform -1 0 29568 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1620_
timestamp 1698431365
transform -1 0 28448 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1621_
timestamp 1698431365
transform 1 0 25200 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1622_
timestamp 1698431365
transform -1 0 27104 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1698431365
transform 1 0 25312 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1624_
timestamp 1698431365
transform -1 0 27664 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1625_
timestamp 1698431365
transform -1 0 26880 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1626_
timestamp 1698431365
transform 1 0 28560 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1627_
timestamp 1698431365
transform 1 0 27664 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1628_
timestamp 1698431365
transform -1 0 30128 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1629_
timestamp 1698431365
transform -1 0 25760 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1630_
timestamp 1698431365
transform 1 0 27888 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1631_
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1632_
timestamp 1698431365
transform 1 0 29568 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1633_
timestamp 1698431365
transform 1 0 31808 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1634_
timestamp 1698431365
transform -1 0 32480 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1635_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31136 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1636_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1637_
timestamp 1698431365
transform -1 0 28336 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1638_
timestamp 1698431365
transform -1 0 28224 0 1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1639_
timestamp 1698431365
transform 1 0 29232 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1640_
timestamp 1698431365
transform 1 0 29456 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1641_
timestamp 1698431365
transform 1 0 30128 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1642_
timestamp 1698431365
transform -1 0 27552 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1643_
timestamp 1698431365
transform 1 0 28560 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1644_
timestamp 1698431365
transform 1 0 30128 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1645_
timestamp 1698431365
transform 1 0 30576 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1646_
timestamp 1698431365
transform -1 0 32704 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1647_
timestamp 1698431365
transform -1 0 33376 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1648_
timestamp 1698431365
transform -1 0 29120 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1649_
timestamp 1698431365
transform 1 0 32144 0 1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1650_
timestamp 1698431365
transform -1 0 32704 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1651_
timestamp 1698431365
transform -1 0 32368 0 1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1652_
timestamp 1698431365
transform 1 0 31136 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1653_
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1654_
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1655_
timestamp 1698431365
transform -1 0 32144 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1656_
timestamp 1698431365
transform 1 0 15568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1657_
timestamp 1698431365
transform 1 0 15456 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1658_
timestamp 1698431365
transform -1 0 17920 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1659_
timestamp 1698431365
transform -1 0 16912 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1660_
timestamp 1698431365
transform 1 0 15456 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1661_
timestamp 1698431365
transform 1 0 16128 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1662_
timestamp 1698431365
transform 1 0 34608 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1663_
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1664_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16464 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1665_
timestamp 1698431365
transform -1 0 20944 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1666_
timestamp 1698431365
transform -1 0 20384 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1667_
timestamp 1698431365
transform 1 0 18928 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1668_
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1669_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1670_
timestamp 1698431365
transform 1 0 18816 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1671_
timestamp 1698431365
transform 1 0 15120 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1672_
timestamp 1698431365
transform -1 0 6496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1673_
timestamp 1698431365
transform 1 0 18480 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1674_
timestamp 1698431365
transform 1 0 13664 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1675_
timestamp 1698431365
transform -1 0 19712 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1676_
timestamp 1698431365
transform 1 0 15904 0 1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1677_
timestamp 1698431365
transform -1 0 17696 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1678_
timestamp 1698431365
transform 1 0 18144 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1679_
timestamp 1698431365
transform -1 0 18816 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1680_
timestamp 1698431365
transform -1 0 17696 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1681_
timestamp 1698431365
transform 1 0 10752 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1682_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11984 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1683_
timestamp 1698431365
transform -1 0 13664 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1684_
timestamp 1698431365
transform 1 0 15792 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1685_
timestamp 1698431365
transform -1 0 16912 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1686_
timestamp 1698431365
transform 1 0 30352 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1687_
timestamp 1698431365
transform 1 0 30912 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1688_
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1689_
timestamp 1698431365
transform 1 0 10976 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1690_
timestamp 1698431365
transform -1 0 14224 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1691_
timestamp 1698431365
transform 1 0 14224 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1692_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1693_
timestamp 1698431365
transform 1 0 16352 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1694_
timestamp 1698431365
transform -1 0 17024 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1695_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18816 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1696_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1697_
timestamp 1698431365
transform 1 0 18928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1698_
timestamp 1698431365
transform 1 0 20048 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1699_
timestamp 1698431365
transform 1 0 17584 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1700_
timestamp 1698431365
transform 1 0 37968 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1701_
timestamp 1698431365
transform 1 0 41888 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1702_
timestamp 1698431365
transform -1 0 42560 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1703_
timestamp 1698431365
transform 1 0 31248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1704_
timestamp 1698431365
transform -1 0 32032 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1705_
timestamp 1698431365
transform 1 0 38640 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1706_
timestamp 1698431365
transform 1 0 41664 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1707_
timestamp 1698431365
transform 1 0 41216 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1708_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1709_
timestamp 1698431365
transform 1 0 18816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1710_
timestamp 1698431365
transform 1 0 21840 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1711_
timestamp 1698431365
transform 1 0 21168 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1712_
timestamp 1698431365
transform 1 0 38864 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1713_
timestamp 1698431365
transform -1 0 45248 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1714_
timestamp 1698431365
transform 1 0 43792 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1715_
timestamp 1698431365
transform -1 0 45024 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1716_
timestamp 1698431365
transform 1 0 43680 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1717_
timestamp 1698431365
transform 1 0 31136 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1718_
timestamp 1698431365
transform -1 0 21840 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1719_
timestamp 1698431365
transform 1 0 16240 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1720_
timestamp 1698431365
transform 1 0 13888 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1721_
timestamp 1698431365
transform -1 0 14000 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1722_
timestamp 1698431365
transform 1 0 31808 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1723_
timestamp 1698431365
transform -1 0 18032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1724_
timestamp 1698431365
transform 1 0 14112 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1725_
timestamp 1698431365
transform -1 0 14112 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1726_
timestamp 1698431365
transform 1 0 17360 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1727_
timestamp 1698431365
transform 1 0 19264 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1728_
timestamp 1698431365
transform 1 0 21840 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1729_
timestamp 1698431365
transform 1 0 37744 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1730_
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1731_
timestamp 1698431365
transform 1 0 38192 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1732_
timestamp 1698431365
transform -1 0 40208 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1733_
timestamp 1698431365
transform 1 0 39200 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1734_
timestamp 1698431365
transform 1 0 15568 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1735_
timestamp 1698431365
transform 1 0 17584 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1736_
timestamp 1698431365
transform 1 0 38304 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1737_
timestamp 1698431365
transform -1 0 40544 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1738_
timestamp 1698431365
transform 1 0 39536 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1739_
timestamp 1698431365
transform 1 0 38752 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1740_
timestamp 1698431365
transform 1 0 39312 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1741_
timestamp 1698431365
transform 1 0 20608 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1742_
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1743_
timestamp 1698431365
transform 1 0 33376 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1744_
timestamp 1698431365
transform 1 0 38528 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1745_
timestamp 1698431365
transform 1 0 33600 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1746_
timestamp 1698431365
transform 1 0 39872 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1747_
timestamp 1698431365
transform 1 0 39648 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1748_
timestamp 1698431365
transform 1 0 34944 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1749_
timestamp 1698431365
transform 1 0 38976 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1750_
timestamp 1698431365
transform 1 0 38752 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1751_
timestamp 1698431365
transform -1 0 36288 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1752_
timestamp 1698431365
transform -1 0 36736 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1753_
timestamp 1698431365
transform -1 0 36848 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1754_
timestamp 1698431365
transform 1 0 36848 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1755_
timestamp 1698431365
transform -1 0 29680 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1756_
timestamp 1698431365
transform 1 0 34384 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1757_
timestamp 1698431365
transform 1 0 34272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1758_
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1759_
timestamp 1698431365
transform -1 0 20608 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1760_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1761_
timestamp 1698431365
transform 1 0 20496 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1762_
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1763_
timestamp 1698431365
transform -1 0 32256 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1764_
timestamp 1698431365
transform 1 0 34048 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1765_
timestamp 1698431365
transform 1 0 31808 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1766_
timestamp 1698431365
transform 1 0 32032 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1767_
timestamp 1698431365
transform -1 0 18032 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1768_
timestamp 1698431365
transform 1 0 17360 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1769_
timestamp 1698431365
transform 1 0 21392 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1770_
timestamp 1698431365
transform -1 0 34048 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1771_
timestamp 1698431365
transform 1 0 31696 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1772_
timestamp 1698431365
transform -1 0 31472 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1773_
timestamp 1698431365
transform 1 0 31808 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1774_
timestamp 1698431365
transform -1 0 31472 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1775_
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1776_
timestamp 1698431365
transform 1 0 38976 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1777_
timestamp 1698431365
transform -1 0 40544 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1778_
timestamp 1698431365
transform -1 0 39984 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1779_
timestamp 1698431365
transform -1 0 40880 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1780_
timestamp 1698431365
transform -1 0 33488 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1781_
timestamp 1698431365
transform 1 0 31024 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1782_
timestamp 1698431365
transform -1 0 30800 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1783_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1784_
timestamp 1698431365
transform 1 0 29904 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1785_
timestamp 1698431365
transform 1 0 11872 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1786_
timestamp 1698431365
transform -1 0 17248 0 1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1787_
timestamp 1698431365
transform 1 0 26320 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1788_
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1789_
timestamp 1698431365
transform -1 0 26096 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1790_
timestamp 1698431365
transform 1 0 27104 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1791_
timestamp 1698431365
transform -1 0 27552 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1792_
timestamp 1698431365
transform -1 0 22400 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1793_
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1794_
timestamp 1698431365
transform 1 0 17136 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1795_
timestamp 1698431365
transform -1 0 17696 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1796_
timestamp 1698431365
transform 1 0 13776 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1797_
timestamp 1698431365
transform -1 0 11872 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1798_
timestamp 1698431365
transform -1 0 23184 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1799_
timestamp 1698431365
transform 1 0 14560 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1800_
timestamp 1698431365
transform -1 0 14000 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1801_
timestamp 1698431365
transform -1 0 14672 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1802_
timestamp 1698431365
transform 1 0 15904 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1803_
timestamp 1698431365
transform 1 0 17696 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1804_
timestamp 1698431365
transform -1 0 15344 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1805_
timestamp 1698431365
transform -1 0 14896 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1806_
timestamp 1698431365
transform -1 0 13776 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1807_
timestamp 1698431365
transform 1 0 14224 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1808_
timestamp 1698431365
transform 1 0 14896 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1809_
timestamp 1698431365
transform -1 0 10752 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1810_
timestamp 1698431365
transform -1 0 8176 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1811_
timestamp 1698431365
transform -1 0 8512 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1812_
timestamp 1698431365
transform -1 0 8064 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1813_
timestamp 1698431365
transform -1 0 7728 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1814_
timestamp 1698431365
transform -1 0 10416 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1815_
timestamp 1698431365
transform 1 0 6160 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1816_
timestamp 1698431365
transform -1 0 7728 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1817_
timestamp 1698431365
transform 1 0 6384 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1818_
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1819_
timestamp 1698431365
transform 1 0 7728 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1820_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8176 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1821_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1822_
timestamp 1698431365
transform 1 0 14896 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1823_
timestamp 1698431365
transform 1 0 15680 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1824_
timestamp 1698431365
transform -1 0 22736 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1825_
timestamp 1698431365
transform -1 0 20944 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1826_
timestamp 1698431365
transform 1 0 20160 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1827_
timestamp 1698431365
transform -1 0 22064 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1828_
timestamp 1698431365
transform -1 0 21840 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1829_
timestamp 1698431365
transform -1 0 22736 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1830_
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1831_
timestamp 1698431365
transform 1 0 20384 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1832_
timestamp 1698431365
transform -1 0 20272 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1833_
timestamp 1698431365
transform 1 0 19264 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1834_
timestamp 1698431365
transform -1 0 19264 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1835_
timestamp 1698431365
transform -1 0 22624 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1836_
timestamp 1698431365
transform 1 0 20608 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1837_
timestamp 1698431365
transform -1 0 20608 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1838_
timestamp 1698431365
transform -1 0 19376 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1839_
timestamp 1698431365
transform -1 0 17024 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1840_
timestamp 1698431365
transform -1 0 18144 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1841_
timestamp 1698431365
transform -1 0 17920 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1842_
timestamp 1698431365
transform -1 0 16800 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1843_
timestamp 1698431365
transform -1 0 17248 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1844_
timestamp 1698431365
transform -1 0 18704 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1845_
timestamp 1698431365
transform -1 0 17024 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1846_
timestamp 1698431365
transform 1 0 15904 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1847_
timestamp 1698431365
transform 1 0 15680 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1848_
timestamp 1698431365
transform 1 0 17696 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1849_
timestamp 1698431365
transform 1 0 17584 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1850_
timestamp 1698431365
transform 1 0 19264 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1851_
timestamp 1698431365
transform -1 0 15904 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1852_
timestamp 1698431365
transform 1 0 16912 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1853_
timestamp 1698431365
transform -1 0 18592 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1854_
timestamp 1698431365
transform 1 0 16128 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1855_
timestamp 1698431365
transform -1 0 37744 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1856_
timestamp 1698431365
transform -1 0 40320 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1857_
timestamp 1698431365
transform -1 0 38752 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1858_
timestamp 1698431365
transform -1 0 37520 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1859_
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1860_
timestamp 1698431365
transform 1 0 40320 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1861_
timestamp 1698431365
transform 1 0 35728 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1862_
timestamp 1698431365
transform -1 0 41664 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1863_
timestamp 1698431365
transform 1 0 41776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1864_
timestamp 1698431365
transform -1 0 39648 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1865_
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1866_
timestamp 1698431365
transform 1 0 36960 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1867_
timestamp 1698431365
transform -1 0 39088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1868_
timestamp 1698431365
transform -1 0 39312 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1869_
timestamp 1698431365
transform -1 0 38528 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1870_
timestamp 1698431365
transform 1 0 39200 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform 1 0 41104 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1872_
timestamp 1698431365
transform -1 0 37520 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1873_
timestamp 1698431365
transform 1 0 38640 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1874_
timestamp 1698431365
transform 1 0 37520 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1875_
timestamp 1698431365
transform 1 0 37520 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1876_
timestamp 1698431365
transform 1 0 39536 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1877_
timestamp 1698431365
transform -1 0 36624 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1878_
timestamp 1698431365
transform 1 0 39312 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1879_
timestamp 1698431365
transform 1 0 39984 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1880_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1881_
timestamp 1698431365
transform -1 0 42672 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1882_
timestamp 1698431365
transform -1 0 41328 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1883_
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1884_
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1885_
timestamp 1698431365
transform 1 0 43456 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1886_
timestamp 1698431365
transform -1 0 38192 0 -1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1887_
timestamp 1698431365
transform -1 0 31696 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1888_
timestamp 1698431365
transform 1 0 34608 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1889_
timestamp 1698431365
transform -1 0 35616 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1890_
timestamp 1698431365
transform -1 0 37856 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1891_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37072 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1892_
timestamp 1698431365
transform 1 0 35504 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1893_
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1894_
timestamp 1698431365
transform -1 0 45360 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1895_
timestamp 1698431365
transform -1 0 57904 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1896_
timestamp 1698431365
transform -1 0 43792 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1897_
timestamp 1698431365
transform 1 0 42224 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1898_
timestamp 1698431365
transform 1 0 45584 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1899_
timestamp 1698431365
transform 1 0 47040 0 1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1900_
timestamp 1698431365
transform -1 0 57344 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1901_
timestamp 1698431365
transform 1 0 56896 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1902_
timestamp 1698431365
transform 1 0 39872 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1903_
timestamp 1698431365
transform 1 0 43120 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1904_
timestamp 1698431365
transform 1 0 46816 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1905_
timestamp 1698431365
transform 1 0 44016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1906_
timestamp 1698431365
transform 1 0 44800 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1907_
timestamp 1698431365
transform 1 0 44688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1908_
timestamp 1698431365
transform 1 0 43792 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1909_
timestamp 1698431365
transform -1 0 45472 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1910_
timestamp 1698431365
transform -1 0 43344 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1911_
timestamp 1698431365
transform 1 0 42224 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1912_
timestamp 1698431365
transform 1 0 42896 0 -1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1913_
timestamp 1698431365
transform -1 0 37296 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1914_
timestamp 1698431365
transform 1 0 42896 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1915_
timestamp 1698431365
transform -1 0 43456 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1916_
timestamp 1698431365
transform 1 0 35952 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1917_
timestamp 1698431365
transform -1 0 42336 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1918_
timestamp 1698431365
transform 1 0 33040 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1919_
timestamp 1698431365
transform 1 0 36400 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1920_
timestamp 1698431365
transform 1 0 35728 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1921_
timestamp 1698431365
transform -1 0 43120 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1922_
timestamp 1698431365
transform 1 0 41776 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1923_
timestamp 1698431365
transform 1 0 42896 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1924_
timestamp 1698431365
transform 1 0 42000 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1925_
timestamp 1698431365
transform 1 0 44576 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1926_
timestamp 1698431365
transform 1 0 44016 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1927_
timestamp 1698431365
transform -1 0 49168 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1928_
timestamp 1698431365
transform -1 0 50400 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1929_
timestamp 1698431365
transform 1 0 49168 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1930_
timestamp 1698431365
transform -1 0 46144 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1931_
timestamp 1698431365
transform -1 0 51968 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1932_
timestamp 1698431365
transform 1 0 46816 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1933_
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1934_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45584 0 1 43904
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1935_
timestamp 1698431365
transform -1 0 57680 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1936_
timestamp 1698431365
transform -1 0 55664 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1937_
timestamp 1698431365
transform 1 0 49952 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1698431365
transform -1 0 50624 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1939_
timestamp 1698431365
transform 1 0 41552 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1940_
timestamp 1698431365
transform -1 0 44128 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1941_
timestamp 1698431365
transform 1 0 41776 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1942_
timestamp 1698431365
transform -1 0 43232 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1943_
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1944_
timestamp 1698431365
transform -1 0 44464 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1945_
timestamp 1698431365
transform 1 0 42672 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1946_
timestamp 1698431365
transform 1 0 43232 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1947_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47040 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1948_
timestamp 1698431365
transform -1 0 49280 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1949_
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1950_
timestamp 1698431365
transform 1 0 42336 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1951_
timestamp 1698431365
transform 1 0 45360 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1952_
timestamp 1698431365
transform -1 0 42784 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1953_
timestamp 1698431365
transform 1 0 39648 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1954_
timestamp 1698431365
transform 1 0 38416 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1955_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37968 0 -1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1956_
timestamp 1698431365
transform -1 0 40544 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1957_
timestamp 1698431365
transform 1 0 39536 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1958_
timestamp 1698431365
transform 1 0 39200 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1959_
timestamp 1698431365
transform -1 0 46256 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1960_
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1961_
timestamp 1698431365
transform 1 0 44240 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1962_
timestamp 1698431365
transform 1 0 43456 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1963_
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1964_
timestamp 1698431365
transform 1 0 46032 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1965_
timestamp 1698431365
transform -1 0 46928 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1966_
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1967_
timestamp 1698431365
transform 1 0 42784 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1968_
timestamp 1698431365
transform -1 0 41440 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1969_
timestamp 1698431365
transform 1 0 42448 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1970_
timestamp 1698431365
transform -1 0 39200 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1971_
timestamp 1698431365
transform 1 0 40880 0 -1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1972_
timestamp 1698431365
transform 1 0 42784 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1973_
timestamp 1698431365
transform -1 0 46032 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1974_
timestamp 1698431365
transform 1 0 44128 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1975_
timestamp 1698431365
transform -1 0 43904 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1976_
timestamp 1698431365
transform 1 0 40992 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1977_
timestamp 1698431365
transform 1 0 45472 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1978_
timestamp 1698431365
transform 1 0 41104 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1979_
timestamp 1698431365
transform 1 0 43344 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1980_
timestamp 1698431365
transform 1 0 37856 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1981_
timestamp 1698431365
transform 1 0 37184 0 -1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1982_
timestamp 1698431365
transform 1 0 37184 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1983_
timestamp 1698431365
transform 1 0 38640 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1984_
timestamp 1698431365
transform -1 0 40992 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1985_
timestamp 1698431365
transform -1 0 39648 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1986_
timestamp 1698431365
transform 1 0 38976 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1987_
timestamp 1698431365
transform 1 0 39088 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1988_
timestamp 1698431365
transform 1 0 38080 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1989_
timestamp 1698431365
transform 1 0 39984 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1990_
timestamp 1698431365
transform 1 0 46256 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1991_
timestamp 1698431365
transform -1 0 42448 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1992_
timestamp 1698431365
transform 1 0 42336 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1993_
timestamp 1698431365
transform 1 0 41216 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1994_
timestamp 1698431365
transform -1 0 41216 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1995_
timestamp 1698431365
transform 1 0 45360 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1996_
timestamp 1698431365
transform -1 0 43568 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1997_
timestamp 1698431365
transform -1 0 41664 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1998_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42784 0 1 39200
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1999_
timestamp 1698431365
transform 1 0 35392 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2000_
timestamp 1698431365
transform -1 0 37520 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2001_
timestamp 1698431365
transform 1 0 37856 0 1 37632
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2002_
timestamp 1698431365
transform 1 0 37072 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2003_
timestamp 1698431365
transform 1 0 38304 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2004_
timestamp 1698431365
transform 1 0 39312 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2005_
timestamp 1698431365
transform -1 0 41104 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2006_
timestamp 1698431365
transform 1 0 37520 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2007_
timestamp 1698431365
transform 1 0 44912 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2008_
timestamp 1698431365
transform 1 0 46480 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2009_
timestamp 1698431365
transform 1 0 39424 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2010_
timestamp 1698431365
transform 1 0 31808 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2011_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39312 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2012_
timestamp 1698431365
transform 1 0 45584 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2013_
timestamp 1698431365
transform -1 0 35392 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2014_
timestamp 1698431365
transform 1 0 46704 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2015_
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2016_
timestamp 1698431365
transform 1 0 39648 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2017_
timestamp 1698431365
transform -1 0 34944 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2018_
timestamp 1698431365
transform 1 0 37184 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2019_
timestamp 1698431365
transform 1 0 37744 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2020_
timestamp 1698431365
transform 1 0 36288 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2021_
timestamp 1698431365
transform 1 0 36064 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2022_
timestamp 1698431365
transform 1 0 37520 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2023_
timestamp 1698431365
transform -1 0 39648 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2024_
timestamp 1698431365
transform -1 0 38752 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2025_
timestamp 1698431365
transform 1 0 38304 0 -1 36064
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2026_
timestamp 1698431365
transform 1 0 35168 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2027_
timestamp 1698431365
transform 1 0 39760 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2028_
timestamp 1698431365
transform -1 0 40432 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2029_
timestamp 1698431365
transform 1 0 30688 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2030_
timestamp 1698431365
transform -1 0 33824 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2031_
timestamp 1698431365
transform 1 0 40544 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2032_
timestamp 1698431365
transform 1 0 34160 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2033_
timestamp 1698431365
transform -1 0 36400 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2034_
timestamp 1698431365
transform 1 0 31696 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2035_
timestamp 1698431365
transform 1 0 34160 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2036_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39536 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2037_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37856 0 1 42336
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2038_
timestamp 1698431365
transform -1 0 37856 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2039_
timestamp 1698431365
transform 1 0 37744 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2040_
timestamp 1698431365
transform -1 0 37968 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2041_
timestamp 1698431365
transform 1 0 37968 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2042_
timestamp 1698431365
transform 1 0 27776 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2043_
timestamp 1698431365
transform 1 0 28560 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2044_
timestamp 1698431365
transform 1 0 38528 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2045_
timestamp 1698431365
transform 1 0 33264 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2046_
timestamp 1698431365
transform 1 0 34272 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2047_
timestamp 1698431365
transform 1 0 35168 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2048_
timestamp 1698431365
transform -1 0 36624 0 1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2049_
timestamp 1698431365
transform 1 0 35728 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2050_
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2051_
timestamp 1698431365
transform -1 0 38864 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2052_
timestamp 1698431365
transform 1 0 37632 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2053_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37968 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2054_
timestamp 1698431365
transform -1 0 32592 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2055_
timestamp 1698431365
transform 1 0 36176 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2056_
timestamp 1698431365
transform 1 0 36176 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2057_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2058_
timestamp 1698431365
transform -1 0 49280 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2059_
timestamp 1698431365
transform 1 0 38864 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2060_
timestamp 1698431365
transform 1 0 39424 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2061_
timestamp 1698431365
transform 1 0 38528 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2062_
timestamp 1698431365
transform 1 0 31248 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2063_
timestamp 1698431365
transform -1 0 38528 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2064_
timestamp 1698431365
transform 1 0 40656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2065_
timestamp 1698431365
transform 1 0 45360 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2066_
timestamp 1698431365
transform 1 0 36064 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2067_
timestamp 1698431365
transform 1 0 36400 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2068_
timestamp 1698431365
transform 1 0 38304 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2069_
timestamp 1698431365
transform 1 0 38304 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2070_
timestamp 1698431365
transform 1 0 38752 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2071_
timestamp 1698431365
transform 1 0 37408 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2072_
timestamp 1698431365
transform 1 0 38864 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2073_
timestamp 1698431365
transform -1 0 42224 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2074_
timestamp 1698431365
transform -1 0 42224 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2075_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2076_
timestamp 1698431365
transform 1 0 38752 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2077_
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2078_
timestamp 1698431365
transform -1 0 40544 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2079_
timestamp 1698431365
transform -1 0 40544 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2080_
timestamp 1698431365
transform 1 0 39312 0 -1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2081_
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2082_
timestamp 1698431365
transform -1 0 42000 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2083_
timestamp 1698431365
transform -1 0 42336 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2084_
timestamp 1698431365
transform 1 0 42000 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2085_
timestamp 1698431365
transform -1 0 42560 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2086_
timestamp 1698431365
transform 1 0 42448 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2087_
timestamp 1698431365
transform -1 0 44352 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2088_
timestamp 1698431365
transform -1 0 40544 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2089_
timestamp 1698431365
transform 1 0 39872 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2090_
timestamp 1698431365
transform -1 0 46480 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2091_
timestamp 1698431365
transform 1 0 40544 0 1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2092_
timestamp 1698431365
transform -1 0 46480 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2093_
timestamp 1698431365
transform 1 0 16464 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2094_
timestamp 1698431365
transform 1 0 42784 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2095_
timestamp 1698431365
transform 1 0 42224 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2096_
timestamp 1698431365
transform -1 0 41776 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2097_
timestamp 1698431365
transform -1 0 43456 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2098_
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2099_
timestamp 1698431365
transform -1 0 45808 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2100_
timestamp 1698431365
transform 1 0 40544 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2101_
timestamp 1698431365
transform -1 0 45472 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2102_
timestamp 1698431365
transform 1 0 44464 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2103_
timestamp 1698431365
transform 1 0 45920 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2104_
timestamp 1698431365
transform -1 0 44464 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2105_
timestamp 1698431365
transform -1 0 44800 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2106_
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2107_
timestamp 1698431365
transform -1 0 44688 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _2108_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37296 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2109_
timestamp 1698431365
transform -1 0 54096 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2110_
timestamp 1698431365
transform -1 0 47824 0 1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2111_
timestamp 1698431365
transform 1 0 46368 0 -1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2112_
timestamp 1698431365
transform 1 0 46704 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2113_
timestamp 1698431365
transform -1 0 50960 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2114_
timestamp 1698431365
transform -1 0 47488 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2115_
timestamp 1698431365
transform -1 0 46368 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2116_
timestamp 1698431365
transform -1 0 46704 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2117_
timestamp 1698431365
transform 1 0 44800 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2118_
timestamp 1698431365
transform 1 0 43456 0 -1 51744
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2119_
timestamp 1698431365
transform 1 0 47824 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2120_
timestamp 1698431365
transform -1 0 49728 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2121_
timestamp 1698431365
transform -1 0 51296 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2122_
timestamp 1698431365
transform 1 0 49728 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2123_
timestamp 1698431365
transform -1 0 49504 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2124_
timestamp 1698431365
transform 1 0 46256 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2125_
timestamp 1698431365
transform -1 0 49728 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2126_
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2127_
timestamp 1698431365
transform -1 0 48384 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2128_
timestamp 1698431365
transform 1 0 51744 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2129_
timestamp 1698431365
transform -1 0 53648 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2130_
timestamp 1698431365
transform 1 0 49168 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2131_
timestamp 1698431365
transform 1 0 49504 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2132_
timestamp 1698431365
transform 1 0 49504 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2133_
timestamp 1698431365
transform -1 0 48384 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2134_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47488 0 1 48608
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2135_
timestamp 1698431365
transform 1 0 50960 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2136_
timestamp 1698431365
transform -1 0 51520 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2137_
timestamp 1698431365
transform 1 0 51072 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2138_
timestamp 1698431365
transform -1 0 51072 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2139_
timestamp 1698431365
transform 1 0 51856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2140_
timestamp 1698431365
transform -1 0 52080 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2141_
timestamp 1698431365
transform 1 0 50736 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2142_
timestamp 1698431365
transform 1 0 51632 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2143_
timestamp 1698431365
transform 1 0 53424 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2144_
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2145_
timestamp 1698431365
transform -1 0 53648 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2146_
timestamp 1698431365
transform 1 0 51968 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2147_
timestamp 1698431365
transform 1 0 52080 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2148_
timestamp 1698431365
transform -1 0 53984 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2149_
timestamp 1698431365
transform -1 0 53200 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2150_
timestamp 1698431365
transform -1 0 51520 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2151_
timestamp 1698431365
transform -1 0 50176 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2152_
timestamp 1698431365
transform -1 0 57008 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2153_
timestamp 1698431365
transform 1 0 52416 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2154_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 55888 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2155_
timestamp 1698431365
transform 1 0 49056 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2156_
timestamp 1698431365
transform 1 0 49056 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2157_
timestamp 1698431365
transform -1 0 46592 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2158_
timestamp 1698431365
transform -1 0 52416 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2159_
timestamp 1698431365
transform -1 0 54656 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2160_
timestamp 1698431365
transform 1 0 54096 0 1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2161_
timestamp 1698431365
transform 1 0 54544 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2162_
timestamp 1698431365
transform -1 0 57792 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2163_
timestamp 1698431365
transform -1 0 53312 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2164_
timestamp 1698431365
transform -1 0 51520 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2165_
timestamp 1698431365
transform -1 0 50624 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2166_
timestamp 1698431365
transform 1 0 50624 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2167_
timestamp 1698431365
transform 1 0 53984 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2168_
timestamp 1698431365
transform -1 0 55776 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2169_
timestamp 1698431365
transform -1 0 54208 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2170_
timestamp 1698431365
transform 1 0 53312 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2171_
timestamp 1698431365
transform 1 0 55216 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2172_
timestamp 1698431365
transform 1 0 57008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2173_
timestamp 1698431365
transform 1 0 56112 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2174_
timestamp 1698431365
transform -1 0 53984 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2175_
timestamp 1698431365
transform 1 0 52640 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2176_
timestamp 1698431365
transform -1 0 54096 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2177_
timestamp 1698431365
transform 1 0 34496 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2178_
timestamp 1698431365
transform -1 0 53424 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2179_
timestamp 1698431365
transform 1 0 53424 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2180_
timestamp 1698431365
transform -1 0 56224 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _2181_
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2182_
timestamp 1698431365
transform -1 0 56224 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2183_
timestamp 1698431365
transform -1 0 52080 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2184_
timestamp 1698431365
transform 1 0 50176 0 -1 45472
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2185_
timestamp 1698431365
transform -1 0 50400 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2186_
timestamp 1698431365
transform 1 0 50400 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2187_
timestamp 1698431365
transform -1 0 49728 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2188_
timestamp 1698431365
transform 1 0 47488 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2189_
timestamp 1698431365
transform 1 0 47488 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2190_
timestamp 1698431365
transform -1 0 53760 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2191_
timestamp 1698431365
transform 1 0 50176 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2192_
timestamp 1698431365
transform -1 0 56224 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2193_
timestamp 1698431365
transform -1 0 52080 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2194_
timestamp 1698431365
transform 1 0 51296 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2195_
timestamp 1698431365
transform 1 0 53536 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2196_
timestamp 1698431365
transform 1 0 52080 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2197_
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2198_
timestamp 1698431365
transform -1 0 58016 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2199_
timestamp 1698431365
transform 1 0 51184 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2200_
timestamp 1698431365
transform 1 0 50624 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2201_
timestamp 1698431365
transform -1 0 53536 0 -1 40768
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2202_
timestamp 1698431365
transform -1 0 51184 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2203_
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2204_
timestamp 1698431365
transform -1 0 54544 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2205_
timestamp 1698431365
transform 1 0 52752 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2206_
timestamp 1698431365
transform 1 0 54208 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2207_
timestamp 1698431365
transform -1 0 56896 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2208_
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2209_
timestamp 1698431365
transform -1 0 57568 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2210_
timestamp 1698431365
transform 1 0 56672 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2211_
timestamp 1698431365
transform 1 0 55664 0 1 36064
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2212_
timestamp 1698431365
transform 1 0 50064 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2213_
timestamp 1698431365
transform 1 0 51632 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2214_
timestamp 1698431365
transform 1 0 55440 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2215_
timestamp 1698431365
transform 1 0 31024 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2216_
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2217_
timestamp 1698431365
transform -1 0 58240 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2218_
timestamp 1698431365
transform -1 0 57792 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2219_
timestamp 1698431365
transform -1 0 54544 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2220_
timestamp 1698431365
transform -1 0 55440 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2221_
timestamp 1698431365
transform -1 0 31136 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2222_
timestamp 1698431365
transform 1 0 53088 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2223_
timestamp 1698431365
transform -1 0 56224 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2224_
timestamp 1698431365
transform -1 0 51856 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2225_
timestamp 1698431365
transform -1 0 53424 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2226_
timestamp 1698431365
transform -1 0 53648 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2227_
timestamp 1698431365
transform -1 0 52304 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2228_
timestamp 1698431365
transform 1 0 50624 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2229_
timestamp 1698431365
transform 1 0 51856 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2230_
timestamp 1698431365
transform -1 0 55104 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2231_
timestamp 1698431365
transform -1 0 54096 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2232_
timestamp 1698431365
transform 1 0 48720 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2233_
timestamp 1698431365
transform -1 0 50064 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2234_
timestamp 1698431365
transform -1 0 48384 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2235_
timestamp 1698431365
transform -1 0 48608 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2236_
timestamp 1698431365
transform 1 0 47264 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2237_
timestamp 1698431365
transform 1 0 49504 0 -1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2238_
timestamp 1698431365
transform -1 0 49952 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2239_
timestamp 1698431365
transform -1 0 49616 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2240_
timestamp 1698431365
transform 1 0 49952 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2241_
timestamp 1698431365
transform -1 0 48384 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2242_
timestamp 1698431365
transform 1 0 47600 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2243_
timestamp 1698431365
transform -1 0 49840 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2244_
timestamp 1698431365
transform -1 0 51744 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2245_
timestamp 1698431365
transform 1 0 49840 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2246_
timestamp 1698431365
transform 1 0 50064 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2247_
timestamp 1698431365
transform 1 0 51408 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2248_
timestamp 1698431365
transform -1 0 50064 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2249_
timestamp 1698431365
transform 1 0 50064 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2250_
timestamp 1698431365
transform 1 0 51072 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2251_
timestamp 1698431365
transform -1 0 52976 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2252_
timestamp 1698431365
transform -1 0 51968 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2253_
timestamp 1698431365
transform 1 0 30576 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2254_
timestamp 1698431365
transform -1 0 31584 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2255_
timestamp 1698431365
transform -1 0 31360 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2256_
timestamp 1698431365
transform 1 0 19712 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2257_
timestamp 1698431365
transform 1 0 25536 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2258_
timestamp 1698431365
transform 1 0 25312 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2259_
timestamp 1698431365
transform -1 0 25872 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2260_
timestamp 1698431365
transform 1 0 23184 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2261_
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2262_
timestamp 1698431365
transform 1 0 25648 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2263_
timestamp 1698431365
transform 1 0 26656 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2264_
timestamp 1698431365
transform -1 0 19712 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2265_
timestamp 1698431365
transform 1 0 18816 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2266_
timestamp 1698431365
transform -1 0 30352 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2267_
timestamp 1698431365
transform 1 0 29456 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2268_
timestamp 1698431365
transform 1 0 29792 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2269_
timestamp 1698431365
transform -1 0 31024 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2270_
timestamp 1698431365
transform -1 0 28112 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2271_
timestamp 1698431365
transform 1 0 19264 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2272_
timestamp 1698431365
transform 1 0 22848 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2273_
timestamp 1698431365
transform -1 0 20944 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2274_
timestamp 1698431365
transform 1 0 14112 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2275_
timestamp 1698431365
transform 1 0 11648 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2276_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20832 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2277_
timestamp 1698431365
transform -1 0 19712 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2278_
timestamp 1698431365
transform -1 0 19264 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2279_
timestamp 1698431365
transform 1 0 18032 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2280_
timestamp 1698431365
transform 1 0 22064 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2281_
timestamp 1698431365
transform -1 0 28672 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2282_
timestamp 1698431365
transform -1 0 29456 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2283_
timestamp 1698431365
transform 1 0 26320 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2284_
timestamp 1698431365
transform 1 0 26208 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2285_
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2286_
timestamp 1698431365
transform 1 0 19936 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2287_
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2288_
timestamp 1698431365
transform 1 0 26096 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2289_
timestamp 1698431365
transform -1 0 28000 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2290_
timestamp 1698431365
transform -1 0 27888 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2291_
timestamp 1698431365
transform 1 0 23520 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2292_
timestamp 1698431365
transform 1 0 23744 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2293_
timestamp 1698431365
transform 1 0 19936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2294_
timestamp 1698431365
transform 1 0 25424 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2295_
timestamp 1698431365
transform 1 0 21392 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2296_
timestamp 1698431365
transform 1 0 27888 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2297_
timestamp 1698431365
transform 1 0 27328 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2298_
timestamp 1698431365
transform -1 0 28784 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2299_
timestamp 1698431365
transform -1 0 27104 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2300_
timestamp 1698431365
transform 1 0 19936 0 -1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2301_
timestamp 1698431365
transform 1 0 17808 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2302_
timestamp 1698431365
transform -1 0 19488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2303_
timestamp 1698431365
transform 1 0 13888 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2304_
timestamp 1698431365
transform 1 0 19600 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2305_
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2306_
timestamp 1698431365
transform 1 0 31360 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2307_
timestamp 1698431365
transform 1 0 25648 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2308_
timestamp 1698431365
transform -1 0 30464 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2309_
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2310_
timestamp 1698431365
transform -1 0 23968 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2311_
timestamp 1698431365
transform 1 0 24528 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2312_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28112 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2313_
timestamp 1698431365
transform -1 0 33824 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2314_
timestamp 1698431365
transform 1 0 34608 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2315_
timestamp 1698431365
transform 1 0 24080 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2316_
timestamp 1698431365
transform -1 0 28000 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2317_
timestamp 1698431365
transform -1 0 27216 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2318_
timestamp 1698431365
transform -1 0 25088 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2319_
timestamp 1698431365
transform -1 0 24752 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2320_
timestamp 1698431365
transform 1 0 23856 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2321_
timestamp 1698431365
transform -1 0 29456 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2322_
timestamp 1698431365
transform -1 0 26432 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2323_
timestamp 1698431365
transform -1 0 25536 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2324_
timestamp 1698431365
transform 1 0 10416 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2325_
timestamp 1698431365
transform 1 0 11088 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2326_
timestamp 1698431365
transform 1 0 12544 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2327_
timestamp 1698431365
transform -1 0 22736 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2328_
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2329_
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2330_
timestamp 1698431365
transform 1 0 26992 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2331_
timestamp 1698431365
transform -1 0 32704 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2332_
timestamp 1698431365
transform 1 0 32256 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2333_
timestamp 1698431365
transform -1 0 19936 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2334_
timestamp 1698431365
transform -1 0 22848 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2335_
timestamp 1698431365
transform 1 0 10528 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2336_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2337_
timestamp 1698431365
transform 1 0 22736 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2338_
timestamp 1698431365
transform 1 0 25648 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2339_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2340_
timestamp 1698431365
transform 1 0 19712 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2341_
timestamp 1698431365
transform 1 0 30464 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2342_
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2343_
timestamp 1698431365
transform -1 0 33824 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2344_
timestamp 1698431365
transform 1 0 26208 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2345_
timestamp 1698431365
transform 1 0 6496 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2346_
timestamp 1698431365
transform 1 0 20944 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2347_
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2348_
timestamp 1698431365
transform 1 0 21952 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2349_
timestamp 1698431365
transform -1 0 27104 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2350_
timestamp 1698431365
transform -1 0 23856 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2351_
timestamp 1698431365
transform -1 0 21728 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2352_
timestamp 1698431365
transform 1 0 21280 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2353_
timestamp 1698431365
transform -1 0 25872 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2354_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2355_
timestamp 1698431365
transform 1 0 25648 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2356_
timestamp 1698431365
transform 1 0 30912 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2357_
timestamp 1698431365
transform 1 0 34048 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2358_
timestamp 1698431365
transform 1 0 32480 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2359_
timestamp 1698431365
transform 1 0 23072 0 1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2360_
timestamp 1698431365
transform 1 0 21840 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2361_
timestamp 1698431365
transform 1 0 25088 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2362_
timestamp 1698431365
transform 1 0 23296 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2363_
timestamp 1698431365
transform -1 0 30240 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2364_
timestamp 1698431365
transform -1 0 32592 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2365_
timestamp 1698431365
transform -1 0 30688 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2366_
timestamp 1698431365
transform 1 0 22176 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2367_
timestamp 1698431365
transform -1 0 23856 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2368_
timestamp 1698431365
transform 1 0 30128 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2369_
timestamp 1698431365
transform 1 0 31136 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2370_
timestamp 1698431365
transform 1 0 31808 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2371_
timestamp 1698431365
transform -1 0 26544 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2372_
timestamp 1698431365
transform -1 0 31360 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2373_
timestamp 1698431365
transform -1 0 29904 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2374_
timestamp 1698431365
transform -1 0 30240 0 -1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2375_
timestamp 1698431365
transform 1 0 34720 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2376_
timestamp 1698431365
transform -1 0 32704 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2377_
timestamp 1698431365
transform -1 0 19712 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2378_
timestamp 1698431365
transform -1 0 27888 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2379_
timestamp 1698431365
transform 1 0 23408 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2380_
timestamp 1698431365
transform -1 0 27552 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2381_
timestamp 1698431365
transform 1 0 26544 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2382_
timestamp 1698431365
transform 1 0 30464 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2383_
timestamp 1698431365
transform 1 0 33488 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2384_
timestamp 1698431365
transform 1 0 32144 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2385_
timestamp 1698431365
transform -1 0 33376 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2386_
timestamp 1698431365
transform -1 0 26208 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2387_
timestamp 1698431365
transform -1 0 28112 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2388_
timestamp 1698431365
transform 1 0 28112 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2389_
timestamp 1698431365
transform 1 0 30800 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2390_
timestamp 1698431365
transform -1 0 27776 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2391_
timestamp 1698431365
transform 1 0 22512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2392_
timestamp 1698431365
transform -1 0 24752 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2393_
timestamp 1698431365
transform 1 0 28112 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2394_
timestamp 1698431365
transform 1 0 27664 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2395_
timestamp 1698431365
transform 1 0 29456 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2396_
timestamp 1698431365
transform -1 0 29120 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2397_
timestamp 1698431365
transform 1 0 9744 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2398_
timestamp 1698431365
transform -1 0 15680 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2399_
timestamp 1698431365
transform -1 0 20160 0 1 36064
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2400_
timestamp 1698431365
transform 1 0 14448 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2401_
timestamp 1698431365
transform -1 0 15232 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2402_
timestamp 1698431365
transform -1 0 9856 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2403_
timestamp 1698431365
transform -1 0 11312 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2404_
timestamp 1698431365
transform -1 0 8064 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2405_
timestamp 1698431365
transform 1 0 5824 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2406_
timestamp 1698431365
transform 1 0 6720 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2407_
timestamp 1698431365
transform 1 0 7840 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2408_
timestamp 1698431365
transform -1 0 8960 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2409_
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2410_
timestamp 1698431365
transform -1 0 10976 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2411_
timestamp 1698431365
transform 1 0 6608 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2412_
timestamp 1698431365
transform 1 0 7168 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2413_
timestamp 1698431365
transform -1 0 11648 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2414_
timestamp 1698431365
transform 1 0 10640 0 -1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2415_
timestamp 1698431365
transform -1 0 4928 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2416_
timestamp 1698431365
transform 1 0 4704 0 -1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2417_
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2418_
timestamp 1698431365
transform -1 0 8064 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2419_
timestamp 1698431365
transform 1 0 7616 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2420_
timestamp 1698431365
transform -1 0 9184 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2421_
timestamp 1698431365
transform -1 0 10416 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2422_
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2423_
timestamp 1698431365
transform -1 0 7616 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2424_
timestamp 1698431365
transform 1 0 15232 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2425_
timestamp 1698431365
transform -1 0 19712 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2426_
timestamp 1698431365
transform 1 0 15456 0 1 37632
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2427_
timestamp 1698431365
transform -1 0 10752 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2428_
timestamp 1698431365
transform -1 0 11984 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2429_
timestamp 1698431365
transform -1 0 10304 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2430_
timestamp 1698431365
transform -1 0 9184 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2431_
timestamp 1698431365
transform 1 0 6944 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2432_
timestamp 1698431365
transform 1 0 8064 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2433_
timestamp 1698431365
transform 1 0 7616 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2434_
timestamp 1698431365
transform 1 0 12544 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2435_
timestamp 1698431365
transform -1 0 14560 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2436_
timestamp 1698431365
transform 1 0 7168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2437_
timestamp 1698431365
transform -1 0 8400 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2438_
timestamp 1698431365
transform -1 0 5712 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2439_
timestamp 1698431365
transform 1 0 9632 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2440_
timestamp 1698431365
transform 1 0 10304 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2441_
timestamp 1698431365
transform -1 0 4928 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2442_
timestamp 1698431365
transform 1 0 4592 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2443_
timestamp 1698431365
transform 1 0 1904 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2444_
timestamp 1698431365
transform 1 0 3248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2445_
timestamp 1698431365
transform -1 0 3248 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2446_
timestamp 1698431365
transform 1 0 2016 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2447_
timestamp 1698431365
transform -1 0 3360 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2448_
timestamp 1698431365
transform 1 0 3696 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2449_
timestamp 1698431365
transform -1 0 13104 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2450_
timestamp 1698431365
transform -1 0 13328 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2451_
timestamp 1698431365
transform 1 0 2576 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2452_
timestamp 1698431365
transform -1 0 3696 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2453_
timestamp 1698431365
transform 1 0 3360 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2454_
timestamp 1698431365
transform 1 0 5936 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2455_
timestamp 1698431365
transform -1 0 7728 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2456_
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2457_
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2458_
timestamp 1698431365
transform -1 0 24864 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2459_
timestamp 1698431365
transform -1 0 14672 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2460_
timestamp 1698431365
transform 1 0 13328 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2461_
timestamp 1698431365
transform -1 0 12992 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2462_
timestamp 1698431365
transform 1 0 12544 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2463_
timestamp 1698431365
transform 1 0 14224 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2464_
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2465_
timestamp 1698431365
transform -1 0 12992 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2466_
timestamp 1698431365
transform -1 0 12544 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2467_
timestamp 1698431365
transform -1 0 11200 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2468_
timestamp 1698431365
transform -1 0 4032 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2469_
timestamp 1698431365
transform 1 0 2576 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2470_
timestamp 1698431365
transform -1 0 3920 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2471_
timestamp 1698431365
transform -1 0 2464 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2472_
timestamp 1698431365
transform -1 0 10304 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2473_
timestamp 1698431365
transform 1 0 6720 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2474_
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2475_
timestamp 1698431365
transform 1 0 5488 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2476_
timestamp 1698431365
transform -1 0 4256 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2477_
timestamp 1698431365
transform -1 0 2800 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2478_
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2479_
timestamp 1698431365
transform -1 0 5376 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2480_
timestamp 1698431365
transform 1 0 4816 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2481_
timestamp 1698431365
transform -1 0 6720 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2482_
timestamp 1698431365
transform -1 0 3696 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2483_
timestamp 1698431365
transform 1 0 5712 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2484_
timestamp 1698431365
transform 1 0 6832 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2485_
timestamp 1698431365
transform -1 0 7616 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2486_
timestamp 1698431365
transform -1 0 7168 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2487_
timestamp 1698431365
transform -1 0 5264 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2488_
timestamp 1698431365
transform 1 0 5488 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2489_
timestamp 1698431365
transform -1 0 6384 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2490_
timestamp 1698431365
transform -1 0 5264 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2491_
timestamp 1698431365
transform 1 0 6160 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2492_
timestamp 1698431365
transform -1 0 6160 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2493_
timestamp 1698431365
transform 1 0 8288 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2494_
timestamp 1698431365
transform 1 0 10528 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2495_
timestamp 1698431365
transform 1 0 10640 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2496_
timestamp 1698431365
transform 1 0 12432 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2497_
timestamp 1698431365
transform 1 0 10416 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2498_
timestamp 1698431365
transform -1 0 13104 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2499_
timestamp 1698431365
transform -1 0 12432 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2500_
timestamp 1698431365
transform 1 0 11984 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2501_
timestamp 1698431365
transform 1 0 10640 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2502_
timestamp 1698431365
transform 1 0 11088 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2503_
timestamp 1698431365
transform 1 0 9744 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2504_
timestamp 1698431365
transform -1 0 12432 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2505_
timestamp 1698431365
transform 1 0 12208 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2506_
timestamp 1698431365
transform -1 0 12208 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2507_
timestamp 1698431365
transform -1 0 9184 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2508_
timestamp 1698431365
transform 1 0 9632 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2509_
timestamp 1698431365
transform -1 0 10304 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2510_
timestamp 1698431365
transform 1 0 11536 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2511_
timestamp 1698431365
transform 1 0 11312 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2512_
timestamp 1698431365
transform -1 0 10976 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2513_
timestamp 1698431365
transform -1 0 11312 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2514_
timestamp 1698431365
transform -1 0 10304 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2515_
timestamp 1698431365
transform -1 0 18928 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2516_
timestamp 1698431365
transform -1 0 16912 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2517_
timestamp 1698431365
transform -1 0 18144 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2518_
timestamp 1698431365
transform 1 0 17808 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2519_
timestamp 1698431365
transform 1 0 18480 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2520_
timestamp 1698431365
transform 1 0 18032 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2521_
timestamp 1698431365
transform 1 0 15344 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2522_
timestamp 1698431365
transform -1 0 16352 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2523_
timestamp 1698431365
transform -1 0 15232 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2524_
timestamp 1698431365
transform 1 0 15008 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2525_
timestamp 1698431365
transform -1 0 15344 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2526_
timestamp 1698431365
transform -1 0 17024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2527_
timestamp 1698431365
transform -1 0 13104 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2528_
timestamp 1698431365
transform -1 0 11648 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2529_
timestamp 1698431365
transform -1 0 13664 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2530_
timestamp 1698431365
transform 1 0 11760 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2531_
timestamp 1698431365
transform -1 0 12656 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2532_
timestamp 1698431365
transform 1 0 14336 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2533_
timestamp 1698431365
transform -1 0 6720 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2534_
timestamp 1698431365
transform -1 0 6160 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2535_
timestamp 1698431365
transform -1 0 6160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2536_
timestamp 1698431365
transform -1 0 6160 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2537_
timestamp 1698431365
transform -1 0 6272 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2538_
timestamp 1698431365
transform -1 0 19152 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2539_
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2540_
timestamp 1698431365
transform 1 0 19488 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2541_
timestamp 1698431365
transform -1 0 21840 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2542_
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2543_
timestamp 1698431365
transform -1 0 19376 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2544_
timestamp 1698431365
transform -1 0 20832 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2545_
timestamp 1698431365
transform 1 0 14896 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2546_
timestamp 1698431365
transform 1 0 16128 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2547_
timestamp 1698431365
transform -1 0 19152 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2548_
timestamp 1698431365
transform 1 0 17472 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2549_
timestamp 1698431365
transform 1 0 17248 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2550_
timestamp 1698431365
transform -1 0 19712 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2551_
timestamp 1698431365
transform -1 0 22848 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2552_
timestamp 1698431365
transform 1 0 21952 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2553_
timestamp 1698431365
transform -1 0 23520 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2554_
timestamp 1698431365
transform -1 0 23184 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2555_
timestamp 1698431365
transform 1 0 19712 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2556_
timestamp 1698431365
transform 1 0 15792 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2557_
timestamp 1698431365
transform 1 0 18928 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2558_
timestamp 1698431365
transform -1 0 21616 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2559_
timestamp 1698431365
transform 1 0 21952 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2560_
timestamp 1698431365
transform -1 0 22848 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2561_
timestamp 1698431365
transform 1 0 20048 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2562_
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2563_
timestamp 1698431365
transform 1 0 14000 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2564_
timestamp 1698431365
transform 1 0 17696 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2565_
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2566_
timestamp 1698431365
transform 1 0 22176 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2567_
timestamp 1698431365
transform -1 0 21280 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2568_
timestamp 1698431365
transform 1 0 16576 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2569_
timestamp 1698431365
transform 1 0 18592 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2570_
timestamp 1698431365
transform 1 0 20832 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2571_
timestamp 1698431365
transform 1 0 22848 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2572_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2573_
timestamp 1698431365
transform -1 0 18928 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2574_
timestamp 1698431365
transform -1 0 19936 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2575_
timestamp 1698431365
transform -1 0 19600 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2576_
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2577_
timestamp 1698431365
transform -1 0 17920 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2578_
timestamp 1698431365
transform -1 0 22960 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2579_
timestamp 1698431365
transform 1 0 20832 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2580_
timestamp 1698431365
transform 1 0 20160 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2581_
timestamp 1698431365
transform -1 0 22960 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2582_
timestamp 1698431365
transform 1 0 23408 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2583_
timestamp 1698431365
transform 1 0 22400 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2584_
timestamp 1698431365
transform 1 0 22736 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2585_
timestamp 1698431365
transform -1 0 34944 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2586_
timestamp 1698431365
transform 1 0 32816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2587_
timestamp 1698431365
transform 1 0 35952 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2588_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2589_
timestamp 1698431365
transform 1 0 22288 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2590_
timestamp 1698431365
transform 1 0 25312 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2591_
timestamp 1698431365
transform -1 0 25312 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2592_
timestamp 1698431365
transform 1 0 27104 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2593_
timestamp 1698431365
transform -1 0 28112 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2594_
timestamp 1698431365
transform -1 0 17024 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2595_
timestamp 1698431365
transform 1 0 17248 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2596_
timestamp 1698431365
transform 1 0 26544 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2597_
timestamp 1698431365
transform 1 0 27776 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2598_
timestamp 1698431365
transform 1 0 27440 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2599_
timestamp 1698431365
transform 1 0 29232 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2600_
timestamp 1698431365
transform 1 0 29232 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2601_
timestamp 1698431365
transform -1 0 19824 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2602_
timestamp 1698431365
transform -1 0 18256 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2603_
timestamp 1698431365
transform 1 0 13664 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2604_
timestamp 1698431365
transform -1 0 12096 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2605_
timestamp 1698431365
transform 1 0 14896 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2606_
timestamp 1698431365
transform -1 0 14784 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2607_
timestamp 1698431365
transform -1 0 21728 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2608_
timestamp 1698431365
transform -1 0 19488 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2609_
timestamp 1698431365
transform -1 0 20832 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2610_
timestamp 1698431365
transform 1 0 19712 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2611_
timestamp 1698431365
transform -1 0 22848 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2612_
timestamp 1698431365
transform 1 0 17584 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2613_
timestamp 1698431365
transform -1 0 18144 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2614_
timestamp 1698431365
transform 1 0 22848 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2615_
timestamp 1698431365
transform 1 0 19376 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2616_
timestamp 1698431365
transform -1 0 19152 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2617_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2618_
timestamp 1698431365
transform -1 0 21840 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2619_
timestamp 1698431365
transform -1 0 17024 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2620_
timestamp 1698431365
transform -1 0 17024 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2621_
timestamp 1698431365
transform 1 0 14000 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2622_
timestamp 1698431365
transform -1 0 12656 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2623_
timestamp 1698431365
transform 1 0 17472 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2624_
timestamp 1698431365
transform -1 0 16016 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2625_
timestamp 1698431365
transform 1 0 21728 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2626_
timestamp 1698431365
transform -1 0 32928 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2627_
timestamp 1698431365
transform 1 0 24192 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2628_
timestamp 1698431365
transform 1 0 23968 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2629_
timestamp 1698431365
transform -1 0 35616 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2630_
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2631_
timestamp 1698431365
transform 1 0 21840 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2632_
timestamp 1698431365
transform 1 0 22960 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2633_
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2634_
timestamp 1698431365
transform 1 0 23520 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2635_
timestamp 1698431365
transform 1 0 24640 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2636_
timestamp 1698431365
transform -1 0 25984 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2637_
timestamp 1698431365
transform -1 0 22400 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2638_
timestamp 1698431365
transform 1 0 19488 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2639_
timestamp 1698431365
transform -1 0 18928 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2640_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2641_
timestamp 1698431365
transform -1 0 21840 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2642_
timestamp 1698431365
transform -1 0 20048 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2643_
timestamp 1698431365
transform 1 0 10976 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2644_
timestamp 1698431365
transform -1 0 10080 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2645_
timestamp 1698431365
transform 1 0 10528 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2646_
timestamp 1698431365
transform 1 0 7616 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2647_
timestamp 1698431365
transform -1 0 19488 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2648_
timestamp 1698431365
transform 1 0 19040 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2649_
timestamp 1698431365
transform 1 0 18032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2650_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2651_
timestamp 1698431365
transform -1 0 17024 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2652_
timestamp 1698431365
transform 1 0 34496 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2653_
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2654_
timestamp 1698431365
transform 1 0 35728 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2655_
timestamp 1698431365
transform 1 0 35168 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2656_
timestamp 1698431365
transform -1 0 37744 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2657_
timestamp 1698431365
transform -1 0 17248 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2658_
timestamp 1698431365
transform 1 0 10864 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2659_
timestamp 1698431365
transform -1 0 10080 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2660_
timestamp 1698431365
transform 1 0 10752 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2661_
timestamp 1698431365
transform -1 0 10752 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2662_
timestamp 1698431365
transform -1 0 36624 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2663_
timestamp 1698431365
transform -1 0 36288 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2664_
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2665_
timestamp 1698431365
transform -1 0 36288 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2666_
timestamp 1698431365
transform -1 0 36960 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2667_
timestamp 1698431365
transform 1 0 33264 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2668_
timestamp 1698431365
transform 1 0 33600 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2669_
timestamp 1698431365
transform 1 0 33376 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2670_
timestamp 1698431365
transform 1 0 34496 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2671_
timestamp 1698431365
transform 1 0 34720 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2672_
timestamp 1698431365
transform 1 0 21392 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2673_
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2674_
timestamp 1698431365
transform -1 0 28224 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2675_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2676_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2677_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41216 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2678_
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2679_
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2680_
timestamp 1698431365
transform 1 0 44016 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2681_
timestamp 1698431365
transform 1 0 12208 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2682_
timestamp 1698431365
transform 1 0 12544 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2683_
timestamp 1698431365
transform -1 0 40768 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2684_
timestamp 1698431365
transform -1 0 40992 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2685_
timestamp 1698431365
transform -1 0 42560 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2686_
timestamp 1698431365
transform -1 0 41328 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2687_
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2688_
timestamp 1698431365
transform 1 0 39648 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2689_
timestamp 1698431365
transform -1 0 40096 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2690_
timestamp 1698431365
transform -1 0 36848 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2691_
timestamp 1698431365
transform 1 0 30800 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2692_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2693_
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2694_
timestamp 1698431365
transform 1 0 29456 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2695_
timestamp 1698431365
transform 1 0 29456 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2696_
timestamp 1698431365
transform 1 0 39424 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2697_
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2698_
timestamp 1698431365
transform 1 0 4816 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2699_
timestamp 1698431365
transform 1 0 8064 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2700_
timestamp 1698431365
transform 1 0 7616 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2701_
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2702_
timestamp 1698431365
transform 1 0 14896 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2703_
timestamp 1698431365
transform -1 0 23744 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2704_
timestamp 1698431365
transform 1 0 5936 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2705_
timestamp 1698431365
transform 1 0 15008 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2706_
timestamp 1698431365
transform 1 0 29008 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2707_
timestamp 1698431365
transform 1 0 30576 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2708_
timestamp 1698431365
transform 1 0 24192 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2709_
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2710_
timestamp 1698431365
transform 1 0 10192 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2711_
timestamp 1698431365
transform 1 0 11984 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2712_
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2713_
timestamp 1698431365
transform 1 0 5824 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2714_
timestamp 1698431365
transform 1 0 5488 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2715_
timestamp 1698431365
transform 1 0 5824 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2716_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2717_
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2718_
timestamp 1698431365
transform 1 0 25536 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2719_
timestamp 1698431365
transform -1 0 32032 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2720_
timestamp 1698431365
transform 1 0 31248 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2721_
timestamp 1698431365
transform 1 0 31696 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2722_
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2723_
timestamp 1698431365
transform 1 0 33376 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2724_
timestamp 1698431365
transform 1 0 35504 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2725_
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2726_
timestamp 1698431365
transform 1 0 13888 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2727_
timestamp 1698431365
transform -1 0 24640 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2728_
timestamp 1698431365
transform 1 0 21616 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2729_
timestamp 1698431365
transform 1 0 16352 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2730_
timestamp 1698431365
transform 1 0 19040 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2731_
timestamp 1698431365
transform 1 0 14112 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2732_
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2733_
timestamp 1698431365
transform 1 0 18928 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2734_
timestamp 1698431365
transform 1 0 12992 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2735_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2736_
timestamp 1698431365
transform -1 0 42560 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2737_
timestamp 1698431365
transform -1 0 44352 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2738_
timestamp 1698431365
transform -1 0 44464 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2739_
timestamp 1698431365
transform -1 0 47824 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2740_
timestamp 1698431365
transform -1 0 45584 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2741_
timestamp 1698431365
transform -1 0 43680 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2742_
timestamp 1698431365
transform -1 0 37520 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2743_
timestamp 1698431365
transform 1 0 31584 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2744_
timestamp 1698431365
transform 1 0 29456 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2745_
timestamp 1698431365
transform 1 0 31696 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2746_
timestamp 1698431365
transform 1 0 33264 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2747_
timestamp 1698431365
transform 1 0 38640 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2748_
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2749_
timestamp 1698431365
transform -1 0 47264 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2750_
timestamp 1698431365
transform -1 0 47936 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2751_
timestamp 1698431365
transform 1 0 47936 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2752_
timestamp 1698431365
transform -1 0 53984 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2753_
timestamp 1698431365
transform 1 0 53648 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2754_
timestamp 1698431365
transform 1 0 54544 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2755_
timestamp 1698431365
transform 1 0 54768 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2756_
timestamp 1698431365
transform 1 0 54768 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2757_
timestamp 1698431365
transform -1 0 49280 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2758_
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2759_
timestamp 1698431365
transform 1 0 54880 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2760_
timestamp 1698431365
transform 1 0 53760 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2761_
timestamp 1698431365
transform 1 0 54208 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2762_
timestamp 1698431365
transform 1 0 52976 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2763_
timestamp 1698431365
transform 1 0 46928 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2764_
timestamp 1698431365
transform 1 0 45584 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2765_
timestamp 1698431365
transform 1 0 49056 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2766_
timestamp 1698431365
transform -1 0 55216 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2767_
timestamp 1698431365
transform -1 0 32256 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2768_
timestamp 1698431365
transform -1 0 28560 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2769_
timestamp 1698431365
transform -1 0 28336 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2770_
timestamp 1698431365
transform 1 0 22624 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2771_
timestamp 1698431365
transform 1 0 17808 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2772_
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2773_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2774_
timestamp 1698431365
transform 1 0 25760 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2775_
timestamp 1698431365
transform -1 0 25536 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2776_
timestamp 1698431365
transform -1 0 28784 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2777_
timestamp 1698431365
transform 1 0 32480 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2778_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2779_
timestamp 1698431365
transform 1 0 32928 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2780_
timestamp 1698431365
transform 1 0 33376 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2781_
timestamp 1698431365
transform 1 0 29232 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2782_
timestamp 1698431365
transform 1 0 34272 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2783_
timestamp 1698431365
transform 1 0 31472 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2784_
timestamp 1698431365
transform 1 0 31696 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2785_
timestamp 1698431365
transform 1 0 30688 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2786_
timestamp 1698431365
transform 1 0 26208 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2787_
timestamp 1698431365
transform 1 0 6496 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2788_
timestamp 1698431365
transform 1 0 5936 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2789_
timestamp 1698431365
transform -1 0 9072 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2790_
timestamp 1698431365
transform 1 0 3024 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2791_
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2792_
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2793_
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2794_
timestamp 1698431365
transform 1 0 3920 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2795_
timestamp 1698431365
transform 1 0 11984 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2796_
timestamp 1698431365
transform 1 0 10976 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2797_
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2798_
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2799_
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2800_
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2801_
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2802_
timestamp 1698431365
transform 1 0 2016 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2803_
timestamp 1698431365
transform -1 0 9072 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2804_
timestamp 1698431365
transform 1 0 2016 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2805_
timestamp 1698431365
transform 1 0 4144 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2806_
timestamp 1698431365
transform -1 0 14336 0 -1 45472
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2807_
timestamp 1698431365
transform -1 0 15008 0 -1 47040
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2808_
timestamp 1698431365
transform 1 0 8288 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2809_
timestamp 1698431365
transform -1 0 14560 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2810_
timestamp 1698431365
transform 1 0 6832 0 1 47040
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2811_
timestamp 1698431365
transform -1 0 13104 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2812_
timestamp 1698431365
transform 1 0 8624 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2813_
timestamp 1698431365
transform 1 0 17696 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2814_
timestamp 1698431365
transform 1 0 9856 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2815_
timestamp 1698431365
transform -1 0 16128 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2816_
timestamp 1698431365
transform 1 0 7168 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2817_
timestamp 1698431365
transform 1 0 7728 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2818_
timestamp 1698431365
transform -1 0 14448 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2819_
timestamp 1698431365
transform 1 0 3024 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2820_
timestamp 1698431365
transform 1 0 3248 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2821_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2822_
timestamp 1698431365
transform 1 0 4704 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2823_
timestamp 1698431365
transform 1 0 16464 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2824_
timestamp 1698431365
transform 1 0 21056 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2825_
timestamp 1698431365
transform -1 0 24864 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2826_
timestamp 1698431365
transform 1 0 23408 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2827_
timestamp 1698431365
transform 1 0 17584 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2828_
timestamp 1698431365
transform 1 0 13776 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2829_
timestamp 1698431365
transform 1 0 20160 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2830_
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2831_
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2832_
timestamp 1698431365
transform 1 0 36176 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2833_
timestamp 1698431365
transform 1 0 23744 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2834_
timestamp 1698431365
transform 1 0 26208 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2835_
timestamp 1698431365
transform 1 0 25536 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2836_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2837_
timestamp 1698431365
transform 1 0 10416 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2838_
timestamp 1698431365
transform 1 0 13104 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2839_
timestamp 1698431365
transform 1 0 19264 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2840_
timestamp 1698431365
transform 1 0 16464 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2841_
timestamp 1698431365
transform 1 0 17136 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2842_
timestamp 1698431365
transform 1 0 19712 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2843_
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2844_
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2845_
timestamp 1698431365
transform 1 0 22288 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2846_
timestamp 1698431365
transform 1 0 20160 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2847_
timestamp 1698431365
transform -1 0 24864 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2848_
timestamp 1698431365
transform 1 0 23856 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2849_
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2850_
timestamp 1698431365
transform 1 0 19824 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2851_
timestamp 1698431365
transform 1 0 8288 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2852_
timestamp 1698431365
transform 1 0 7728 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2853_
timestamp 1698431365
transform 1 0 18704 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2854_
timestamp 1698431365
transform 1 0 15232 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2855_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2856_
timestamp 1698431365
transform 1 0 35616 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2857_
timestamp 1698431365
transform 1 0 8288 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2858_
timestamp 1698431365
transform 1 0 8064 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2859_
timestamp 1698431365
transform 1 0 35616 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2860_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2861_
timestamp 1698431365
transform 1 0 32928 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2862_
timestamp 1698431365
transform 1 0 34384 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2863_
timestamp 1698431365
transform 1 0 25536 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2864_
timestamp 1698431365
transform 1 0 27552 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__A2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__I
timestamp 1698431365
transform -1 0 25424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__I
timestamp 1698431365
transform -1 0 24304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1352__I
timestamp 1698431365
transform 1 0 30688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__I
timestamp 1698431365
transform -1 0 25984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__I
timestamp 1698431365
transform 1 0 30240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1374__I
timestamp 1698431365
transform -1 0 27328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1377__I
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__I
timestamp 1698431365
transform 1 0 30576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__I
timestamp 1698431365
transform -1 0 25984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1397__I
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A1
timestamp 1698431365
transform -1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1498__I
timestamp 1698431365
transform 1 0 14784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__B
timestamp 1698431365
transform 1 0 17472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__I
timestamp 1698431365
transform -1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__I
timestamp 1698431365
transform 1 0 18480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__B
timestamp 1698431365
transform -1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__A4
timestamp 1698431365
transform 1 0 19264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__I
timestamp 1698431365
transform 1 0 20496 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__A1
timestamp 1698431365
transform 1 0 24416 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__A1
timestamp 1698431365
transform 1 0 8624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__B
timestamp 1698431365
transform 1 0 14784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__I
timestamp 1698431365
transform -1 0 14448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__B
timestamp 1698431365
transform 1 0 14896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__I
timestamp 1698431365
transform -1 0 15568 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__I
timestamp 1698431365
transform 1 0 34384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A2
timestamp 1698431365
transform 1 0 19488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A1
timestamp 1698431365
transform 1 0 16464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A2
timestamp 1698431365
transform 1 0 18592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__B
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__B
timestamp 1698431365
transform 1 0 13776 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A2
timestamp 1698431365
transform 1 0 11760 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A1
timestamp 1698431365
transform 1 0 15568 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__I
timestamp 1698431365
transform 1 0 37968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__I
timestamp 1698431365
transform -1 0 18704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A1
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A2
timestamp 1698431365
transform 1 0 37632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__I
timestamp 1698431365
transform 1 0 38416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__A1
timestamp 1698431365
transform 1 0 39648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__A2
timestamp 1698431365
transform 1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__A1
timestamp 1698431365
transform 1 0 20272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__I
timestamp 1698431365
transform -1 0 18928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__A1
timestamp 1698431365
transform 1 0 38192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__A2
timestamp 1698431365
transform 1 0 37296 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__A1
timestamp 1698431365
transform 1 0 37408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__A2
timestamp 1698431365
transform -1 0 38080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1744__A1
timestamp 1698431365
transform 1 0 38304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__I
timestamp 1698431365
transform 1 0 33376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__I
timestamp 1698431365
transform 1 0 34496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__A1
timestamp 1698431365
transform 1 0 36960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__A2
timestamp 1698431365
transform 1 0 35728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__I
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__A3
timestamp 1698431365
transform -1 0 22288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__I1
timestamp 1698431365
transform 1 0 35280 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__I
timestamp 1698431365
transform 1 0 35840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__I1
timestamp 1698431365
transform -1 0 33712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A1
timestamp 1698431365
transform -1 0 33488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A2
timestamp 1698431365
transform -1 0 34272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A2
timestamp 1698431365
transform 1 0 38976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A1
timestamp 1698431365
transform -1 0 33824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A2
timestamp 1698431365
transform 1 0 34272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__A1
timestamp 1698431365
transform 1 0 26096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__A2
timestamp 1698431365
transform 1 0 25872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__I
timestamp 1698431365
transform 1 0 23184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__A1
timestamp 1698431365
transform -1 0 17136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__I
timestamp 1698431365
transform 1 0 23184 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__C
timestamp 1698431365
transform 1 0 16016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__I
timestamp 1698431365
transform 1 0 17024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__A1
timestamp 1698431365
transform -1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__A2
timestamp 1698431365
transform -1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A1
timestamp 1698431365
transform 1 0 15568 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__A1
timestamp 1698431365
transform -1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__I
timestamp 1698431365
transform 1 0 35504 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__B
timestamp 1698431365
transform -1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A1
timestamp 1698431365
transform 1 0 40880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__A1
timestamp 1698431365
transform 1 0 41440 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__I
timestamp 1698431365
transform -1 0 45360 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__C
timestamp 1698431365
transform -1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__I
timestamp 1698431365
transform 1 0 48384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A2
timestamp 1698431365
transform -1 0 45472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__B
timestamp 1698431365
transform 1 0 43904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A1
timestamp 1698431365
transform 1 0 44128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__B
timestamp 1698431365
transform 1 0 43792 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__C
timestamp 1698431365
transform 1 0 40992 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2009__B
timestamp 1698431365
transform 1 0 40992 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__A2
timestamp 1698431365
transform 1 0 41888 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__C
timestamp 1698431365
transform -1 0 39312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A2
timestamp 1698431365
transform 1 0 36064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__A1
timestamp 1698431365
transform 1 0 41440 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__B
timestamp 1698431365
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__A2
timestamp 1698431365
transform 1 0 37968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__B
timestamp 1698431365
transform 1 0 36848 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A1
timestamp 1698431365
transform 1 0 39088 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__I
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__B
timestamp 1698431365
transform 1 0 39424 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__A2
timestamp 1698431365
transform 1 0 39984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2054__A1
timestamp 1698431365
transform 1 0 31024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2060__B
timestamp 1698431365
transform 1 0 40432 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__C
timestamp 1698431365
transform -1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__B
timestamp 1698431365
transform -1 0 39648 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__A2
timestamp 1698431365
transform -1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__C
timestamp 1698431365
transform -1 0 39312 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__C
timestamp 1698431365
transform -1 0 43344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2094__I
timestamp 1698431365
transform -1 0 42784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__A2
timestamp 1698431365
transform -1 0 43568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__B
timestamp 1698431365
transform -1 0 44016 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2103__B
timestamp 1698431365
transform 1 0 49280 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2105__C
timestamp 1698431365
transform 1 0 43792 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__B
timestamp 1698431365
transform 1 0 48832 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A2
timestamp 1698431365
transform -1 0 48048 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__C
timestamp 1698431365
transform -1 0 44016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__C
timestamp 1698431365
transform -1 0 51744 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__A2
timestamp 1698431365
transform 1 0 47040 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__B
timestamp 1698431365
transform 1 0 47488 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2136__A1
timestamp 1698431365
transform 1 0 51744 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A2
timestamp 1698431365
transform -1 0 51632 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__B
timestamp 1698431365
transform 1 0 52752 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2143__B
timestamp 1698431365
transform 1 0 54544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__A2
timestamp 1698431365
transform 1 0 50512 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__C
timestamp 1698431365
transform 1 0 51632 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__A2
timestamp 1698431365
transform 1 0 46368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__B
timestamp 1698431365
transform 1 0 44240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2158__A1
timestamp 1698431365
transform 1 0 51744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2169__B
timestamp 1698431365
transform 1 0 55328 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__A2
timestamp 1698431365
transform 1 0 54880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__C
timestamp 1698431365
transform 1 0 54208 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2176__C
timestamp 1698431365
transform 1 0 54320 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2177__I
timestamp 1698431365
transform 1 0 34272 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2178__A2
timestamp 1698431365
transform -1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2178__B
timestamp 1698431365
transform -1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2187__C
timestamp 1698431365
transform 1 0 48384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__A2
timestamp 1698431365
transform 1 0 47264 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__B
timestamp 1698431365
transform 1 0 46592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A1
timestamp 1698431365
transform 1 0 51408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__A1
timestamp 1698431365
transform 1 0 54096 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__A2
timestamp 1698431365
transform 1 0 53648 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__C
timestamp 1698431365
transform 1 0 54880 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__C
timestamp 1698431365
transform 1 0 50400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2204__A2
timestamp 1698431365
transform 1 0 53984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2205__A1
timestamp 1698431365
transform -1 0 50512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__A1
timestamp 1698431365
transform 1 0 55440 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__A2
timestamp 1698431365
transform 1 0 54096 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__C
timestamp 1698431365
transform 1 0 49840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2219__B
timestamp 1698431365
transform 1 0 54544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2222__A2
timestamp 1698431365
transform -1 0 51856 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2222__C
timestamp 1698431365
transform 1 0 52080 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2229__A1
timestamp 1698431365
transform 1 0 50960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2230__A2
timestamp 1698431365
transform 1 0 54880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2230__B
timestamp 1698431365
transform -1 0 54656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2234__A2
timestamp 1698431365
transform -1 0 47264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2234__B
timestamp 1698431365
transform -1 0 47488 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A1
timestamp 1698431365
transform 1 0 48832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2242__A1
timestamp 1698431365
transform 1 0 47376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__A2
timestamp 1698431365
transform 1 0 48832 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__C
timestamp 1698431365
transform 1 0 48160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__B
timestamp 1698431365
transform -1 0 49504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__A2
timestamp 1698431365
transform 1 0 51968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__C
timestamp 1698431365
transform 1 0 49728 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2252__A1
timestamp 1698431365
transform 1 0 52752 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2252__C
timestamp 1698431365
transform 1 0 50736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__I
timestamp 1698431365
transform -1 0 30576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2254__B
timestamp 1698431365
transform 1 0 32032 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2254__C
timestamp 1698431365
transform 1 0 31584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__A1
timestamp 1698431365
transform 1 0 26208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__A1
timestamp 1698431365
transform 1 0 26656 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__A2
timestamp 1698431365
transform 1 0 25088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__A1
timestamp 1698431365
transform 1 0 22064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2262__I
timestamp 1698431365
transform 1 0 25088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2264__B
timestamp 1698431365
transform -1 0 16464 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A1
timestamp 1698431365
transform -1 0 20160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A2
timestamp 1698431365
transform 1 0 18592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2266__A1
timestamp 1698431365
transform -1 0 29680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2267__I
timestamp 1698431365
transform 1 0 28336 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2322__A2
timestamp 1698431365
transform -1 0 25536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2343__B
timestamp 1698431365
transform 1 0 34160 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2357__B
timestamp 1698431365
transform -1 0 35392 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2359__A2
timestamp 1698431365
transform -1 0 27776 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A1
timestamp 1698431365
transform 1 0 21616 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2365__B
timestamp 1698431365
transform 1 0 30576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2366__A1
timestamp 1698431365
transform 1 0 21168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2375__B
timestamp 1698431365
transform 1 0 35952 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__A1
timestamp 1698431365
transform 1 0 27776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2383__B
timestamp 1698431365
transform 1 0 34608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2389__C
timestamp 1698431365
transform 1 0 33600 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__I
timestamp 1698431365
transform 1 0 27776 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2408__A1
timestamp 1698431365
transform -1 0 10304 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2413__A1
timestamp 1698431365
transform 1 0 12768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2420__C
timestamp 1698431365
transform 1 0 9184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2421__A1
timestamp 1698431365
transform -1 0 9856 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2433__C
timestamp 1698431365
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__B
timestamp 1698431365
transform 1 0 14784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2440__A1
timestamp 1698431365
transform 1 0 11536 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A1
timestamp 1698431365
transform -1 0 4592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2450__B
timestamp 1698431365
transform 1 0 11872 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__B
timestamp 1698431365
transform 1 0 15904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2515__I
timestamp 1698431365
transform -1 0 19376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2517__B
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__C
timestamp 1698431365
transform 1 0 19824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2521__B
timestamp 1698431365
transform 1 0 17472 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__C
timestamp 1698431365
transform 1 0 15120 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__I
timestamp 1698431365
transform 1 0 6944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__A2
timestamp 1698431365
transform 1 0 6496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__B2
timestamp 1698431365
transform 1 0 21952 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__C
timestamp 1698431365
transform 1 0 17024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__A1
timestamp 1698431365
transform 1 0 19712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__A2
timestamp 1698431365
transform -1 0 19152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__A1
timestamp 1698431365
transform 1 0 21952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__A2
timestamp 1698431365
transform 1 0 23632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__A2
timestamp 1698431365
transform 1 0 22512 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A2
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__I1
timestamp 1698431365
transform 1 0 26992 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__I1
timestamp 1698431365
transform 1 0 28784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__A1
timestamp 1698431365
transform 1 0 26096 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__A2
timestamp 1698431365
transform 1 0 26320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__A1
timestamp 1698431365
transform 1 0 28560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2599__A1
timestamp 1698431365
transform 1 0 30016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__I
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__A2
timestamp 1698431365
transform 1 0 20160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__I
timestamp 1698431365
transform 1 0 23072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__A1
timestamp 1698431365
transform 1 0 22736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2620__A1
timestamp 1698431365
transform 1 0 19152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__I
timestamp 1698431365
transform 1 0 35392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__A2
timestamp 1698431365
transform -1 0 22960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__A2
timestamp 1698431365
transform 1 0 20944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__A2
timestamp 1698431365
transform 1 0 18704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__A2
timestamp 1698431365
transform -1 0 34496 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__A1
timestamp 1698431365
transform 1 0 37632 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2667__A1
timestamp 1698431365
transform 1 0 32368 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2667__A2
timestamp 1698431365
transform 1 0 32816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__I1
timestamp 1698431365
transform 1 0 33376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2670__I1
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2677__CLK
timestamp 1698431365
transform 1 0 44912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__CLK
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2679__CLK
timestamp 1698431365
transform 1 0 45248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__CLK
timestamp 1698431365
transform 1 0 43792 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__CLK
timestamp 1698431365
transform 1 0 11984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__CLK
timestamp 1698431365
transform 1 0 16016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__CLK
timestamp 1698431365
transform 1 0 40992 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__CLK
timestamp 1698431365
transform 1 0 42784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2686__CLK
timestamp 1698431365
transform 1 0 41552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2687__CLK
timestamp 1698431365
transform 1 0 44240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__CLK
timestamp 1698431365
transform 1 0 43120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__CLK
timestamp 1698431365
transform 1 0 40320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__CLK
timestamp 1698431365
transform 1 0 37744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__CLK
timestamp 1698431365
transform 1 0 34272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__CLK
timestamp 1698431365
transform 1 0 21952 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__CLK
timestamp 1698431365
transform 1 0 31920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__CLK
timestamp 1698431365
transform 1 0 33712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__CLK
timestamp 1698431365
transform 1 0 43344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__CLK
timestamp 1698431365
transform 1 0 44240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__CLK
timestamp 1698431365
transform -1 0 11312 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__CLK
timestamp 1698431365
transform 1 0 10864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__CLK
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__CLK
timestamp 1698431365
transform 1 0 14224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__CLK
timestamp 1698431365
transform -1 0 24192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__CLK
timestamp 1698431365
transform -1 0 9856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__CLK
timestamp 1698431365
transform -1 0 18704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__CLK
timestamp 1698431365
transform 1 0 34048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__CLK
timestamp 1698431365
transform 1 0 23968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2709__CLK
timestamp 1698431365
transform 1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__CLK
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__CLK
timestamp 1698431365
transform 1 0 15456 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__CLK
timestamp 1698431365
transform 1 0 24640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2714__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2715__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2716__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__CLK
timestamp 1698431365
transform 1 0 22624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2718__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__CLK
timestamp 1698431365
transform -1 0 21392 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2728__CLK
timestamp 1698431365
transform 1 0 20720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2729__CLK
timestamp 1698431365
transform 1 0 19824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2730__CLK
timestamp 1698431365
transform 1 0 22512 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__CLK
timestamp 1698431365
transform 1 0 18144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__CLK
timestamp 1698431365
transform 1 0 15792 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__CLK
timestamp 1698431365
transform 1 0 22400 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__CLK
timestamp 1698431365
transform 1 0 15904 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__CLK
timestamp 1698431365
transform 1 0 42784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__CLK
timestamp 1698431365
transform 1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2738__CLK
timestamp 1698431365
transform 1 0 44912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2739__CLK
timestamp 1698431365
transform 1 0 48048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2740__CLK
timestamp 1698431365
transform 1 0 46704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__CLK
timestamp 1698431365
transform 1 0 43680 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2742__CLK
timestamp 1698431365
transform 1 0 37520 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__CLK
timestamp 1698431365
transform 1 0 35616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2744__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__CLK
timestamp 1698431365
transform 1 0 35168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2746__CLK
timestamp 1698431365
transform 1 0 35504 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2756__CLK
timestamp 1698431365
transform 1 0 54544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2757__CLK
timestamp 1698431365
transform 1 0 49504 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2758__CLK
timestamp 1698431365
transform 1 0 54432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2759__CLK
timestamp 1698431365
transform 1 0 55888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__CLK
timestamp 1698431365
transform 1 0 54992 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2761__CLK
timestamp 1698431365
transform 1 0 53984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2762__CLK
timestamp 1698431365
transform 1 0 52752 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2763__CLK
timestamp 1698431365
transform 1 0 50400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2764__CLK
timestamp 1698431365
transform 1 0 45360 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2765__CLK
timestamp 1698431365
transform 1 0 48832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2766__CLK
timestamp 1698431365
transform 1 0 52192 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2767__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2768__CLK
timestamp 1698431365
transform 1 0 29232 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2769__CLK
timestamp 1698431365
transform 1 0 28560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2770__CLK
timestamp 1698431365
transform 1 0 22400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2771__CLK
timestamp 1698431365
transform 1 0 21392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2772__CLK
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2773__CLK
timestamp 1698431365
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2774__CLK
timestamp 1698431365
transform 1 0 25536 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2775__CLK
timestamp 1698431365
transform 1 0 22064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2776__CLK
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2777__CLK
timestamp 1698431365
transform 1 0 35952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2778__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2779__CLK
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2780__CLK
timestamp 1698431365
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2781__CLK
timestamp 1698431365
transform 1 0 34608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2782__CLK
timestamp 1698431365
transform 1 0 37520 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2783__CLK
timestamp 1698431365
transform 1 0 35504 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2784__CLK
timestamp 1698431365
transform 1 0 35840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2785__CLK
timestamp 1698431365
transform 1 0 34608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2786__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2787__CLK
timestamp 1698431365
transform 1 0 9968 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2788__CLK
timestamp 1698431365
transform 1 0 9184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2789__CLK
timestamp 1698431365
transform 1 0 9296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2790__CLK
timestamp 1698431365
transform 1 0 6496 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2791__CLK
timestamp 1698431365
transform 1 0 4816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2792__CLK
timestamp 1698431365
transform 1 0 4816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2793__CLK
timestamp 1698431365
transform 1 0 5040 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2794__CLK
timestamp 1698431365
transform 1 0 8064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2795__CLK
timestamp 1698431365
transform 1 0 11760 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2796__CLK
timestamp 1698431365
transform 1 0 10752 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2806__CLK
timestamp 1698431365
transform 1 0 14560 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2807__CLK
timestamp 1698431365
transform 1 0 15232 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2809__CLK
timestamp 1698431365
transform 1 0 14784 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2811__CLK
timestamp 1698431365
transform 1 0 13104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2813__CLK
timestamp 1698431365
transform 1 0 20944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2814__CLK
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2815__CLK
timestamp 1698431365
transform 1 0 16128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2816__CLK
timestamp 1698431365
transform 1 0 10640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2817__CLK
timestamp 1698431365
transform 1 0 10976 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2818__CLK
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2819__CLK
timestamp 1698431365
transform 1 0 6496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2820__CLK
timestamp 1698431365
transform 1 0 6720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2821__CLK
timestamp 1698431365
transform 1 0 8960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2822__CLK
timestamp 1698431365
transform 1 0 8176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2823__CLK
timestamp 1698431365
transform 1 0 19712 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2824__CLK
timestamp 1698431365
transform 1 0 21840 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2825__CLK
timestamp 1698431365
transform 1 0 21392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2826__CLK
timestamp 1698431365
transform 1 0 23184 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2827__CLK
timestamp 1698431365
transform -1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2828__CLK
timestamp 1698431365
transform -1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2829__CLK
timestamp 1698431365
transform 1 0 24304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2830__CLK
timestamp 1698431365
transform -1 0 22960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2831__CLK
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2832__CLK
timestamp 1698431365
transform 1 0 39648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2833__CLK
timestamp 1698431365
transform 1 0 23520 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2834__CLK
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2835__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2836__CLK
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2837__CLK
timestamp 1698431365
transform 1 0 13664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2838__CLK
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2839__CLK
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2840__CLK
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2841__CLK
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2842__CLK
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2843__CLK
timestamp 1698431365
transform 1 0 14000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2844__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2845__CLK
timestamp 1698431365
transform 1 0 21504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2846__CLK
timestamp 1698431365
transform 1 0 23968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2847__CLK
timestamp 1698431365
transform 1 0 25536 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2848__CLK
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2849__CLK
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2850__CLK
timestamp 1698431365
transform 1 0 23296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2851__CLK
timestamp 1698431365
transform 1 0 12432 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2852__CLK
timestamp 1698431365
transform 1 0 10528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2853__CLK
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2854__CLK
timestamp 1698431365
transform 1 0 15680 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2855__CLK
timestamp 1698431365
transform 1 0 36848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__CLK
timestamp 1698431365
transform -1 0 35168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2857__CLK
timestamp 1698431365
transform 1 0 11760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2858__CLK
timestamp 1698431365
transform 1 0 11536 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2859__CLK
timestamp 1698431365
transform 1 0 37184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2860__CLK
timestamp 1698431365
transform -1 0 41328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2861__CLK
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2862__CLK
timestamp 1698431365
transform 1 0 37856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2863__CLK
timestamp 1698431365
transform 1 0 25312 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2864__CLK
timestamp 1698431365
transform 1 0 27328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 16688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 24304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 24416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 9632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 8064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 22960 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 32928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 38752 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 39648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 35616 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 35840 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 44352 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 45920 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 18928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 20608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 41216 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 41664 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 15568 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 14784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 4704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_wb_clk_i asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16240 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1698431365
transform -1 0 13328 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1698431365
transform -1 0 24080 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1698431365
transform -1 0 24080 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1698431365
transform 1 0 6272 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1698431365
transform -1 0 8960 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1698431365
transform 1 0 33152 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1698431365
transform 1 0 33488 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1698431365
transform 1 0 40320 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1698431365
transform 1 0 40992 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1698431365
transform -1 0 38752 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1698431365
transform -1 0 39760 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1698431365
transform 1 0 45472 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1698431365
transform 1 0 46144 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_142 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_158 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19040 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_166 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_176
timestamp 1698431365
transform 1 0 21056 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_184
timestamp 1698431365
transform 1 0 21952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_188
timestamp 1698431365
transform 1 0 22400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_190 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22624 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_193
timestamp 1698431365
transform 1 0 22960 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_222
timestamp 1698431365
transform 1 0 26208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_226
timestamp 1698431365
transform 1 0 26656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_234
timestamp 1698431365
transform 1 0 27552 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_290
timestamp 1698431365
transform 1 0 33824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_300
timestamp 1698431365
transform 1 0 34944 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_304
timestamp 1698431365
transform 1 0 35392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494
timestamp 1698431365
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698431365
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_104
timestamp 1698431365
transform 1 0 12992 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_108
timestamp 1698431365
transform 1 0 13440 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_110
timestamp 1698431365
transform 1 0 13664 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_148
timestamp 1698431365
transform 1 0 17920 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_166
timestamp 1698431365
transform 1 0 19936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_203
timestamp 1698431365
transform 1 0 24080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698431365
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_286
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_323
timestamp 1698431365
transform 1 0 37520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_327
timestamp 1698431365
transform 1 0 37968 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_343
timestamp 1698431365
transform 1 0 39760 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_347
timestamp 1698431365
transform 1 0 40208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_111
timestamp 1698431365
transform 1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_113
timestamp 1698431365
transform 1 0 14000 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_120
timestamp 1698431365
transform 1 0 14784 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_136
timestamp 1698431365
transform 1 0 16576 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_144
timestamp 1698431365
transform 1 0 17472 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_222
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_290
timestamp 1698431365
transform 1 0 33824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_294
timestamp 1698431365
transform 1 0 34272 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_310
timestamp 1698431365
transform 1 0 36064 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698431365
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_346
timestamp 1698431365
transform 1 0 40096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_350
timestamp 1698431365
transform 1 0 40544 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_382
timestamp 1698431365
transform 1 0 44128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_384
timestamp 1698431365
transform 1 0 44352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698431365
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_104
timestamp 1698431365
transform 1 0 12992 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_134
timestamp 1698431365
transform 1 0 16352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_138
timestamp 1698431365
transform 1 0 16800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_163
timestamp 1698431365
transform 1 0 19600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_167
timestamp 1698431365
transform 1 0 20048 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_204
timestamp 1698431365
transform 1 0 24192 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_208
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_214
timestamp 1698431365
transform 1 0 25312 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_221
timestamp 1698431365
transform 1 0 26096 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_252
timestamp 1698431365
transform 1 0 29568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_256
timestamp 1698431365
transform 1 0 30016 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_263
timestamp 1698431365
transform 1 0 30800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_297
timestamp 1698431365
transform 1 0 34608 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_301
timestamp 1698431365
transform 1 0 35056 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_317
timestamp 1698431365
transform 1 0 36848 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_113
timestamp 1698431365
transform 1 0 14000 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_136
timestamp 1698431365
transform 1 0 16576 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_168
timestamp 1698431365
transform 1 0 20160 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_185
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_191
timestamp 1698431365
transform 1 0 22736 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_197
timestamp 1698431365
transform 1 0 23408 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_201
timestamp 1698431365
transform 1 0 23856 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_233
timestamp 1698431365
transform 1 0 27440 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_253
timestamp 1698431365
transform 1 0 29680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_257
timestamp 1698431365
transform 1 0 30128 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_261
timestamp 1698431365
transform 1 0 30576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_269
timestamp 1698431365
transform 1 0 31472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_271
timestamp 1698431365
transform 1 0 31696 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_287
timestamp 1698431365
transform 1 0 33488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_303
timestamp 1698431365
transform 1 0 35280 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_325
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_327
timestamp 1698431365
transform 1 0 37968 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_357
timestamp 1698431365
transform 1 0 41328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_361
timestamp 1698431365
transform 1 0 41776 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_377
timestamp 1698431365
transform 1 0 43568 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_88
timestamp 1698431365
transform 1 0 11200 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_92
timestamp 1698431365
transform 1 0 11648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_94
timestamp 1698431365
transform 1 0 11872 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_124
timestamp 1698431365
transform 1 0 15232 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_128
timestamp 1698431365
transform 1 0 15680 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_144
timestamp 1698431365
transform 1 0 17472 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_228
timestamp 1698431365
transform 1 0 26880 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_232
timestamp 1698431365
transform 1 0 27328 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_248
timestamp 1698431365
transform 1 0 29120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_250
timestamp 1698431365
transform 1 0 29344 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_284
timestamp 1698431365
transform 1 0 33152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_287
timestamp 1698431365
transform 1 0 33488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_291
timestamp 1698431365
transform 1 0 33936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_324
timestamp 1698431365
transform 1 0 37632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_328
timestamp 1698431365
transform 1 0 38080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_330
timestamp 1698431365
transform 1 0 38304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_345
timestamp 1698431365
transform 1 0 39984 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_349
timestamp 1698431365
transform 1 0 40432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698431365
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_85
timestamp 1698431365
transform 1 0 10864 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_89
timestamp 1698431365
transform 1 0 11312 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_96
timestamp 1698431365
transform 1 0 12096 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_109
timestamp 1698431365
transform 1 0 13552 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_112
timestamp 1698431365
transform 1 0 13888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_116
timestamp 1698431365
transform 1 0 14336 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_133
timestamp 1698431365
transform 1 0 16240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_170
timestamp 1698431365
transform 1 0 20384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_183
timestamp 1698431365
transform 1 0 21840 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_192
timestamp 1698431365
transform 1 0 22848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_196
timestamp 1698431365
transform 1 0 23296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_229
timestamp 1698431365
transform 1 0 26992 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_269
timestamp 1698431365
transform 1 0 31472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_286
timestamp 1698431365
transform 1 0 33376 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_290
timestamp 1698431365
transform 1 0 33824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_294
timestamp 1698431365
transform 1 0 34272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_304
timestamp 1698431365
transform 1 0 35392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_312
timestamp 1698431365
transform 1 0 36288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_332
timestamp 1698431365
transform 1 0 38528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_349
timestamp 1698431365
transform 1 0 40432 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_489
timestamp 1698431365
transform 1 0 56112 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_505
timestamp 1698431365
transform 1 0 57904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_80
timestamp 1698431365
transform 1 0 10304 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_152
timestamp 1698431365
transform 1 0 18368 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_155
timestamp 1698431365
transform 1 0 18704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_174
timestamp 1698431365
transform 1 0 20832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_193
timestamp 1698431365
transform 1 0 22960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_197
timestamp 1698431365
transform 1 0 23408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_201
timestamp 1698431365
transform 1 0 23856 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_292
timestamp 1698431365
transform 1 0 34048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_316
timestamp 1698431365
transform 1 0 36736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_320
timestamp 1698431365
transform 1 0 37184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_324
timestamp 1698431365
transform 1 0 37632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_328
timestamp 1698431365
transform 1 0 38080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_85
timestamp 1698431365
transform 1 0 10864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_87
timestamp 1698431365
transform 1 0 11088 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_94
timestamp 1698431365
transform 1 0 11872 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_102
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_126
timestamp 1698431365
transform 1 0 15456 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_134
timestamp 1698431365
transform 1 0 16352 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_138
timestamp 1698431365
transform 1 0 16800 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_151
timestamp 1698431365
transform 1 0 18256 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_162
timestamp 1698431365
transform 1 0 19488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_166
timestamp 1698431365
transform 1 0 19936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_170
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_183
timestamp 1698431365
transform 1 0 21840 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_195
timestamp 1698431365
transform 1 0 23184 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_199
timestamp 1698431365
transform 1 0 23632 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_229
timestamp 1698431365
transform 1 0 26992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_253
timestamp 1698431365
transform 1 0 29680 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_269
timestamp 1698431365
transform 1 0 31472 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_275
timestamp 1698431365
transform 1 0 32144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_279
timestamp 1698431365
transform 1 0 32592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_283
timestamp 1698431365
transform 1 0 33040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_293
timestamp 1698431365
transform 1 0 34160 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_301
timestamp 1698431365
transform 1 0 35056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_305
timestamp 1698431365
transform 1 0 35504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_309
timestamp 1698431365
transform 1 0 35952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_335
timestamp 1698431365
transform 1 0 38864 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_368
timestamp 1698431365
transform 1 0 42560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_372
timestamp 1698431365
transform 1 0 43008 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_380
timestamp 1698431365
transform 1 0 43904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698431365
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_489
timestamp 1698431365
transform 1 0 56112 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_505
timestamp 1698431365
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_76
timestamp 1698431365
transform 1 0 9856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_78
timestamp 1698431365
transform 1 0 10080 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_108
timestamp 1698431365
transform 1 0 13440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_125
timestamp 1698431365
transform 1 0 15344 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_133
timestamp 1698431365
transform 1 0 16240 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_144
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_159
timestamp 1698431365
transform 1 0 19152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_176
timestamp 1698431365
transform 1 0 21056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_180
timestamp 1698431365
transform 1 0 21504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_182
timestamp 1698431365
transform 1 0 21728 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_189
timestamp 1698431365
transform 1 0 22512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_201
timestamp 1698431365
transform 1 0 23856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_205
timestamp 1698431365
transform 1 0 24304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_218
timestamp 1698431365
transform 1 0 25760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_232
timestamp 1698431365
transform 1 0 27328 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_239
timestamp 1698431365
transform 1 0 28112 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_243
timestamp 1698431365
transform 1 0 28560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_247
timestamp 1698431365
transform 1 0 29008 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_263
timestamp 1698431365
transform 1 0 30800 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_270
timestamp 1698431365
transform 1 0 31584 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_278
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_303
timestamp 1698431365
transform 1 0 35280 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_305
timestamp 1698431365
transform 1 0 35504 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_321
timestamp 1698431365
transform 1 0 37296 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_335
timestamp 1698431365
transform 1 0 38864 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_339
timestamp 1698431365
transform 1 0 39312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_347
timestamp 1698431365
transform 1 0 40208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_360
timestamp 1698431365
transform 1 0 41664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_368
timestamp 1698431365
transform 1 0 42560 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_400
timestamp 1698431365
transform 1 0 46144 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698431365
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_85
timestamp 1698431365
transform 1 0 10864 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_93
timestamp 1698431365
transform 1 0 11760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_111
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_115
timestamp 1698431365
transform 1 0 14224 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_123
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_135
timestamp 1698431365
transform 1 0 16464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_139
timestamp 1698431365
transform 1 0 16912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_170
timestamp 1698431365
transform 1 0 20384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_217
timestamp 1698431365
transform 1 0 25648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_221
timestamp 1698431365
transform 1 0 26096 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_231
timestamp 1698431365
transform 1 0 27216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_255
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_257
timestamp 1698431365
transform 1 0 30128 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_274
timestamp 1698431365
transform 1 0 32032 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_352
timestamp 1698431365
transform 1 0 40768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_391
timestamp 1698431365
transform 1 0 45136 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_489
timestamp 1698431365
transform 1 0 56112 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_505
timestamp 1698431365
transform 1 0 57904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_128
timestamp 1698431365
transform 1 0 15680 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_162
timestamp 1698431365
transform 1 0 19488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_193
timestamp 1698431365
transform 1 0 22960 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_216
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_228
timestamp 1698431365
transform 1 0 26880 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_292
timestamp 1698431365
transform 1 0 34048 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_317
timestamp 1698431365
transform 1 0 36848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_345
timestamp 1698431365
transform 1 0 39984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_360
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_392
timestamp 1698431365
transform 1 0 45248 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_408
timestamp 1698431365
transform 1 0 47040 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_53
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_57
timestamp 1698431365
transform 1 0 7728 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_59
timestamp 1698431365
transform 1 0 7952 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_89
timestamp 1698431365
transform 1 0 11312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_93
timestamp 1698431365
transform 1 0 11760 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_159
timestamp 1698431365
transform 1 0 19152 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_183
timestamp 1698431365
transform 1 0 21840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_191
timestamp 1698431365
transform 1 0 22736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_211
timestamp 1698431365
transform 1 0 24976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_221
timestamp 1698431365
transform 1 0 26096 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_228
timestamp 1698431365
transform 1 0 26880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_230
timestamp 1698431365
transform 1 0 27104 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_253
timestamp 1698431365
transform 1 0 29680 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_277
timestamp 1698431365
transform 1 0 32368 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_288
timestamp 1698431365
transform 1 0 33600 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_292
timestamp 1698431365
transform 1 0 34048 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_294
timestamp 1698431365
transform 1 0 34272 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_327
timestamp 1698431365
transform 1 0 37968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_331
timestamp 1698431365
transform 1 0 38416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_340
timestamp 1698431365
transform 1 0 39424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_344
timestamp 1698431365
transform 1 0 39872 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_360
timestamp 1698431365
transform 1 0 41664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_377
timestamp 1698431365
transform 1 0 43568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_416
timestamp 1698431365
transform 1 0 47936 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_448
timestamp 1698431365
transform 1 0 51520 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_452
timestamp 1698431365
transform 1 0 51968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_454
timestamp 1698431365
transform 1 0 52192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_489
timestamp 1698431365
transform 1 0 56112 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_505
timestamp 1698431365
transform 1 0 57904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_34
timestamp 1698431365
transform 1 0 5152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_36
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_84
timestamp 1698431365
transform 1 0 10752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_100
timestamp 1698431365
transform 1 0 12544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_104
timestamp 1698431365
transform 1 0 12992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_106
timestamp 1698431365
transform 1 0 13216 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_122
timestamp 1698431365
transform 1 0 15008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_124
timestamp 1698431365
transform 1 0 15232 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_157
timestamp 1698431365
transform 1 0 18928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_161
timestamp 1698431365
transform 1 0 19376 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_185
timestamp 1698431365
transform 1 0 22064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_187
timestamp 1698431365
transform 1 0 22288 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_227
timestamp 1698431365
transform 1 0 26768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_229
timestamp 1698431365
transform 1 0 26992 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_268
timestamp 1698431365
transform 1 0 31360 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_300
timestamp 1698431365
transform 1 0 34944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_322
timestamp 1698431365
transform 1 0 37408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_326
timestamp 1698431365
transform 1 0 37856 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_356
timestamp 1698431365
transform 1 0 41216 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_390
timestamp 1698431365
transform 1 0 45024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_394
timestamp 1698431365
transform 1 0 45472 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_410
timestamp 1698431365
transform 1 0 47264 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_418
timestamp 1698431365
transform 1 0 48160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698431365
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_53
timestamp 1698431365
transform 1 0 7280 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_61
timestamp 1698431365
transform 1 0 8176 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_91
timestamp 1698431365
transform 1 0 11536 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_95
timestamp 1698431365
transform 1 0 11984 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698431365
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698431365
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_131
timestamp 1698431365
transform 1 0 16016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_192
timestamp 1698431365
transform 1 0 22848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_210
timestamp 1698431365
transform 1 0 24864 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_270
timestamp 1698431365
transform 1 0 31584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_286
timestamp 1698431365
transform 1 0 33376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_294
timestamp 1698431365
transform 1 0 34272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_296
timestamp 1698431365
transform 1 0 34496 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_354
timestamp 1698431365
transform 1 0 40992 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_377
timestamp 1698431365
transform 1 0 43568 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_489
timestamp 1698431365
transform 1 0 56112 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_505
timestamp 1698431365
transform 1 0 57904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_34
timestamp 1698431365
transform 1 0 5152 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_38
timestamp 1698431365
transform 1 0 5600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_76
timestamp 1698431365
transform 1 0 9856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_99
timestamp 1698431365
transform 1 0 12432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_129
timestamp 1698431365
transform 1 0 15792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_148
timestamp 1698431365
transform 1 0 17920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_157
timestamp 1698431365
transform 1 0 18928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_194
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_198
timestamp 1698431365
transform 1 0 23520 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_202
timestamp 1698431365
transform 1 0 23968 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698431365
transform 1 0 24304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_226
timestamp 1698431365
transform 1 0 26656 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_234
timestamp 1698431365
transform 1 0 27552 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_236
timestamp 1698431365
transform 1 0 27776 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_247
timestamp 1698431365
transform 1 0 29008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_259
timestamp 1698431365
transform 1 0 30352 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_275
timestamp 1698431365
transform 1 0 32144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_298
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_306
timestamp 1698431365
transform 1 0 35616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_310
timestamp 1698431365
transform 1 0 36064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_312
timestamp 1698431365
transform 1 0 36288 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_323
timestamp 1698431365
transform 1 0 37520 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_331
timestamp 1698431365
transform 1 0 38416 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_344
timestamp 1698431365
transform 1 0 39872 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_348
timestamp 1698431365
transform 1 0 40320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_410
timestamp 1698431365
transform 1 0 47264 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_418
timestamp 1698431365
transform 1 0 48160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698431365
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_53
timestamp 1698431365
transform 1 0 7280 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_135
timestamp 1698431365
transform 1 0 16464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_139
timestamp 1698431365
transform 1 0 16912 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_162
timestamp 1698431365
transform 1 0 19488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_170
timestamp 1698431365
transform 1 0 20384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_213
timestamp 1698431365
transform 1 0 25200 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_217
timestamp 1698431365
transform 1 0 25648 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_220
timestamp 1698431365
transform 1 0 25984 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_236
timestamp 1698431365
transform 1 0 27776 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_257
timestamp 1698431365
transform 1 0 30128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_261
timestamp 1698431365
transform 1 0 30576 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_264
timestamp 1698431365
transform 1 0 30912 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_268
timestamp 1698431365
transform 1 0 31360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_276
timestamp 1698431365
transform 1 0 32256 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_292
timestamp 1698431365
transform 1 0 34048 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_301
timestamp 1698431365
transform 1 0 35056 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_309
timestamp 1698431365
transform 1 0 35952 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_313
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_325
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_331
timestamp 1698431365
transform 1 0 38416 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_363
timestamp 1698431365
transform 1 0 42000 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_489
timestamp 1698431365
transform 1 0 56112 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_505
timestamp 1698431365
transform 1 0 57904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_78
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_80
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_133
timestamp 1698431365
transform 1 0 16240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_157
timestamp 1698431365
transform 1 0 18928 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_167
timestamp 1698431365
transform 1 0 20048 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698431365
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_242
timestamp 1698431365
transform 1 0 28448 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_250
timestamp 1698431365
transform 1 0 29344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_270
timestamp 1698431365
transform 1 0 31584 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_340
timestamp 1698431365
transform 1 0 39424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_344
timestamp 1698431365
transform 1 0 39872 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_348
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_360
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_365
timestamp 1698431365
transform 1 0 42224 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_397
timestamp 1698431365
transform 1 0 45808 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_413
timestamp 1698431365
transform 1 0 47600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_417
timestamp 1698431365
transform 1 0 48048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698431365
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_53
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_55
timestamp 1698431365
transform 1 0 7504 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_91
timestamp 1698431365
transform 1 0 11536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_97
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_113
timestamp 1698431365
transform 1 0 14000 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_115
timestamp 1698431365
transform 1 0 14224 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_122
timestamp 1698431365
transform 1 0 15008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_153
timestamp 1698431365
transform 1 0 18480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_157
timestamp 1698431365
transform 1 0 18928 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_203
timestamp 1698431365
transform 1 0 24080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_211
timestamp 1698431365
transform 1 0 24976 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_238
timestamp 1698431365
transform 1 0 28000 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_249
timestamp 1698431365
transform 1 0 29232 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_256
timestamp 1698431365
transform 1 0 30016 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_276
timestamp 1698431365
transform 1 0 32256 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_280
timestamp 1698431365
transform 1 0 32704 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_298
timestamp 1698431365
transform 1 0 34720 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_307
timestamp 1698431365
transform 1 0 35728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_333
timestamp 1698431365
transform 1 0 38640 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_371
timestamp 1698431365
transform 1 0 42896 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_375
timestamp 1698431365
transform 1 0 43344 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_383
timestamp 1698431365
transform 1 0 44240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_489
timestamp 1698431365
transform 1 0 56112 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_505
timestamp 1698431365
transform 1 0 57904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_34
timestamp 1698431365
transform 1 0 5152 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_38
timestamp 1698431365
transform 1 0 5600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_80
timestamp 1698431365
transform 1 0 10304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_126
timestamp 1698431365
transform 1 0 15456 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_130
timestamp 1698431365
transform 1 0 15904 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_184
timestamp 1698431365
transform 1 0 21952 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_188
timestamp 1698431365
transform 1 0 22400 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_191
timestamp 1698431365
transform 1 0 22736 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_267
timestamp 1698431365
transform 1 0 31248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_290
timestamp 1698431365
transform 1 0 33824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_302
timestamp 1698431365
transform 1 0 35168 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_312
timestamp 1698431365
transform 1 0 36288 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_320
timestamp 1698431365
transform 1 0 37184 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_324
timestamp 1698431365
transform 1 0 37632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_330
timestamp 1698431365
transform 1 0 38304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_381
timestamp 1698431365
transform 1 0 44016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_385
timestamp 1698431365
transform 1 0 44464 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_417
timestamp 1698431365
transform 1 0 48048 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_419
timestamp 1698431365
transform 1 0 48272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698431365
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_45
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_49
timestamp 1698431365
transform 1 0 6832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_51
timestamp 1698431365
transform 1 0 7056 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_81
timestamp 1698431365
transform 1 0 10416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_85
timestamp 1698431365
transform 1 0 10864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_93
timestamp 1698431365
transform 1 0 11760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_111
timestamp 1698431365
transform 1 0 13776 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_127
timestamp 1698431365
transform 1 0 15568 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_131
timestamp 1698431365
transform 1 0 16016 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_134
timestamp 1698431365
transform 1 0 16352 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_142
timestamp 1698431365
transform 1 0 17248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_144
timestamp 1698431365
transform 1 0 17472 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_200
timestamp 1698431365
transform 1 0 23744 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_204
timestamp 1698431365
transform 1 0 24192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_208
timestamp 1698431365
transform 1 0 24640 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_216
timestamp 1698431365
transform 1 0 25536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_220
timestamp 1698431365
transform 1 0 25984 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_223
timestamp 1698431365
transform 1 0 26320 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_237
timestamp 1698431365
transform 1 0 27888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_257
timestamp 1698431365
transform 1 0 30128 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_273
timestamp 1698431365
transform 1 0 31920 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_281
timestamp 1698431365
transform 1 0 32816 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_284
timestamp 1698431365
transform 1 0 33152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698431365
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_346
timestamp 1698431365
transform 1 0 40096 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_378
timestamp 1698431365
transform 1 0 43680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_382
timestamp 1698431365
transform 1 0 44128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_384
timestamp 1698431365
transform 1 0 44352 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698431365
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_489
timestamp 1698431365
transform 1 0 56112 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_505
timestamp 1698431365
transform 1 0 57904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_84
timestamp 1698431365
transform 1 0 10752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_92
timestamp 1698431365
transform 1 0 11648 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_110
timestamp 1698431365
transform 1 0 13664 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_201
timestamp 1698431365
transform 1 0 23856 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_218
timestamp 1698431365
transform 1 0 25760 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_222
timestamp 1698431365
transform 1 0 26208 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_245
timestamp 1698431365
transform 1 0 28784 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_257
timestamp 1698431365
transform 1 0 30128 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_261
timestamp 1698431365
transform 1 0 30576 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698431365
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_290
timestamp 1698431365
transform 1 0 33824 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_306
timestamp 1698431365
transform 1 0 35616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_318
timestamp 1698431365
transform 1 0 36960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_322
timestamp 1698431365
transform 1 0 37408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_326
timestamp 1698431365
transform 1 0 37856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_337
timestamp 1698431365
transform 1 0 39088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_341
timestamp 1698431365
transform 1 0 39536 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_380
timestamp 1698431365
transform 1 0 43904 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_412
timestamp 1698431365
transform 1 0 47488 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_41
timestamp 1698431365
transform 1 0 5936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_49
timestamp 1698431365
transform 1 0 6832 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698431365
transform 1 0 21392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_282
timestamp 1698431365
transform 1 0 32928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_334
timestamp 1698431365
transform 1 0 38752 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_338
timestamp 1698431365
transform 1 0 39200 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_353
timestamp 1698431365
transform 1 0 40880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_357
timestamp 1698431365
transform 1 0 41328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_361
timestamp 1698431365
transform 1 0 41776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_363
timestamp 1698431365
transform 1 0 42000 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_368
timestamp 1698431365
transform 1 0 42560 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698431365
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_489
timestamp 1698431365
transform 1 0 56112 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_505
timestamp 1698431365
transform 1 0 57904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_34
timestamp 1698431365
transform 1 0 5152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_36
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_43
timestamp 1698431365
transform 1 0 6160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_57
timestamp 1698431365
transform 1 0 7728 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_65
timestamp 1698431365
transform 1 0 8624 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_76
timestamp 1698431365
transform 1 0 9856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_92
timestamp 1698431365
transform 1 0 11648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_102
timestamp 1698431365
transform 1 0 12768 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_196
timestamp 1698431365
transform 1 0 23296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_216
timestamp 1698431365
transform 1 0 25536 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_232
timestamp 1698431365
transform 1 0 27328 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_241
timestamp 1698431365
transform 1 0 28336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_245
timestamp 1698431365
transform 1 0 28784 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_254
timestamp 1698431365
transform 1 0 29792 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_258
timestamp 1698431365
transform 1 0 30240 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_274
timestamp 1698431365
transform 1 0 32032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698431365
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_292
timestamp 1698431365
transform 1 0 34048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_304
timestamp 1698431365
transform 1 0 35392 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_335
timestamp 1698431365
transform 1 0 38864 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_381
timestamp 1698431365
transform 1 0 44016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_385
timestamp 1698431365
transform 1 0 44464 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_417
timestamp 1698431365
transform 1 0 48048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_419
timestamp 1698431365
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698431365
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1698431365
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_66
timestamp 1698431365
transform 1 0 8736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_70
timestamp 1698431365
transform 1 0 9184 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_94
timestamp 1698431365
transform 1 0 11872 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_102
timestamp 1698431365
transform 1 0 12768 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_125
timestamp 1698431365
transform 1 0 15344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_189
timestamp 1698431365
transform 1 0 22512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_206
timestamp 1698431365
transform 1 0 24416 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698431365
transform 1 0 25312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_218
timestamp 1698431365
transform 1 0 25760 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_226
timestamp 1698431365
transform 1 0 26656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_230
timestamp 1698431365
transform 1 0 27104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_234
timestamp 1698431365
transform 1 0 27552 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698431365
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_255
timestamp 1698431365
transform 1 0 29904 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_292
timestamp 1698431365
transform 1 0 34048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_296
timestamp 1698431365
transform 1 0 34496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_330
timestamp 1698431365
transform 1 0 38304 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_338
timestamp 1698431365
transform 1 0 39200 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_373
timestamp 1698431365
transform 1 0 43120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_377
timestamp 1698431365
transform 1 0 43568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_451
timestamp 1698431365
transform 1 0 51856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_489
timestamp 1698431365
transform 1 0 56112 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_505
timestamp 1698431365
transform 1 0 57904 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_10
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_14
timestamp 1698431365
transform 1 0 2912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_44
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_48
timestamp 1698431365
transform 1 0 6720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_50
timestamp 1698431365
transform 1 0 6944 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_64
timestamp 1698431365
transform 1 0 8512 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_128
timestamp 1698431365
transform 1 0 15680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_130
timestamp 1698431365
transform 1 0 15904 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_168
timestamp 1698431365
transform 1 0 20160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_170
timestamp 1698431365
transform 1 0 20384 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_226
timestamp 1698431365
transform 1 0 26656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_267
timestamp 1698431365
transform 1 0 31248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_269
timestamp 1698431365
transform 1 0 31472 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_301
timestamp 1698431365
transform 1 0 35056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_305
timestamp 1698431365
transform 1 0 35504 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_335
timestamp 1698431365
transform 1 0 38864 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_343
timestamp 1698431365
transform 1 0 39760 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_347
timestamp 1698431365
transform 1 0 40208 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698431365
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_43
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_47
timestamp 1698431365
transform 1 0 6608 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_73
timestamp 1698431365
transform 1 0 9520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_75
timestamp 1698431365
transform 1 0 9744 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_115
timestamp 1698431365
transform 1 0 14224 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_183
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_187
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_230
timestamp 1698431365
transform 1 0 27104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_240
timestamp 1698431365
transform 1 0 28224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_253
timestamp 1698431365
transform 1 0 29680 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_269
timestamp 1698431365
transform 1 0 31472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_271
timestamp 1698431365
transform 1 0 31696 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_346
timestamp 1698431365
transform 1 0 40096 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_378
timestamp 1698431365
transform 1 0 43680 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_382
timestamp 1698431365
transform 1 0 44128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_451
timestamp 1698431365
transform 1 0 51856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_489
timestamp 1698431365
transform 1 0 56112 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_505
timestamp 1698431365
transform 1 0 57904 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_34
timestamp 1698431365
transform 1 0 5152 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_50
timestamp 1698431365
transform 1 0 6944 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_87
timestamp 1698431365
transform 1 0 11088 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_129
timestamp 1698431365
transform 1 0 15792 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_131
timestamp 1698431365
transform 1 0 16016 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_165
timestamp 1698431365
transform 1 0 19824 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_177
timestamp 1698431365
transform 1 0 21168 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_224
timestamp 1698431365
transform 1 0 26432 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_230
timestamp 1698431365
transform 1 0 27104 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_238
timestamp 1698431365
transform 1 0 28000 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_242
timestamp 1698431365
transform 1 0 28448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_248
timestamp 1698431365
transform 1 0 29120 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_264
timestamp 1698431365
transform 1 0 30912 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_272
timestamp 1698431365
transform 1 0 31808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_311
timestamp 1698431365
transform 1 0 36176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_315
timestamp 1698431365
transform 1 0 36624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_319
timestamp 1698431365
transform 1 0 37072 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_335
timestamp 1698431365
transform 1 0 38864 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_343
timestamp 1698431365
transform 1 0 39760 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698431365
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698431365
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_43
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_59
timestamp 1698431365
transform 1 0 7952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_61
timestamp 1698431365
transform 1 0 8176 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_75
timestamp 1698431365
transform 1 0 9744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_77
timestamp 1698431365
transform 1 0 9968 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_109
timestamp 1698431365
transform 1 0 13552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_126
timestamp 1698431365
transform 1 0 15456 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_128
timestamp 1698431365
transform 1 0 15680 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_206
timestamp 1698431365
transform 1 0 24416 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_210
timestamp 1698431365
transform 1 0 24864 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_255
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_267
timestamp 1698431365
transform 1 0 31248 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_283
timestamp 1698431365
transform 1 0 33040 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_289
timestamp 1698431365
transform 1 0 33712 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_305
timestamp 1698431365
transform 1 0 35504 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_333
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_337
timestamp 1698431365
transform 1 0 39088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_368
timestamp 1698431365
transform 1 0 42560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_372
timestamp 1698431365
transform 1 0 43008 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_380
timestamp 1698431365
transform 1 0 43904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698431365
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_489
timestamp 1698431365
transform 1 0 56112 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_505
timestamp 1698431365
transform 1 0 57904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_10
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_14
timestamp 1698431365
transform 1 0 2912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_16
timestamp 1698431365
transform 1 0 3136 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_46
timestamp 1698431365
transform 1 0 6496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_55
timestamp 1698431365
transform 1 0 7504 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_81
timestamp 1698431365
transform 1 0 10416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_163
timestamp 1698431365
transform 1 0 19600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_167
timestamp 1698431365
transform 1 0 20048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_171
timestamp 1698431365
transform 1 0 20496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_177
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_193
timestamp 1698431365
transform 1 0 22960 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_201
timestamp 1698431365
transform 1 0 23856 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_205
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_243
timestamp 1698431365
transform 1 0 28560 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_251
timestamp 1698431365
transform 1 0 29456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_253
timestamp 1698431365
transform 1 0 29680 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_275
timestamp 1698431365
transform 1 0 32144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_302
timestamp 1698431365
transform 1 0 35168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_304
timestamp 1698431365
transform 1 0 35392 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_307
timestamp 1698431365
transform 1 0 35728 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_311
timestamp 1698431365
transform 1 0 36176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_323
timestamp 1698431365
transform 1 0 37520 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_339
timestamp 1698431365
transform 1 0 39312 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_345
timestamp 1698431365
transform 1 0 39984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_347
timestamp 1698431365
transform 1 0 40208 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_366
timestamp 1698431365
transform 1 0 42336 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_398
timestamp 1698431365
transform 1 0 45920 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_414
timestamp 1698431365
transform 1 0 47712 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_418
timestamp 1698431365
transform 1 0 48160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698431365
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_508
timestamp 1698431365
transform 1 0 58240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_44
timestamp 1698431365
transform 1 0 6272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_48
timestamp 1698431365
transform 1 0 6720 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_52
timestamp 1698431365
transform 1 0 7168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_54
timestamp 1698431365
transform 1 0 7392 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_100
timestamp 1698431365
transform 1 0 12544 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_150
timestamp 1698431365
transform 1 0 18144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_152
timestamp 1698431365
transform 1 0 18368 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_157
timestamp 1698431365
transform 1 0 18928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_161
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_169
timestamp 1698431365
transform 1 0 20272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_185
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_187
timestamp 1698431365
transform 1 0 22288 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_219
timestamp 1698431365
transform 1 0 25872 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_235
timestamp 1698431365
transform 1 0 27664 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_276
timestamp 1698431365
transform 1 0 32256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_346
timestamp 1698431365
transform 1 0 40096 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_369
timestamp 1698431365
transform 1 0 42672 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698431365
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_489
timestamp 1698431365
transform 1 0 56112 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_505
timestamp 1698431365
transform 1 0 57904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_26
timestamp 1698431365
transform 1 0 4256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_59
timestamp 1698431365
transform 1 0 7952 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_63
timestamp 1698431365
transform 1 0 8400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_67
timestamp 1698431365
transform 1 0 8848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_84
timestamp 1698431365
transform 1 0 10752 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_100
timestamp 1698431365
transform 1 0 12544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_102
timestamp 1698431365
transform 1 0 12768 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_111
timestamp 1698431365
transform 1 0 13776 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_119
timestamp 1698431365
transform 1 0 14672 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_125
timestamp 1698431365
transform 1 0 15344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_129
timestamp 1698431365
transform 1 0 15792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_133
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_200
timestamp 1698431365
transform 1 0 23744 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_218
timestamp 1698431365
transform 1 0 25760 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_250
timestamp 1698431365
transform 1 0 29344 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_265
timestamp 1698431365
transform 1 0 31024 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_273
timestamp 1698431365
transform 1 0 31920 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_275
timestamp 1698431365
transform 1 0 32144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_278
timestamp 1698431365
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_311
timestamp 1698431365
transform 1 0 36176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_315
timestamp 1698431365
transform 1 0 36624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_317
timestamp 1698431365
transform 1 0 36848 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_348
timestamp 1698431365
transform 1 0 40320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_367
timestamp 1698431365
transform 1 0 42448 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_399
timestamp 1698431365
transform 1 0 46032 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_415
timestamp 1698431365
transform 1 0 47824 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_419
timestamp 1698431365
transform 1 0 48272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_48
timestamp 1698431365
transform 1 0 6720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_52
timestamp 1698431365
transform 1 0 7168 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_84
timestamp 1698431365
transform 1 0 10752 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_100
timestamp 1698431365
transform 1 0 12544 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_115
timestamp 1698431365
transform 1 0 14224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_117
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_122
timestamp 1698431365
transform 1 0 15008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_135
timestamp 1698431365
transform 1 0 16464 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_164
timestamp 1698431365
transform 1 0 19712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_200
timestamp 1698431365
transform 1 0 23744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_204
timestamp 1698431365
transform 1 0 24192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_208
timestamp 1698431365
transform 1 0 24640 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_212
timestamp 1698431365
transform 1 0 25088 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_237
timestamp 1698431365
transform 1 0 27888 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698431365
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_344
timestamp 1698431365
transform 1 0 39872 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_350
timestamp 1698431365
transform 1 0 40544 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_358
timestamp 1698431365
transform 1 0 41440 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_367
timestamp 1698431365
transform 1 0 42448 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_383
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698431365
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_489
timestamp 1698431365
transform 1 0 56112 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_505
timestamp 1698431365
transform 1 0 57904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_34
timestamp 1698431365
transform 1 0 5152 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_38
timestamp 1698431365
transform 1 0 5600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_40
timestamp 1698431365
transform 1 0 5824 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_76
timestamp 1698431365
transform 1 0 9856 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_84
timestamp 1698431365
transform 1 0 10752 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_86
timestamp 1698431365
transform 1 0 10976 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_97
timestamp 1698431365
transform 1 0 12208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_146
timestamp 1698431365
transform 1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_150
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_156
timestamp 1698431365
transform 1 0 18816 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_161
timestamp 1698431365
transform 1 0 19376 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_169
timestamp 1698431365
transform 1 0 20272 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_177
timestamp 1698431365
transform 1 0 21168 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_187
timestamp 1698431365
transform 1 0 22288 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_194
timestamp 1698431365
transform 1 0 23072 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_196
timestamp 1698431365
transform 1 0 23296 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_201
timestamp 1698431365
transform 1 0 23856 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_216
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_238
timestamp 1698431365
transform 1 0 28000 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_240
timestamp 1698431365
transform 1 0 28224 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_257
timestamp 1698431365
transform 1 0 30128 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_265
timestamp 1698431365
transform 1 0 31024 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_269
timestamp 1698431365
transform 1 0 31472 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_271
timestamp 1698431365
transform 1 0 31696 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_290
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_337
timestamp 1698431365
transform 1 0 39088 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_354
timestamp 1698431365
transform 1 0 40992 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_384
timestamp 1698431365
transform 1 0 44352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_388
timestamp 1698431365
transform 1 0 44800 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_508
timestamp 1698431365
transform 1 0 58240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_45
timestamp 1698431365
transform 1 0 6384 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_55
timestamp 1698431365
transform 1 0 7504 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_59
timestamp 1698431365
transform 1 0 7952 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_89
timestamp 1698431365
transform 1 0 11312 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_132
timestamp 1698431365
transform 1 0 16128 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_140
timestamp 1698431365
transform 1 0 17024 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_164
timestamp 1698431365
transform 1 0 19712 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_172
timestamp 1698431365
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_182
timestamp 1698431365
transform 1 0 21728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_186
timestamp 1698431365
transform 1 0 22176 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_198
timestamp 1698431365
transform 1 0 23520 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_200
timestamp 1698431365
transform 1 0 23744 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_206
timestamp 1698431365
transform 1 0 24416 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_224
timestamp 1698431365
transform 1 0 26432 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_231
timestamp 1698431365
transform 1 0 27216 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_239
timestamp 1698431365
transform 1 0 28112 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_303
timestamp 1698431365
transform 1 0 35280 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_319
timestamp 1698431365
transform 1 0 37072 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_332
timestamp 1698431365
transform 1 0 38528 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_351
timestamp 1698431365
transform 1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_361
timestamp 1698431365
transform 1 0 41776 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_377
timestamp 1698431365
transform 1 0 43568 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_419
timestamp 1698431365
transform 1 0 48272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_423
timestamp 1698431365
transform 1 0 48720 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_489
timestamp 1698431365
transform 1 0 56112 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_505
timestamp 1698431365
transform 1 0 57904 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_18
timestamp 1698431365
transform 1 0 3360 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_26
timestamp 1698431365
transform 1 0 4256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_30
timestamp 1698431365
transform 1 0 4704 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_76
timestamp 1698431365
transform 1 0 9856 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_102
timestamp 1698431365
transform 1 0 12768 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_110
timestamp 1698431365
transform 1 0 13664 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_119
timestamp 1698431365
transform 1 0 14672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_130
timestamp 1698431365
transform 1 0 15904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_138
timestamp 1698431365
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_183
timestamp 1698431365
transform 1 0 21840 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_199
timestamp 1698431365
transform 1 0 23632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_232
timestamp 1698431365
transform 1 0 27328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_236
timestamp 1698431365
transform 1 0 27776 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_244
timestamp 1698431365
transform 1 0 28672 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_248
timestamp 1698431365
transform 1 0 29120 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_278
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_295
timestamp 1698431365
transform 1 0 34384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_299
timestamp 1698431365
transform 1 0 34832 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_315
timestamp 1698431365
transform 1 0 36624 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_319
timestamp 1698431365
transform 1 0 37072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_369
timestamp 1698431365
transform 1 0 42672 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_401
timestamp 1698431365
transform 1 0 46256 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_417
timestamp 1698431365
transform 1 0 48048 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_426
timestamp 1698431365
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_430
timestamp 1698431365
transform 1 0 49504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_434
timestamp 1698431365
transform 1 0 49952 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_450
timestamp 1698431365
transform 1 0 51744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_454
timestamp 1698431365
transform 1 0 52192 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698431365
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_508
timestamp 1698431365
transform 1 0 58240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_41
timestamp 1698431365
transform 1 0 5936 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_46
timestamp 1698431365
transform 1 0 6496 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_54
timestamp 1698431365
transform 1 0 7392 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_116
timestamp 1698431365
transform 1 0 14336 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_125
timestamp 1698431365
transform 1 0 15344 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_129
timestamp 1698431365
transform 1 0 15792 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_192
timestamp 1698431365
transform 1 0 22848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_239
timestamp 1698431365
transform 1 0 28112 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_252
timestamp 1698431365
transform 1 0 29568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_291
timestamp 1698431365
transform 1 0 33936 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_295
timestamp 1698431365
transform 1 0 34384 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_299
timestamp 1698431365
transform 1 0 34832 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_354
timestamp 1698431365
transform 1 0 40992 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_391
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_424
timestamp 1698431365
transform 1 0 48832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_426
timestamp 1698431365
transform 1 0 49056 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_461
timestamp 1698431365
transform 1 0 52976 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_493
timestamp 1698431365
transform 1 0 56560 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_10
timestamp 1698431365
transform 1 0 2464 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_14
timestamp 1698431365
transform 1 0 2912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_44
timestamp 1698431365
transform 1 0 6272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_48
timestamp 1698431365
transform 1 0 6720 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_64
timestamp 1698431365
transform 1 0 8512 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_68
timestamp 1698431365
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_80
timestamp 1698431365
transform 1 0 10304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_84
timestamp 1698431365
transform 1 0 10752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_87
timestamp 1698431365
transform 1 0 11088 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_103
timestamp 1698431365
transform 1 0 12880 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_113
timestamp 1698431365
transform 1 0 14000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_121
timestamp 1698431365
transform 1 0 14896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_150
timestamp 1698431365
transform 1 0 18144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_152
timestamp 1698431365
transform 1 0 18368 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_195
timestamp 1698431365
transform 1 0 23184 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698431365
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_216
timestamp 1698431365
transform 1 0 25536 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_223
timestamp 1698431365
transform 1 0 26320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_225
timestamp 1698431365
transform 1 0 26544 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_237
timestamp 1698431365
transform 1 0 27888 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_258
timestamp 1698431365
transform 1 0 30240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_260
timestamp 1698431365
transform 1 0 30464 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_286
timestamp 1698431365
transform 1 0 33376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_290
timestamp 1698431365
transform 1 0 33824 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_331
timestamp 1698431365
transform 1 0 38416 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_339
timestamp 1698431365
transform 1 0 39312 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_357
timestamp 1698431365
transform 1 0 41328 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_359
timestamp 1698431365
transform 1 0 41552 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_403
timestamp 1698431365
transform 1 0 46480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_407
timestamp 1698431365
transform 1 0 46928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_409
timestamp 1698431365
transform 1 0 47152 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_441
timestamp 1698431365
transform 1 0 50736 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_481
timestamp 1698431365
transform 1 0 55216 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_489
timestamp 1698431365
transform 1 0 56112 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_508
timestamp 1698431365
transform 1 0 58240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_18
timestamp 1698431365
transform 1 0 3360 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_26
timestamp 1698431365
transform 1 0 4256 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_30
timestamp 1698431365
transform 1 0 4704 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_33
timestamp 1698431365
transform 1 0 5040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_39
timestamp 1698431365
transform 1 0 5712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_69
timestamp 1698431365
transform 1 0 9072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_73
timestamp 1698431365
transform 1 0 9520 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_109
timestamp 1698431365
transform 1 0 13552 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_118
timestamp 1698431365
transform 1 0 14560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_122
timestamp 1698431365
transform 1 0 15008 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_126
timestamp 1698431365
transform 1 0 15456 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_129
timestamp 1698431365
transform 1 0 15792 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_133
timestamp 1698431365
transform 1 0 16240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_137
timestamp 1698431365
transform 1 0 16688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_139
timestamp 1698431365
transform 1 0 16912 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_142
timestamp 1698431365
transform 1 0 17248 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_146
timestamp 1698431365
transform 1 0 17696 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_153
timestamp 1698431365
transform 1 0 18480 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_162
timestamp 1698431365
transform 1 0 19488 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_191
timestamp 1698431365
transform 1 0 22736 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_207
timestamp 1698431365
transform 1 0 24528 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_211
timestamp 1698431365
transform 1 0 24976 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_234
timestamp 1698431365
transform 1 0 27552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_238
timestamp 1698431365
transform 1 0 28000 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_242
timestamp 1698431365
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_253
timestamp 1698431365
transform 1 0 29680 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_257
timestamp 1698431365
transform 1 0 30128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_259
timestamp 1698431365
transform 1 0 30352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_265
timestamp 1698431365
transform 1 0 31024 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_269
timestamp 1698431365
transform 1 0 31472 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_271
timestamp 1698431365
transform 1 0 31696 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_321
timestamp 1698431365
transform 1 0 37296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_333
timestamp 1698431365
transform 1 0 38640 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_346
timestamp 1698431365
transform 1 0 40096 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_354
timestamp 1698431365
transform 1 0 40992 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_360
timestamp 1698431365
transform 1 0 41664 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_376
timestamp 1698431365
transform 1 0 43456 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_384
timestamp 1698431365
transform 1 0 44352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_411
timestamp 1698431365
transform 1 0 47376 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_431
timestamp 1698431365
transform 1 0 49616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_433
timestamp 1698431365
transform 1 0 49840 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_452
timestamp 1698431365
transform 1 0 51968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_454
timestamp 1698431365
transform 1 0 52192 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_461
timestamp 1698431365
transform 1 0 52976 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_469
timestamp 1698431365
transform 1 0 53872 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_472
timestamp 1698431365
transform 1 0 54208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_476
timestamp 1698431365
transform 1 0 54656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_480
timestamp 1698431365
transform 1 0 55104 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_496
timestamp 1698431365
transform 1 0 56896 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_504
timestamp 1698431365
transform 1 0 57792 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_508
timestamp 1698431365
transform 1 0 58240 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_39
timestamp 1698431365
transform 1 0 5712 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_47
timestamp 1698431365
transform 1 0 6608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_49
timestamp 1698431365
transform 1 0 6832 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_74
timestamp 1698431365
transform 1 0 9632 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_99
timestamp 1698431365
transform 1 0 12432 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_120
timestamp 1698431365
transform 1 0 14784 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_127
timestamp 1698431365
transform 1 0 15568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_137
timestamp 1698431365
transform 1 0 16688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_146
timestamp 1698431365
transform 1 0 17696 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_161
timestamp 1698431365
transform 1 0 19376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_163
timestamp 1698431365
transform 1 0 19600 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_174
timestamp 1698431365
transform 1 0 20832 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_183
timestamp 1698431365
transform 1 0 21840 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_187
timestamp 1698431365
transform 1 0 22288 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_197
timestamp 1698431365
transform 1 0 23408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_201
timestamp 1698431365
transform 1 0 23856 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_258
timestamp 1698431365
transform 1 0 30240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_275
timestamp 1698431365
transform 1 0 32144 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_290
timestamp 1698431365
transform 1 0 33824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_300
timestamp 1698431365
transform 1 0 34944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_304
timestamp 1698431365
transform 1 0 35392 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_312
timestamp 1698431365
transform 1 0 36288 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_316
timestamp 1698431365
transform 1 0 36736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_377
timestamp 1698431365
transform 1 0 43568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_409
timestamp 1698431365
transform 1 0 47152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_413
timestamp 1698431365
transform 1 0 47600 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_417
timestamp 1698431365
transform 1 0 48048 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_419
timestamp 1698431365
transform 1 0 48272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_439
timestamp 1698431365
transform 1 0 50512 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_443
timestamp 1698431365
transform 1 0 50960 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_452
timestamp 1698431365
transform 1 0 51968 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_456
timestamp 1698431365
transform 1 0 52416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_458
timestamp 1698431365
transform 1 0 52640 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_508
timestamp 1698431365
transform 1 0 58240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_10
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_18
timestamp 1698431365
transform 1 0 3360 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_26
timestamp 1698431365
transform 1 0 4256 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_30
timestamp 1698431365
transform 1 0 4704 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_33
timestamp 1698431365
transform 1 0 5040 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_70
timestamp 1698431365
transform 1 0 9184 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_87
timestamp 1698431365
transform 1 0 11088 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_95
timestamp 1698431365
transform 1 0 11984 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_99
timestamp 1698431365
transform 1 0 12432 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_118
timestamp 1698431365
transform 1 0 14560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_151
timestamp 1698431365
transform 1 0 18256 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_155
timestamp 1698431365
transform 1 0 18704 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_170
timestamp 1698431365
transform 1 0 20384 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_174
timestamp 1698431365
transform 1 0 20832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_182
timestamp 1698431365
transform 1 0 21728 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_195
timestamp 1698431365
transform 1 0 23184 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_208
timestamp 1698431365
transform 1 0 24640 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_255
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_274
timestamp 1698431365
transform 1 0 32032 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_283
timestamp 1698431365
transform 1 0 33040 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_291
timestamp 1698431365
transform 1 0 33936 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_325
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_375
timestamp 1698431365
transform 1 0 43344 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_379
timestamp 1698431365
transform 1 0 43792 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_382
timestamp 1698431365
transform 1 0 44128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_395
timestamp 1698431365
transform 1 0 45584 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_399
timestamp 1698431365
transform 1 0 46032 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_436
timestamp 1698431365
transform 1 0 50176 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_440
timestamp 1698431365
transform 1 0 50624 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_448
timestamp 1698431365
transform 1 0 51520 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_451
timestamp 1698431365
transform 1 0 51856 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_471
timestamp 1698431365
transform 1 0 54096 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_501
timestamp 1698431365
transform 1 0 57456 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_19
timestamp 1698431365
transform 1 0 3472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_45
timestamp 1698431365
transform 1 0 6384 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_63
timestamp 1698431365
transform 1 0 8400 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_67
timestamp 1698431365
transform 1 0 8848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_116
timestamp 1698431365
transform 1 0 14336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_160
timestamp 1698431365
transform 1 0 19264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_164
timestamp 1698431365
transform 1 0 19712 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_172
timestamp 1698431365
transform 1 0 20608 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_176
timestamp 1698431365
transform 1 0 21056 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_179
timestamp 1698431365
transform 1 0 21392 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_183
timestamp 1698431365
transform 1 0 21840 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_185
timestamp 1698431365
transform 1 0 22064 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_192
timestamp 1698431365
transform 1 0 22848 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_196
timestamp 1698431365
transform 1 0 23296 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_204
timestamp 1698431365
transform 1 0 24192 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_208
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_262
timestamp 1698431365
transform 1 0 30688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_270
timestamp 1698431365
transform 1 0 31584 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_295
timestamp 1698431365
transform 1 0 34384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_299
timestamp 1698431365
transform 1 0 34832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_319
timestamp 1698431365
transform 1 0 37072 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_323
timestamp 1698431365
transform 1 0 37520 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_390
timestamp 1698431365
transform 1 0 45024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_394
timestamp 1698431365
transform 1 0 45472 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_403
timestamp 1698431365
transform 1 0 46480 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_407
timestamp 1698431365
transform 1 0 46928 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_410
timestamp 1698431365
transform 1 0 47264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_435
timestamp 1698431365
transform 1 0 50064 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_459
timestamp 1698431365
transform 1 0 52752 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_461
timestamp 1698431365
transform 1 0 52976 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_480
timestamp 1698431365
transform 1 0 55104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_39
timestamp 1698431365
transform 1 0 5712 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_51
timestamp 1698431365
transform 1 0 7056 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_98
timestamp 1698431365
transform 1 0 12320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_168
timestamp 1698431365
transform 1 0 20160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_209
timestamp 1698431365
transform 1 0 24752 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_217
timestamp 1698431365
transform 1 0 25648 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_219
timestamp 1698431365
transform 1 0 25872 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_230
timestamp 1698431365
transform 1 0 27104 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_234
timestamp 1698431365
transform 1 0 27552 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_261
timestamp 1698431365
transform 1 0 30576 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_342
timestamp 1698431365
transform 1 0 39648 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_358
timestamp 1698431365
transform 1 0 41440 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_366
timestamp 1698431365
transform 1 0 42336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_370
timestamp 1698431365
transform 1 0 42784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_380
timestamp 1698431365
transform 1 0 43904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_384
timestamp 1698431365
transform 1 0 44352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_413
timestamp 1698431365
transform 1 0 47600 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_4
timestamp 1698431365
transform 1 0 1792 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_25
timestamp 1698431365
transform 1 0 4144 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_32
timestamp 1698431365
transform 1 0 4928 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_76
timestamp 1698431365
transform 1 0 9856 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_124
timestamp 1698431365
transform 1 0 15232 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_198
timestamp 1698431365
transform 1 0 23520 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698431365
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_237
timestamp 1698431365
transform 1 0 27888 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_247
timestamp 1698431365
transform 1 0 29008 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_263
timestamp 1698431365
transform 1 0 30800 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698431365
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_290
timestamp 1698431365
transform 1 0 33824 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_294
timestamp 1698431365
transform 1 0 34272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_296
timestamp 1698431365
transform 1 0 34496 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_303
timestamp 1698431365
transform 1 0 35280 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_307
timestamp 1698431365
transform 1 0 35728 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_311
timestamp 1698431365
transform 1 0 36176 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_347
timestamp 1698431365
transform 1 0 40208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_360
timestamp 1698431365
transform 1 0 41664 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_371
timestamp 1698431365
transform 1 0 42896 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_375
timestamp 1698431365
transform 1 0 43344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_377
timestamp 1698431365
transform 1 0 43568 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_380
timestamp 1698431365
transform 1 0 43904 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_384
timestamp 1698431365
transform 1 0 44352 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_407
timestamp 1698431365
transform 1 0 46928 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_409
timestamp 1698431365
transform 1 0 47152 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_412
timestamp 1698431365
transform 1 0 47488 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_426
timestamp 1698431365
transform 1 0 49056 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_489
timestamp 1698431365
transform 1 0 56112 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_504
timestamp 1698431365
transform 1 0 57792 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1698431365
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_25
timestamp 1698431365
transform 1 0 4144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_65
timestamp 1698431365
transform 1 0 8624 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_69
timestamp 1698431365
transform 1 0 9072 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_72
timestamp 1698431365
transform 1 0 9408 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_76
timestamp 1698431365
transform 1 0 9856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_78
timestamp 1698431365
transform 1 0 10080 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_94
timestamp 1698431365
transform 1 0 11872 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_98
timestamp 1698431365
transform 1 0 12320 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_109
timestamp 1698431365
transform 1 0 13552 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_119
timestamp 1698431365
transform 1 0 14672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698431365
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_183
timestamp 1698431365
transform 1 0 21840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_191
timestamp 1698431365
transform 1 0 22736 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_195
timestamp 1698431365
transform 1 0 23184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_197
timestamp 1698431365
transform 1 0 23408 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_206
timestamp 1698431365
transform 1 0 24416 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_226
timestamp 1698431365
transform 1 0 26656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_230
timestamp 1698431365
transform 1 0 27104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_232
timestamp 1698431365
transform 1 0 27328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_238
timestamp 1698431365
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_260
timestamp 1698431365
transform 1 0 30464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_264
timestamp 1698431365
transform 1 0 30912 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_306
timestamp 1698431365
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_319
timestamp 1698431365
transform 1 0 37072 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_345
timestamp 1698431365
transform 1 0 39984 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_382
timestamp 1698431365
transform 1 0 44128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_407
timestamp 1698431365
transform 1 0 46928 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_415
timestamp 1698431365
transform 1 0 47824 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_419
timestamp 1698431365
transform 1 0 48272 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_422
timestamp 1698431365
transform 1 0 48608 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_430
timestamp 1698431365
transform 1 0 49504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_432
timestamp 1698431365
transform 1 0 49728 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_454
timestamp 1698431365
transform 1 0 52192 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_502
timestamp 1698431365
transform 1 0 57568 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_506
timestamp 1698431365
transform 1 0 58016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_508
timestamp 1698431365
transform 1 0 58240 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_10
timestamp 1698431365
transform 1 0 2464 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_57
timestamp 1698431365
transform 1 0 7728 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_59
timestamp 1698431365
transform 1 0 7952 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_92
timestamp 1698431365
transform 1 0 11648 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_128
timestamp 1698431365
transform 1 0 15680 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_148
timestamp 1698431365
transform 1 0 17920 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_216
timestamp 1698431365
transform 1 0 25536 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_220
timestamp 1698431365
transform 1 0 25984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_222
timestamp 1698431365
transform 1 0 26208 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_231
timestamp 1698431365
transform 1 0 27216 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_243
timestamp 1698431365
transform 1 0 28560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_251
timestamp 1698431365
transform 1 0 29456 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_274
timestamp 1698431365
transform 1 0 32032 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_278
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_290
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_317
timestamp 1698431365
transform 1 0 36848 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_343
timestamp 1698431365
transform 1 0 39760 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_374
timestamp 1698431365
transform 1 0 43232 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_415
timestamp 1698431365
transform 1 0 47824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_419
timestamp 1698431365
transform 1 0 48272 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_430
timestamp 1698431365
transform 1 0 49504 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_434
timestamp 1698431365
transform 1 0 49952 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_436
timestamp 1698431365
transform 1 0 50176 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_469
timestamp 1698431365
transform 1 0 53872 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_473
timestamp 1698431365
transform 1 0 54320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_477
timestamp 1698431365
transform 1 0 54768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_481
timestamp 1698431365
transform 1 0 55216 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_485
timestamp 1698431365
transform 1 0 55664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_489
timestamp 1698431365
transform 1 0 56112 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_496
timestamp 1698431365
transform 1 0 56896 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_503
timestamp 1698431365
transform 1 0 57680 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_507
timestamp 1698431365
transform 1 0 58128 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_33
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_47
timestamp 1698431365
transform 1 0 6608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_49
timestamp 1698431365
transform 1 0 6832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_89
timestamp 1698431365
transform 1 0 11312 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_93
timestamp 1698431365
transform 1 0 11760 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_115
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_123
timestamp 1698431365
transform 1 0 15120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_154
timestamp 1698431365
transform 1 0 18592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_158
timestamp 1698431365
transform 1 0 19040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_162
timestamp 1698431365
transform 1 0 19488 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_170
timestamp 1698431365
transform 1 0 20384 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698431365
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_187
timestamp 1698431365
transform 1 0 22288 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_195
timestamp 1698431365
transform 1 0 23184 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_202
timestamp 1698431365
transform 1 0 23968 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_218
timestamp 1698431365
transform 1 0 25760 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_230
timestamp 1698431365
transform 1 0 27104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_232
timestamp 1698431365
transform 1 0 27328 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_255
timestamp 1698431365
transform 1 0 29904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_267
timestamp 1698431365
transform 1 0 31248 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_299
timestamp 1698431365
transform 1 0 34832 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_307
timestamp 1698431365
transform 1 0 35728 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_331
timestamp 1698431365
transform 1 0 38416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_335
timestamp 1698431365
transform 1 0 38864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_378
timestamp 1698431365
transform 1 0 43680 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_382
timestamp 1698431365
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_395
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_411
timestamp 1698431365
transform 1 0 47376 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_419
timestamp 1698431365
transform 1 0 48272 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_422
timestamp 1698431365
transform 1 0 48608 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_454
timestamp 1698431365
transform 1 0 52192 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_475
timestamp 1698431365
transform 1 0 54544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_477
timestamp 1698431365
transform 1 0 54768 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_507
timestamp 1698431365
transform 1 0 58128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_10
timestamp 1698431365
transform 1 0 2464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_12
timestamp 1698431365
transform 1 0 2688 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_21
timestamp 1698431365
transform 1 0 3696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_58
timestamp 1698431365
transform 1 0 7840 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_92
timestamp 1698431365
transform 1 0 11648 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_104
timestamp 1698431365
transform 1 0 12992 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_122
timestamp 1698431365
transform 1 0 15008 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_150
timestamp 1698431365
transform 1 0 18144 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_164
timestamp 1698431365
transform 1 0 19712 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_168
timestamp 1698431365
transform 1 0 20160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_178
timestamp 1698431365
transform 1 0 21280 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_198
timestamp 1698431365
transform 1 0 23520 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_202
timestamp 1698431365
transform 1 0 23968 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_220
timestamp 1698431365
transform 1 0 25984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_230
timestamp 1698431365
transform 1 0 27104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_232
timestamp 1698431365
transform 1 0 27328 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_239
timestamp 1698431365
transform 1 0 28112 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_255
timestamp 1698431365
transform 1 0 29904 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_259
timestamp 1698431365
transform 1 0 30352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_261
timestamp 1698431365
transform 1 0 30576 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_268
timestamp 1698431365
transform 1 0 31360 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_272
timestamp 1698431365
transform 1 0 31808 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_290
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_336
timestamp 1698431365
transform 1 0 38976 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_348
timestamp 1698431365
transform 1 0 40320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_356
timestamp 1698431365
transform 1 0 41216 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_358
timestamp 1698431365
transform 1 0 41440 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_367
timestamp 1698431365
transform 1 0 42448 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_369
timestamp 1698431365
transform 1 0 42672 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_401
timestamp 1698431365
transform 1 0 46256 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_409
timestamp 1698431365
transform 1 0 47152 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_418
timestamp 1698431365
transform 1 0 48160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_428
timestamp 1698431365
transform 1 0 49280 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_432
timestamp 1698431365
transform 1 0 49728 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_505
timestamp 1698431365
transform 1 0 57904 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_18
timestamp 1698431365
transform 1 0 3360 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_26
timestamp 1698431365
transform 1 0 4256 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_30
timestamp 1698431365
transform 1 0 4704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_32
timestamp 1698431365
transform 1 0 4928 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_69
timestamp 1698431365
transform 1 0 9072 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_72
timestamp 1698431365
transform 1 0 9408 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_74
timestamp 1698431365
transform 1 0 9632 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_83
timestamp 1698431365
transform 1 0 10640 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_99
timestamp 1698431365
transform 1 0 12432 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_103
timestamp 1698431365
transform 1 0 12880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_134
timestamp 1698431365
transform 1 0 16352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_155
timestamp 1698431365
transform 1 0 18704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_185
timestamp 1698431365
transform 1 0 22064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_251
timestamp 1698431365
transform 1 0 29456 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_259
timestamp 1698431365
transform 1 0 30352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_304
timestamp 1698431365
transform 1 0 35392 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_308
timestamp 1698431365
transform 1 0 35840 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_312
timestamp 1698431365
transform 1 0 36288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_321
timestamp 1698431365
transform 1 0 37296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_333
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_360
timestamp 1698431365
transform 1 0 41664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_364
timestamp 1698431365
transform 1 0 42112 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_370
timestamp 1698431365
transform 1 0 42784 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_377
timestamp 1698431365
transform 1 0 43568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_393
timestamp 1698431365
transform 1 0 45360 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_397
timestamp 1698431365
transform 1 0 45808 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_428
timestamp 1698431365
transform 1 0 49280 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_454
timestamp 1698431365
transform 1 0 52192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_486
timestamp 1698431365
transform 1 0 55776 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_490
timestamp 1698431365
transform 1 0 56224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_492
timestamp 1698431365
transform 1 0 56448 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_506
timestamp 1698431365
transform 1 0 58016 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_508
timestamp 1698431365
transform 1 0 58240 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_34
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_38
timestamp 1698431365
transform 1 0 5600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_40
timestamp 1698431365
transform 1 0 5824 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_74
timestamp 1698431365
transform 1 0 9632 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_134
timestamp 1698431365
transform 1 0 16352 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_138
timestamp 1698431365
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_168
timestamp 1698431365
transform 1 0 20160 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_172
timestamp 1698431365
transform 1 0 20608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_183
timestamp 1698431365
transform 1 0 21840 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_187
timestamp 1698431365
transform 1 0 22288 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_203
timestamp 1698431365
transform 1 0 24080 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_207
timestamp 1698431365
transform 1 0 24528 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_290
timestamp 1698431365
transform 1 0 33824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_292
timestamp 1698431365
transform 1 0 34048 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_301
timestamp 1698431365
transform 1 0 35056 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_317
timestamp 1698431365
transform 1 0 36848 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_338
timestamp 1698431365
transform 1 0 39200 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_349
timestamp 1698431365
transform 1 0 40432 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_356
timestamp 1698431365
transform 1 0 41216 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_380
timestamp 1698431365
transform 1 0 43904 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_388
timestamp 1698431365
transform 1 0 44800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_390
timestamp 1698431365
transform 1 0 45024 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_399
timestamp 1698431365
transform 1 0 46032 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_403
timestamp 1698431365
transform 1 0 46480 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_432
timestamp 1698431365
transform 1 0 49728 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_434
timestamp 1698431365
transform 1 0 49952 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_468
timestamp 1698431365
transform 1 0 53760 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_472
timestamp 1698431365
transform 1 0 54208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_476
timestamp 1698431365
transform 1 0 54656 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_480
timestamp 1698431365
transform 1 0 55104 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_501
timestamp 1698431365
transform 1 0 57456 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_45
timestamp 1698431365
transform 1 0 6384 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_75
timestamp 1698431365
transform 1 0 9744 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_79
timestamp 1698431365
transform 1 0 10192 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_83
timestamp 1698431365
transform 1 0 10640 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_86
timestamp 1698431365
transform 1 0 10976 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_90
timestamp 1698431365
transform 1 0 11424 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_92
timestamp 1698431365
transform 1 0 11648 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_95
timestamp 1698431365
transform 1 0 11984 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_103
timestamp 1698431365
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_115
timestamp 1698431365
transform 1 0 14224 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_123
timestamp 1698431365
transform 1 0 15120 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_131
timestamp 1698431365
transform 1 0 16016 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_136
timestamp 1698431365
transform 1 0 16576 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_159
timestamp 1698431365
transform 1 0 19152 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_192
timestamp 1698431365
transform 1 0 22848 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_194
timestamp 1698431365
transform 1 0 23072 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_226
timestamp 1698431365
transform 1 0 26656 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_234
timestamp 1698431365
transform 1 0 27552 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_238
timestamp 1698431365
transform 1 0 28000 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_242
timestamp 1698431365
transform 1 0 28448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_255
timestamp 1698431365
transform 1 0 29904 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_259
timestamp 1698431365
transform 1 0 30352 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_268
timestamp 1698431365
transform 1 0 31360 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_280
timestamp 1698431365
transform 1 0 32704 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_300
timestamp 1698431365
transform 1 0 34944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_356
timestamp 1698431365
transform 1 0 41216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_360
timestamp 1698431365
transform 1 0 41664 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_364
timestamp 1698431365
transform 1 0 42112 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_393
timestamp 1698431365
transform 1 0 45360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_407
timestamp 1698431365
transform 1 0 46928 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_453
timestamp 1698431365
transform 1 0 52080 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_465
timestamp 1698431365
transform 1 0 53424 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_469
timestamp 1698431365
transform 1 0 53872 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_473
timestamp 1698431365
transform 1 0 54320 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_506
timestamp 1698431365
transform 1 0 58016 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_508
timestamp 1698431365
transform 1 0 58240 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_34
timestamp 1698431365
transform 1 0 5152 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_42
timestamp 1698431365
transform 1 0 6048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_124
timestamp 1698431365
transform 1 0 15232 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_144
timestamp 1698431365
transform 1 0 17472 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_151
timestamp 1698431365
transform 1 0 18256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_159
timestamp 1698431365
transform 1 0 19152 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_163
timestamp 1698431365
transform 1 0 19600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_166
timestamp 1698431365
transform 1 0 19936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_170
timestamp 1698431365
transform 1 0 20384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_172
timestamp 1698431365
transform 1 0 20608 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_228
timestamp 1698431365
transform 1 0 26880 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_248
timestamp 1698431365
transform 1 0 29120 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_262
timestamp 1698431365
transform 1 0 30688 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_278
timestamp 1698431365
transform 1 0 32480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_284
timestamp 1698431365
transform 1 0 33152 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_318
timestamp 1698431365
transform 1 0 36960 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_326
timestamp 1698431365
transform 1 0 37856 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_329
timestamp 1698431365
transform 1 0 38192 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_341
timestamp 1698431365
transform 1 0 39536 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_348
timestamp 1698431365
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_360
timestamp 1698431365
transform 1 0 41664 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_364
timestamp 1698431365
transform 1 0 42112 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_374
timestamp 1698431365
transform 1 0 43232 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_390
timestamp 1698431365
transform 1 0 45024 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_464
timestamp 1698431365
transform 1 0 53312 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_471
timestamp 1698431365
transform 1 0 54096 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_479
timestamp 1698431365
transform 1 0 54992 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_481
timestamp 1698431365
transform 1 0 55216 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_503
timestamp 1698431365
transform 1 0 57680 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_507
timestamp 1698431365
transform 1 0 58128 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_45
timestamp 1698431365
transform 1 0 6384 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_100
timestamp 1698431365
transform 1 0 12544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_115
timestamp 1698431365
transform 1 0 14224 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_119
timestamp 1698431365
transform 1 0 14672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_128
timestamp 1698431365
transform 1 0 15680 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_172
timestamp 1698431365
transform 1 0 20608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_181
timestamp 1698431365
transform 1 0 21616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_183
timestamp 1698431365
transform 1 0 21840 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_190
timestamp 1698431365
transform 1 0 22624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_198
timestamp 1698431365
transform 1 0 23520 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_243
timestamp 1698431365
transform 1 0 28560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_251
timestamp 1698431365
transform 1 0 29456 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_259
timestamp 1698431365
transform 1 0 30352 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_289
timestamp 1698431365
transform 1 0 33712 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_291
timestamp 1698431365
transform 1 0 33936 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_335
timestamp 1698431365
transform 1 0 38864 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_339
timestamp 1698431365
transform 1 0 39312 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_347
timestamp 1698431365
transform 1 0 40208 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_349
timestamp 1698431365
transform 1 0 40432 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_356
timestamp 1698431365
transform 1 0 41216 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_364
timestamp 1698431365
transform 1 0 42112 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_445
timestamp 1698431365
transform 1 0 51184 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_449
timestamp 1698431365
transform 1 0 51632 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_471
timestamp 1698431365
transform 1 0 54096 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_505
timestamp 1698431365
transform 1 0 57904 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_18
timestamp 1698431365
transform 1 0 3360 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_22
timestamp 1698431365
transform 1 0 3808 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_24
timestamp 1698431365
transform 1 0 4032 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_76
timestamp 1698431365
transform 1 0 9856 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_80
timestamp 1698431365
transform 1 0 10304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_84
timestamp 1698431365
transform 1 0 10752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_116
timestamp 1698431365
transform 1 0 14336 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_120
timestamp 1698431365
transform 1 0 14784 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_146
timestamp 1698431365
transform 1 0 17696 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_205
timestamp 1698431365
transform 1 0 24304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_286
timestamp 1698431365
transform 1 0 33376 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_306
timestamp 1698431365
transform 1 0 35616 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_314
timestamp 1698431365
transform 1 0 36512 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_316
timestamp 1698431365
transform 1 0 36736 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_319
timestamp 1698431365
transform 1 0 37072 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_323
timestamp 1698431365
transform 1 0 37520 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_338
timestamp 1698431365
transform 1 0 39200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_342
timestamp 1698431365
transform 1 0 39648 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_358
timestamp 1698431365
transform 1 0 41440 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_362
timestamp 1698431365
transform 1 0 41888 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_379
timestamp 1698431365
transform 1 0 43792 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_395
timestamp 1698431365
transform 1 0 45584 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_397
timestamp 1698431365
transform 1 0 45808 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_400
timestamp 1698431365
transform 1 0 46144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_404
timestamp 1698431365
transform 1 0 46592 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_428
timestamp 1698431365
transform 1 0 49280 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_486
timestamp 1698431365
transform 1 0 55776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_504
timestamp 1698431365
transform 1 0 57792 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698431365
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_18
timestamp 1698431365
transform 1 0 3360 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_26
timestamp 1698431365
transform 1 0 4256 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_28
timestamp 1698431365
transform 1 0 4480 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_41
timestamp 1698431365
transform 1 0 5936 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_100
timestamp 1698431365
transform 1 0 12544 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_111
timestamp 1698431365
transform 1 0 13776 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_149
timestamp 1698431365
transform 1 0 18032 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_153
timestamp 1698431365
transform 1 0 18480 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_164
timestamp 1698431365
transform 1 0 19712 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_168
timestamp 1698431365
transform 1 0 20160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_172
timestamp 1698431365
transform 1 0 20608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_174
timestamp 1698431365
transform 1 0 20832 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_181
timestamp 1698431365
transform 1 0 21616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_185
timestamp 1698431365
transform 1 0 22064 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_201
timestamp 1698431365
transform 1 0 23856 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_209
timestamp 1698431365
transform 1 0 24752 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_211
timestamp 1698431365
transform 1 0 24976 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_220
timestamp 1698431365
transform 1 0 25984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_224
timestamp 1698431365
transform 1 0 26432 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_228
timestamp 1698431365
transform 1 0 26880 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_244
timestamp 1698431365
transform 1 0 28672 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_251
timestamp 1698431365
transform 1 0 29456 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_259
timestamp 1698431365
transform 1 0 30352 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_267
timestamp 1698431365
transform 1 0 31248 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_300
timestamp 1698431365
transform 1 0 34944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_304
timestamp 1698431365
transform 1 0 35392 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_312
timestamp 1698431365
transform 1 0 36288 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_343
timestamp 1698431365
transform 1 0 39760 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_347
timestamp 1698431365
transform 1 0 40208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_351
timestamp 1698431365
transform 1 0 40656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_375
timestamp 1698431365
transform 1 0 43344 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_381
timestamp 1698431365
transform 1 0 44016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_389
timestamp 1698431365
transform 1 0 44912 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_448
timestamp 1698431365
transform 1 0 51520 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_452
timestamp 1698431365
transform 1 0 51968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_454
timestamp 1698431365
transform 1 0 52192 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_463
timestamp 1698431365
transform 1 0 53200 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_475
timestamp 1698431365
transform 1 0 54544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_506
timestamp 1698431365
transform 1 0 58016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_508
timestamp 1698431365
transform 1 0 58240 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_51
timestamp 1698431365
transform 1 0 7056 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_58
timestamp 1698431365
transform 1 0 7840 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_86
timestamp 1698431365
transform 1 0 10976 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_90
timestamp 1698431365
transform 1 0 11424 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_122
timestamp 1698431365
transform 1 0 15008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_126
timestamp 1698431365
transform 1 0 15456 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_134
timestamp 1698431365
transform 1 0 16352 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_138
timestamp 1698431365
transform 1 0 16800 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_174
timestamp 1698431365
transform 1 0 20832 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_176
timestamp 1698431365
transform 1 0 21056 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_208
timestamp 1698431365
transform 1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_241
timestamp 1698431365
transform 1 0 28336 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_245
timestamp 1698431365
transform 1 0 28784 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_261
timestamp 1698431365
transform 1 0 30576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_279
timestamp 1698431365
transform 1 0 32592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_298
timestamp 1698431365
transform 1 0 34720 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_302
timestamp 1698431365
transform 1 0 35168 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_304
timestamp 1698431365
transform 1 0 35392 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_321
timestamp 1698431365
transform 1 0 37296 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_348
timestamp 1698431365
transform 1 0 40320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_381
timestamp 1698431365
transform 1 0 44016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_383
timestamp 1698431365
transform 1 0 44240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_422
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_476
timestamp 1698431365
transform 1 0 54656 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_480
timestamp 1698431365
transform 1 0 55104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_484
timestamp 1698431365
transform 1 0 55552 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_488
timestamp 1698431365
transform 1 0 56000 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_496
timestamp 1698431365
transform 1 0 56896 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_505
timestamp 1698431365
transform 1 0 57904 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_18
timestamp 1698431365
transform 1 0 3360 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_26
timestamp 1698431365
transform 1 0 4256 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_28
timestamp 1698431365
transform 1 0 4480 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_45
timestamp 1698431365
transform 1 0 6384 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_80
timestamp 1698431365
transform 1 0 10304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_82
timestamp 1698431365
transform 1 0 10528 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_123
timestamp 1698431365
transform 1 0 15120 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_127
timestamp 1698431365
transform 1 0 15568 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_163
timestamp 1698431365
transform 1 0 19600 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_191
timestamp 1698431365
transform 1 0 22736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_195
timestamp 1698431365
transform 1 0 23184 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_227
timestamp 1698431365
transform 1 0 26768 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_235
timestamp 1698431365
transform 1 0 27664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_269
timestamp 1698431365
transform 1 0 31472 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_314
timestamp 1698431365
transform 1 0 36512 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_350
timestamp 1698431365
transform 1 0 40544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_377
timestamp 1698431365
transform 1 0 43568 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_404
timestamp 1698431365
transform 1 0 46592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_470
timestamp 1698431365
transform 1 0 53984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_474
timestamp 1698431365
transform 1 0 54432 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_504
timestamp 1698431365
transform 1 0 57792 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_508
timestamp 1698431365
transform 1 0 58240 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_31
timestamp 1698431365
transform 1 0 4816 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_35
timestamp 1698431365
transform 1 0 5264 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_45
timestamp 1698431365
transform 1 0 6384 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_52
timestamp 1698431365
transform 1 0 7168 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_56
timestamp 1698431365
transform 1 0 7616 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_63
timestamp 1698431365
transform 1 0 8400 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_80
timestamp 1698431365
transform 1 0 10304 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_118
timestamp 1698431365
transform 1 0 14560 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_122
timestamp 1698431365
transform 1 0 15008 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_138
timestamp 1698431365
transform 1 0 16800 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_168
timestamp 1698431365
transform 1 0 20160 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_180
timestamp 1698431365
transform 1 0 21504 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_220
timestamp 1698431365
transform 1 0 25984 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_227
timestamp 1698431365
transform 1 0 26768 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_234
timestamp 1698431365
transform 1 0 27552 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_277
timestamp 1698431365
transform 1 0 32368 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698431365
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_298
timestamp 1698431365
transform 1 0 34720 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_376
timestamp 1698431365
transform 1 0 43456 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_426
timestamp 1698431365
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_436
timestamp 1698431365
transform 1 0 50176 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_438
timestamp 1698431365
transform 1 0 50400 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_473
timestamp 1698431365
transform 1 0 54320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_477
timestamp 1698431365
transform 1 0 54768 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_485
timestamp 1698431365
transform 1 0 55664 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_489
timestamp 1698431365
transform 1 0 56112 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_500
timestamp 1698431365
transform 1 0 57344 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698431365
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_10
timestamp 1698431365
transform 1 0 2464 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_17
timestamp 1698431365
transform 1 0 3248 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_24
timestamp 1698431365
transform 1 0 4032 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_32
timestamp 1698431365
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_45
timestamp 1698431365
transform 1 0 6384 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_61
timestamp 1698431365
transform 1 0 8176 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_69
timestamp 1698431365
transform 1 0 9072 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_73
timestamp 1698431365
transform 1 0 9520 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_88
timestamp 1698431365
transform 1 0 11200 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_111
timestamp 1698431365
transform 1 0 13776 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_113
timestamp 1698431365
transform 1 0 14000 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_149
timestamp 1698431365
transform 1 0 18032 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_151
timestamp 1698431365
transform 1 0 18256 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_170
timestamp 1698431365
transform 1 0 20384 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_172
timestamp 1698431365
transform 1 0 20608 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_205
timestamp 1698431365
transform 1 0 24304 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_213
timestamp 1698431365
transform 1 0 25200 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_215
timestamp 1698431365
transform 1 0 25424 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_244
timestamp 1698431365
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_284
timestamp 1698431365
transform 1 0 33152 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_300
timestamp 1698431365
transform 1 0 34944 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_343
timestamp 1698431365
transform 1 0 39760 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_376
timestamp 1698431365
transform 1 0 43456 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_447
timestamp 1698431365
transform 1 0 51408 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_504
timestamp 1698431365
transform 1 0 57792 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_508
timestamp 1698431365
transform 1 0 58240 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_23
timestamp 1698431365
transform 1 0 3920 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_27
timestamp 1698431365
transform 1 0 4368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_29
timestamp 1698431365
transform 1 0 4592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_58
timestamp 1698431365
transform 1 0 7840 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1698431365
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_77
timestamp 1698431365
transform 1 0 9968 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_81
timestamp 1698431365
transform 1 0 10416 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_88
timestamp 1698431365
transform 1 0 11200 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_105
timestamp 1698431365
transform 1 0 13104 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_121
timestamp 1698431365
transform 1 0 14896 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_129
timestamp 1698431365
transform 1 0 15792 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_133
timestamp 1698431365
transform 1 0 16240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_150
timestamp 1698431365
transform 1 0 18144 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_152
timestamp 1698431365
transform 1 0 18368 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_169
timestamp 1698431365
transform 1 0 20272 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_171
timestamp 1698431365
transform 1 0 20496 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_191
timestamp 1698431365
transform 1 0 22736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_195
timestamp 1698431365
transform 1 0 23184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_248
timestamp 1698431365
transform 1 0 29120 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_298
timestamp 1698431365
transform 1 0 34720 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_306
timestamp 1698431365
transform 1 0 35616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_310
timestamp 1698431365
transform 1 0 36064 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_340
timestamp 1698431365
transform 1 0 39424 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_366
timestamp 1698431365
transform 1 0 42336 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_389
timestamp 1698431365
transform 1 0 44912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_413
timestamp 1698431365
transform 1 0 47600 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_438
timestamp 1698431365
transform 1 0 50400 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_440
timestamp 1698431365
transform 1 0 50624 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_453
timestamp 1698431365
transform 1 0 52080 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_455
timestamp 1698431365
transform 1 0 52304 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_487
timestamp 1698431365
transform 1 0 55888 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_489
timestamp 1698431365
transform 1 0 56112 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_497
timestamp 1698431365
transform 1 0 57008 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_505
timestamp 1698431365
transform 1 0 57904 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_31
timestamp 1698431365
transform 1 0 4816 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_68
timestamp 1698431365
transform 1 0 8960 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_72
timestamp 1698431365
transform 1 0 9408 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_80
timestamp 1698431365
transform 1 0 10304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_82
timestamp 1698431365
transform 1 0 10528 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_123
timestamp 1698431365
transform 1 0 15120 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_127
timestamp 1698431365
transform 1 0 15568 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_129
timestamp 1698431365
transform 1 0 15792 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_148
timestamp 1698431365
transform 1 0 17920 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_152
timestamp 1698431365
transform 1 0 18368 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_154
timestamp 1698431365
transform 1 0 18592 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_172
timestamp 1698431365
transform 1 0 20608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_174
timestamp 1698431365
transform 1 0 20832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_183
timestamp 1698431365
transform 1 0 21840 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_185
timestamp 1698431365
transform 1 0 22064 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_194
timestamp 1698431365
transform 1 0 23072 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_198
timestamp 1698431365
transform 1 0 23520 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_209
timestamp 1698431365
transform 1 0 24752 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_235
timestamp 1698431365
transform 1 0 27664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_321
timestamp 1698431365
transform 1 0 37296 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_338
timestamp 1698431365
transform 1 0 39200 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698431365
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_448
timestamp 1698431365
transform 1 0 51520 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_452
timestamp 1698431365
transform 1 0 51968 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_454
timestamp 1698431365
transform 1 0 52192 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_467
timestamp 1698431365
transform 1 0 53648 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_485
timestamp 1698431365
transform 1 0 55664 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_501
timestamp 1698431365
transform 1 0 57456 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_18
timestamp 1698431365
transform 1 0 3360 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_26
timestamp 1698431365
transform 1 0 4256 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_36
timestamp 1698431365
transform 1 0 5376 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_45
timestamp 1698431365
transform 1 0 6384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_54
timestamp 1698431365
transform 1 0 7392 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_74
timestamp 1698431365
transform 1 0 9632 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_101
timestamp 1698431365
transform 1 0 12656 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_103
timestamp 1698431365
transform 1 0 12880 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_133
timestamp 1698431365
transform 1 0 16240 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_154
timestamp 1698431365
transform 1 0 18592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_187
timestamp 1698431365
transform 1 0 22288 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_191
timestamp 1698431365
transform 1 0 22736 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_193
timestamp 1698431365
transform 1 0 22960 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_204
timestamp 1698431365
transform 1 0 24192 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_208
timestamp 1698431365
transform 1 0 24640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_219
timestamp 1698431365
transform 1 0 25872 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_221
timestamp 1698431365
transform 1 0 26096 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_242
timestamp 1698431365
transform 1 0 28448 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_249
timestamp 1698431365
transform 1 0 29232 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_265
timestamp 1698431365
transform 1 0 31024 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_269
timestamp 1698431365
transform 1 0 31472 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_287
timestamp 1698431365
transform 1 0 33488 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_295
timestamp 1698431365
transform 1 0 34384 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_303
timestamp 1698431365
transform 1 0 35280 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_335
timestamp 1698431365
transform 1 0 38864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_357
timestamp 1698431365
transform 1 0 41328 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_368
timestamp 1698431365
transform 1 0 42560 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_413
timestamp 1698431365
transform 1 0 47600 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_417
timestamp 1698431365
transform 1 0 48048 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_419
timestamp 1698431365
transform 1 0 48272 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_432
timestamp 1698431365
transform 1 0 49728 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_446
timestamp 1698431365
transform 1 0 51296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_459
timestamp 1698431365
transform 1 0 52752 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_471
timestamp 1698431365
transform 1 0 54096 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_487
timestamp 1698431365
transform 1 0 55888 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_489
timestamp 1698431365
transform 1 0 56112 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698431365
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_31
timestamp 1698431365
transform 1 0 4816 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_47
timestamp 1698431365
transform 1 0 6608 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_60
timestamp 1698431365
transform 1 0 8064 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_99
timestamp 1698431365
transform 1 0 12432 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_103
timestamp 1698431365
transform 1 0 12880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_123
timestamp 1698431365
transform 1 0 15120 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_138
timestamp 1698431365
transform 1 0 16800 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_155
timestamp 1698431365
transform 1 0 18704 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_159
timestamp 1698431365
transform 1 0 19152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_166
timestamp 1698431365
transform 1 0 19936 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_174
timestamp 1698431365
transform 1 0 20832 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_194
timestamp 1698431365
transform 1 0 23072 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_198
timestamp 1698431365
transform 1 0 23520 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_213
timestamp 1698431365
transform 1 0 25200 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_217
timestamp 1698431365
transform 1 0 25648 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_240
timestamp 1698431365
transform 1 0 28224 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_244
timestamp 1698431365
transform 1 0 28672 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_261
timestamp 1698431365
transform 1 0 30576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_277
timestamp 1698431365
transform 1 0 32368 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_281
timestamp 1698431365
transform 1 0 32816 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_283
timestamp 1698431365
transform 1 0 33040 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_302
timestamp 1698431365
transform 1 0 35168 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_310
timestamp 1698431365
transform 1 0 36064 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_314
timestamp 1698431365
transform 1 0 36512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_325
timestamp 1698431365
transform 1 0 37744 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_329
timestamp 1698431365
transform 1 0 38192 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_350
timestamp 1698431365
transform 1 0 40544 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_371
timestamp 1698431365
transform 1 0 42896 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_375
timestamp 1698431365
transform 1 0 43344 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_399
timestamp 1698431365
transform 1 0 46032 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_435
timestamp 1698431365
transform 1 0 50064 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_437
timestamp 1698431365
transform 1 0 50288 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_452
timestamp 1698431365
transform 1 0 51968 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_454
timestamp 1698431365
transform 1 0 52192 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_461
timestamp 1698431365
transform 1 0 52976 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_493
timestamp 1698431365
transform 1 0 56560 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_10
timestamp 1698431365
transform 1 0 2464 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_14
timestamp 1698431365
transform 1 0 2912 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_21
timestamp 1698431365
transform 1 0 3696 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_29
timestamp 1698431365
transform 1 0 4592 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_57
timestamp 1698431365
transform 1 0 7728 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_65
timestamp 1698431365
transform 1 0 8624 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_69
timestamp 1698431365
transform 1 0 9072 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_76
timestamp 1698431365
transform 1 0 9856 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_97
timestamp 1698431365
transform 1 0 12208 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_107
timestamp 1698431365
transform 1 0 13328 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_123
timestamp 1698431365
transform 1 0 15120 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_127
timestamp 1698431365
transform 1 0 15568 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_138
timestamp 1698431365
transform 1 0 16800 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_144
timestamp 1698431365
transform 1 0 17472 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_186
timestamp 1698431365
transform 1 0 22176 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_190
timestamp 1698431365
transform 1 0 22624 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_228
timestamp 1698431365
transform 1 0 26880 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_232
timestamp 1698431365
transform 1 0 27328 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_234
timestamp 1698431365
transform 1 0 27552 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_269
timestamp 1698431365
transform 1 0 31472 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_277
timestamp 1698431365
transform 1 0 32368 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_279
timestamp 1698431365
transform 1 0 32592 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_311
timestamp 1698431365
transform 1 0 36176 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_327
timestamp 1698431365
transform 1 0 37968 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_331
timestamp 1698431365
transform 1 0 38416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_333
timestamp 1698431365
transform 1 0 38640 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_342
timestamp 1698431365
transform 1 0 39648 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_346
timestamp 1698431365
transform 1 0 40096 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_354
timestamp 1698431365
transform 1 0 40992 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_366
timestamp 1698431365
transform 1 0 42336 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_391
timestamp 1698431365
transform 1 0 45136 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_407
timestamp 1698431365
transform 1 0 46928 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_410
timestamp 1698431365
transform 1 0 47264 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_430
timestamp 1698431365
transform 1 0 49504 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_438
timestamp 1698431365
transform 1 0 50400 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_440
timestamp 1698431365
transform 1 0 50624 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_470
timestamp 1698431365
transform 1 0 53984 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_486
timestamp 1698431365
transform 1 0 55776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_508
timestamp 1698431365
transform 1 0 58240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_6
timestamp 1698431365
transform 1 0 2016 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_26
timestamp 1698431365
transform 1 0 4256 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_39
timestamp 1698431365
transform 1 0 5712 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_69
timestamp 1698431365
transform 1 0 9072 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_73
timestamp 1698431365
transform 1 0 9520 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_75
timestamp 1698431365
transform 1 0 9744 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_142
timestamp 1698431365
transform 1 0 17248 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_144
timestamp 1698431365
transform 1 0 17472 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_153
timestamp 1698431365
transform 1 0 18480 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_161
timestamp 1698431365
transform 1 0 19376 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_163
timestamp 1698431365
transform 1 0 19600 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_168
timestamp 1698431365
transform 1 0 20160 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_172
timestamp 1698431365
transform 1 0 20608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_174
timestamp 1698431365
transform 1 0 20832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_185
timestamp 1698431365
transform 1 0 22064 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_189
timestamp 1698431365
transform 1 0 22512 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_212
timestamp 1698431365
transform 1 0 25088 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_228
timestamp 1698431365
transform 1 0 26880 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_233
timestamp 1698431365
transform 1 0 27440 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_263
timestamp 1698431365
transform 1 0 30800 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_300
timestamp 1698431365
transform 1 0 34944 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_304
timestamp 1698431365
transform 1 0 35392 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698431365
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_321
timestamp 1698431365
transform 1 0 37296 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_329
timestamp 1698431365
transform 1 0 38192 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_362
timestamp 1698431365
transform 1 0 41888 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_364
timestamp 1698431365
transform 1 0 42112 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_373
timestamp 1698431365
transform 1 0 43120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_377
timestamp 1698431365
transform 1 0 43568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_381
timestamp 1698431365
transform 1 0 44016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_445
timestamp 1698431365
transform 1 0 51184 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_449
timestamp 1698431365
transform 1 0 51632 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_453
timestamp 1698431365
transform 1 0 52080 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_489
timestamp 1698431365
transform 1 0 56112 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_505
timestamp 1698431365
transform 1 0 57904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_31
timestamp 1698431365
transform 1 0 4816 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_56
timestamp 1698431365
transform 1 0 7616 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_64
timestamp 1698431365
transform 1 0 8512 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_68
timestamp 1698431365
transform 1 0 8960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_80
timestamp 1698431365
transform 1 0 10304 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_86
timestamp 1698431365
transform 1 0 10976 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_118
timestamp 1698431365
transform 1 0 14560 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_122
timestamp 1698431365
transform 1 0 15008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_124
timestamp 1698431365
transform 1 0 15232 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_127
timestamp 1698431365
transform 1 0 15568 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_131
timestamp 1698431365
transform 1 0 16016 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_155
timestamp 1698431365
transform 1 0 18704 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_182
timestamp 1698431365
transform 1 0 21728 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_186
timestamp 1698431365
transform 1 0 22176 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_206
timestamp 1698431365
transform 1 0 24416 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_218
timestamp 1698431365
transform 1 0 25760 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_220
timestamp 1698431365
transform 1 0 25984 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_231
timestamp 1698431365
transform 1 0 27216 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_286
timestamp 1698431365
transform 1 0 33376 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_302
timestamp 1698431365
transform 1 0 35168 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_304
timestamp 1698431365
transform 1 0 35392 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_342
timestamp 1698431365
transform 1 0 39648 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_410
timestamp 1698431365
transform 1 0 47264 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_418
timestamp 1698431365
transform 1 0 48160 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698431365
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_39
timestamp 1698431365
transform 1 0 5712 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_46
timestamp 1698431365
transform 1 0 6496 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_62
timestamp 1698431365
transform 1 0 8288 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_64
timestamp 1698431365
transform 1 0 8512 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_94
timestamp 1698431365
transform 1 0 11872 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_102
timestamp 1698431365
transform 1 0 12768 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_104
timestamp 1698431365
transform 1 0 12992 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_112
timestamp 1698431365
transform 1 0 13888 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_116
timestamp 1698431365
transform 1 0 14336 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_210
timestamp 1698431365
transform 1 0 24864 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_261
timestamp 1698431365
transform 1 0 30576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_306
timestamp 1698431365
transform 1 0 35616 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_314
timestamp 1698431365
transform 1 0 36512 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_356
timestamp 1698431365
transform 1 0 41216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_372
timestamp 1698431365
transform 1 0 43008 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_380
timestamp 1698431365
transform 1 0 43904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_384
timestamp 1698431365
transform 1 0 44352 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_451
timestamp 1698431365
transform 1 0 51856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_489
timestamp 1698431365
transform 1 0 56112 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_505
timestamp 1698431365
transform 1 0 57904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_18
timestamp 1698431365
transform 1 0 3360 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_26
timestamp 1698431365
transform 1 0 4256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_46
timestamp 1698431365
transform 1 0 6496 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_48
timestamp 1698431365
transform 1 0 6720 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_57
timestamp 1698431365
transform 1 0 7728 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_59
timestamp 1698431365
transform 1 0 7952 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_81
timestamp 1698431365
transform 1 0 10416 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_104
timestamp 1698431365
transform 1 0 12992 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_132
timestamp 1698431365
transform 1 0 16128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_140
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_167
timestamp 1698431365
transform 1 0 20048 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_169
timestamp 1698431365
transform 1 0 20272 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_235
timestamp 1698431365
transform 1 0 27664 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_237
timestamp 1698431365
transform 1 0 27888 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_240
timestamp 1698431365
transform 1 0 28224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_242
timestamp 1698431365
transform 1 0 28448 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_267
timestamp 1698431365
transform 1 0 31248 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_271
timestamp 1698431365
transform 1 0 31696 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_284
timestamp 1698431365
transform 1 0 33152 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_318
timestamp 1698431365
transform 1 0 36960 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_332
timestamp 1698431365
transform 1 0 38528 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_372
timestamp 1698431365
transform 1 0 43008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_384
timestamp 1698431365
transform 1 0 44352 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_393
timestamp 1698431365
transform 1 0 45360 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_405
timestamp 1698431365
transform 1 0 46704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_407
timestamp 1698431365
transform 1 0 46928 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_418
timestamp 1698431365
transform 1 0 48160 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_420
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_429
timestamp 1698431365
transform 1 0 49392 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_441
timestamp 1698431365
transform 1 0 50736 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_444
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_453
timestamp 1698431365
transform 1 0 52080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_465
timestamp 1698431365
transform 1 0 53424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_473
timestamp 1698431365
transform 1 0 54320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_475
timestamp 1698431365
transform 1 0 54544 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_490
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_506
timestamp 1698431365
transform 1 0 58016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1698431365
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input1
timestamp 1698431365
transform 1 0 19712 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 21280 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 41888 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 41888 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input5
timestamp 1698431365
transform 1 0 15232 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 14560 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output8 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21056 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output9 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24416 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output10
timestamp 1698431365
transform 1 0 22624 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output11
timestamp 1698431365
transform 1 0 26096 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output12
timestamp 1698431365
transform -1 0 30576 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output13
timestamp 1698431365
transform 1 0 28560 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output14
timestamp 1698431365
transform 1 0 30128 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output15
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output16
timestamp 1698431365
transform 1 0 34048 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output17
timestamp 1698431365
transform 1 0 34496 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output18
timestamp 1698431365
transform 1 0 35840 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output19
timestamp 1698431365
transform 1 0 37408 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output20
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output21
timestamp 1698431365
transform 1 0 40096 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_153
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_154
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_155
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_159
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_160
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_161
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_162
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_164
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_165
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_166
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_167
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_168
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_169
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_171
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_172
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_173
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_174
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_175
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_176
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_178
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_179
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_180
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_181
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_182
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_183
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_185
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_186
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_187
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_188
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_189
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_190
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_192
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_193
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_194
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_195
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_196
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_197
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_199
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_200
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_201
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_202
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_203
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_204
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_206
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_207
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_208
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_209
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_210
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_211
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_213
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_214
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_215
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_216
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_217
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_218
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_220
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_221
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_222
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_223
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_224
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_225
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_227
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_228
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_229
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_230
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_231
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_232
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_234
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_235
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_236
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_237
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_238
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_239
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_241
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_242
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_243
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_244
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_245
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_246
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_248
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_249
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_250
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_251
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_252
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_253
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_258
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_259
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_260
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_267
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_276
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_283
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_284
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_285
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_290
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_291
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_292
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_293
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_294
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_295
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_297
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_298
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_299
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_300
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_301
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_302
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_304
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_305
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_306
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_307
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_308
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_309
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_311
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_312
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_313
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_314
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_315
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_316
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_318
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_319
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_320
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_321
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_322
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_323
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_325
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_326
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_327
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_328
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_329
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_330
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_332
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_333
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_334
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_335
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_336
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_337
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_339
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_340
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_341
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_342
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_343
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_344
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_346
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_347
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_348
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_349
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_350
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_351
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_353
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_354
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_355
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_356
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_357
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_358
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_360
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_361
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_362
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_363
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_364
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_367
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_368
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_369
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_374
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_375
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_392
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_393
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_398
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_399
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_403
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_404
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_405
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_409
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_410
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_416
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_428
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_433
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_434
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_448
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_449
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_453
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_454
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_455
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_456
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_458
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_459
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_460
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_461
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_462
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_463
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_465
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_466
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_467
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_468
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_469
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_470
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_472
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_473
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_474
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_475
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_476
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_477
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_479
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_480
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_481
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_482
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_483
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_484
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_486
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_487
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_488
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_489
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_490
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_491
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_493
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_494
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_495
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_496
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_497
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_498
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_500
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_501
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_502
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_503
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_504
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_505
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_507
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_508
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_509
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_510
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_511
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_512
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_514
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_515
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_516
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_517
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_518
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_519
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_521
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_522
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_523
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_524
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_525
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_526
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_528
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_529
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_530
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_531
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_532
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_533
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_535
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_536
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_537
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_538
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_539
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_540
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_542
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_543
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_544
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_545
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_546
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_547
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_549
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_550
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_551
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_552
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_553
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_554
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_556
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_557
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_558
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_559
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_560
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_561
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_563
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_564
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_565
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_566
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_567
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_568
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_570
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_571
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_572
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_573
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_574
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_575
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_577
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_578
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_579
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_580
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_581
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_582
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_584
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_585
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_586
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_587
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_588
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_589
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_591
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_592
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_593
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_594
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_595
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_596
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_598
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_599
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_600
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_601
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_602
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_603
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_605
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_606
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_607
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_608
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_609
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_610
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_612
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_613
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_614
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_615
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_616
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_617
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_625
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_22 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_23
timestamp 1698431365
transform -1 0 23296 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_24
timestamp 1698431365
transform -1 0 24864 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_25
timestamp 1698431365
transform 1 0 25088 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_26
timestamp 1698431365
transform -1 0 27440 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_27
timestamp 1698431365
transform -1 0 28784 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_28
timestamp 1698431365
transform 1 0 28336 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_29
timestamp 1698431365
transform -1 0 31248 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_30
timestamp 1698431365
transform -1 0 33376 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_31
timestamp 1698431365
transform -1 0 35616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_32
timestamp 1698431365
transform -1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_33
timestamp 1698431365
transform -1 0 39424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_34
timestamp 1698431365
transform -1 0 39200 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_35
timestamp 1698431365
transform -1 0 39648 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_36
timestamp 1698431365
transform -1 0 6496 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_37
timestamp 1698431365
transform -1 0 7728 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_38
timestamp 1698431365
transform -1 0 8960 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_39
timestamp 1698431365
transform -1 0 10416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_40
timestamp 1698431365
transform 1 0 10976 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_41
timestamp 1698431365
transform 1 0 11872 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_42
timestamp 1698431365
transform 1 0 13440 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_43
timestamp 1698431365
transform 1 0 14784 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_44
timestamp 1698431365
transform 1 0 14112 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_45
timestamp 1698431365
transform -1 0 18480 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_46
timestamp 1698431365
transform -1 0 20160 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_47
timestamp 1698431365
transform -1 0 20944 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_48
timestamp 1698431365
transform -1 0 42112 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_49
timestamp 1698431365
transform -1 0 43008 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_50
timestamp 1698431365
transform -1 0 44352 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_51
timestamp 1698431365
transform -1 0 45360 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_52
timestamp 1698431365
transform -1 0 46704 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_53
timestamp 1698431365
transform -1 0 48160 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_54
timestamp 1698431365
transform -1 0 49392 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_55
timestamp 1698431365
transform -1 0 50736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_56
timestamp 1698431365
transform -1 0 52080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_57
timestamp 1698431365
transform -1 0 53424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_58
timestamp 1698431365
transform -1 0 55328 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_59
timestamp 1698431365
transform -1 0 56224 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_60 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_61
timestamp 1698431365
transform -1 0 7280 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_62
timestamp 1698431365
transform -1 0 8512 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_63
timestamp 1698431365
transform -1 0 9968 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_64
timestamp 1698431365
transform 1 0 10528 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_65
timestamp 1698431365
transform 1 0 11424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_66
timestamp 1698431365
transform 1 0 12320 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_67
timestamp 1698431365
transform 1 0 13216 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_68
timestamp 1698431365
transform 1 0 13664 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_69
timestamp 1698431365
transform -1 0 18032 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_70
timestamp 1698431365
transform -1 0 19376 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_71
timestamp 1698431365
transform -1 0 21056 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_72
timestamp 1698431365
transform -1 0 43008 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_73
timestamp 1698431365
transform -1 0 42560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_74
timestamp 1698431365
transform -1 0 43904 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_75
timestamp 1698431365
transform -1 0 44912 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_76
timestamp 1698431365
transform -1 0 46256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_77
timestamp 1698431365
transform -1 0 47712 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_78
timestamp 1698431365
transform -1 0 48944 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_79
timestamp 1698431365
transform -1 0 50288 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_80
timestamp 1698431365
transform -1 0 51632 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_81
timestamp 1698431365
transform -1 0 52976 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_82
timestamp 1698431365
transform -1 0 54320 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_83
timestamp 1698431365
transform -1 0 55776 0 -1 56448
box -86 -86 534 870
<< labels >>
flabel metal2 s 4928 59200 5040 60000 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 18368 59200 18480 60000 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 19712 59200 19824 60000 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 21056 59200 21168 60000 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 22400 59200 22512 60000 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 23744 59200 23856 60000 0 FreeSans 448 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 25088 59200 25200 60000 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 26432 59200 26544 60000 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 27776 59200 27888 60000 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 29120 59200 29232 60000 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 30464 59200 30576 60000 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 6272 59200 6384 60000 0 FreeSans 448 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 31808 59200 31920 60000 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 33152 59200 33264 60000 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 34496 59200 34608 60000 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 35840 59200 35952 60000 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 37184 59200 37296 60000 0 FreeSans 448 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 38528 59200 38640 60000 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 39872 59200 39984 60000 0 FreeSans 448 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 41216 59200 41328 60000 0 FreeSans 448 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 42560 59200 42672 60000 0 FreeSans 448 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 43904 59200 44016 60000 0 FreeSans 448 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 7616 59200 7728 60000 0 FreeSans 448 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 45248 59200 45360 60000 0 FreeSans 448 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 46592 59200 46704 60000 0 FreeSans 448 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 47936 59200 48048 60000 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 49280 59200 49392 60000 0 FreeSans 448 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 50624 59200 50736 60000 0 FreeSans 448 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 51968 59200 52080 60000 0 FreeSans 448 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 53312 59200 53424 60000 0 FreeSans 448 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 54656 59200 54768 60000 0 FreeSans 448 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 8960 59200 9072 60000 0 FreeSans 448 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 10304 59200 10416 60000 0 FreeSans 448 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 11648 59200 11760 60000 0 FreeSans 448 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 12992 59200 13104 60000 0 FreeSans 448 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 14336 59200 14448 60000 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 15680 59200 15792 60000 0 FreeSans 448 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 17024 59200 17136 60000 0 FreeSans 448 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 5376 59200 5488 60000 0 FreeSans 448 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 18816 59200 18928 60000 0 FreeSans 448 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 20160 59200 20272 60000 0 FreeSans 448 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 21504 59200 21616 60000 0 FreeSans 448 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 22848 59200 22960 60000 0 FreeSans 448 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 24192 59200 24304 60000 0 FreeSans 448 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 25536 59200 25648 60000 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 26880 59200 26992 60000 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 28224 59200 28336 60000 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 29568 59200 29680 60000 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 30912 59200 31024 60000 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 6720 59200 6832 60000 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 32256 59200 32368 60000 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 33600 59200 33712 60000 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 34944 59200 35056 60000 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 36288 59200 36400 60000 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 37632 59200 37744 60000 0 FreeSans 448 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 38976 59200 39088 60000 0 FreeSans 448 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 40320 59200 40432 60000 0 FreeSans 448 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 41664 59200 41776 60000 0 FreeSans 448 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 43008 59200 43120 60000 0 FreeSans 448 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 44352 59200 44464 60000 0 FreeSans 448 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 8064 59200 8176 60000 0 FreeSans 448 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 45696 59200 45808 60000 0 FreeSans 448 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 47040 59200 47152 60000 0 FreeSans 448 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 48384 59200 48496 60000 0 FreeSans 448 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 49728 59200 49840 60000 0 FreeSans 448 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 51072 59200 51184 60000 0 FreeSans 448 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 52416 59200 52528 60000 0 FreeSans 448 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 53760 59200 53872 60000 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 55104 59200 55216 60000 0 FreeSans 448 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 9408 59200 9520 60000 0 FreeSans 448 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 10752 59200 10864 60000 0 FreeSans 448 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 12096 59200 12208 60000 0 FreeSans 448 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 13440 59200 13552 60000 0 FreeSans 448 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 14784 59200 14896 60000 0 FreeSans 448 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 16128 59200 16240 60000 0 FreeSans 448 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 17472 59200 17584 60000 0 FreeSans 448 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 5824 59200 5936 60000 0 FreeSans 448 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 19264 59200 19376 60000 0 FreeSans 448 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 20608 59200 20720 60000 0 FreeSans 448 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 21952 59200 22064 60000 0 FreeSans 448 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 23296 59200 23408 60000 0 FreeSans 448 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 24640 59200 24752 60000 0 FreeSans 448 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 25984 59200 26096 60000 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 27328 59200 27440 60000 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 28672 59200 28784 60000 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 30016 59200 30128 60000 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 31360 59200 31472 60000 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 7168 59200 7280 60000 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 32704 59200 32816 60000 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 34048 59200 34160 60000 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 35392 59200 35504 60000 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 36736 59200 36848 60000 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 38080 59200 38192 60000 0 FreeSans 448 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 39424 59200 39536 60000 0 FreeSans 448 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 40768 59200 40880 60000 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 42112 59200 42224 60000 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 43456 59200 43568 60000 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 44800 59200 44912 60000 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 8512 59200 8624 60000 0 FreeSans 448 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 46144 59200 46256 60000 0 FreeSans 448 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 47488 59200 47600 60000 0 FreeSans 448 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 48832 59200 48944 60000 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 50176 59200 50288 60000 0 FreeSans 448 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 51520 59200 51632 60000 0 FreeSans 448 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 52864 59200 52976 60000 0 FreeSans 448 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 54208 59200 54320 60000 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 55552 59200 55664 60000 0 FreeSans 448 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 9856 59200 9968 60000 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 11200 59200 11312 60000 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 12544 59200 12656 60000 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 13888 59200 14000 60000 0 FreeSans 448 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 15232 59200 15344 60000 0 FreeSans 448 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 16576 59200 16688 60000 0 FreeSans 448 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 17920 59200 18032 60000 0 FreeSans 448 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 114 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 114 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 115 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 115 nsew ground bidirectional
flabel metal2 s 4032 59200 4144 60000 0 FreeSans 448 90 0 0 wb_clk_i
port 116 nsew signal input
flabel metal2 s 4480 59200 4592 60000 0 FreeSans 448 90 0 0 wb_rst_i
port 117 nsew signal input
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal3 25368 17248 25368 17248 0 _0000_
rlabel metal2 24024 18256 24024 18256 0 _0001_
rlabel metal2 8568 13160 8568 13160 0 _0002_
rlabel metal3 19880 15456 19880 15456 0 _0003_
rlabel metal2 27832 18872 27832 18872 0 _0004_
rlabel metal2 5768 31304 5768 31304 0 _0005_
rlabel metal2 9016 30520 9016 30520 0 _0006_
rlabel metal2 8568 32480 8568 32480 0 _0007_
rlabel metal2 18200 28280 18200 28280 0 _0008_
rlabel metal2 15456 35560 15456 35560 0 _0009_
rlabel metal2 22792 28000 22792 28000 0 _0010_
rlabel metal2 6888 29904 6888 29904 0 _0011_
rlabel metal2 16072 34552 16072 34552 0 _0012_
rlabel metal2 36960 53704 36960 53704 0 _0013_
rlabel metal3 37464 53816 37464 53816 0 _0014_
rlabel metal2 42112 10808 42112 10808 0 _0015_
rlabel metal2 41720 14784 41720 14784 0 _0016_
rlabel metal3 44968 12824 44968 12824 0 _0017_
rlabel metal2 44184 14560 44184 14560 0 _0018_
rlabel metal2 13496 17920 13496 17920 0 _0019_
rlabel metal2 13496 15624 13496 15624 0 _0020_
rlabel metal2 38808 10808 38808 10808 0 _0021_
rlabel metal2 40040 15008 40040 15008 0 _0022_
rlabel metal3 40824 9912 40824 9912 0 _0023_
rlabel metal3 40096 6552 40096 6552 0 _0024_
rlabel metal3 40824 18312 40824 18312 0 _0025_
rlabel metal3 39816 17752 39816 17752 0 _0026_
rlabel metal2 37352 4816 37352 4816 0 _0027_
rlabel metal2 34776 3808 34776 3808 0 _0028_
rlabel metal2 31752 22848 31752 22848 0 _0029_
rlabel metal3 33208 24808 33208 24808 0 _0030_
rlabel metal2 21896 54544 21896 54544 0 _0031_
rlabel metal2 30968 8512 30968 8512 0 _0032_
rlabel metal2 30968 6944 30968 6944 0 _0033_
rlabel metal2 40264 22008 40264 22008 0 _0034_
rlabel metal2 40712 20888 40712 20888 0 _0035_
rlabel metal2 29960 5208 29960 5208 0 _0036_
rlabel metal2 30408 5208 30408 5208 0 _0037_
rlabel metal2 25592 6328 25592 6328 0 _0038_
rlabel metal2 27048 3808 27048 3808 0 _0039_
rlabel metal2 11368 10080 11368 10080 0 _0040_
rlabel metal2 13496 6944 13496 6944 0 _0041_
rlabel metal2 22120 26040 22120 26040 0 _0042_
rlabel metal2 6776 19992 6776 19992 0 _0043_
rlabel metal2 6440 17192 6440 17192 0 _0044_
rlabel metal2 6832 15400 6832 15400 0 _0045_
rlabel metal2 26040 26628 26040 26628 0 _0046_
rlabel metal2 15400 42896 15400 42896 0 _0047_
rlabel metal3 22736 46760 22736 46760 0 _0048_
rlabel metal2 22568 48384 22568 48384 0 _0049_
rlabel metal2 17304 48216 17304 48216 0 _0050_
rlabel metal2 19152 51240 19152 51240 0 _0051_
rlabel metal2 15064 48608 15064 48608 0 _0052_
rlabel metal2 14280 53368 14280 53368 0 _0053_
rlabel metal2 19824 52360 19824 52360 0 _0054_
rlabel metal2 13944 50792 13944 50792 0 _0055_
rlabel metal2 36792 26628 36792 26628 0 _0056_
rlabel metal2 41608 26152 41608 26152 0 _0057_
rlabel metal2 43400 29736 43400 29736 0 _0058_
rlabel metal2 43288 31752 43288 31752 0 _0059_
rlabel metal2 46872 38976 46872 38976 0 _0060_
rlabel metal2 44632 33264 44632 33264 0 _0061_
rlabel metal3 42112 38136 42112 38136 0 _0062_
rlabel metal2 36568 40712 36568 40712 0 _0063_
rlabel metal2 33544 40824 33544 40824 0 _0064_
rlabel metal3 34328 44408 34328 44408 0 _0065_
rlabel metal2 32648 46032 32648 46032 0 _0066_
rlabel metal2 34216 47152 34216 47152 0 _0067_
rlabel metal2 39928 52584 39928 52584 0 _0068_
rlabel metal2 41496 53760 41496 53760 0 _0069_
rlabel metal3 44912 48440 44912 48440 0 _0070_
rlabel metal2 45752 48944 45752 48944 0 _0071_
rlabel metal3 48496 53144 48496 53144 0 _0072_
rlabel metal2 50792 52528 50792 52528 0 _0073_
rlabel metal3 53984 48888 53984 48888 0 _0074_
rlabel metal2 52136 46984 52136 46984 0 _0075_
rlabel metal2 54488 45696 54488 45696 0 _0076_
rlabel metal2 55720 43064 55720 43064 0 _0077_
rlabel metal2 47992 40656 47992 40656 0 _0078_
rlabel metal2 53480 41328 53480 41328 0 _0079_
rlabel metal3 55272 39704 55272 39704 0 _0080_
rlabel metal2 53704 37856 53704 37856 0 _0081_
rlabel metal3 54264 35000 54264 35000 0 _0082_
rlabel metal2 53872 34216 53872 34216 0 _0083_
rlabel metal2 47880 35616 47880 35616 0 _0084_
rlabel metal3 47712 32424 47712 32424 0 _0085_
rlabel metal2 50008 30520 50008 30520 0 _0086_
rlabel metal3 52976 32536 52976 32536 0 _0087_
rlabel metal2 31304 42112 31304 42112 0 _0088_
rlabel metal2 27608 44632 27608 44632 0 _0089_
rlabel metal2 25816 46312 25816 46312 0 _0090_
rlabel metal2 23464 27048 23464 27048 0 _0091_
rlabel metal2 18760 45248 18760 45248 0 _0092_
rlabel metal2 30072 28280 30072 28280 0 _0093_
rlabel metal2 29960 27216 29960 27216 0 _0094_
rlabel metal2 26488 41216 26488 41216 0 _0095_
rlabel metal2 24472 40040 24472 40040 0 _0096_
rlabel metal2 26432 39704 26432 39704 0 _0097_
rlabel metal2 33376 27160 33376 27160 0 _0098_
rlabel metal2 33880 28168 33880 28168 0 _0099_
rlabel metal2 33880 29288 33880 29288 0 _0100_
rlabel metal3 33544 33208 33544 33208 0 _0101_
rlabel metal2 30240 31080 30240 31080 0 _0102_
rlabel metal2 35224 32704 35224 32704 0 _0103_
rlabel metal2 32424 36120 32424 36120 0 _0104_
rlabel metal2 32424 35336 32424 35336 0 _0105_
rlabel metal2 31696 31864 31696 31864 0 _0106_
rlabel metal2 28616 43456 28616 43456 0 _0107_
rlabel metal2 7448 41496 7448 41496 0 _0108_
rlabel metal2 8904 41216 8904 41216 0 _0109_
rlabel metal2 8120 33880 8120 33880 0 _0110_
rlabel metal2 3976 33096 3976 33096 0 _0111_
rlabel metal2 2520 36792 2520 36792 0 _0112_
rlabel metal2 2520 34608 2520 34608 0 _0113_
rlabel metal2 2520 39928 2520 39928 0 _0114_
rlabel metal2 4872 40040 4872 40040 0 _0115_
rlabel metal2 14672 40488 14672 40488 0 _0116_
rlabel metal2 11984 41832 11984 41832 0 _0117_
rlabel metal2 2520 48384 2520 48384 0 _0118_
rlabel metal2 2184 50232 2184 50232 0 _0119_
rlabel metal2 6440 50904 6440 50904 0 _0120_
rlabel metal2 2520 54096 2520 54096 0 _0121_
rlabel metal2 2520 52472 2520 52472 0 _0122_
rlabel metal2 3136 52808 3136 52808 0 _0123_
rlabel metal2 8120 54264 8120 54264 0 _0124_
rlabel metal2 2968 46928 2968 46928 0 _0125_
rlabel metal2 5152 45192 5152 45192 0 _0126_
rlabel metal2 11368 46704 11368 46704 0 _0127_
rlabel metal3 12880 46760 12880 46760 0 _0128_
rlabel metal2 10024 51800 10024 51800 0 _0129_
rlabel metal3 12600 48328 12600 48328 0 _0130_
rlabel metal2 7784 47768 7784 47768 0 _0131_
rlabel metal2 11704 53368 11704 53368 0 _0132_
rlabel metal2 9800 54768 9800 54768 0 _0133_
rlabel metal2 18704 25592 18704 25592 0 _0134_
rlabel metal3 12656 23800 12656 23800 0 _0135_
rlabel metal2 15176 21336 15176 21336 0 _0136_
rlabel metal2 8120 19936 8120 19936 0 _0137_
rlabel metal3 10416 19432 10416 19432 0 _0138_
rlabel metal2 13496 25032 13496 25032 0 _0139_
rlabel metal2 3976 23464 3976 23464 0 _0140_
rlabel metal2 5656 25928 5656 25928 0 _0141_
rlabel metal2 5880 21896 5880 21896 0 _0142_
rlabel metal2 5768 27496 5768 27496 0 _0143_
rlabel metal2 17416 43680 17416 43680 0 _0144_
rlabel metal2 22232 44688 22232 44688 0 _0145_
rlabel metal2 22680 43176 22680 43176 0 _0146_
rlabel metal3 23744 42840 23744 42840 0 _0147_
rlabel metal2 18536 5600 18536 5600 0 _0148_
rlabel metal3 16072 4424 16072 4424 0 _0149_
rlabel metal2 21168 4424 21168 4424 0 _0150_
rlabel metal2 23912 4760 23912 4760 0 _0151_
rlabel metal2 33880 17192 33880 17192 0 _0152_
rlabel metal2 37128 17192 37128 17192 0 _0153_
rlabel metal2 24696 8960 24696 8960 0 _0154_
rlabel metal2 27160 9912 27160 9912 0 _0155_
rlabel metal2 26488 20384 26488 20384 0 _0156_
rlabel metal2 29512 20440 29512 20440 0 _0157_
rlabel metal2 11592 8260 11592 8260 0 _0158_
rlabel metal2 14280 5376 14280 5376 0 _0159_
rlabel metal2 20216 7784 20216 7784 0 _0160_
rlabel metal2 17416 8736 17416 8736 0 _0161_
rlabel metal2 18648 11032 18648 11032 0 _0162_
rlabel metal2 20664 12488 20664 12488 0 _0163_
rlabel metal2 11928 11256 11928 11256 0 _0164_
rlabel metal2 15176 13440 15176 13440 0 _0165_
rlabel metal3 23688 20104 23688 20104 0 _0166_
rlabel metal2 22120 19600 22120 19600 0 _0167_
rlabel metal2 23912 22568 23912 22568 0 _0168_
rlabel metal3 25200 23352 25200 23352 0 _0169_
rlabel metal2 18424 15260 18424 15260 0 _0170_
rlabel metal2 20776 15736 20776 15736 0 _0171_
rlabel metal2 9576 17304 9576 17304 0 _0172_
rlabel metal2 8680 16464 8680 16464 0 _0173_
rlabel metal3 19096 18312 19096 18312 0 _0174_
rlabel metal2 16520 17304 16520 17304 0 _0175_
rlabel metal2 36064 22456 36064 22456 0 _0176_
rlabel metal2 37464 22736 37464 22736 0 _0177_
rlabel metal2 9576 14168 9576 14168 0 _0178_
rlabel metal2 9016 13272 9016 13272 0 _0179_
rlabel metal2 37128 21168 37128 21168 0 _0180_
rlabel metal3 37240 19320 37240 19320 0 _0181_
rlabel metal2 33880 11872 33880 11872 0 _0182_
rlabel metal2 35336 7784 35336 7784 0 _0183_
rlabel metal2 26488 24696 26488 24696 0 _0184_
rlabel metal2 29288 22736 29288 22736 0 _0185_
rlabel metal2 25256 55328 25256 55328 0 _0186_
rlabel metal2 27832 54936 27832 54936 0 _0187_
rlabel metal2 30632 53984 30632 53984 0 _0188_
rlabel metal2 32200 54936 32200 54936 0 _0189_
rlabel metal2 32200 52584 32200 52584 0 _0190_
rlabel metal2 33432 51856 33432 51856 0 _0191_
rlabel metal3 33824 50456 33824 50456 0 _0192_
rlabel metal2 48888 37856 48888 37856 0 _0193_
rlabel metal2 43288 38024 43288 38024 0 _0194_
rlabel metal2 40936 36120 40936 36120 0 _0195_
rlabel metal3 42280 34888 42280 34888 0 _0196_
rlabel metal2 41160 34048 41160 34048 0 _0197_
rlabel metal2 43064 36344 43064 36344 0 _0198_
rlabel metal2 43960 36120 43960 36120 0 _0199_
rlabel metal2 45528 36624 45528 36624 0 _0200_
rlabel metal2 44408 36120 44408 36120 0 _0201_
rlabel metal3 42840 37576 42840 37576 0 _0202_
rlabel metal2 41048 44968 41048 44968 0 _0203_
rlabel metal3 46872 48328 46872 48328 0 _0204_
rlabel metal3 42840 40600 42840 40600 0 _0205_
rlabel metal2 38864 36344 38864 36344 0 _0206_
rlabel metal3 39144 37240 39144 37240 0 _0207_
rlabel metal2 37912 30464 37912 30464 0 _0208_
rlabel metal2 40152 32592 40152 32592 0 _0209_
rlabel metal2 40488 35000 40488 35000 0 _0210_
rlabel metal2 39368 34216 39368 34216 0 _0211_
rlabel metal2 39704 36008 39704 36008 0 _0212_
rlabel metal2 40208 37464 40208 37464 0 _0213_
rlabel metal2 40096 38920 40096 38920 0 _0214_
rlabel metal2 42336 38808 42336 38808 0 _0215_
rlabel metal2 43904 40936 43904 40936 0 _0216_
rlabel metal2 42896 38808 42896 38808 0 _0217_
rlabel metal3 42224 38696 42224 38696 0 _0218_
rlabel metal2 40376 41440 40376 41440 0 _0219_
rlabel via2 46088 37800 46088 37800 0 _0220_
rlabel metal2 31304 42616 31304 42616 0 _0221_
rlabel metal2 41160 40264 41160 40264 0 _0222_
rlabel metal2 40936 40432 40936 40432 0 _0223_
rlabel metal2 37800 39984 37800 39984 0 _0224_
rlabel metal3 37408 39032 37408 39032 0 _0225_
rlabel metal2 38136 39928 38136 39928 0 _0226_
rlabel metal2 38584 40712 38584 40712 0 _0227_
rlabel metal2 38808 43568 38808 43568 0 _0228_
rlabel metal2 39816 41552 39816 41552 0 _0229_
rlabel metal3 40264 40488 40264 40488 0 _0230_
rlabel metal2 39144 40376 39144 40376 0 _0231_
rlabel metal2 46424 34720 46424 34720 0 _0232_
rlabel metal2 49448 31472 49448 31472 0 _0233_
rlabel metal2 39704 40824 39704 40824 0 _0234_
rlabel metal3 44240 41160 44240 41160 0 _0235_
rlabel metal2 48944 31192 48944 31192 0 _0236_
rlabel metal2 33432 40656 33432 40656 0 _0237_
rlabel metal2 47432 36232 47432 36232 0 _0238_
rlabel metal2 50792 46088 50792 46088 0 _0239_
rlabel metal2 40152 43008 40152 43008 0 _0240_
rlabel metal2 35896 43120 35896 43120 0 _0241_
rlabel metal2 38472 37352 38472 37352 0 _0242_
rlabel metal2 38080 35448 38080 35448 0 _0243_
rlabel metal2 37576 36232 37576 36232 0 _0244_
rlabel metal3 37016 38808 37016 38808 0 _0245_
rlabel metal2 38024 37632 38024 37632 0 _0246_
rlabel metal3 38808 36232 38808 36232 0 _0247_
rlabel metal2 38304 35672 38304 35672 0 _0248_
rlabel metal2 38808 37016 38808 37016 0 _0249_
rlabel metal3 39704 42840 39704 42840 0 _0250_
rlabel metal2 40264 42504 40264 42504 0 _0251_
rlabel metal2 33768 41048 33768 41048 0 _0252_
rlabel metal3 19432 39592 19432 39592 0 _0253_
rlabel metal2 47096 48720 47096 48720 0 _0254_
rlabel metal3 35224 43624 35224 43624 0 _0255_
rlabel metal3 35504 43512 35504 43512 0 _0256_
rlabel metal3 34048 43512 34048 43512 0 _0257_
rlabel metal2 39312 42728 39312 42728 0 _0258_
rlabel metal2 39032 42784 39032 42784 0 _0259_
rlabel metal2 38696 45416 38696 45416 0 _0260_
rlabel metal2 37912 42504 37912 42504 0 _0261_
rlabel metal2 38248 42448 38248 42448 0 _0262_
rlabel metal3 38192 44296 38192 44296 0 _0263_
rlabel metal2 27776 42504 27776 42504 0 _0264_
rlabel metal3 26488 45640 26488 45640 0 _0265_
rlabel metal2 38808 45584 38808 45584 0 _0266_
rlabel metal2 33992 43960 33992 43960 0 _0267_
rlabel metal3 34944 45080 34944 45080 0 _0268_
rlabel metal3 35504 44184 35504 44184 0 _0269_
rlabel metal3 35504 51352 35504 51352 0 _0270_
rlabel metal3 36960 50456 36960 50456 0 _0271_
rlabel metal3 40040 48216 40040 48216 0 _0272_
rlabel metal2 37576 45808 37576 45808 0 _0273_
rlabel metal2 37856 45304 37856 45304 0 _0274_
rlabel metal2 37240 46200 37240 46200 0 _0275_
rlabel metal2 38920 47208 38920 47208 0 _0276_
rlabel metal3 38668 49784 38668 49784 0 _0277_
rlabel metal2 39256 49000 39256 49000 0 _0278_
rlabel metal2 48776 45192 48776 45192 0 _0279_
rlabel metal2 39592 46536 39592 46536 0 _0280_
rlabel metal2 39256 46816 39256 46816 0 _0281_
rlabel metal3 38360 46536 38360 46536 0 _0282_
rlabel metal2 45640 49168 45640 49168 0 _0283_
rlabel metal2 41160 52136 41160 52136 0 _0284_
rlabel metal2 45976 38304 45976 38304 0 _0285_
rlabel metal2 36568 50904 36568 50904 0 _0286_
rlabel metal2 37128 51576 37128 51576 0 _0287_
rlabel metal2 39032 52584 39032 52584 0 _0288_
rlabel metal2 40040 50624 40040 50624 0 _0289_
rlabel metal2 41272 47712 41272 47712 0 _0290_
rlabel metal2 38024 51240 38024 51240 0 _0291_
rlabel metal2 41048 47376 41048 47376 0 _0292_
rlabel metal2 42168 47880 42168 47880 0 _0293_
rlabel metal2 41944 47544 41944 47544 0 _0294_
rlabel metal2 42504 48664 42504 48664 0 _0295_
rlabel metal2 42056 49000 42056 49000 0 _0296_
rlabel metal2 40824 50204 40824 50204 0 _0297_
rlabel metal2 39760 51464 39760 51464 0 _0298_
rlabel metal2 40264 50792 40264 50792 0 _0299_
rlabel metal2 41272 50960 41272 50960 0 _0300_
rlabel metal2 41720 51744 41720 51744 0 _0301_
rlabel metal2 37912 51744 37912 51744 0 _0302_
rlabel metal2 45360 51352 45360 51352 0 _0303_
rlabel metal3 42224 51240 42224 51240 0 _0304_
rlabel metal2 42728 50232 42728 50232 0 _0305_
rlabel metal2 41328 48888 41328 48888 0 _0306_
rlabel metal2 40264 50204 40264 50204 0 _0307_
rlabel metal2 40264 49448 40264 49448 0 _0308_
rlabel metal2 45696 32648 45696 32648 0 _0309_
rlabel metal2 41832 50372 41832 50372 0 _0310_
rlabel metal2 45752 36176 45752 36176 0 _0311_
rlabel metal2 42952 39648 42952 39648 0 _0312_
rlabel metal2 43512 39928 43512 39928 0 _0313_
rlabel metal2 41608 53424 41608 53424 0 _0314_
rlabel metal2 43176 51856 43176 51856 0 _0315_
rlabel metal2 48440 49336 48440 49336 0 _0316_
rlabel metal2 50344 47880 50344 47880 0 _0317_
rlabel metal2 45304 48160 45304 48160 0 _0318_
rlabel metal2 45248 48440 45248 48440 0 _0319_
rlabel metal3 45920 37240 45920 37240 0 _0320_
rlabel metal2 43848 48944 43848 48944 0 _0321_
rlabel metal2 44184 48496 44184 48496 0 _0322_
rlabel metal2 46760 51464 46760 51464 0 _0323_
rlabel metal2 38136 51408 38136 51408 0 _0324_
rlabel metal2 53032 50848 53032 50848 0 _0325_
rlabel metal2 47768 51744 47768 51744 0 _0326_
rlabel metal2 46200 48552 46200 48552 0 _0327_
rlabel metal2 48104 47880 48104 47880 0 _0328_
rlabel metal3 46648 49784 46648 49784 0 _0329_
rlabel metal3 49672 49560 49672 49560 0 _0330_
rlabel metal2 46648 50064 46648 50064 0 _0331_
rlabel metal2 46032 48440 46032 48440 0 _0332_
rlabel metal2 45528 49336 45528 49336 0 _0333_
rlabel metal3 47488 52136 47488 52136 0 _0334_
rlabel metal2 49224 51688 49224 51688 0 _0335_
rlabel metal2 49504 50680 49504 50680 0 _0336_
rlabel metal2 50344 50848 50344 50848 0 _0337_
rlabel metal2 49392 49784 49392 49784 0 _0338_
rlabel metal3 49616 49672 49616 49672 0 _0339_
rlabel metal2 46760 35112 46760 35112 0 _0340_
rlabel metal2 47992 52304 47992 52304 0 _0341_
rlabel metal3 48552 52808 48552 52808 0 _0342_
rlabel metal2 54600 50092 54600 50092 0 _0343_
rlabel metal2 49896 49000 49896 49000 0 _0344_
rlabel metal2 49672 49056 49672 49056 0 _0345_
rlabel metal3 50680 49896 50680 49896 0 _0346_
rlabel metal3 49112 47992 49112 47992 0 _0347_
rlabel metal2 48104 49336 48104 49336 0 _0348_
rlabel metal2 50344 44632 50344 44632 0 _0349_
rlabel metal2 51632 47656 51632 47656 0 _0350_
rlabel metal2 50792 50960 50792 50960 0 _0351_
rlabel metal2 51128 52136 51128 52136 0 _0352_
rlabel metal2 53088 49000 53088 49000 0 _0353_
rlabel metal2 50960 49672 50960 49672 0 _0354_
rlabel metal2 51912 47600 51912 47600 0 _0355_
rlabel metal2 52696 47824 52696 47824 0 _0356_
rlabel metal2 53480 47432 53480 47432 0 _0357_
rlabel metal2 52920 48216 52920 48216 0 _0358_
rlabel metal2 52472 43064 52472 43064 0 _0359_
rlabel metal2 52920 46200 52920 46200 0 _0360_
rlabel metal2 51408 45864 51408 45864 0 _0361_
rlabel metal2 52696 45920 52696 45920 0 _0362_
rlabel metal2 50008 45248 50008 45248 0 _0363_
rlabel metal2 49672 45808 49672 45808 0 _0364_
rlabel metal3 55888 49784 55888 49784 0 _0365_
rlabel metal3 53480 49784 53480 49784 0 _0366_
rlabel metal2 50120 46144 50120 46144 0 _0367_
rlabel metal2 50288 45976 50288 45976 0 _0368_
rlabel metal3 51240 46648 51240 46648 0 _0369_
rlabel metal2 46536 47152 46536 47152 0 _0370_
rlabel metal2 54376 46144 54376 46144 0 _0371_
rlabel metal2 54880 44296 54880 44296 0 _0372_
rlabel metal2 57288 44184 57288 44184 0 _0373_
rlabel metal2 53816 45528 53816 45528 0 _0374_
rlabel metal2 53480 45080 53480 45080 0 _0375_
rlabel metal2 50848 45192 50848 45192 0 _0376_
rlabel metal3 50456 44072 50456 44072 0 _0377_
rlabel metal2 53032 44240 53032 44240 0 _0378_
rlabel metal2 54656 44968 54656 44968 0 _0379_
rlabel metal2 53704 45024 53704 45024 0 _0380_
rlabel metal2 53536 45864 53536 45864 0 _0381_
rlabel metal3 56560 43624 56560 43624 0 _0382_
rlabel metal2 57176 44408 57176 44408 0 _0383_
rlabel metal3 55160 44296 55160 44296 0 _0384_
rlabel metal2 52864 44856 52864 44856 0 _0385_
rlabel metal2 53200 43400 53200 43400 0 _0386_
rlabel metal2 53704 43624 53704 43624 0 _0387_
rlabel metal3 43456 41832 43456 41832 0 _0388_
rlabel metal2 53200 42840 53200 42840 0 _0389_
rlabel metal2 55888 42168 55888 42168 0 _0390_
rlabel metal2 57064 42616 57064 42616 0 _0391_
rlabel metal3 53424 41832 53424 41832 0 _0392_
rlabel metal2 50008 41496 50008 41496 0 _0393_
rlabel metal2 50568 41384 50568 41384 0 _0394_
rlabel metal2 51800 41384 51800 41384 0 _0395_
rlabel metal2 50680 41496 50680 41496 0 _0396_
rlabel metal2 47880 41272 47880 41272 0 _0397_
rlabel metal2 47712 40488 47712 40488 0 _0398_
rlabel metal2 53312 41944 53312 41944 0 _0399_
rlabel metal2 51688 42840 51688 42840 0 _0400_
rlabel metal3 53312 41272 53312 41272 0 _0401_
rlabel metal3 52136 41944 52136 41944 0 _0402_
rlabel metal3 52864 40264 52864 40264 0 _0403_
rlabel metal2 53928 40208 53928 40208 0 _0404_
rlabel metal2 57288 40040 57288 40040 0 _0405_
rlabel metal2 51352 40376 51352 40376 0 _0406_
rlabel metal2 51464 39200 51464 39200 0 _0407_
rlabel metal2 50904 40152 50904 40152 0 _0408_
rlabel metal2 51016 39592 51016 39592 0 _0409_
rlabel metal2 50344 38192 50344 38192 0 _0410_
rlabel metal2 53144 39032 53144 39032 0 _0411_
rlabel metal2 53256 39144 53256 39144 0 _0412_
rlabel metal2 53704 39480 53704 39480 0 _0413_
rlabel metal3 55104 38024 55104 38024 0 _0414_
rlabel metal2 57008 36456 57008 36456 0 _0415_
rlabel metal2 57176 37464 57176 37464 0 _0416_
rlabel metal2 57624 36792 57624 36792 0 _0417_
rlabel metal2 50232 37688 50232 37688 0 _0418_
rlabel metal3 51744 37912 51744 37912 0 _0419_
rlabel metal2 53256 37520 53256 37520 0 _0420_
rlabel metal3 54208 37464 54208 37464 0 _0421_
rlabel metal3 47376 31864 47376 31864 0 _0422_
rlabel metal3 54600 35672 54600 35672 0 _0423_
rlabel metal2 55272 36512 55272 36512 0 _0424_
rlabel metal3 54488 37240 54488 37240 0 _0425_
rlabel metal3 54488 35448 54488 35448 0 _0426_
rlabel metal2 41944 36288 41944 36288 0 _0427_
rlabel metal2 53032 35224 53032 35224 0 _0428_
rlabel metal3 52248 36456 52248 36456 0 _0429_
rlabel metal2 49560 34832 49560 34832 0 _0430_
rlabel metal2 52416 35672 52416 35672 0 _0431_
rlabel metal2 51352 37688 51352 37688 0 _0432_
rlabel metal2 49672 36400 49672 36400 0 _0433_
rlabel metal2 53592 34776 53592 34776 0 _0434_
rlabel metal2 53928 35336 53928 35336 0 _0435_
rlabel metal2 49560 36624 49560 36624 0 _0436_
rlabel metal2 48664 36456 48664 36456 0 _0437_
rlabel metal2 48048 35896 48048 35896 0 _0438_
rlabel metal2 48776 32984 48776 32984 0 _0439_
rlabel metal2 48048 32760 48048 32760 0 _0440_
rlabel metal2 49560 33320 49560 33320 0 _0441_
rlabel metal2 48440 33768 48440 33768 0 _0442_
rlabel metal2 49672 31696 49672 31696 0 _0443_
rlabel metal2 47824 32424 47824 32424 0 _0444_
rlabel metal2 49672 32872 49672 32872 0 _0445_
rlabel metal2 51296 30968 51296 30968 0 _0446_
rlabel metal2 50512 32760 50512 32760 0 _0447_
rlabel metal3 51520 31752 51520 31752 0 _0448_
rlabel metal2 50456 31304 50456 31304 0 _0449_
rlabel metal2 50120 31136 50120 31136 0 _0450_
rlabel metal2 51800 33264 51800 33264 0 _0451_
rlabel metal3 52024 31864 52024 31864 0 _0452_
rlabel metal2 13160 39032 13160 39032 0 _0453_
rlabel metal2 30632 41944 30632 41944 0 _0454_
rlabel metal2 20104 44464 20104 44464 0 _0455_
rlabel metal2 25816 30576 25816 30576 0 _0456_
rlabel metal2 23128 28728 23128 28728 0 _0457_
rlabel metal2 25872 32760 25872 32760 0 _0458_
rlabel metal2 20160 45640 20160 45640 0 _0459_
rlabel metal2 19544 46452 19544 46452 0 _0460_
rlabel metal2 32648 30632 32648 30632 0 _0461_
rlabel metal2 31080 26628 31080 26628 0 _0462_
rlabel metal2 26600 40320 26600 40320 0 _0463_
rlabel metal3 20832 39480 20832 39480 0 _0464_
rlabel metal3 21784 38808 21784 38808 0 _0465_
rlabel metal2 20552 38304 20552 38304 0 _0466_
rlabel metal2 16968 40880 16968 40880 0 _0467_
rlabel metal2 24920 38136 24920 38136 0 _0468_
rlabel metal3 19096 38136 19096 38136 0 _0469_
rlabel metal2 18984 35392 18984 35392 0 _0470_
rlabel metal2 18760 36176 18760 36176 0 _0471_
rlabel metal2 22120 38864 22120 38864 0 _0472_
rlabel metal2 24136 38864 24136 38864 0 _0473_
rlabel metal3 28840 37912 28840 37912 0 _0474_
rlabel metal2 26488 38668 26488 38668 0 _0475_
rlabel metal2 26824 39704 26824 39704 0 _0476_
rlabel metal3 24864 38808 24864 38808 0 _0477_
rlabel metal4 21336 38192 21336 38192 0 _0478_
rlabel metal3 23800 35616 23800 35616 0 _0479_
rlabel metal2 26656 37800 26656 37800 0 _0480_
rlabel metal3 25872 34888 25872 34888 0 _0481_
rlabel metal2 24248 37520 24248 37520 0 _0482_
rlabel metal2 23912 38192 23912 38192 0 _0483_
rlabel metal2 25704 37800 25704 37800 0 _0484_
rlabel metal2 26208 39032 26208 39032 0 _0485_
rlabel metal2 22232 39592 22232 39592 0 _0486_
rlabel metal2 28392 38780 28392 38780 0 _0487_
rlabel metal2 27832 39312 27832 39312 0 _0488_
rlabel metal2 27272 39704 27272 39704 0 _0489_
rlabel metal2 20104 34104 20104 34104 0 _0490_
rlabel metal3 24584 32536 24584 32536 0 _0491_
rlabel metal2 19992 33712 19992 33712 0 _0492_
rlabel metal2 17640 34944 17640 34944 0 _0493_
rlabel metal3 28448 33208 28448 33208 0 _0494_
rlabel metal2 31248 35672 31248 35672 0 _0495_
rlabel metal3 33096 29400 33096 29400 0 _0496_
rlabel metal2 26824 36848 26824 36848 0 _0497_
rlabel metal2 29960 35616 29960 35616 0 _0498_
rlabel metal3 23184 37912 23184 37912 0 _0499_
rlabel metal2 24584 38304 24584 38304 0 _0500_
rlabel metal2 24920 36736 24920 36736 0 _0501_
rlabel metal2 33096 29792 33096 29792 0 _0502_
rlabel metal2 33544 29512 33544 29512 0 _0503_
rlabel metal2 25928 31920 25928 31920 0 _0504_
rlabel metal2 25816 31584 25816 31584 0 _0505_
rlabel metal2 26712 30520 26712 30520 0 _0506_
rlabel metal2 24752 30408 24752 30408 0 _0507_
rlabel metal3 20328 30968 20328 30968 0 _0508_
rlabel metal2 24416 30184 24416 30184 0 _0509_
rlabel metal2 29176 36120 29176 36120 0 _0510_
rlabel metal3 25816 30184 25816 30184 0 _0511_
rlabel metal2 24696 34608 24696 34608 0 _0512_
rlabel metal2 10976 42168 10976 42168 0 _0513_
rlabel metal3 12040 39144 12040 39144 0 _0514_
rlabel metal2 13048 37576 13048 37576 0 _0515_
rlabel metal3 24640 35784 24640 35784 0 _0516_
rlabel metal2 27496 32368 27496 32368 0 _0517_
rlabel metal2 28280 32088 28280 32088 0 _0518_
rlabel metal2 31976 29512 31976 29512 0 _0519_
rlabel metal2 32424 29064 32424 29064 0 _0520_
rlabel metal3 20720 40376 20720 40376 0 _0521_
rlabel metal2 22344 40936 22344 40936 0 _0522_
rlabel metal3 20496 36232 20496 36232 0 _0523_
rlabel metal3 22120 36568 22120 36568 0 _0524_
rlabel metal3 24584 31640 24584 31640 0 _0525_
rlabel metal3 26740 31528 26740 31528 0 _0526_
rlabel metal2 33320 31304 33320 31304 0 _0527_
rlabel metal2 28560 34216 28560 34216 0 _0528_
rlabel metal2 32424 31808 32424 31808 0 _0529_
rlabel metal2 33768 30856 33768 30856 0 _0530_
rlabel metal2 27608 34048 27608 34048 0 _0531_
rlabel metal2 21112 34496 21112 34496 0 _0532_
rlabel metal2 22288 35000 22288 35000 0 _0533_
rlabel metal2 22008 33936 22008 33936 0 _0534_
rlabel metal2 26824 33936 26824 33936 0 _0535_
rlabel metal2 25424 34328 25424 34328 0 _0536_
rlabel metal2 23632 31752 23632 31752 0 _0537_
rlabel metal2 21448 31360 21448 31360 0 _0538_
rlabel metal2 25704 33152 25704 33152 0 _0539_
rlabel metal2 25312 33320 25312 33320 0 _0540_
rlabel metal2 25592 34160 25592 34160 0 _0541_
rlabel metal2 32536 33376 32536 33376 0 _0542_
rlabel metal2 31416 36064 31416 36064 0 _0543_
rlabel metal2 33208 33656 33208 33656 0 _0544_
rlabel metal2 25032 32200 25032 32200 0 _0545_
rlabel metal2 23240 34888 23240 34888 0 _0546_
rlabel metal3 24752 34664 24752 34664 0 _0547_
rlabel metal2 24248 34552 24248 34552 0 _0548_
rlabel metal2 30240 31752 30240 31752 0 _0549_
rlabel metal2 30632 31864 30632 31864 0 _0550_
rlabel metal2 22680 35952 22680 35952 0 _0551_
rlabel metal2 23464 35616 23464 35616 0 _0552_
rlabel metal2 31528 33936 31528 33936 0 _0553_
rlabel metal2 31808 33544 31808 33544 0 _0554_
rlabel metal2 26040 33936 26040 33936 0 _0555_
rlabel metal3 30128 34888 30128 34888 0 _0556_
rlabel metal2 29792 34216 29792 34216 0 _0557_
rlabel metal2 32200 35504 32200 35504 0 _0558_
rlabel metal3 33768 35448 33768 35448 0 _0559_
rlabel metal2 31192 32368 31192 32368 0 _0560_
rlabel metal2 27328 32760 27328 32760 0 _0561_
rlabel metal2 24024 34272 24024 34272 0 _0562_
rlabel metal2 26712 33992 26712 33992 0 _0563_
rlabel metal3 29064 33320 29064 33320 0 _0564_
rlabel metal2 30968 33600 30968 33600 0 _0565_
rlabel metal2 32872 35224 32872 35224 0 _0566_
rlabel metal3 32480 32536 32480 32536 0 _0567_
rlabel metal2 26040 30968 26040 30968 0 _0568_
rlabel metal2 27664 34664 27664 34664 0 _0569_
rlabel metal3 30072 32536 30072 32536 0 _0570_
rlabel metal2 23352 43904 23352 43904 0 _0571_
rlabel metal3 23688 36344 23688 36344 0 _0572_
rlabel metal3 26152 36232 26152 36232 0 _0573_
rlabel metal2 28168 36512 28168 36512 0 _0574_
rlabel metal2 28616 36512 28616 36512 0 _0575_
rlabel metal2 29624 40936 29624 40936 0 _0576_
rlabel metal3 9408 38808 9408 38808 0 _0577_
rlabel metal2 15400 37744 15400 37744 0 _0578_
rlabel metal3 14840 36400 14840 36400 0 _0579_
rlabel metal2 15064 36120 15064 36120 0 _0580_
rlabel metal2 9688 36960 9688 36960 0 _0581_
rlabel metal2 9016 38724 9016 38724 0 _0582_
rlabel metal3 10360 39592 10360 39592 0 _0583_
rlabel metal2 7560 52136 7560 52136 0 _0584_
rlabel metal2 6328 54768 6328 54768 0 _0585_
rlabel metal2 7728 52360 7728 52360 0 _0586_
rlabel metal2 8568 45304 8568 45304 0 _0587_
rlabel metal2 8904 45528 8904 45528 0 _0588_
rlabel metal2 9800 44464 9800 44464 0 _0589_
rlabel metal2 10360 45360 10360 45360 0 _0590_
rlabel metal2 7336 48944 7336 48944 0 _0591_
rlabel metal2 10584 44744 10584 44744 0 _0592_
rlabel metal2 9576 43960 9576 43960 0 _0593_
rlabel metal3 10360 51576 10360 51576 0 _0594_
rlabel metal2 5768 48888 5768 48888 0 _0595_
rlabel metal2 9576 49952 9576 49952 0 _0596_
rlabel metal2 10584 43736 10584 43736 0 _0597_
rlabel metal3 9800 44408 9800 44408 0 _0598_
rlabel metal2 8624 38808 8624 38808 0 _0599_
rlabel metal2 9800 40488 9800 40488 0 _0600_
rlabel metal2 7504 39592 7504 39592 0 _0601_
rlabel metal2 7112 39592 7112 39592 0 _0602_
rlabel metal2 15512 37128 15512 37128 0 _0603_
rlabel metal2 18984 30240 18984 30240 0 _0604_
rlabel metal2 10584 38080 10584 38080 0 _0605_
rlabel metal2 9632 39368 9632 39368 0 _0606_
rlabel metal3 9576 39368 9576 39368 0 _0607_
rlabel metal2 9352 39928 9352 39928 0 _0608_
rlabel metal2 8120 35112 8120 35112 0 _0609_
rlabel metal2 8568 33880 8568 33880 0 _0610_
rlabel metal2 13496 35112 13496 35112 0 _0611_
rlabel metal2 2968 34272 2968 34272 0 _0612_
rlabel metal2 5320 34384 5320 34384 0 _0613_
rlabel metal2 4984 35784 4984 35784 0 _0614_
rlabel metal2 10360 39256 10360 39256 0 _0615_
rlabel metal2 6440 39424 6440 39424 0 _0616_
rlabel metal2 3640 37184 3640 37184 0 _0617_
rlabel metal2 3080 35840 3080 35840 0 _0618_
rlabel via2 3416 38808 3416 38808 0 _0619_
rlabel metal2 2744 36512 2744 36512 0 _0620_
rlabel metal2 3192 35280 3192 35280 0 _0621_
rlabel metal2 3976 39592 3976 39592 0 _0622_
rlabel metal2 12376 39088 12376 39088 0 _0623_
rlabel metal2 12040 40320 12040 40320 0 _0624_
rlabel metal2 3528 39592 3528 39592 0 _0625_
rlabel metal3 4872 39480 4872 39480 0 _0626_
rlabel metal3 10696 38024 10696 38024 0 _0627_
rlabel metal2 7224 39312 7224 39312 0 _0628_
rlabel metal2 14000 40936 14000 40936 0 _0629_
rlabel metal2 24584 34720 24584 34720 0 _0630_
rlabel metal2 14168 38472 14168 38472 0 _0631_
rlabel metal2 14616 38864 14616 38864 0 _0632_
rlabel metal2 12712 34160 12712 34160 0 _0633_
rlabel metal3 13384 38808 13384 38808 0 _0634_
rlabel metal3 12992 39704 12992 39704 0 _0635_
rlabel metal3 10472 50456 10472 50456 0 _0636_
rlabel metal3 5432 48440 5432 48440 0 _0637_
rlabel metal2 3304 53312 3304 53312 0 _0638_
rlabel metal2 2464 49784 2464 49784 0 _0639_
rlabel metal2 5432 52024 5432 52024 0 _0640_
rlabel metal2 5208 51912 5208 51912 0 _0641_
rlabel metal2 5712 49112 5712 49112 0 _0642_
rlabel metal2 2800 53592 2800 53592 0 _0643_
rlabel metal2 6216 53704 6216 53704 0 _0644_
rlabel metal2 5096 52136 5096 52136 0 _0645_
rlabel metal2 3528 53648 3528 53648 0 _0646_
rlabel metal2 6664 53536 6664 53536 0 _0647_
rlabel metal2 7280 53144 7280 53144 0 _0648_
rlabel metal2 11536 47544 11536 47544 0 _0649_
rlabel metal3 5488 47432 5488 47432 0 _0650_
rlabel metal2 6552 46256 6552 46256 0 _0651_
rlabel metal2 4984 46200 4984 46200 0 _0652_
rlabel metal2 8680 46704 8680 46704 0 _0653_
rlabel metal3 10024 47432 10024 47432 0 _0654_
rlabel metal2 10920 47936 10920 47936 0 _0655_
rlabel metal2 12040 47320 12040 47320 0 _0656_
rlabel metal3 11536 48888 11536 48888 0 _0657_
rlabel metal2 11256 50624 11256 50624 0 _0658_
rlabel metal2 11480 50792 11480 50792 0 _0659_
rlabel metal2 11984 50568 11984 50568 0 _0660_
rlabel metal2 11368 50736 11368 50736 0 _0661_
rlabel metal3 9520 49000 9520 49000 0 _0662_
rlabel metal3 12208 49784 12208 49784 0 _0663_
rlabel metal3 9408 48104 9408 48104 0 _0664_
rlabel metal2 11480 52584 11480 52584 0 _0665_
rlabel metal2 11872 52248 11872 52248 0 _0666_
rlabel metal2 10472 53648 10472 53648 0 _0667_
rlabel metal2 10136 53648 10136 53648 0 _0668_
rlabel metal2 18648 26600 18648 26600 0 _0669_
rlabel metal2 16576 28056 16576 28056 0 _0670_
rlabel metal2 18088 24304 18088 24304 0 _0671_
rlabel metal3 18704 26040 18704 26040 0 _0672_
rlabel metal2 14672 24136 14672 24136 0 _0673_
rlabel metal2 15176 24752 15176 24752 0 _0674_
rlabel metal2 15288 23464 15288 23464 0 _0675_
rlabel metal2 16632 21840 16632 21840 0 _0676_
rlabel metal2 14616 21728 14616 21728 0 _0677_
rlabel metal2 11648 20664 11648 20664 0 _0678_
rlabel metal2 13160 20132 13160 20132 0 _0679_
rlabel metal2 12488 19656 12488 19656 0 _0680_
rlabel metal2 5656 22736 5656 22736 0 _0681_
rlabel metal2 18480 42728 18480 42728 0 _0682_
rlabel metal2 18872 42616 18872 42616 0 _0683_
rlabel via2 19992 41832 19992 41832 0 _0684_
rlabel metal2 21112 31416 21112 31416 0 _0685_
rlabel metal2 17360 40040 17360 40040 0 _0686_
rlabel metal2 19544 40712 19544 40712 0 _0687_
rlabel metal2 19096 40992 19096 40992 0 _0688_
rlabel metal2 16296 40656 16296 40656 0 _0689_
rlabel metal2 16408 40824 16408 40824 0 _0690_
rlabel metal2 19320 41720 19320 41720 0 _0691_
rlabel metal2 17416 42168 17416 42168 0 _0692_
rlabel metal3 21224 40600 21224 40600 0 _0693_
rlabel metal2 22344 30576 22344 30576 0 _0694_
rlabel metal2 20944 32648 20944 32648 0 _0695_
rlabel metal2 23016 31472 23016 31472 0 _0696_
rlabel metal2 21504 40936 21504 40936 0 _0697_
rlabel metal3 20888 41160 20888 41160 0 _0698_
rlabel metal3 17808 41160 17808 41160 0 _0699_
rlabel metal2 19880 41664 19880 41664 0 _0700_
rlabel metal2 21336 43904 21336 43904 0 _0701_
rlabel metal3 21672 31752 21672 31752 0 _0702_
rlabel metal2 20328 32536 20328 32536 0 _0703_
rlabel metal2 21448 41496 21448 41496 0 _0704_
rlabel metal3 17752 41888 17752 41888 0 _0705_
rlabel metal2 17976 42168 17976 42168 0 _0706_
rlabel metal2 22064 42840 22064 42840 0 _0707_
rlabel metal2 21000 40432 21000 40432 0 _0708_
rlabel metal3 18032 41384 18032 41384 0 _0709_
rlabel metal3 19936 41944 19936 41944 0 _0710_
rlabel metal2 21336 42168 21336 42168 0 _0711_
rlabel metal2 22624 9800 22624 9800 0 _0712_
rlabel metal2 18312 6216 18312 6216 0 _0713_
rlabel metal2 19656 5208 19656 5208 0 _0714_
rlabel metal2 17640 4984 17640 4984 0 _0715_
rlabel metal2 22344 5880 22344 5880 0 _0716_
rlabel metal2 20440 5824 20440 5824 0 _0717_
rlabel metal2 23576 4648 23576 4648 0 _0718_
rlabel metal3 22512 20664 22512 20664 0 _0719_
rlabel metal3 23464 18928 23464 18928 0 _0720_
rlabel metal2 33544 17864 33544 17864 0 _0721_
rlabel metal2 37464 17696 37464 17696 0 _0722_
rlabel metal3 24584 9688 24584 9688 0 _0723_
rlabel metal2 25368 9688 25368 9688 0 _0724_
rlabel metal2 27384 10080 27384 10080 0 _0725_
rlabel metal2 15848 20832 15848 20832 0 _0726_
rlabel metal2 22344 16856 22344 16856 0 _0727_
rlabel metal2 29400 20888 29400 20888 0 _0728_
rlabel metal2 28056 20776 28056 20776 0 _0729_
rlabel metal2 30072 20440 30072 20440 0 _0730_
rlabel metal3 18144 15400 18144 15400 0 _0731_
rlabel metal2 17752 9296 17752 9296 0 _0732_
rlabel metal3 12936 8792 12936 8792 0 _0733_
rlabel metal2 15176 5768 15176 5768 0 _0734_
rlabel metal2 20552 10360 20552 10360 0 _0735_
rlabel metal2 19376 9016 19376 9016 0 _0736_
rlabel metal2 19992 8512 19992 8512 0 _0737_
rlabel metal2 18760 12292 18760 12292 0 _0738_
rlabel metal2 17920 7672 17920 7672 0 _0739_
rlabel metal2 22008 10920 22008 10920 0 _0740_
rlabel metal3 19320 10584 19320 10584 0 _0741_
rlabel metal2 21448 12264 21448 12264 0 _0742_
rlabel metal2 16744 20328 16744 20328 0 _0743_
rlabel metal2 16744 13328 16744 13328 0 _0744_
rlabel metal2 12488 11648 12488 11648 0 _0745_
rlabel metal3 16800 12936 16800 12936 0 _0746_
rlabel metal2 22232 20440 22232 20440 0 _0747_
rlabel metal2 24696 21728 24696 21728 0 _0748_
rlabel metal2 24696 20720 24696 20720 0 _0749_
rlabel metal2 24080 21560 24080 21560 0 _0750_
rlabel metal2 22568 19712 22568 19712 0 _0751_
rlabel metal2 26040 23128 26040 23128 0 _0752_
rlabel metal2 24248 22680 24248 22680 0 _0753_
rlabel metal2 25144 22848 25144 22848 0 _0754_
rlabel metal2 22120 15876 22120 15876 0 _0755_
rlabel metal2 18760 15204 18760 15204 0 _0756_
rlabel metal2 21504 14728 21504 14728 0 _0757_
rlabel metal2 19208 17080 19208 17080 0 _0758_
rlabel metal3 10584 16296 10584 16296 0 _0759_
rlabel metal2 7896 17920 7896 17920 0 _0760_
rlabel metal2 18648 17192 18648 17192 0 _0761_
rlabel metal2 19320 17920 19320 17920 0 _0762_
rlabel metal3 17192 16968 17192 16968 0 _0763_
rlabel metal2 37744 22232 37744 22232 0 _0764_
rlabel metal3 37296 22120 37296 22120 0 _0765_
rlabel metal3 36344 22344 36344 22344 0 _0766_
rlabel metal2 12264 14056 12264 14056 0 _0767_
rlabel metal3 10528 13720 10528 13720 0 _0768_
rlabel metal2 10584 14448 10584 14448 0 _0769_
rlabel metal2 36120 18760 36120 18760 0 _0770_
rlabel metal2 36008 19992 36008 19992 0 _0771_
rlabel metal2 36008 18256 36008 18256 0 _0772_
rlabel metal2 33992 9352 33992 9352 0 _0773_
rlabel metal2 33824 10808 33824 10808 0 _0774_
rlabel metal2 34888 8512 34888 8512 0 _0775_
rlabel metal2 22008 21896 22008 21896 0 _0776_
rlabel metal2 27384 23408 27384 23408 0 _0777_
rlabel metal2 29624 23184 29624 23184 0 _0778_
rlabel metal2 17528 55216 17528 55216 0 _0779_
rlabel metal2 18480 43624 18480 43624 0 _0780_
rlabel metal3 21672 37240 21672 37240 0 _0781_
rlabel metal2 23912 34832 23912 34832 0 _0782_
rlabel metal2 20664 28616 20664 28616 0 _0783_
rlabel metal2 20440 32144 20440 32144 0 _0784_
rlabel metal3 17136 31080 17136 31080 0 _0785_
rlabel metal3 26152 13720 26152 13720 0 _0786_
rlabel metal2 23240 10864 23240 10864 0 _0787_
rlabel metal2 24864 17640 24864 17640 0 _0788_
rlabel metal2 32256 13944 32256 13944 0 _0789_
rlabel metal2 31864 16464 31864 16464 0 _0790_
rlabel metal2 29848 18816 29848 18816 0 _0791_
rlabel metal2 29400 22064 29400 22064 0 _0792_
rlabel metal2 27440 19208 27440 19208 0 _0793_
rlabel metal3 30128 18424 30128 18424 0 _0794_
rlabel metal2 27720 13552 27720 13552 0 _0795_
rlabel metal2 27832 11480 27832 11480 0 _0796_
rlabel metal2 23128 17864 23128 17864 0 _0797_
rlabel metal3 23016 12376 23016 12376 0 _0798_
rlabel metal2 17752 13608 17752 13608 0 _0799_
rlabel metal2 16744 10248 16744 10248 0 _0800_
rlabel metal3 24920 12152 24920 12152 0 _0801_
rlabel metal3 25928 11368 25928 11368 0 _0802_
rlabel metal3 35560 12152 35560 12152 0 _0803_
rlabel metal2 31080 8792 31080 8792 0 _0804_
rlabel metal2 29176 6104 29176 6104 0 _0805_
rlabel metal2 24472 16576 24472 16576 0 _0806_
rlabel metal3 34160 15848 34160 15848 0 _0807_
rlabel metal2 23408 7448 23408 7448 0 _0808_
rlabel metal2 29568 10024 29568 10024 0 _0809_
rlabel metal3 33096 15288 33096 15288 0 _0810_
rlabel metal2 30016 11928 30016 11928 0 _0811_
rlabel metal2 35448 13776 35448 13776 0 _0812_
rlabel metal2 28168 11592 28168 11592 0 _0813_
rlabel metal2 27552 11144 27552 11144 0 _0814_
rlabel metal2 28616 15736 28616 15736 0 _0815_
rlabel metal2 26152 17136 26152 17136 0 _0816_
rlabel metal2 38752 15512 38752 15512 0 _0817_
rlabel metal3 27720 18424 27720 18424 0 _0818_
rlabel metal2 37352 22008 37352 22008 0 _0819_
rlabel metal2 27608 17248 27608 17248 0 _0820_
rlabel metal2 27048 17024 27048 17024 0 _0821_
rlabel metal3 30240 19992 30240 19992 0 _0822_
rlabel metal2 27384 17752 27384 17752 0 _0823_
rlabel metal3 24864 17528 24864 17528 0 _0824_
rlabel metal2 27832 17360 27832 17360 0 _0825_
rlabel metal2 26712 15008 26712 15008 0 _0826_
rlabel metal2 26488 15260 26488 15260 0 _0827_
rlabel metal3 20608 13720 20608 13720 0 _0828_
rlabel metal2 24808 16240 24808 16240 0 _0829_
rlabel metal2 22344 19488 22344 19488 0 _0830_
rlabel metal2 13552 13720 13552 13720 0 _0831_
rlabel metal2 18312 17080 18312 17080 0 _0832_
rlabel metal2 24136 16632 24136 16632 0 _0833_
rlabel metal2 22848 15960 22848 15960 0 _0834_
rlabel metal2 24472 14112 24472 14112 0 _0835_
rlabel metal2 25368 13888 25368 13888 0 _0836_
rlabel metal3 26096 13496 26096 13496 0 _0837_
rlabel metal2 27048 14560 27048 14560 0 _0838_
rlabel metal2 32872 12544 32872 12544 0 _0839_
rlabel metal2 39144 17248 39144 17248 0 _0840_
rlabel metal2 34664 14336 34664 14336 0 _0841_
rlabel metal3 35392 12936 35392 12936 0 _0842_
rlabel metal2 37128 10080 37128 10080 0 _0843_
rlabel metal2 34776 12600 34776 12600 0 _0844_
rlabel metal2 35896 14168 35896 14168 0 _0845_
rlabel metal3 39312 14392 39312 14392 0 _0846_
rlabel metal3 37296 18312 37296 18312 0 _0847_
rlabel metal3 37800 15176 37800 15176 0 _0848_
rlabel metal2 36512 15512 36512 15512 0 _0849_
rlabel metal2 36008 13608 36008 13608 0 _0850_
rlabel metal2 30856 13440 30856 13440 0 _0851_
rlabel metal2 25592 18200 25592 18200 0 _0852_
rlabel metal2 40488 20720 40488 20720 0 _0853_
rlabel metal2 26040 18256 26040 18256 0 _0854_
rlabel metal2 34832 18312 34832 18312 0 _0855_
rlabel metal2 34328 14112 34328 14112 0 _0856_
rlabel metal2 34104 18200 34104 18200 0 _0857_
rlabel metal3 33544 16968 33544 16968 0 _0858_
rlabel metal2 33320 13048 33320 13048 0 _0859_
rlabel metal2 29960 14000 29960 14000 0 _0860_
rlabel metal2 28896 7672 28896 7672 0 _0861_
rlabel metal2 25592 22736 25592 22736 0 _0862_
rlabel metal3 23184 15064 23184 15064 0 _0863_
rlabel metal2 28504 13832 28504 13832 0 _0864_
rlabel metal2 28840 12600 28840 12600 0 _0865_
rlabel metal2 29288 13384 29288 13384 0 _0866_
rlabel metal2 28336 14504 28336 14504 0 _0867_
rlabel metal2 28224 18200 28224 18200 0 _0868_
rlabel metal2 27720 28952 27720 28952 0 _0869_
rlabel metal3 27440 23800 27440 23800 0 _0870_
rlabel metal2 25816 17136 25816 17136 0 _0871_
rlabel metal2 25480 15344 25480 15344 0 _0872_
rlabel metal2 15176 11312 15176 11312 0 _0873_
rlabel metal2 23968 12376 23968 12376 0 _0874_
rlabel metal2 23912 6384 23912 6384 0 _0875_
rlabel metal2 25032 16408 25032 16408 0 _0876_
rlabel metal2 24640 16072 24640 16072 0 _0877_
rlabel metal3 24416 13496 24416 13496 0 _0878_
rlabel metal3 25032 15288 25032 15288 0 _0879_
rlabel metal2 25368 15148 25368 15148 0 _0880_
rlabel metal3 33208 22120 33208 22120 0 _0881_
rlabel metal2 27048 18368 27048 18368 0 _0882_
rlabel metal2 26432 17080 26432 17080 0 _0883_
rlabel metal2 27832 19488 27832 19488 0 _0884_
rlabel metal2 26264 17864 26264 17864 0 _0885_
rlabel metal2 26040 17136 26040 17136 0 _0886_
rlabel metal2 26152 16632 26152 16632 0 _0887_
rlabel metal2 24024 13160 24024 13160 0 _0888_
rlabel metal3 24976 19992 24976 19992 0 _0889_
rlabel metal2 24808 18032 24808 18032 0 _0890_
rlabel metal2 25536 17080 25536 17080 0 _0891_
rlabel metal2 24808 12768 24808 12768 0 _0892_
rlabel metal2 25816 13552 25816 13552 0 _0893_
rlabel metal2 27496 14000 27496 14000 0 _0894_
rlabel metal2 40040 18312 40040 18312 0 _0895_
rlabel metal2 35168 16632 35168 16632 0 _0896_
rlabel metal2 35392 12264 35392 12264 0 _0897_
rlabel metal2 35896 11256 35896 11256 0 _0898_
rlabel metal2 35896 12264 35896 12264 0 _0899_
rlabel metal2 42168 13440 42168 13440 0 _0900_
rlabel metal2 37352 20104 37352 20104 0 _0901_
rlabel metal2 37072 12040 37072 12040 0 _0902_
rlabel metal3 36064 13496 36064 13496 0 _0903_
rlabel metal2 35224 12656 35224 12656 0 _0904_
rlabel metal2 35560 12488 35560 12488 0 _0905_
rlabel metal2 40152 21672 40152 21672 0 _0906_
rlabel metal2 33488 16184 33488 16184 0 _0907_
rlabel metal2 32088 14112 32088 14112 0 _0908_
rlabel metal2 32536 19936 32536 19936 0 _0909_
rlabel metal3 32928 15960 32928 15960 0 _0910_
rlabel metal2 32424 14000 32424 14000 0 _0911_
rlabel metal2 30184 14560 30184 14560 0 _0912_
rlabel metal2 24584 10024 24584 10024 0 _0913_
rlabel metal2 24024 22008 24024 22008 0 _0914_
rlabel metal3 18256 16296 18256 16296 0 _0915_
rlabel metal2 24360 15792 24360 15792 0 _0916_
rlabel metal2 26376 13216 26376 13216 0 _0917_
rlabel metal2 26768 13160 26768 13160 0 _0918_
rlabel metal2 28392 14000 28392 14000 0 _0919_
rlabel metal2 26992 23800 26992 23800 0 _0920_
rlabel metal2 27216 28616 27216 28616 0 _0921_
rlabel metal2 14728 28784 14728 28784 0 _0922_
rlabel metal2 15960 29960 15960 29960 0 _0923_
rlabel metal2 6216 36904 6216 36904 0 _0924_
rlabel metal3 10136 35672 10136 35672 0 _0925_
rlabel metal2 11144 37856 11144 37856 0 _0926_
rlabel metal2 14672 42056 14672 42056 0 _0927_
rlabel metal2 15960 40880 15960 40880 0 _0928_
rlabel metal2 11760 35672 11760 35672 0 _0929_
rlabel metal2 7672 37352 7672 37352 0 _0930_
rlabel metal2 12152 36176 12152 36176 0 _0931_
rlabel metal2 13384 29904 13384 29904 0 _0932_
rlabel metal2 14840 37520 14840 37520 0 _0933_
rlabel metal2 15344 38920 15344 38920 0 _0934_
rlabel metal2 15904 31192 15904 31192 0 _0935_
rlabel metal2 16072 43512 16072 43512 0 _0936_
rlabel metal2 16296 44688 16296 44688 0 _0937_
rlabel metal2 30184 46200 30184 46200 0 _0938_
rlabel metal3 31024 38920 31024 38920 0 _0939_
rlabel metal3 17248 32760 17248 32760 0 _0940_
rlabel metal2 6832 21784 6832 21784 0 _0941_
rlabel metal2 18648 31808 18648 31808 0 _0942_
rlabel metal3 18816 31528 18816 31528 0 _0943_
rlabel metal2 3080 37184 3080 37184 0 _0944_
rlabel metal2 18536 40600 18536 40600 0 _0945_
rlabel metal2 5544 39032 5544 39032 0 _0946_
rlabel metal3 9520 38360 9520 38360 0 _0947_
rlabel metal2 21560 36568 21560 36568 0 _0948_
rlabel metal3 10472 34776 10472 34776 0 _0949_
rlabel metal2 10192 34328 10192 34328 0 _0950_
rlabel metal2 18424 30464 18424 30464 0 _0951_
rlabel metal2 7336 30576 7336 30576 0 _0952_
rlabel metal2 31976 43176 31976 43176 0 _0953_
rlabel metal2 15904 26264 15904 26264 0 _0954_
rlabel metal2 19880 30520 19880 30520 0 _0955_
rlabel metal2 20216 30800 20216 30800 0 _0956_
rlabel metal2 20552 30800 20552 30800 0 _0957_
rlabel metal2 16632 41048 16632 41048 0 _0958_
rlabel metal2 19040 34104 19040 34104 0 _0959_
rlabel metal2 18144 43624 18144 43624 0 _0960_
rlabel metal2 18424 54936 18424 54936 0 _0961_
rlabel metal2 17360 55496 17360 55496 0 _0962_
rlabel metal2 17192 54600 17192 54600 0 _0963_
rlabel metal2 23800 44520 23800 44520 0 _0964_
rlabel metal2 19320 39816 19320 39816 0 _0965_
rlabel metal2 18704 45976 18704 45976 0 _0966_
rlabel metal2 21448 28952 21448 28952 0 _0967_
rlabel metal3 17080 35560 17080 35560 0 _0968_
rlabel metal2 10976 37240 10976 37240 0 _0969_
rlabel metal3 21056 35560 21056 35560 0 _0970_
rlabel metal2 4312 38864 4312 38864 0 _0971_
rlabel metal2 9912 36736 9912 36736 0 _0972_
rlabel metal2 10864 38808 10864 38808 0 _0973_
rlabel metal2 10304 37128 10304 37128 0 _0974_
rlabel metal2 14728 36400 14728 36400 0 _0975_
rlabel metal3 14616 33320 14616 33320 0 _0976_
rlabel metal2 9352 24192 9352 24192 0 _0977_
rlabel metal2 9688 24976 9688 24976 0 _0978_
rlabel metal3 9128 26264 9128 26264 0 _0979_
rlabel metal2 11200 24920 11200 24920 0 _0980_
rlabel metal2 14168 22960 14168 22960 0 _0981_
rlabel metal2 7224 25816 7224 25816 0 _0982_
rlabel metal3 9016 25592 9016 25592 0 _0983_
rlabel metal2 11424 27272 11424 27272 0 _0984_
rlabel metal3 18368 24696 18368 24696 0 _0985_
rlabel metal2 12376 24640 12376 24640 0 _0986_
rlabel metal2 14560 26488 14560 26488 0 _0987_
rlabel metal3 13832 24808 13832 24808 0 _0988_
rlabel metal2 12880 23128 12880 23128 0 _0989_
rlabel metal2 7896 23632 7896 23632 0 _0990_
rlabel metal2 10808 22960 10808 22960 0 _0991_
rlabel metal2 13384 25424 13384 25424 0 _0992_
rlabel metal2 10248 27384 10248 27384 0 _0993_
rlabel metal3 12712 27048 12712 27048 0 _0994_
rlabel metal3 13384 28616 13384 28616 0 _0995_
rlabel metal3 12936 34664 12936 34664 0 _0996_
rlabel metal2 12152 33656 12152 33656 0 _0997_
rlabel metal2 12264 32424 12264 32424 0 _0998_
rlabel metal2 25256 39200 25256 39200 0 _0999_
rlabel metal3 15568 41160 15568 41160 0 _1000_
rlabel metal2 15064 41832 15064 41832 0 _1001_
rlabel metal2 23464 39872 23464 39872 0 _1002_
rlabel metal2 11424 38808 11424 38808 0 _1003_
rlabel metal2 21112 38920 21112 38920 0 _1004_
rlabel metal2 20664 38808 20664 38808 0 _1005_
rlabel metal2 23128 33656 23128 33656 0 _1006_
rlabel metal3 20552 34104 20552 34104 0 _1007_
rlabel metal2 13552 33320 13552 33320 0 _1008_
rlabel metal2 15624 30464 15624 30464 0 _1009_
rlabel metal3 15512 30184 15512 30184 0 _1010_
rlabel metal3 14616 30408 14616 30408 0 _1011_
rlabel metal2 14168 32032 14168 32032 0 _1012_
rlabel metal2 13832 31248 13832 31248 0 _1013_
rlabel metal2 34328 52360 34328 52360 0 _1014_
rlabel metal2 29736 51072 29736 51072 0 _1015_
rlabel metal2 28952 52584 28952 52584 0 _1016_
rlabel metal3 35336 52248 35336 52248 0 _1017_
rlabel metal2 29960 50568 29960 50568 0 _1018_
rlabel metal2 22960 50344 22960 50344 0 _1019_
rlabel metal2 23912 50148 23912 50148 0 _1020_
rlabel metal2 23240 51968 23240 51968 0 _1021_
rlabel metal2 23632 51352 23632 51352 0 _1022_
rlabel metal2 24808 50148 24808 50148 0 _1023_
rlabel metal2 22568 50148 22568 50148 0 _1024_
rlabel metal2 22792 51408 22792 51408 0 _1025_
rlabel metal2 25592 51408 25592 51408 0 _1026_
rlabel metal3 26572 49000 26572 49000 0 _1027_
rlabel metal3 28896 48776 28896 48776 0 _1028_
rlabel metal2 26208 48440 26208 48440 0 _1029_
rlabel metal2 26712 48440 26712 48440 0 _1030_
rlabel metal2 24024 52808 24024 52808 0 _1031_
rlabel metal2 26712 49784 26712 49784 0 _1032_
rlabel metal2 28000 51128 28000 51128 0 _1033_
rlabel metal3 29624 49112 29624 49112 0 _1034_
rlabel metal2 32760 49336 32760 49336 0 _1035_
rlabel metal2 31976 51464 31976 51464 0 _1036_
rlabel metal2 27160 50512 27160 50512 0 _1037_
rlabel metal3 28000 50568 28000 50568 0 _1038_
rlabel metal2 26936 52472 26936 52472 0 _1039_
rlabel metal3 29400 49672 29400 49672 0 _1040_
rlabel metal2 31696 51352 31696 51352 0 _1041_
rlabel metal2 31920 51128 31920 51128 0 _1042_
rlabel metal2 26824 49448 26824 49448 0 _1043_
rlabel metal3 30296 48328 30296 48328 0 _1044_
rlabel metal2 31192 49840 31192 49840 0 _1045_
rlabel metal2 29624 49616 29624 49616 0 _1046_
rlabel metal2 31472 52136 31472 52136 0 _1047_
rlabel metal2 32648 50064 32648 50064 0 _1048_
rlabel metal3 30856 53032 30856 53032 0 _1049_
rlabel metal2 28336 51352 28336 51352 0 _1050_
rlabel metal2 27776 51464 27776 51464 0 _1051_
rlabel metal2 26208 50120 26208 50120 0 _1052_
rlabel metal2 26600 49728 26600 49728 0 _1053_
rlabel metal2 27496 50960 27496 50960 0 _1054_
rlabel metal2 27048 50792 27048 50792 0 _1055_
rlabel metal3 27804 51464 27804 51464 0 _1056_
rlabel metal3 28616 52920 28616 52920 0 _1057_
rlabel metal2 29624 53312 29624 53312 0 _1058_
rlabel metal2 29400 53592 29400 53592 0 _1059_
rlabel metal2 28616 50904 28616 50904 0 _1060_
rlabel metal2 29344 50344 29344 50344 0 _1061_
rlabel metal3 30184 50456 30184 50456 0 _1062_
rlabel metal2 31976 47992 31976 47992 0 _1063_
rlabel metal2 30072 49728 30072 49728 0 _1064_
rlabel metal2 30408 51016 30408 51016 0 _1065_
rlabel metal3 29120 52360 29120 52360 0 _1066_
rlabel metal3 28896 52696 28896 52696 0 _1067_
rlabel metal2 29736 52360 29736 52360 0 _1068_
rlabel metal2 30520 53424 30520 53424 0 _1069_
rlabel metal2 27384 51576 27384 51576 0 _1070_
rlabel metal2 30296 52528 30296 52528 0 _1071_
rlabel metal2 31024 52696 31024 52696 0 _1072_
rlabel metal2 31304 53816 31304 53816 0 _1073_
rlabel metal2 33096 50176 33096 50176 0 _1074_
rlabel metal3 30520 50568 30520 50568 0 _1075_
rlabel metal2 32536 51016 32536 51016 0 _1076_
rlabel metal2 33208 51744 33208 51744 0 _1077_
rlabel metal2 33096 51016 33096 51016 0 _1078_
rlabel metal2 19208 26320 19208 26320 0 _1079_
rlabel metal2 15736 40152 15736 40152 0 _1080_
rlabel metal3 16016 34552 16016 34552 0 _1081_
rlabel metal3 16688 37464 16688 37464 0 _1082_
rlabel metal3 16296 32648 16296 32648 0 _1083_
rlabel metal2 15568 36456 15568 36456 0 _1084_
rlabel metal3 18928 25368 18928 25368 0 _1085_
rlabel metal2 47488 37128 47488 37128 0 _1086_
rlabel metal3 16072 35672 16072 35672 0 _1087_
rlabel metal2 19992 34832 19992 34832 0 _1088_
rlabel metal2 18648 30800 18648 30800 0 _1089_
rlabel metal2 19208 28896 19208 28896 0 _1090_
rlabel metal2 13832 30464 13832 30464 0 _1091_
rlabel metal2 25480 45696 25480 45696 0 _1092_
rlabel metal2 6552 31640 6552 31640 0 _1093_
rlabel metal2 19376 32648 19376 32648 0 _1094_
rlabel metal2 17864 29960 17864 29960 0 _1095_
rlabel metal3 17584 33096 17584 33096 0 _1096_
rlabel metal2 17528 26628 17528 26628 0 _1097_
rlabel metal2 17416 25760 17416 25760 0 _1098_
rlabel metal2 18424 35504 18424 35504 0 _1099_
rlabel metal2 18312 30184 18312 30184 0 _1100_
rlabel metal3 18088 38808 18088 38808 0 _1101_
rlabel metal2 12264 30576 12264 30576 0 _1102_
rlabel metal2 12712 29680 12712 29680 0 _1103_
rlabel metal2 15848 25480 15848 25480 0 _1104_
rlabel metal3 16912 21672 16912 21672 0 _1105_
rlabel metal2 30744 25928 30744 25928 0 _1106_
rlabel metal2 31304 22680 31304 22680 0 _1107_
rlabel metal2 22232 8960 22232 8960 0 _1108_
rlabel metal3 41440 12264 41440 12264 0 _1109_
rlabel metal2 16520 22008 16520 22008 0 _1110_
rlabel metal2 19208 19600 19208 19600 0 _1111_
rlabel metal2 15400 22568 15400 22568 0 _1112_
rlabel metal2 19208 21224 19208 21224 0 _1113_
rlabel metal3 20048 24696 20048 24696 0 _1114_
rlabel metal2 16800 23128 16800 23128 0 _1115_
rlabel metal2 18368 20104 18368 20104 0 _1116_
rlabel metal3 39424 12824 39424 12824 0 _1117_
rlabel metal2 18984 23184 18984 23184 0 _1118_
rlabel metal2 20776 18648 20776 18648 0 _1119_
rlabel metal2 26712 19432 26712 19432 0 _1120_
rlabel metal2 42672 12264 42672 12264 0 _1121_
rlabel metal2 42280 11256 42280 11256 0 _1122_
rlabel metal2 31976 23072 31976 23072 0 _1123_
rlabel metal2 38808 7392 38808 7392 0 _1124_
rlabel metal2 39928 8064 39928 8064 0 _1125_
rlabel metal2 41944 14000 41944 14000 0 _1126_
rlabel metal2 21672 23016 21672 23016 0 _1127_
rlabel metal2 22008 22736 22008 22736 0 _1128_
rlabel metal2 21336 14952 21336 14952 0 _1129_
rlabel metal2 38696 12040 38696 12040 0 _1130_
rlabel via2 43848 12936 43848 12936 0 _1131_
rlabel metal3 44520 12376 44520 12376 0 _1132_
rlabel metal2 44744 14000 44744 14000 0 _1133_
rlabel metal2 31640 19656 31640 19656 0 _1134_
rlabel metal2 12040 14224 12040 14224 0 _1135_
rlabel metal3 16464 19544 16464 19544 0 _1136_
rlabel metal2 13832 18312 13832 18312 0 _1137_
rlabel metal3 19712 17752 19712 17752 0 _1138_
rlabel metal2 17528 17920 17528 17920 0 _1139_
rlabel metal2 14168 15960 14168 15960 0 _1140_
rlabel metal2 20776 23408 20776 23408 0 _1141_
rlabel metal2 19656 17192 19656 17192 0 _1142_
rlabel metal2 22848 10472 22848 10472 0 _1143_
rlabel metal2 39256 12656 39256 12656 0 _1144_
rlabel metal2 38472 11256 38472 11256 0 _1145_
rlabel metal2 39928 14168 39928 14168 0 _1146_
rlabel metal2 17528 19992 17528 19992 0 _1147_
rlabel metal2 38808 19992 38808 19992 0 _1148_
rlabel metal2 39592 8260 39592 8260 0 _1149_
rlabel metal2 40264 9464 40264 9464 0 _1150_
rlabel metal2 39480 7784 39480 7784 0 _1151_
rlabel metal2 21280 22568 21280 22568 0 _1152_
rlabel metal2 22680 21504 22680 21504 0 _1153_
rlabel metal2 38696 20132 38696 20132 0 _1154_
rlabel metal2 39032 20048 39032 20048 0 _1155_
rlabel metal2 39368 21616 39368 21616 0 _1156_
rlabel metal2 40320 18424 40320 18424 0 _1157_
rlabel metal2 39592 20356 39592 20356 0 _1158_
rlabel metal2 39480 17920 39480 17920 0 _1159_
rlabel metal3 29904 5992 29904 5992 0 _1160_
rlabel metal2 36008 7504 36008 7504 0 _1161_
rlabel metal2 36960 4424 36960 4424 0 _1162_
rlabel metal2 34328 5880 34328 5880 0 _1163_
rlabel metal2 34608 3528 34608 3528 0 _1164_
rlabel metal2 25928 10080 25928 10080 0 _1165_
rlabel metal2 20104 24528 20104 24528 0 _1166_
rlabel metal2 21112 21280 21112 21280 0 _1167_
rlabel metal2 21448 23408 21448 23408 0 _1168_
rlabel metal3 32648 23240 32648 23240 0 _1169_
rlabel metal2 34664 19768 34664 19768 0 _1170_
rlabel metal2 32144 24136 32144 24136 0 _1171_
rlabel metal3 16856 48216 16856 48216 0 _1172_
rlabel metal3 19488 48776 19488 48776 0 _1173_
rlabel metal2 33096 8400 33096 8400 0 _1174_
rlabel metal3 31640 8120 31640 8120 0 _1175_
rlabel metal3 31696 6552 31696 6552 0 _1176_
rlabel metal2 39144 21168 39144 21168 0 _1177_
rlabel metal2 39816 21504 39816 21504 0 _1178_
rlabel metal2 40152 20832 40152 20832 0 _1179_
rlabel metal3 33544 5992 33544 5992 0 _1180_
rlabel metal2 30968 5880 30968 5880 0 _1181_
rlabel metal2 30184 5376 30184 5376 0 _1182_
rlabel metal2 15176 20524 15176 20524 0 _1183_
rlabel metal3 17640 20664 17640 20664 0 _1184_
rlabel metal2 27048 8232 27048 8232 0 _1185_
rlabel metal2 26208 5880 26208 5880 0 _1186_
rlabel metal2 27384 4200 27384 4200 0 _1187_
rlabel metal2 14952 9408 14952 9408 0 _1188_
rlabel metal2 19096 21616 19096 21616 0 _1189_
rlabel metal2 18088 9856 18088 9856 0 _1190_
rlabel metal2 14840 9744 14840 9744 0 _1191_
rlabel metal3 12880 9688 12880 9688 0 _1192_
rlabel metal2 21784 5824 21784 5824 0 _1193_
rlabel metal2 13832 7336 13832 7336 0 _1194_
rlabel metal2 14392 29064 14392 29064 0 _1195_
rlabel metal2 16184 29176 16184 29176 0 _1196_
rlabel metal2 15176 29568 15176 29568 0 _1197_
rlabel metal2 14728 27496 14728 27496 0 _1198_
rlabel metal2 14840 26264 14840 26264 0 _1199_
rlabel metal3 10528 27608 10528 27608 0 _1200_
rlabel metal2 14952 25872 14952 25872 0 _1201_
rlabel metal2 7000 24920 7000 24920 0 _1202_
rlabel metal2 7336 24136 7336 24136 0 _1203_
rlabel metal2 8064 23128 8064 23128 0 _1204_
rlabel metal3 6776 23352 6776 23352 0 _1205_
rlabel metal2 5992 25928 5992 25928 0 _1206_
rlabel metal2 6552 22064 6552 22064 0 _1207_
rlabel metal3 41216 30072 41216 30072 0 _1208_
rlabel metal2 8904 26712 8904 26712 0 _1209_
rlabel metal2 24360 27552 24360 27552 0 _1210_
rlabel metal2 18648 48216 18648 48216 0 _1211_
rlabel metal2 21952 47656 21952 47656 0 _1212_
rlabel metal2 20272 47656 20272 47656 0 _1213_
rlabel metal2 20552 48832 20552 48832 0 _1214_
rlabel metal3 21672 49000 21672 49000 0 _1215_
rlabel metal2 22064 49784 22064 49784 0 _1216_
rlabel metal2 21168 47992 21168 47992 0 _1217_
rlabel metal2 18928 49224 18928 49224 0 _1218_
rlabel metal2 19096 49056 19096 49056 0 _1219_
rlabel metal2 22120 49112 22120 49112 0 _1220_
rlabel metal3 19824 49784 19824 49784 0 _1221_
rlabel metal2 19208 50092 19208 50092 0 _1222_
rlabel metal2 16464 48216 16464 48216 0 _1223_
rlabel metal2 17472 50008 17472 50008 0 _1224_
rlabel metal2 16688 48216 16688 48216 0 _1225_
rlabel metal2 16632 52080 16632 52080 0 _1226_
rlabel metal2 16856 51688 16856 51688 0 _1227_
rlabel metal2 16128 52024 16128 52024 0 _1228_
rlabel metal2 16184 52472 16184 52472 0 _1229_
rlabel metal2 17976 52584 17976 52584 0 _1230_
rlabel metal2 19432 52584 19432 52584 0 _1231_
rlabel metal2 16296 50680 16296 50680 0 _1232_
rlabel metal2 17640 51632 17640 51632 0 _1233_
rlabel metal2 16912 50792 16912 50792 0 _1234_
rlabel metal2 39816 27944 39816 27944 0 _1235_
rlabel metal2 37184 26264 37184 26264 0 _1236_
rlabel metal2 37352 26376 37352 26376 0 _1237_
rlabel metal2 41216 26264 41216 26264 0 _1238_
rlabel metal2 41496 27496 41496 27496 0 _1239_
rlabel metal2 43960 35056 43960 35056 0 _1240_
rlabel metal2 41328 26488 41328 26488 0 _1241_
rlabel metal2 38920 29400 38920 29400 0 _1242_
rlabel metal2 42000 28616 42000 28616 0 _1243_
rlabel metal2 37688 28336 37688 28336 0 _1244_
rlabel metal2 38920 28728 38920 28728 0 _1245_
rlabel metal2 39704 29064 39704 29064 0 _1246_
rlabel metal3 41384 29400 41384 29400 0 _1247_
rlabel metal2 40376 29904 40376 29904 0 _1248_
rlabel metal2 38808 32144 38808 32144 0 _1249_
rlabel metal2 40264 30688 40264 30688 0 _1250_
rlabel metal2 34384 29512 34384 29512 0 _1251_
rlabel metal2 38920 31360 38920 31360 0 _1252_
rlabel metal3 40544 31416 40544 31416 0 _1253_
rlabel metal2 39480 30464 39480 30464 0 _1254_
rlabel metal2 39872 28616 39872 28616 0 _1255_
rlabel metal2 40824 28112 40824 28112 0 _1256_
rlabel metal3 42056 31080 42056 31080 0 _1257_
rlabel metal3 41664 31192 41664 31192 0 _1258_
rlabel metal2 41048 31640 41048 31640 0 _1259_
rlabel metal2 41888 31080 41888 31080 0 _1260_
rlabel metal2 42504 36848 42504 36848 0 _1261_
rlabel metal2 35784 32200 35784 32200 0 _1262_
rlabel metal2 34272 44296 34272 44296 0 _1263_
rlabel metal3 35560 36456 35560 36456 0 _1264_
rlabel metal3 34608 35784 34608 35784 0 _1265_
rlabel metal2 40712 34832 40712 34832 0 _1266_
rlabel metal2 35784 36120 35784 36120 0 _1267_
rlabel metal2 45080 34944 45080 34944 0 _1268_
rlabel metal2 45304 38024 45304 38024 0 _1269_
rlabel metal2 44632 47600 44632 47600 0 _1270_
rlabel metal2 47208 44464 47208 44464 0 _1271_
rlabel metal2 43064 48972 43064 48972 0 _1272_
rlabel metal2 44968 42784 44968 42784 0 _1273_
rlabel metal3 47040 42616 47040 42616 0 _1274_
rlabel metal2 49000 43512 49000 43512 0 _1275_
rlabel metal2 48776 47768 48776 47768 0 _1276_
rlabel metal2 49000 47880 49000 47880 0 _1277_
rlabel metal3 41160 46648 41160 46648 0 _1278_
rlabel metal2 44912 47208 44912 47208 0 _1279_
rlabel metal2 49336 45864 49336 45864 0 _1280_
rlabel metal2 45080 47152 45080 47152 0 _1281_
rlabel metal2 49560 44632 49560 44632 0 _1282_
rlabel metal2 44968 52528 44968 52528 0 _1283_
rlabel metal2 44464 48216 44464 48216 0 _1284_
rlabel metal2 44296 45360 44296 45360 0 _1285_
rlabel metal2 48552 46200 48552 46200 0 _1286_
rlabel metal2 43400 48720 43400 48720 0 _1287_
rlabel metal3 44968 45136 44968 45136 0 _1288_
rlabel metal2 42168 46032 42168 46032 0 _1289_
rlabel metal2 42168 36904 42168 36904 0 _1290_
rlabel metal2 42280 41944 42280 41944 0 _1291_
rlabel metal2 42616 37856 42616 37856 0 _1292_
rlabel metal2 42056 43232 42056 43232 0 _1293_
rlabel metal2 36680 43848 36680 43848 0 _1294_
rlabel metal2 43008 45080 43008 45080 0 _1295_
rlabel metal2 40040 47152 40040 47152 0 _1296_
rlabel metal2 42672 45864 42672 45864 0 _1297_
rlabel metal2 43512 45472 43512 45472 0 _1298_
rlabel metal2 43008 45304 43008 45304 0 _1299_
rlabel metal3 43512 45080 43512 45080 0 _1300_
rlabel metal2 44184 45024 44184 45024 0 _1301_
rlabel metal2 44520 44632 44520 44632 0 _1302_
rlabel metal2 45752 46536 45752 46536 0 _1303_
rlabel metal2 49672 47656 49672 47656 0 _1304_
rlabel metal2 45640 46144 45640 46144 0 _1305_
rlabel metal2 46088 44800 46088 44800 0 _1306_
rlabel metal3 49448 43456 49448 43456 0 _1307_
rlabel metal3 48776 42168 48776 42168 0 _1308_
rlabel metal2 48104 44016 48104 44016 0 _1309_
rlabel metal2 46200 43792 46200 43792 0 _1310_
rlabel metal3 54880 39480 54880 39480 0 _1311_
rlabel metal3 52192 36232 52192 36232 0 _1312_
rlabel metal2 50456 35728 50456 35728 0 _1313_
rlabel metal2 50064 36456 50064 36456 0 _1314_
rlabel metal3 42560 42728 42560 42728 0 _1315_
rlabel metal2 43848 37520 43848 37520 0 _1316_
rlabel metal3 42840 42616 42840 42616 0 _1317_
rlabel metal2 43176 42840 43176 42840 0 _1318_
rlabel metal2 45192 42896 45192 42896 0 _1319_
rlabel metal2 43792 42728 43792 42728 0 _1320_
rlabel metal2 43904 42952 43904 42952 0 _1321_
rlabel metal2 45864 43456 45864 43456 0 _1322_
rlabel metal3 49672 40488 49672 40488 0 _1323_
rlabel metal2 48776 40768 48776 40768 0 _1324_
rlabel metal2 45192 41384 45192 41384 0 _1325_
rlabel metal2 43064 44576 43064 44576 0 _1326_
rlabel metal2 48888 45360 48888 45360 0 _1327_
rlabel metal2 40096 35784 40096 35784 0 _1328_
rlabel metal2 39816 34440 39816 34440 0 _1329_
rlabel metal3 39816 31752 39816 31752 0 _1330_
rlabel metal2 39816 30520 39816 30520 0 _1331_
rlabel metal2 39984 31192 39984 31192 0 _1332_
rlabel metal2 40376 31892 40376 31892 0 _1333_
rlabel metal2 41496 40432 41496 40432 0 _1334_
rlabel metal3 44968 40376 44968 40376 0 _1335_
rlabel metal2 44968 40040 44968 40040 0 _1336_
rlabel metal2 44352 38584 44352 38584 0 _1337_
rlabel metal2 46368 37800 46368 37800 0 _1338_
rlabel metal2 46872 36848 46872 36848 0 _1339_
rlabel metal2 48440 38360 48440 38360 0 _1340_
rlabel metal3 39312 20328 39312 20328 0 clknet_0_wb_clk_i
rlabel metal2 5880 13720 5880 13720 0 clknet_4_0_0_wb_clk_i
rlabel metal2 44912 11144 44912 11144 0 clknet_4_10_0_wb_clk_i
rlabel metal2 44072 29120 44072 29120 0 clknet_4_11_0_wb_clk_i
rlabel metal2 35224 46032 35224 46032 0 clknet_4_12_0_wb_clk_i
rlabel metal2 31864 54096 31864 54096 0 clknet_4_13_0_wb_clk_i
rlabel metal3 46088 32536 46088 32536 0 clknet_4_14_0_wb_clk_i
rlabel metal2 48664 46704 48664 46704 0 clknet_4_15_0_wb_clk_i
rlabel metal2 15512 17976 15512 17976 0 clknet_4_1_0_wb_clk_i
rlabel metal2 23352 15848 23352 15848 0 clknet_4_2_0_wb_clk_i
rlabel metal2 15960 20440 15960 20440 0 clknet_4_3_0_wb_clk_i
rlabel metal2 1848 39984 1848 39984 0 clknet_4_4_0_wb_clk_i
rlabel metal2 2296 46312 2296 46312 0 clknet_4_5_0_wb_clk_i
rlabel metal2 19712 43400 19712 43400 0 clknet_4_6_0_wb_clk_i
rlabel metal2 13608 53648 13608 53648 0 clknet_4_7_0_wb_clk_i
rlabel metal2 36288 15848 36288 15848 0 clknet_4_8_0_wb_clk_i
rlabel metal2 36512 26488 36512 26488 0 clknet_4_9_0_wb_clk_i
rlabel metal3 18536 53816 18536 53816 0 io_in[10]
rlabel metal2 21112 54992 21112 54992 0 io_in[11]
rlabel metal3 40544 56280 40544 56280 0 io_in[26]
rlabel metal3 41664 56056 41664 56056 0 io_in[27]
rlabel metal2 15512 56336 15512 56336 0 io_in[8]
rlabel metal2 14784 55384 14784 55384 0 io_in[9]
rlabel metal2 22008 57610 22008 57610 0 io_out[12]
rlabel metal2 23408 54712 23408 54712 0 io_out[13]
rlabel metal2 23688 56392 23688 56392 0 io_out[14]
rlabel metal2 26712 55664 26712 55664 0 io_out[15]
rlabel metal3 28504 55384 28504 55384 0 io_out[16]
rlabel metal2 29400 56280 29400 56280 0 io_out[17]
rlabel metal3 30576 56280 30576 56280 0 io_out[18]
rlabel metal2 31416 57778 31416 57778 0 io_out[19]
rlabel metal2 34664 56504 34664 56504 0 io_out[20]
rlabel metal2 35112 55412 35112 55412 0 io_out[21]
rlabel metal2 36792 56448 36792 56448 0 io_out[22]
rlabel metal2 38024 56504 38024 56504 0 io_out[23]
rlabel metal2 38136 58114 38136 58114 0 io_out[24]
rlabel metal3 40096 55384 40096 55384 0 io_out[25]
rlabel metal2 20328 54824 20328 54824 0 net1
rlabel metal2 21784 44296 21784 44296 0 net10
rlabel metal2 21448 42224 21448 42224 0 net11
rlabel metal3 30632 55048 30632 55048 0 net12
rlabel metal2 27496 56000 27496 56000 0 net13
rlabel metal3 29456 55720 29456 55720 0 net14
rlabel metal3 30632 54376 30632 54376 0 net15
rlabel metal2 34328 55720 34328 55720 0 net16
rlabel metal2 34776 54544 34776 54544 0 net17
rlabel metal2 36064 52808 36064 52808 0 net18
rlabel metal2 36456 51856 36456 51856 0 net19
rlabel metal2 16632 54656 16632 54656 0 net2
rlabel metal2 38584 55216 38584 55216 0 net20
rlabel metal2 40264 55328 40264 55328 0 net21
rlabel metal2 21560 56994 21560 56994 0 net22
rlabel metal2 22960 54712 22960 54712 0 net23
rlabel metal2 24584 56168 24584 56168 0 net24
rlabel metal2 25368 55328 25368 55328 0 net25
rlabel metal2 27160 54516 27160 54516 0 net26
rlabel metal2 28504 54516 28504 54516 0 net27
rlabel metal2 28672 54712 28672 54712 0 net28
rlabel metal2 30968 57218 30968 57218 0 net29
rlabel metal2 34216 52752 34216 52752 0 net3
rlabel metal2 32704 57400 32704 57400 0 net30
rlabel metal3 34496 56280 34496 56280 0 net31
rlabel metal3 35560 55160 35560 55160 0 net32
rlabel metal2 36344 57778 36344 57778 0 net33
rlabel metal2 37688 56994 37688 56994 0 net34
rlabel metal2 39200 54712 39200 54712 0 net35
rlabel metal2 6216 57008 6216 57008 0 net36
rlabel metal2 7336 56280 7336 56280 0 net37
rlabel metal2 8624 56280 8624 56280 0 net38
rlabel metal2 10024 56280 10024 56280 0 net39
rlabel metal2 40152 48888 40152 48888 0 net4
rlabel metal2 11256 57778 11256 57778 0 net40
rlabel metal2 12152 57008 12152 57008 0 net41
rlabel metal2 13832 57400 13832 57400 0 net42
rlabel metal2 15064 55300 15064 55300 0 net43
rlabel metal2 16632 57778 16632 57778 0 net44
rlabel metal2 18088 53592 18088 53592 0 net45
rlabel metal2 19824 53592 19824 53592 0 net46
rlabel metal2 20664 57218 20664 57218 0 net47
rlabel metal2 41664 55160 41664 55160 0 net48
rlabel metal2 42672 55160 42672 55160 0 net49
rlabel metal3 19488 55944 19488 55944 0 net5
rlabel metal2 44072 56616 44072 56616 0 net50
rlabel metal2 44968 56280 44968 56280 0 net51
rlabel metal2 46312 56280 46312 56280 0 net52
rlabel metal2 47880 57008 47880 57008 0 net53
rlabel metal2 49000 56280 49000 56280 0 net54
rlabel metal2 50232 57778 50232 57778 0 net55
rlabel metal2 51688 56280 51688 56280 0 net56
rlabel metal2 53032 56280 53032 56280 0 net57
rlabel metal2 55048 56560 55048 56560 0 net58
rlabel metal2 55944 57008 55944 57008 0 net59
rlabel metal2 15400 55720 15400 55720 0 net6
rlabel metal2 4984 56392 4984 56392 0 net60
rlabel metal2 6888 55944 6888 55944 0 net61
rlabel metal2 8176 55944 8176 55944 0 net62
rlabel metal2 9576 55944 9576 55944 0 net63
rlabel metal2 10808 57610 10808 57610 0 net64
rlabel metal2 11760 55944 11760 55944 0 net65
rlabel metal2 12600 56392 12600 56392 0 net66
rlabel metal2 13496 56280 13496 56280 0 net67
rlabel metal2 16184 57610 16184 57610 0 net68
rlabel metal2 17752 55216 17752 55216 0 net69
rlabel metal3 7504 56168 7504 56168 0 net7
rlabel metal2 19096 54824 19096 54824 0 net70
rlabel metal2 20776 56280 20776 56280 0 net71
rlabel metal3 41552 55944 41552 55944 0 net72
rlabel metal2 42280 55944 42280 55944 0 net73
rlabel metal2 43624 56280 43624 56280 0 net74
rlabel metal2 44520 55944 44520 55944 0 net75
rlabel metal2 45864 55944 45864 55944 0 net76
rlabel metal2 47264 55944 47264 55944 0 net77
rlabel metal2 48552 55944 48552 55944 0 net78
rlabel metal2 49896 55944 49896 55944 0 net79
rlabel metal2 19544 44800 19544 44800 0 net8
rlabel metal2 51240 55944 51240 55944 0 net80
rlabel metal2 52584 55944 52584 55944 0 net81
rlabel metal2 53928 55944 53928 55944 0 net82
rlabel metal2 55328 55944 55328 55944 0 net83
rlabel metal2 24192 44968 24192 44968 0 net9
rlabel metal2 9912 42504 9912 42504 0 simon1.millis_counter\[0\]
rlabel metal2 9968 39592 9968 39592 0 simon1.millis_counter\[1\]
rlabel metal2 10696 36064 10696 36064 0 simon1.millis_counter\[2\]
rlabel metal3 6440 34888 6440 34888 0 simon1.millis_counter\[3\]
rlabel metal2 4592 35672 4592 35672 0 simon1.millis_counter\[4\]
rlabel metal2 6104 35504 6104 35504 0 simon1.millis_counter\[5\]
rlabel metal2 4704 39368 4704 39368 0 simon1.millis_counter\[6\]
rlabel metal2 7336 40320 7336 40320 0 simon1.millis_counter\[7\]
rlabel metal2 15288 42280 15288 42280 0 simon1.millis_counter\[8\]
rlabel metal2 14056 41888 14056 41888 0 simon1.millis_counter\[9\]
rlabel metal2 30520 25928 30520 25928 0 simon1.next_random\[0\]
rlabel metal2 31136 26152 31136 26152 0 simon1.next_random\[1\]
rlabel metal2 39704 27440 39704 27440 0 simon1.play1.freq\[0\]
rlabel metal2 39368 27776 39368 27776 0 simon1.play1.freq\[1\]
rlabel metal3 37128 30072 37128 30072 0 simon1.play1.freq\[2\]
rlabel metal3 37072 32648 37072 32648 0 simon1.play1.freq\[3\]
rlabel metal2 41160 35672 41160 35672 0 simon1.play1.freq\[4\]
rlabel metal2 37688 33488 37688 33488 0 simon1.play1.freq\[5\]
rlabel metal2 34552 36624 34552 36624 0 simon1.play1.freq\[6\]
rlabel metal3 35616 38024 35616 38024 0 simon1.play1.freq\[7\]
rlabel metal2 34328 41440 34328 41440 0 simon1.play1.freq\[8\]
rlabel metal2 31416 44632 31416 44632 0 simon1.play1.freq\[9\]
rlabel metal3 40992 27944 40992 27944 0 simon1.play1.tick_counter\[0\]
rlabel metal2 35896 46312 35896 46312 0 simon1.play1.tick_counter\[10\]
rlabel metal3 36848 48888 36848 48888 0 simon1.play1.tick_counter\[11\]
rlabel metal2 43568 49784 43568 49784 0 simon1.play1.tick_counter\[12\]
rlabel metal2 44016 50120 44016 50120 0 simon1.play1.tick_counter\[13\]
rlabel metal2 44520 53704 44520 53704 0 simon1.play1.tick_counter\[14\]
rlabel metal2 44184 47768 44184 47768 0 simon1.play1.tick_counter\[15\]
rlabel metal2 50232 52640 50232 52640 0 simon1.play1.tick_counter\[16\]
rlabel metal3 49840 52024 49840 52024 0 simon1.play1.tick_counter\[17\]
rlabel metal2 56784 49112 56784 49112 0 simon1.play1.tick_counter\[18\]
rlabel metal2 57064 48384 57064 48384 0 simon1.play1.tick_counter\[19\]
rlabel metal2 40824 26824 40824 26824 0 simon1.play1.tick_counter\[1\]
rlabel metal2 57848 45752 57848 45752 0 simon1.play1.tick_counter\[20\]
rlabel metal3 52024 42728 52024 42728 0 simon1.play1.tick_counter\[21\]
rlabel metal3 46648 41944 46648 41944 0 simon1.play1.tick_counter\[22\]
rlabel metal2 55608 41720 55608 41720 0 simon1.play1.tick_counter\[23\]
rlabel metal2 57960 40432 57960 40432 0 simon1.play1.tick_counter\[24\]
rlabel metal2 56728 38724 56728 38724 0 simon1.play1.tick_counter\[25\]
rlabel metal2 57288 35728 57288 35728 0 simon1.play1.tick_counter\[26\]
rlabel metal2 54712 34832 54712 34832 0 simon1.play1.tick_counter\[27\]
rlabel metal3 48608 35672 48608 35672 0 simon1.play1.tick_counter\[28\]
rlabel metal2 50008 32368 50008 32368 0 simon1.play1.tick_counter\[29\]
rlabel metal2 41272 29064 41272 29064 0 simon1.play1.tick_counter\[2\]
rlabel metal2 51576 30576 51576 30576 0 simon1.play1.tick_counter\[30\]
rlabel metal3 52472 32424 52472 32424 0 simon1.play1.tick_counter\[31\]
rlabel metal3 42504 31864 42504 31864 0 simon1.play1.tick_counter\[3\]
rlabel metal2 41216 36792 41216 36792 0 simon1.play1.tick_counter\[4\]
rlabel metal2 38752 33992 38752 33992 0 simon1.play1.tick_counter\[5\]
rlabel metal2 43960 38192 43960 38192 0 simon1.play1.tick_counter\[6\]
rlabel metal3 35280 39592 35280 39592 0 simon1.play1.tick_counter\[7\]
rlabel metal2 34664 42896 34664 42896 0 simon1.play1.tick_counter\[8\]
rlabel metal2 32536 44688 32536 44688 0 simon1.play1.tick_counter\[9\]
rlabel metal2 24360 54544 24360 54544 0 simon1.score1.active_digit
rlabel metal2 25480 44352 25480 44352 0 simon1.score1.ena
rlabel metal3 23800 47320 23800 47320 0 simon1.score1.inc
rlabel metal2 22680 48888 22680 48888 0 simon1.score1.ones\[0\]
rlabel metal2 21280 49784 21280 49784 0 simon1.score1.ones\[1\]
rlabel metal2 19544 50176 19544 50176 0 simon1.score1.ones\[2\]
rlabel metal2 22400 50008 22400 50008 0 simon1.score1.ones\[3\]
rlabel metal2 17976 49560 17976 49560 0 simon1.score1.tens\[0\]
rlabel metal2 23464 53200 23464 53200 0 simon1.score1.tens\[1\]
rlabel metal2 22008 52416 22008 52416 0 simon1.score1.tens\[2\]
rlabel metal2 18088 51408 18088 51408 0 simon1.score1.tens\[3\]
rlabel metal3 17304 45976 17304 45976 0 simon1.score_rst
rlabel metal2 15288 17808 15288 17808 0 simon1.seq\[0\]\[0\]
rlabel metal3 16520 15176 16520 15176 0 simon1.seq\[0\]\[1\]
rlabel metal2 44632 12600 44632 12600 0 simon1.seq\[10\]\[0\]
rlabel metal3 45752 13720 45752 13720 0 simon1.seq\[10\]\[1\]
rlabel metal2 44296 11536 44296 11536 0 simon1.seq\[11\]\[0\]
rlabel metal2 42504 14952 42504 14952 0 simon1.seq\[11\]\[1\]
rlabel metal2 36288 5880 36288 5880 0 simon1.seq\[12\]\[0\]
rlabel metal2 35000 7168 35000 7168 0 simon1.seq\[12\]\[1\]
rlabel metal2 43848 18368 43848 18368 0 simon1.seq\[13\]\[0\]
rlabel metal2 42056 17360 42056 17360 0 simon1.seq\[13\]\[1\]
rlabel metal2 39480 9968 39480 9968 0 simon1.seq\[14\]\[0\]
rlabel metal2 38248 8176 38248 8176 0 simon1.seq\[14\]\[1\]
rlabel metal2 36232 10640 36232 10640 0 simon1.seq\[15\]\[0\]
rlabel metal3 36680 8344 36680 8344 0 simon1.seq\[15\]\[1\]
rlabel metal2 24472 17304 24472 17304 0 simon1.seq\[16\]\[0\]
rlabel metal2 11144 18032 11144 18032 0 simon1.seq\[16\]\[1\]
rlabel metal2 25592 20496 25592 20496 0 simon1.seq\[17\]\[0\]
rlabel metal2 23240 19936 23240 19936 0 simon1.seq\[17\]\[1\]
rlabel metal2 11480 13776 11480 13776 0 simon1.seq\[18\]\[0\]
rlabel metal2 11200 13048 11200 13048 0 simon1.seq\[18\]\[1\]
rlabel metal2 14616 12824 14616 12824 0 simon1.seq\[19\]\[0\]
rlabel metal2 18088 13328 18088 13328 0 simon1.seq\[19\]\[1\]
rlabel metal2 21784 23408 21784 23408 0 simon1.seq\[1\]\[0\]
rlabel metal2 26936 24304 26936 24304 0 simon1.seq\[1\]\[1\]
rlabel metal3 23520 16520 23520 16520 0 simon1.seq\[20\]\[0\]
rlabel metal3 22344 15176 22344 15176 0 simon1.seq\[20\]\[1\]
rlabel metal2 39928 24304 39928 24304 0 simon1.seq\[21\]\[0\]
rlabel metal2 38248 23800 38248 23800 0 simon1.seq\[21\]\[1\]
rlabel metal2 21784 17976 21784 17976 0 simon1.seq\[22\]\[0\]
rlabel metal2 18368 17752 18368 17752 0 simon1.seq\[22\]\[1\]
rlabel metal2 28616 20496 28616 20496 0 simon1.seq\[23\]\[0\]
rlabel metal2 30968 20496 30968 20496 0 simon1.seq\[23\]\[1\]
rlabel metal2 26488 10024 26488 10024 0 simon1.seq\[24\]\[0\]
rlabel metal2 29176 9296 29176 9296 0 simon1.seq\[24\]\[1\]
rlabel metal3 35280 16744 35280 16744 0 simon1.seq\[25\]\[0\]
rlabel metal2 38248 16464 38248 16464 0 simon1.seq\[25\]\[1\]
rlabel metal2 23016 5096 23016 5096 0 simon1.seq\[26\]\[0\]
rlabel metal3 24192 5208 24192 5208 0 simon1.seq\[26\]\[1\]
rlabel metal2 20664 5264 20664 5264 0 simon1.seq\[27\]\[0\]
rlabel metal2 16856 4480 16856 4480 0 simon1.seq\[27\]\[1\]
rlabel metal2 25200 16856 25200 16856 0 simon1.seq\[28\]\[0\]
rlabel metal2 21784 11816 21784 11816 0 simon1.seq\[28\]\[1\]
rlabel metal2 28952 25200 28952 25200 0 simon1.seq\[29\]\[0\]
rlabel metal2 30632 23072 30632 23072 0 simon1.seq\[29\]\[1\]
rlabel metal3 21392 7336 21392 7336 0 simon1.seq\[2\]\[0\]
rlabel metal2 19544 8288 19544 8288 0 simon1.seq\[2\]\[1\]
rlabel metal2 14280 9856 14280 9856 0 simon1.seq\[30\]\[0\]
rlabel metal2 15456 6888 15456 6888 0 simon1.seq\[30\]\[1\]
rlabel metal3 14000 10472 14000 10472 0 simon1.seq\[31\]\[0\]
rlabel metal2 15064 7840 15064 7840 0 simon1.seq\[31\]\[1\]
rlabel metal2 26824 6552 26824 6552 0 simon1.seq\[3\]\[0\]
rlabel metal2 27720 5040 27720 5040 0 simon1.seq\[3\]\[1\]
rlabel metal2 31808 5880 31808 5880 0 simon1.seq\[4\]\[0\]
rlabel metal2 33544 6272 33544 6272 0 simon1.seq\[4\]\[1\]
rlabel metal2 42728 22456 42728 22456 0 simon1.seq\[5\]\[0\]
rlabel metal2 42392 21168 42392 21168 0 simon1.seq\[5\]\[1\]
rlabel metal2 32536 9576 32536 9576 0 simon1.seq\[6\]\[0\]
rlabel metal2 32536 7784 32536 7784 0 simon1.seq\[6\]\[1\]
rlabel metal2 33880 22512 33880 22512 0 simon1.seq\[7\]\[0\]
rlabel metal2 34888 23912 34888 23912 0 simon1.seq\[7\]\[1\]
rlabel metal2 37632 11480 37632 11480 0 simon1.seq\[8\]\[0\]
rlabel metal2 39032 14392 39032 14392 0 simon1.seq\[8\]\[1\]
rlabel metal2 38696 21168 38696 21168 0 simon1.seq\[9\]\[0\]
rlabel metal2 38136 18872 38136 18872 0 simon1.seq\[9\]\[1\]
rlabel metal2 11424 24584 11424 24584 0 simon1.seq_counter\[0\]
rlabel metal2 7448 23072 7448 23072 0 simon1.seq_counter\[1\]
rlabel metal2 9352 25592 9352 25592 0 simon1.seq_counter\[2\]
rlabel metal3 8176 23800 8176 23800 0 simon1.seq_counter\[3\]
rlabel metal2 8456 25592 8456 25592 0 simon1.seq_counter\[4\]
rlabel metal2 15960 24248 15960 24248 0 simon1.seq_length\[0\]
rlabel metal2 12936 24192 12936 24192 0 simon1.seq_length\[1\]
rlabel metal2 17416 22848 17416 22848 0 simon1.seq_length\[2\]
rlabel metal2 10248 20440 10248 20440 0 simon1.seq_length\[3\]
rlabel metal2 11144 22568 11144 22568 0 simon1.seq_length\[4\]
rlabel metal2 16632 32144 16632 32144 0 simon1.state\[0\]
rlabel metal3 11592 30968 11592 30968 0 simon1.state\[1\]
rlabel metal2 10920 31752 10920 31752 0 simon1.state\[2\]
rlabel metal2 20272 27720 20272 27720 0 simon1.state\[3\]
rlabel metal2 18312 28728 18312 28728 0 simon1.state\[4\]
rlabel metal2 20328 28952 20328 28952 0 simon1.state\[5\]
rlabel metal2 12824 29792 12824 29792 0 simon1.state\[6\]
rlabel metal2 18144 35000 18144 35000 0 simon1.state\[7\]
rlabel metal3 5936 49000 5936 49000 0 simon1.tick_counter\[0\]
rlabel metal2 11928 46704 11928 46704 0 simon1.tick_counter\[10\]
rlabel metal2 12376 51520 12376 51520 0 simon1.tick_counter\[11\]
rlabel metal2 12656 51352 12656 51352 0 simon1.tick_counter\[12\]
rlabel metal2 9800 46200 9800 46200 0 simon1.tick_counter\[13\]
rlabel metal2 10024 54208 10024 54208 0 simon1.tick_counter\[14\]
rlabel metal2 10584 54152 10584 54152 0 simon1.tick_counter\[15\]
rlabel metal3 4088 49784 4088 49784 0 simon1.tick_counter\[1\]
rlabel metal2 8456 44688 8456 44688 0 simon1.tick_counter\[2\]
rlabel metal2 5656 52192 5656 52192 0 simon1.tick_counter\[3\]
rlabel metal3 6888 52136 6888 52136 0 simon1.tick_counter\[4\]
rlabel metal2 5936 55048 5936 55048 0 simon1.tick_counter\[5\]
rlabel metal2 6048 53032 6048 53032 0 simon1.tick_counter\[6\]
rlabel metal2 5600 48216 5600 48216 0 simon1.tick_counter\[7\]
rlabel metal2 7672 46816 7672 46816 0 simon1.tick_counter\[8\]
rlabel metal2 10360 46648 10360 46648 0 simon1.tick_counter\[9\]
rlabel metal2 23016 39984 23016 39984 0 simon1.tone_sequence_counter\[0\]
rlabel metal2 23240 40936 23240 40936 0 simon1.tone_sequence_counter\[1\]
rlabel metal2 21616 38920 21616 38920 0 simon1.tone_sequence_counter\[2\]
rlabel metal2 26040 28616 26040 28616 0 simon1.user_input\[0\]
rlabel metal2 20832 44968 20832 44968 0 simon1.user_input\[1\]
rlabel metal3 2856 53816 2856 53816 0 wb_clk_i
rlabel metal2 4592 56280 4592 56280 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
