VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_design_mux
  CLASS BLOCK ;
  FOREIGN top_design_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 2400.000 BY 220.000 ;
  PIN diego_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1515.360 0.000 1515.920 4.000 ;
    END
  END diego_clk
  PIN diego_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1528.800 0.000 1529.360 4.000 ;
    END
  END diego_ena
  PIN diego_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1965.600 0.000 1966.160 4.000 ;
    END
  END diego_io_in[0]
  PIN diego_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2032.800 0.000 2033.360 4.000 ;
    END
  END diego_io_in[10]
  PIN diego_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2039.520 0.000 2040.080 4.000 ;
    END
  END diego_io_in[11]
  PIN diego_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2046.240 0.000 2046.800 4.000 ;
    END
  END diego_io_in[12]
  PIN diego_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2052.960 0.000 2053.520 4.000 ;
    END
  END diego_io_in[13]
  PIN diego_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2059.680 0.000 2060.240 4.000 ;
    END
  END diego_io_in[14]
  PIN diego_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2066.400 0.000 2066.960 4.000 ;
    END
  END diego_io_in[15]
  PIN diego_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2073.120 0.000 2073.680 4.000 ;
    END
  END diego_io_in[16]
  PIN diego_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2079.840 0.000 2080.400 4.000 ;
    END
  END diego_io_in[17]
  PIN diego_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2086.560 0.000 2087.120 4.000 ;
    END
  END diego_io_in[18]
  PIN diego_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2093.280 0.000 2093.840 4.000 ;
    END
  END diego_io_in[19]
  PIN diego_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1972.320 0.000 1972.880 4.000 ;
    END
  END diego_io_in[1]
  PIN diego_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2100.000 0.000 2100.560 4.000 ;
    END
  END diego_io_in[20]
  PIN diego_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2106.720 0.000 2107.280 4.000 ;
    END
  END diego_io_in[21]
  PIN diego_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2113.440 0.000 2114.000 4.000 ;
    END
  END diego_io_in[22]
  PIN diego_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2120.160 0.000 2120.720 4.000 ;
    END
  END diego_io_in[23]
  PIN diego_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2126.880 0.000 2127.440 4.000 ;
    END
  END diego_io_in[24]
  PIN diego_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2133.600 0.000 2134.160 4.000 ;
    END
  END diego_io_in[25]
  PIN diego_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2140.320 0.000 2140.880 4.000 ;
    END
  END diego_io_in[26]
  PIN diego_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2147.040 0.000 2147.600 4.000 ;
    END
  END diego_io_in[27]
  PIN diego_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2153.760 0.000 2154.320 4.000 ;
    END
  END diego_io_in[28]
  PIN diego_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2160.480 0.000 2161.040 4.000 ;
    END
  END diego_io_in[29]
  PIN diego_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1979.040 0.000 1979.600 4.000 ;
    END
  END diego_io_in[2]
  PIN diego_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2167.200 0.000 2167.760 4.000 ;
    END
  END diego_io_in[30]
  PIN diego_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2173.920 0.000 2174.480 4.000 ;
    END
  END diego_io_in[31]
  PIN diego_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2180.640 0.000 2181.200 4.000 ;
    END
  END diego_io_in[32]
  PIN diego_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2187.360 0.000 2187.920 4.000 ;
    END
  END diego_io_in[33]
  PIN diego_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2194.080 0.000 2194.640 4.000 ;
    END
  END diego_io_in[34]
  PIN diego_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2200.800 0.000 2201.360 4.000 ;
    END
  END diego_io_in[35]
  PIN diego_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2207.520 0.000 2208.080 4.000 ;
    END
  END diego_io_in[36]
  PIN diego_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2214.240 0.000 2214.800 4.000 ;
    END
  END diego_io_in[37]
  PIN diego_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1985.760 0.000 1986.320 4.000 ;
    END
  END diego_io_in[3]
  PIN diego_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1992.480 0.000 1993.040 4.000 ;
    END
  END diego_io_in[4]
  PIN diego_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1999.200 0.000 1999.760 4.000 ;
    END
  END diego_io_in[5]
  PIN diego_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2005.920 0.000 2006.480 4.000 ;
    END
  END diego_io_in[6]
  PIN diego_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2012.640 0.000 2013.200 4.000 ;
    END
  END diego_io_in[7]
  PIN diego_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2019.360 0.000 2019.920 4.000 ;
    END
  END diego_io_in[8]
  PIN diego_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2026.080 0.000 2026.640 4.000 ;
    END
  END diego_io_in[9]
  PIN diego_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1750.560 0.000 1751.120 4.000 ;
    END
  END diego_io_oeb[0]
  PIN diego_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1817.760 0.000 1818.320 4.000 ;
    END
  END diego_io_oeb[10]
  PIN diego_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1824.480 0.000 1825.040 4.000 ;
    END
  END diego_io_oeb[11]
  PIN diego_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1831.200 0.000 1831.760 4.000 ;
    END
  END diego_io_oeb[12]
  PIN diego_io_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1837.920 0.000 1838.480 4.000 ;
    END
  END diego_io_oeb[13]
  PIN diego_io_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1844.640 0.000 1845.200 4.000 ;
    END
  END diego_io_oeb[14]
  PIN diego_io_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1851.360 0.000 1851.920 4.000 ;
    END
  END diego_io_oeb[15]
  PIN diego_io_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1858.080 0.000 1858.640 4.000 ;
    END
  END diego_io_oeb[16]
  PIN diego_io_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1864.800 0.000 1865.360 4.000 ;
    END
  END diego_io_oeb[17]
  PIN diego_io_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1871.520 0.000 1872.080 4.000 ;
    END
  END diego_io_oeb[18]
  PIN diego_io_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1878.240 0.000 1878.800 4.000 ;
    END
  END diego_io_oeb[19]
  PIN diego_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1757.280 0.000 1757.840 4.000 ;
    END
  END diego_io_oeb[1]
  PIN diego_io_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1884.960 0.000 1885.520 4.000 ;
    END
  END diego_io_oeb[20]
  PIN diego_io_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1891.680 0.000 1892.240 4.000 ;
    END
  END diego_io_oeb[21]
  PIN diego_io_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1898.400 0.000 1898.960 4.000 ;
    END
  END diego_io_oeb[22]
  PIN diego_io_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1905.120 0.000 1905.680 4.000 ;
    END
  END diego_io_oeb[23]
  PIN diego_io_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1911.840 0.000 1912.400 4.000 ;
    END
  END diego_io_oeb[24]
  PIN diego_io_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1918.560 0.000 1919.120 4.000 ;
    END
  END diego_io_oeb[25]
  PIN diego_io_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1925.280 0.000 1925.840 4.000 ;
    END
  END diego_io_oeb[26]
  PIN diego_io_oeb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1932.000 0.000 1932.560 4.000 ;
    END
  END diego_io_oeb[27]
  PIN diego_io_oeb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1938.720 0.000 1939.280 4.000 ;
    END
  END diego_io_oeb[28]
  PIN diego_io_oeb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1945.440 0.000 1946.000 4.000 ;
    END
  END diego_io_oeb[29]
  PIN diego_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1764.000 0.000 1764.560 4.000 ;
    END
  END diego_io_oeb[2]
  PIN diego_io_oeb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1952.160 0.000 1952.720 4.000 ;
    END
  END diego_io_oeb[30]
  PIN diego_io_oeb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1958.880 0.000 1959.440 4.000 ;
    END
  END diego_io_oeb[31]
  PIN diego_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1770.720 0.000 1771.280 4.000 ;
    END
  END diego_io_oeb[3]
  PIN diego_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1777.440 0.000 1778.000 4.000 ;
    END
  END diego_io_oeb[4]
  PIN diego_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1784.160 0.000 1784.720 4.000 ;
    END
  END diego_io_oeb[5]
  PIN diego_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1790.880 0.000 1791.440 4.000 ;
    END
  END diego_io_oeb[6]
  PIN diego_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1797.600 0.000 1798.160 4.000 ;
    END
  END diego_io_oeb[7]
  PIN diego_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1804.320 0.000 1804.880 4.000 ;
    END
  END diego_io_oeb[8]
  PIN diego_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1811.040 0.000 1811.600 4.000 ;
    END
  END diego_io_oeb[9]
  PIN diego_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1535.520 0.000 1536.080 4.000 ;
    END
  END diego_io_out[0]
  PIN diego_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1602.720 0.000 1603.280 4.000 ;
    END
  END diego_io_out[10]
  PIN diego_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1609.440 0.000 1610.000 4.000 ;
    END
  END diego_io_out[11]
  PIN diego_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1616.160 0.000 1616.720 4.000 ;
    END
  END diego_io_out[12]
  PIN diego_io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1622.880 0.000 1623.440 4.000 ;
    END
  END diego_io_out[13]
  PIN diego_io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1629.600 0.000 1630.160 4.000 ;
    END
  END diego_io_out[14]
  PIN diego_io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1636.320 0.000 1636.880 4.000 ;
    END
  END diego_io_out[15]
  PIN diego_io_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1643.040 0.000 1643.600 4.000 ;
    END
  END diego_io_out[16]
  PIN diego_io_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1649.760 0.000 1650.320 4.000 ;
    END
  END diego_io_out[17]
  PIN diego_io_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1656.480 0.000 1657.040 4.000 ;
    END
  END diego_io_out[18]
  PIN diego_io_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1663.200 0.000 1663.760 4.000 ;
    END
  END diego_io_out[19]
  PIN diego_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1542.240 0.000 1542.800 4.000 ;
    END
  END diego_io_out[1]
  PIN diego_io_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1669.920 0.000 1670.480 4.000 ;
    END
  END diego_io_out[20]
  PIN diego_io_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1676.640 0.000 1677.200 4.000 ;
    END
  END diego_io_out[21]
  PIN diego_io_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1683.360 0.000 1683.920 4.000 ;
    END
  END diego_io_out[22]
  PIN diego_io_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1690.080 0.000 1690.640 4.000 ;
    END
  END diego_io_out[23]
  PIN diego_io_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1696.800 0.000 1697.360 4.000 ;
    END
  END diego_io_out[24]
  PIN diego_io_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1703.520 0.000 1704.080 4.000 ;
    END
  END diego_io_out[25]
  PIN diego_io_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1710.240 0.000 1710.800 4.000 ;
    END
  END diego_io_out[26]
  PIN diego_io_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1716.960 0.000 1717.520 4.000 ;
    END
  END diego_io_out[27]
  PIN diego_io_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1723.680 0.000 1724.240 4.000 ;
    END
  END diego_io_out[28]
  PIN diego_io_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1730.400 0.000 1730.960 4.000 ;
    END
  END diego_io_out[29]
  PIN diego_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1548.960 0.000 1549.520 4.000 ;
    END
  END diego_io_out[2]
  PIN diego_io_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1737.120 0.000 1737.680 4.000 ;
    END
  END diego_io_out[30]
  PIN diego_io_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1743.840 0.000 1744.400 4.000 ;
    END
  END diego_io_out[31]
  PIN diego_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1555.680 0.000 1556.240 4.000 ;
    END
  END diego_io_out[3]
  PIN diego_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1562.400 0.000 1562.960 4.000 ;
    END
  END diego_io_out[4]
  PIN diego_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1569.120 0.000 1569.680 4.000 ;
    END
  END diego_io_out[5]
  PIN diego_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1575.840 0.000 1576.400 4.000 ;
    END
  END diego_io_out[6]
  PIN diego_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1582.560 0.000 1583.120 4.000 ;
    END
  END diego_io_out[7]
  PIN diego_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1589.280 0.000 1589.840 4.000 ;
    END
  END diego_io_out[8]
  PIN diego_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1596.000 0.000 1596.560 4.000 ;
    END
  END diego_io_out[9]
  PIN diego_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1522.080 0.000 1522.640 4.000 ;
    END
  END diego_rst
  PIN i_design_reset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 26.880 2400.000 27.440 ;
    END
  END i_design_reset[0]
  PIN i_design_reset[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 30.240 2400.000 30.800 ;
    END
  END i_design_reset[1]
  PIN i_design_reset[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 33.600 2400.000 34.160 ;
    END
  END i_design_reset[2]
  PIN i_design_reset[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 36.960 2400.000 37.520 ;
    END
  END i_design_reset[3]
  PIN i_design_reset[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 40.320 2400.000 40.880 ;
    END
  END i_design_reset[4]
  PIN i_design_reset[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 43.680 2400.000 44.240 ;
    END
  END i_design_reset[5]
  PIN i_design_reset[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 47.040 2400.000 47.600 ;
    END
  END i_design_reset[6]
  PIN i_design_reset[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 50.400 2400.000 50.960 ;
    END
  END i_design_reset[7]
  PIN i_mux_auto_reset_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 23.520 2400.000 24.080 ;
    END
  END i_mux_auto_reset_enb
  PIN i_mux_io5_reset_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 3.360 2400.000 3.920 ;
    END
  END i_mux_io5_reset_enb
  PIN i_mux_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 6.720 2400.000 7.280 ;
    END
  END i_mux_sel[0]
  PIN i_mux_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 10.080 2400.000 10.640 ;
    END
  END i_mux_sel[1]
  PIN i_mux_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 13.440 2400.000 14.000 ;
    END
  END i_mux_sel[2]
  PIN i_mux_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 16.800 2400.000 17.360 ;
    END
  END i_mux_sel[3]
  PIN i_mux_sys_reset_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 20.160 2400.000 20.720 ;
    END
  END i_mux_sys_reset_enb
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 57.120 2400.000 57.680 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 157.920 2400.000 158.480 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 168.000 2400.000 168.560 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 178.080 2400.000 178.640 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 188.160 2400.000 188.720 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 198.240 2400.000 198.800 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 208.320 2400.000 208.880 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1327.200 216.000 1327.760 220.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1307.040 216.000 1307.600 220.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1286.880 216.000 1287.440 220.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 216.000 669.200 220.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 67.200 2400.000 67.760 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 216.000 649.040 220.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 216.000 628.880 220.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 216.000 608.720 220.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.800 4.000 213.360 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 199.360 4.000 199.920 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.920 4.000 186.480 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 172.480 4.000 173.040 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 159.040 4.000 159.600 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.600 4.000 146.160 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.160 4.000 132.720 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 77.280 2400.000 77.840 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.720 4.000 119.280 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.280 4.000 105.840 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 91.840 4.000 92.400 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.960 4.000 65.520 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 4.000 52.080 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.080 4.000 38.640 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.640 4.000 25.200 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 87.360 2400.000 87.920 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 97.440 2400.000 98.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 107.520 2400.000 108.080 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 117.600 2400.000 118.160 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 127.680 2400.000 128.240 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 137.760 2400.000 138.320 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 147.840 2400.000 148.400 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 63.840 2400.000 64.400 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 164.640 2400.000 165.200 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 174.720 2400.000 175.280 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 184.800 2400.000 185.360 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 194.880 2400.000 195.440 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 204.960 2400.000 205.520 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 215.040 2400.000 215.600 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1313.760 216.000 1314.320 220.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1293.600 216.000 1294.160 220.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1273.440 216.000 1274.000 220.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 216.000 655.760 220.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 73.920 2400.000 74.480 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 216.000 635.600 220.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 216.000 615.440 220.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 216.000 595.280 220.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 203.840 4.000 204.400 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.400 4.000 190.960 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 176.960 4.000 177.520 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 163.520 4.000 164.080 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.080 4.000 150.640 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 136.640 4.000 137.200 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.200 4.000 123.760 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 84.000 2400.000 84.560 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.760 4.000 110.320 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.320 4.000 96.880 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 82.880 4.000 83.440 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.440 4.000 70.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.000 4.000 56.560 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 4.000 43.120 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 4.000 29.680 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.680 4.000 16.240 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 94.080 2400.000 94.640 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 104.160 2400.000 104.720 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 114.240 2400.000 114.800 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 124.320 2400.000 124.880 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 134.400 2400.000 134.960 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 144.480 2400.000 145.040 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 154.560 2400.000 155.120 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 60.480 2400.000 61.040 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 161.280 2400.000 161.840 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 171.360 2400.000 171.920 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 181.440 2400.000 182.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 191.520 2400.000 192.080 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 201.600 2400.000 202.160 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 211.680 2400.000 212.240 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1320.480 216.000 1321.040 220.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1300.320 216.000 1300.880 220.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1280.160 216.000 1280.720 220.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 216.000 662.480 220.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 70.560 2400.000 71.120 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 216.000 642.320 220.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 216.000 622.160 220.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 216.000 602.000 220.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.320 4.000 208.880 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 4.000 182.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 80.640 2400.000 81.200 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 4.000 74.480 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.040 4.000 47.600 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 4.000 34.160 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 90.720 2400.000 91.280 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 100.800 2400.000 101.360 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 110.880 2400.000 111.440 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 120.960 2400.000 121.520 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 131.040 2400.000 131.600 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 141.120 2400.000 141.680 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 151.200 2400.000 151.760 ;
    END
  END io_out[9]
  PIN la_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1273.440 0.000 1274.000 4.000 ;
    END
  END la_in[0]
  PIN la_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1340.640 0.000 1341.200 4.000 ;
    END
  END la_in[10]
  PIN la_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1347.360 0.000 1347.920 4.000 ;
    END
  END la_in[11]
  PIN la_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1354.080 0.000 1354.640 4.000 ;
    END
  END la_in[12]
  PIN la_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1360.800 0.000 1361.360 4.000 ;
    END
  END la_in[13]
  PIN la_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1367.520 0.000 1368.080 4.000 ;
    END
  END la_in[14]
  PIN la_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1374.240 0.000 1374.800 4.000 ;
    END
  END la_in[15]
  PIN la_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1280.160 0.000 1280.720 4.000 ;
    END
  END la_in[1]
  PIN la_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1286.880 0.000 1287.440 4.000 ;
    END
  END la_in[2]
  PIN la_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1293.600 0.000 1294.160 4.000 ;
    END
  END la_in[3]
  PIN la_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1300.320 0.000 1300.880 4.000 ;
    END
  END la_in[4]
  PIN la_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1307.040 0.000 1307.600 4.000 ;
    END
  END la_in[5]
  PIN la_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1313.760 0.000 1314.320 4.000 ;
    END
  END la_in[6]
  PIN la_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1320.480 0.000 1321.040 4.000 ;
    END
  END la_in[7]
  PIN la_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1327.200 0.000 1327.760 4.000 ;
    END
  END la_in[8]
  PIN la_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1333.920 0.000 1334.480 4.000 ;
    END
  END la_in[9]
  PIN mux_conf_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 53.760 2400.000 54.320 ;
    END
  END mux_conf_clk
  PIN pawel_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END pawel_clk
  PIN pawel_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END pawel_ena
  PIN pawel_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END pawel_io_in[0]
  PIN pawel_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 0.000 420.560 4.000 ;
    END
  END pawel_io_in[10]
  PIN pawel_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 0.000 427.280 4.000 ;
    END
  END pawel_io_in[11]
  PIN pawel_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 0.000 434.000 4.000 ;
    END
  END pawel_io_in[12]
  PIN pawel_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 0.000 440.720 4.000 ;
    END
  END pawel_io_in[13]
  PIN pawel_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 0.000 447.440 4.000 ;
    END
  END pawel_io_in[14]
  PIN pawel_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 0.000 454.160 4.000 ;
    END
  END pawel_io_in[15]
  PIN pawel_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 0.000 460.880 4.000 ;
    END
  END pawel_io_in[16]
  PIN pawel_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 0.000 467.600 4.000 ;
    END
  END pawel_io_in[17]
  PIN pawel_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 0.000 474.320 4.000 ;
    END
  END pawel_io_in[18]
  PIN pawel_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 0.000 481.040 4.000 ;
    END
  END pawel_io_in[19]
  PIN pawel_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 0.000 360.080 4.000 ;
    END
  END pawel_io_in[1]
  PIN pawel_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 0.000 487.760 4.000 ;
    END
  END pawel_io_in[20]
  PIN pawel_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 0.000 494.480 4.000 ;
    END
  END pawel_io_in[21]
  PIN pawel_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 0.000 501.200 4.000 ;
    END
  END pawel_io_in[22]
  PIN pawel_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 0.000 507.920 4.000 ;
    END
  END pawel_io_in[23]
  PIN pawel_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 0.000 514.640 4.000 ;
    END
  END pawel_io_in[24]
  PIN pawel_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 0.000 521.360 4.000 ;
    END
  END pawel_io_in[25]
  PIN pawel_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 0.000 528.080 4.000 ;
    END
  END pawel_io_in[26]
  PIN pawel_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 0.000 534.800 4.000 ;
    END
  END pawel_io_in[27]
  PIN pawel_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 0.000 541.520 4.000 ;
    END
  END pawel_io_in[28]
  PIN pawel_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 0.000 548.240 4.000 ;
    END
  END pawel_io_in[29]
  PIN pawel_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 0.000 366.800 4.000 ;
    END
  END pawel_io_in[2]
  PIN pawel_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 0.000 554.960 4.000 ;
    END
  END pawel_io_in[30]
  PIN pawel_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 0.000 561.680 4.000 ;
    END
  END pawel_io_in[31]
  PIN pawel_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 0.000 568.400 4.000 ;
    END
  END pawel_io_in[32]
  PIN pawel_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 0.000 575.120 4.000 ;
    END
  END pawel_io_in[33]
  PIN pawel_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 0.000 581.840 4.000 ;
    END
  END pawel_io_in[34]
  PIN pawel_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 0.000 588.560 4.000 ;
    END
  END pawel_io_in[35]
  PIN pawel_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 0.000 595.280 4.000 ;
    END
  END pawel_io_in[36]
  PIN pawel_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 0.000 602.000 4.000 ;
    END
  END pawel_io_in[37]
  PIN pawel_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 0.000 373.520 4.000 ;
    END
  END pawel_io_in[3]
  PIN pawel_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 0.000 380.240 4.000 ;
    END
  END pawel_io_in[4]
  PIN pawel_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END pawel_io_in[5]
  PIN pawel_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 0.000 393.680 4.000 ;
    END
  END pawel_io_in[6]
  PIN pawel_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 0.000 400.400 4.000 ;
    END
  END pawel_io_in[7]
  PIN pawel_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 0.000 407.120 4.000 ;
    END
  END pawel_io_in[8]
  PIN pawel_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 0.000 413.840 4.000 ;
    END
  END pawel_io_in[9]
  PIN pawel_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END pawel_io_oeb[0]
  PIN pawel_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END pawel_io_oeb[10]
  PIN pawel_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 0.000 232.400 4.000 ;
    END
  END pawel_io_oeb[11]
  PIN pawel_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 4.000 ;
    END
  END pawel_io_oeb[12]
  PIN pawel_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END pawel_io_oeb[1]
  PIN pawel_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END pawel_io_oeb[2]
  PIN pawel_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END pawel_io_oeb[3]
  PIN pawel_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END pawel_io_oeb[4]
  PIN pawel_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END pawel_io_oeb[5]
  PIN pawel_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 4.000 ;
    END
  END pawel_io_oeb[6]
  PIN pawel_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END pawel_io_oeb[7]
  PIN pawel_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END pawel_io_oeb[8]
  PIN pawel_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END pawel_io_oeb[9]
  PIN pawel_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END pawel_io_out[0]
  PIN pawel_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 4.000 ;
    END
  END pawel_io_out[10]
  PIN pawel_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END pawel_io_out[11]
  PIN pawel_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END pawel_io_out[12]
  PIN pawel_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END pawel_io_out[1]
  PIN pawel_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END pawel_io_out[2]
  PIN pawel_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END pawel_io_out[3]
  PIN pawel_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END pawel_io_out[4]
  PIN pawel_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END pawel_io_out[5]
  PIN pawel_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END pawel_io_out[6]
  PIN pawel_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END pawel_io_out[7]
  PIN pawel_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END pawel_io_out[8]
  PIN pawel_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END pawel_io_out[9]
  PIN pawel_la_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 0.000 245.840 4.000 ;
    END
  END pawel_la_in[0]
  PIN pawel_la_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 0.000 313.040 4.000 ;
    END
  END pawel_la_in[10]
  PIN pawel_la_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 0.000 319.760 4.000 ;
    END
  END pawel_la_in[11]
  PIN pawel_la_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 0.000 326.480 4.000 ;
    END
  END pawel_la_in[12]
  PIN pawel_la_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 0.000 333.200 4.000 ;
    END
  END pawel_la_in[13]
  PIN pawel_la_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 0.000 339.920 4.000 ;
    END
  END pawel_la_in[14]
  PIN pawel_la_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 0.000 346.640 4.000 ;
    END
  END pawel_la_in[15]
  PIN pawel_la_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 0.000 252.560 4.000 ;
    END
  END pawel_la_in[1]
  PIN pawel_la_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 0.000 259.280 4.000 ;
    END
  END pawel_la_in[2]
  PIN pawel_la_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 0.000 266.000 4.000 ;
    END
  END pawel_la_in[3]
  PIN pawel_la_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 0.000 272.720 4.000 ;
    END
  END pawel_la_in[4]
  PIN pawel_la_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 4.000 ;
    END
  END pawel_la_in[5]
  PIN pawel_la_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 0.000 286.160 4.000 ;
    END
  END pawel_la_in[6]
  PIN pawel_la_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 0.000 292.880 4.000 ;
    END
  END pawel_la_in[7]
  PIN pawel_la_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 0.000 299.600 4.000 ;
    END
  END pawel_la_in[8]
  PIN pawel_la_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 0.000 306.320 4.000 ;
    END
  END pawel_la_in[9]
  PIN pawel_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END pawel_rst
  PIN solos_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1905.120 216.000 1905.680 220.000 ;
    END
  END solos_clk
  PIN solos_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1918.560 216.000 1919.120 220.000 ;
    END
  END solos_ena
  PIN solos_gpio_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1925.280 216.000 1925.840 220.000 ;
    END
  END solos_gpio_ready
  PIN solos_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2180.640 216.000 2181.200 220.000 ;
    END
  END solos_io_in[0]
  PIN solos_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2113.440 216.000 2114.000 220.000 ;
    END
  END solos_io_in[10]
  PIN solos_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2106.720 216.000 2107.280 220.000 ;
    END
  END solos_io_in[11]
  PIN solos_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2100.000 216.000 2100.560 220.000 ;
    END
  END solos_io_in[12]
  PIN solos_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2093.280 216.000 2093.840 220.000 ;
    END
  END solos_io_in[13]
  PIN solos_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2086.560 216.000 2087.120 220.000 ;
    END
  END solos_io_in[14]
  PIN solos_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2079.840 216.000 2080.400 220.000 ;
    END
  END solos_io_in[15]
  PIN solos_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2073.120 216.000 2073.680 220.000 ;
    END
  END solos_io_in[16]
  PIN solos_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2066.400 216.000 2066.960 220.000 ;
    END
  END solos_io_in[17]
  PIN solos_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2059.680 216.000 2060.240 220.000 ;
    END
  END solos_io_in[18]
  PIN solos_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2052.960 216.000 2053.520 220.000 ;
    END
  END solos_io_in[19]
  PIN solos_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2173.920 216.000 2174.480 220.000 ;
    END
  END solos_io_in[1]
  PIN solos_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2046.240 216.000 2046.800 220.000 ;
    END
  END solos_io_in[20]
  PIN solos_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2039.520 216.000 2040.080 220.000 ;
    END
  END solos_io_in[21]
  PIN solos_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2032.800 216.000 2033.360 220.000 ;
    END
  END solos_io_in[22]
  PIN solos_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2026.080 216.000 2026.640 220.000 ;
    END
  END solos_io_in[23]
  PIN solos_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2019.360 216.000 2019.920 220.000 ;
    END
  END solos_io_in[24]
  PIN solos_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2012.640 216.000 2013.200 220.000 ;
    END
  END solos_io_in[25]
  PIN solos_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2005.920 216.000 2006.480 220.000 ;
    END
  END solos_io_in[26]
  PIN solos_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1999.200 216.000 1999.760 220.000 ;
    END
  END solos_io_in[27]
  PIN solos_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1992.480 216.000 1993.040 220.000 ;
    END
  END solos_io_in[28]
  PIN solos_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1985.760 216.000 1986.320 220.000 ;
    END
  END solos_io_in[29]
  PIN solos_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2167.200 216.000 2167.760 220.000 ;
    END
  END solos_io_in[2]
  PIN solos_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1979.040 216.000 1979.600 220.000 ;
    END
  END solos_io_in[30]
  PIN solos_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1972.320 216.000 1972.880 220.000 ;
    END
  END solos_io_in[31]
  PIN solos_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1965.600 216.000 1966.160 220.000 ;
    END
  END solos_io_in[32]
  PIN solos_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1958.880 216.000 1959.440 220.000 ;
    END
  END solos_io_in[33]
  PIN solos_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1952.160 216.000 1952.720 220.000 ;
    END
  END solos_io_in[34]
  PIN solos_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1945.440 216.000 1946.000 220.000 ;
    END
  END solos_io_in[35]
  PIN solos_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1938.720 216.000 1939.280 220.000 ;
    END
  END solos_io_in[36]
  PIN solos_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1932.000 216.000 1932.560 220.000 ;
    END
  END solos_io_in[37]
  PIN solos_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2160.480 216.000 2161.040 220.000 ;
    END
  END solos_io_in[3]
  PIN solos_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2153.760 216.000 2154.320 220.000 ;
    END
  END solos_io_in[4]
  PIN solos_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2147.040 216.000 2147.600 220.000 ;
    END
  END solos_io_in[5]
  PIN solos_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2140.320 216.000 2140.880 220.000 ;
    END
  END solos_io_in[6]
  PIN solos_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2133.600 216.000 2134.160 220.000 ;
    END
  END solos_io_in[7]
  PIN solos_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2126.880 216.000 2127.440 220.000 ;
    END
  END solos_io_in[8]
  PIN solos_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2120.160 216.000 2120.720 220.000 ;
    END
  END solos_io_in[9]
  PIN solos_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2268.000 216.000 2268.560 220.000 ;
    END
  END solos_io_out[0]
  PIN solos_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2200.800 216.000 2201.360 220.000 ;
    END
  END solos_io_out[10]
  PIN solos_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2194.080 216.000 2194.640 220.000 ;
    END
  END solos_io_out[11]
  PIN solos_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2187.360 216.000 2187.920 220.000 ;
    END
  END solos_io_out[12]
  PIN solos_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2261.280 216.000 2261.840 220.000 ;
    END
  END solos_io_out[1]
  PIN solos_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2254.560 216.000 2255.120 220.000 ;
    END
  END solos_io_out[2]
  PIN solos_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2247.840 216.000 2248.400 220.000 ;
    END
  END solos_io_out[3]
  PIN solos_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2241.120 216.000 2241.680 220.000 ;
    END
  END solos_io_out[4]
  PIN solos_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2234.400 216.000 2234.960 220.000 ;
    END
  END solos_io_out[5]
  PIN solos_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2227.680 216.000 2228.240 220.000 ;
    END
  END solos_io_out[6]
  PIN solos_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2220.960 216.000 2221.520 220.000 ;
    END
  END solos_io_out[7]
  PIN solos_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2214.240 216.000 2214.800 220.000 ;
    END
  END solos_io_out[8]
  PIN solos_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2207.520 216.000 2208.080 220.000 ;
    END
  END solos_io_out[9]
  PIN solos_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1911.840 216.000 1912.400 220.000 ;
    END
  END solos_rst
  PIN trzf2_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 216.000 749.840 220.000 ;
    END
  END trzf2_clk
  PIN trzf2_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 216.000 743.120 220.000 ;
    END
  END trzf2_ena
  PIN trzf2_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1199.520 216.000 1200.080 220.000 ;
    END
  END trzf2_io_in[0]
  PIN trzf2_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1132.320 216.000 1132.880 220.000 ;
    END
  END trzf2_io_in[10]
  PIN trzf2_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1125.600 216.000 1126.160 220.000 ;
    END
  END trzf2_io_in[11]
  PIN trzf2_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1118.880 216.000 1119.440 220.000 ;
    END
  END trzf2_io_in[12]
  PIN trzf2_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1112.160 216.000 1112.720 220.000 ;
    END
  END trzf2_io_in[13]
  PIN trzf2_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1105.440 216.000 1106.000 220.000 ;
    END
  END trzf2_io_in[14]
  PIN trzf2_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1098.720 216.000 1099.280 220.000 ;
    END
  END trzf2_io_in[15]
  PIN trzf2_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1092.000 216.000 1092.560 220.000 ;
    END
  END trzf2_io_in[16]
  PIN trzf2_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1085.280 216.000 1085.840 220.000 ;
    END
  END trzf2_io_in[17]
  PIN trzf2_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1078.560 216.000 1079.120 220.000 ;
    END
  END trzf2_io_in[18]
  PIN trzf2_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1071.840 216.000 1072.400 220.000 ;
    END
  END trzf2_io_in[19]
  PIN trzf2_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1192.800 216.000 1193.360 220.000 ;
    END
  END trzf2_io_in[1]
  PIN trzf2_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1065.120 216.000 1065.680 220.000 ;
    END
  END trzf2_io_in[20]
  PIN trzf2_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1058.400 216.000 1058.960 220.000 ;
    END
  END trzf2_io_in[21]
  PIN trzf2_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1051.680 216.000 1052.240 220.000 ;
    END
  END trzf2_io_in[22]
  PIN trzf2_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1044.960 216.000 1045.520 220.000 ;
    END
  END trzf2_io_in[23]
  PIN trzf2_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1038.240 216.000 1038.800 220.000 ;
    END
  END trzf2_io_in[24]
  PIN trzf2_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1031.520 216.000 1032.080 220.000 ;
    END
  END trzf2_io_in[25]
  PIN trzf2_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1024.800 216.000 1025.360 220.000 ;
    END
  END trzf2_io_in[26]
  PIN trzf2_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1018.080 216.000 1018.640 220.000 ;
    END
  END trzf2_io_in[27]
  PIN trzf2_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1011.360 216.000 1011.920 220.000 ;
    END
  END trzf2_io_in[28]
  PIN trzf2_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1004.640 216.000 1005.200 220.000 ;
    END
  END trzf2_io_in[29]
  PIN trzf2_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1186.080 216.000 1186.640 220.000 ;
    END
  END trzf2_io_in[2]
  PIN trzf2_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 997.920 216.000 998.480 220.000 ;
    END
  END trzf2_io_in[30]
  PIN trzf2_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 216.000 991.760 220.000 ;
    END
  END trzf2_io_in[31]
  PIN trzf2_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 216.000 985.040 220.000 ;
    END
  END trzf2_io_in[32]
  PIN trzf2_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 977.760 216.000 978.320 220.000 ;
    END
  END trzf2_io_in[33]
  PIN trzf2_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 216.000 971.600 220.000 ;
    END
  END trzf2_io_in[34]
  PIN trzf2_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 964.320 216.000 964.880 220.000 ;
    END
  END trzf2_io_in[35]
  PIN trzf2_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 216.000 958.160 220.000 ;
    END
  END trzf2_io_in[36]
  PIN trzf2_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 950.880 216.000 951.440 220.000 ;
    END
  END trzf2_io_in[37]
  PIN trzf2_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1179.360 216.000 1179.920 220.000 ;
    END
  END trzf2_io_in[3]
  PIN trzf2_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1172.640 216.000 1173.200 220.000 ;
    END
  END trzf2_io_in[4]
  PIN trzf2_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1165.920 216.000 1166.480 220.000 ;
    END
  END trzf2_io_in[5]
  PIN trzf2_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1159.200 216.000 1159.760 220.000 ;
    END
  END trzf2_io_in[6]
  PIN trzf2_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1152.480 216.000 1153.040 220.000 ;
    END
  END trzf2_io_in[7]
  PIN trzf2_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1145.760 216.000 1146.320 220.000 ;
    END
  END trzf2_io_in[8]
  PIN trzf2_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1139.040 216.000 1139.600 220.000 ;
    END
  END trzf2_io_in[9]
  PIN trzf2_la_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 216.000 843.920 220.000 ;
    END
  END trzf2_la_in[0]
  PIN trzf2_la_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 216.000 776.720 220.000 ;
    END
  END trzf2_la_in[10]
  PIN trzf2_la_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 216.000 770.000 220.000 ;
    END
  END trzf2_la_in[11]
  PIN trzf2_la_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 216.000 763.280 220.000 ;
    END
  END trzf2_la_in[12]
  PIN trzf2_la_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 216.000 837.200 220.000 ;
    END
  END trzf2_la_in[1]
  PIN trzf2_la_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 216.000 830.480 220.000 ;
    END
  END trzf2_la_in[2]
  PIN trzf2_la_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 216.000 823.760 220.000 ;
    END
  END trzf2_la_in[3]
  PIN trzf2_la_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 216.000 817.040 220.000 ;
    END
  END trzf2_la_in[4]
  PIN trzf2_la_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 809.760 216.000 810.320 220.000 ;
    END
  END trzf2_la_in[5]
  PIN trzf2_la_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 216.000 803.600 220.000 ;
    END
  END trzf2_la_in[6]
  PIN trzf2_la_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 796.320 216.000 796.880 220.000 ;
    END
  END trzf2_la_in[7]
  PIN trzf2_la_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 216.000 790.160 220.000 ;
    END
  END trzf2_la_in[8]
  PIN trzf2_la_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 216.000 783.440 220.000 ;
    END
  END trzf2_la_in[9]
  PIN trzf2_o_gpout[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 216.000 864.080 220.000 ;
    END
  END trzf2_o_gpout[0]
  PIN trzf2_o_gpout[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 216.000 857.360 220.000 ;
    END
  END trzf2_o_gpout[1]
  PIN trzf2_o_gpout[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 216.000 850.640 220.000 ;
    END
  END trzf2_o_gpout[2]
  PIN trzf2_o_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 944.160 216.000 944.720 220.000 ;
    END
  END trzf2_o_hsync
  PIN trzf2_o_rgb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 930.720 216.000 931.280 220.000 ;
    END
  END trzf2_o_rgb[0]
  PIN trzf2_o_rgb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 924.000 216.000 924.560 220.000 ;
    END
  END trzf2_o_rgb[1]
  PIN trzf2_o_rgb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 216.000 917.840 220.000 ;
    END
  END trzf2_o_rgb[2]
  PIN trzf2_o_rgb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 910.560 216.000 911.120 220.000 ;
    END
  END trzf2_o_rgb[3]
  PIN trzf2_o_rgb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 216.000 904.400 220.000 ;
    END
  END trzf2_o_rgb[4]
  PIN trzf2_o_rgb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 216.000 897.680 220.000 ;
    END
  END trzf2_o_rgb[5]
  PIN trzf2_o_tex_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 216.000 890.960 220.000 ;
    END
  END trzf2_o_tex_csb
  PIN trzf2_o_tex_oeb0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 216.000 870.800 220.000 ;
    END
  END trzf2_o_tex_oeb0
  PIN trzf2_o_tex_out0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 876.960 216.000 877.520 220.000 ;
    END
  END trzf2_o_tex_out0
  PIN trzf2_o_tex_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 216.000 884.240 220.000 ;
    END
  END trzf2_o_tex_sclk
  PIN trzf2_o_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 216.000 938.000 220.000 ;
    END
  END trzf2_o_vsync
  PIN trzf2_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 216.000 756.560 220.000 ;
    END
  END trzf2_rst
  PIN trzf_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 216.000 71.120 220.000 ;
    END
  END trzf_clk
  PIN trzf_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 216.000 64.400 220.000 ;
    END
  END trzf_ena
  PIN trzf_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 216.000 521.360 220.000 ;
    END
  END trzf_io_in[0]
  PIN trzf_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 216.000 454.160 220.000 ;
    END
  END trzf_io_in[10]
  PIN trzf_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 216.000 447.440 220.000 ;
    END
  END trzf_io_in[11]
  PIN trzf_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 216.000 440.720 220.000 ;
    END
  END trzf_io_in[12]
  PIN trzf_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 216.000 434.000 220.000 ;
    END
  END trzf_io_in[13]
  PIN trzf_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 216.000 427.280 220.000 ;
    END
  END trzf_io_in[14]
  PIN trzf_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 216.000 420.560 220.000 ;
    END
  END trzf_io_in[15]
  PIN trzf_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 216.000 413.840 220.000 ;
    END
  END trzf_io_in[16]
  PIN trzf_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 216.000 407.120 220.000 ;
    END
  END trzf_io_in[17]
  PIN trzf_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 216.000 400.400 220.000 ;
    END
  END trzf_io_in[18]
  PIN trzf_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 216.000 393.680 220.000 ;
    END
  END trzf_io_in[19]
  PIN trzf_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 216.000 514.640 220.000 ;
    END
  END trzf_io_in[1]
  PIN trzf_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 216.000 386.960 220.000 ;
    END
  END trzf_io_in[20]
  PIN trzf_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 216.000 380.240 220.000 ;
    END
  END trzf_io_in[21]
  PIN trzf_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 216.000 373.520 220.000 ;
    END
  END trzf_io_in[22]
  PIN trzf_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 216.000 366.800 220.000 ;
    END
  END trzf_io_in[23]
  PIN trzf_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 216.000 360.080 220.000 ;
    END
  END trzf_io_in[24]
  PIN trzf_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 216.000 353.360 220.000 ;
    END
  END trzf_io_in[25]
  PIN trzf_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 216.000 346.640 220.000 ;
    END
  END trzf_io_in[26]
  PIN trzf_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 216.000 339.920 220.000 ;
    END
  END trzf_io_in[27]
  PIN trzf_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 216.000 333.200 220.000 ;
    END
  END trzf_io_in[28]
  PIN trzf_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 216.000 326.480 220.000 ;
    END
  END trzf_io_in[29]
  PIN trzf_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 216.000 507.920 220.000 ;
    END
  END trzf_io_in[2]
  PIN trzf_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 216.000 319.760 220.000 ;
    END
  END trzf_io_in[30]
  PIN trzf_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 216.000 313.040 220.000 ;
    END
  END trzf_io_in[31]
  PIN trzf_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 216.000 306.320 220.000 ;
    END
  END trzf_io_in[32]
  PIN trzf_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 216.000 299.600 220.000 ;
    END
  END trzf_io_in[33]
  PIN trzf_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 216.000 292.880 220.000 ;
    END
  END trzf_io_in[34]
  PIN trzf_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 216.000 286.160 220.000 ;
    END
  END trzf_io_in[35]
  PIN trzf_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 216.000 279.440 220.000 ;
    END
  END trzf_io_in[36]
  PIN trzf_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 216.000 272.720 220.000 ;
    END
  END trzf_io_in[37]
  PIN trzf_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 216.000 501.200 220.000 ;
    END
  END trzf_io_in[3]
  PIN trzf_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 216.000 494.480 220.000 ;
    END
  END trzf_io_in[4]
  PIN trzf_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 216.000 487.760 220.000 ;
    END
  END trzf_io_in[5]
  PIN trzf_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 216.000 481.040 220.000 ;
    END
  END trzf_io_in[6]
  PIN trzf_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 216.000 474.320 220.000 ;
    END
  END trzf_io_in[7]
  PIN trzf_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 216.000 467.600 220.000 ;
    END
  END trzf_io_in[8]
  PIN trzf_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 216.000 460.880 220.000 ;
    END
  END trzf_io_in[9]
  PIN trzf_la_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 216.000 165.200 220.000 ;
    END
  END trzf_la_in[0]
  PIN trzf_la_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 216.000 98.000 220.000 ;
    END
  END trzf_la_in[10]
  PIN trzf_la_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 216.000 91.280 220.000 ;
    END
  END trzf_la_in[11]
  PIN trzf_la_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 216.000 84.560 220.000 ;
    END
  END trzf_la_in[12]
  PIN trzf_la_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 216.000 158.480 220.000 ;
    END
  END trzf_la_in[1]
  PIN trzf_la_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 216.000 151.760 220.000 ;
    END
  END trzf_la_in[2]
  PIN trzf_la_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 216.000 145.040 220.000 ;
    END
  END trzf_la_in[3]
  PIN trzf_la_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 216.000 138.320 220.000 ;
    END
  END trzf_la_in[4]
  PIN trzf_la_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 216.000 131.600 220.000 ;
    END
  END trzf_la_in[5]
  PIN trzf_la_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 216.000 124.880 220.000 ;
    END
  END trzf_la_in[6]
  PIN trzf_la_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 216.000 118.160 220.000 ;
    END
  END trzf_la_in[7]
  PIN trzf_la_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 216.000 111.440 220.000 ;
    END
  END trzf_la_in[8]
  PIN trzf_la_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 216.000 104.720 220.000 ;
    END
  END trzf_la_in[9]
  PIN trzf_o_gpout[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 216.000 185.360 220.000 ;
    END
  END trzf_o_gpout[0]
  PIN trzf_o_gpout[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 216.000 178.640 220.000 ;
    END
  END trzf_o_gpout[1]
  PIN trzf_o_gpout[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 216.000 171.920 220.000 ;
    END
  END trzf_o_gpout[2]
  PIN trzf_o_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 216.000 266.000 220.000 ;
    END
  END trzf_o_hsync
  PIN trzf_o_rgb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 216.000 252.560 220.000 ;
    END
  END trzf_o_rgb[0]
  PIN trzf_o_rgb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 216.000 245.840 220.000 ;
    END
  END trzf_o_rgb[1]
  PIN trzf_o_rgb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 216.000 239.120 220.000 ;
    END
  END trzf_o_rgb[2]
  PIN trzf_o_rgb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 216.000 232.400 220.000 ;
    END
  END trzf_o_rgb[3]
  PIN trzf_o_rgb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 216.000 225.680 220.000 ;
    END
  END trzf_o_rgb[4]
  PIN trzf_o_rgb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 216.000 218.960 220.000 ;
    END
  END trzf_o_rgb[5]
  PIN trzf_o_tex_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 216.000 212.240 220.000 ;
    END
  END trzf_o_tex_csb
  PIN trzf_o_tex_oeb0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 216.000 192.080 220.000 ;
    END
  END trzf_o_tex_oeb0
  PIN trzf_o_tex_out0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 216.000 198.800 220.000 ;
    END
  END trzf_o_tex_out0
  PIN trzf_o_tex_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 216.000 205.520 220.000 ;
    END
  END trzf_o_tex_sclk
  PIN trzf_o_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 216.000 259.280 220.000 ;
    END
  END trzf_o_vsync
  PIN trzf_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 216.000 77.840 220.000 ;
    END
  END trzf_rst
  PIN uri_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 0.000 675.920 4.000 ;
    END
  END uri_clk
  PIN uri_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 0.000 689.360 4.000 ;
    END
  END uri_ena
  PIN uri_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 950.880 0.000 951.440 4.000 ;
    END
  END uri_io_in[0]
  PIN uri_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1018.080 0.000 1018.640 4.000 ;
    END
  END uri_io_in[10]
  PIN uri_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1024.800 0.000 1025.360 4.000 ;
    END
  END uri_io_in[11]
  PIN uri_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1031.520 0.000 1032.080 4.000 ;
    END
  END uri_io_in[12]
  PIN uri_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1038.240 0.000 1038.800 4.000 ;
    END
  END uri_io_in[13]
  PIN uri_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1044.960 0.000 1045.520 4.000 ;
    END
  END uri_io_in[14]
  PIN uri_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1051.680 0.000 1052.240 4.000 ;
    END
  END uri_io_in[15]
  PIN uri_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1058.400 0.000 1058.960 4.000 ;
    END
  END uri_io_in[16]
  PIN uri_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1065.120 0.000 1065.680 4.000 ;
    END
  END uri_io_in[17]
  PIN uri_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1071.840 0.000 1072.400 4.000 ;
    END
  END uri_io_in[18]
  PIN uri_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1078.560 0.000 1079.120 4.000 ;
    END
  END uri_io_in[19]
  PIN uri_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 0.000 958.160 4.000 ;
    END
  END uri_io_in[1]
  PIN uri_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1085.280 0.000 1085.840 4.000 ;
    END
  END uri_io_in[20]
  PIN uri_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1092.000 0.000 1092.560 4.000 ;
    END
  END uri_io_in[21]
  PIN uri_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1098.720 0.000 1099.280 4.000 ;
    END
  END uri_io_in[22]
  PIN uri_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1105.440 0.000 1106.000 4.000 ;
    END
  END uri_io_in[23]
  PIN uri_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1112.160 0.000 1112.720 4.000 ;
    END
  END uri_io_in[24]
  PIN uri_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1118.880 0.000 1119.440 4.000 ;
    END
  END uri_io_in[25]
  PIN uri_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1125.600 0.000 1126.160 4.000 ;
    END
  END uri_io_in[26]
  PIN uri_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1132.320 0.000 1132.880 4.000 ;
    END
  END uri_io_in[27]
  PIN uri_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1139.040 0.000 1139.600 4.000 ;
    END
  END uri_io_in[28]
  PIN uri_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1145.760 0.000 1146.320 4.000 ;
    END
  END uri_io_in[29]
  PIN uri_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 964.320 0.000 964.880 4.000 ;
    END
  END uri_io_in[2]
  PIN uri_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1152.480 0.000 1153.040 4.000 ;
    END
  END uri_io_in[30]
  PIN uri_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1159.200 0.000 1159.760 4.000 ;
    END
  END uri_io_in[31]
  PIN uri_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1165.920 0.000 1166.480 4.000 ;
    END
  END uri_io_in[32]
  PIN uri_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1172.640 0.000 1173.200 4.000 ;
    END
  END uri_io_in[33]
  PIN uri_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1179.360 0.000 1179.920 4.000 ;
    END
  END uri_io_in[34]
  PIN uri_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1186.080 0.000 1186.640 4.000 ;
    END
  END uri_io_in[35]
  PIN uri_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1192.800 0.000 1193.360 4.000 ;
    END
  END uri_io_in[36]
  PIN uri_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1199.520 0.000 1200.080 4.000 ;
    END
  END uri_io_in[37]
  PIN uri_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 0.000 971.600 4.000 ;
    END
  END uri_io_in[3]
  PIN uri_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 977.760 0.000 978.320 4.000 ;
    END
  END uri_io_in[4]
  PIN uri_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 0.000 985.040 4.000 ;
    END
  END uri_io_in[5]
  PIN uri_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 0.000 991.760 4.000 ;
    END
  END uri_io_in[6]
  PIN uri_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 997.920 0.000 998.480 4.000 ;
    END
  END uri_io_in[7]
  PIN uri_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1004.640 0.000 1005.200 4.000 ;
    END
  END uri_io_in[8]
  PIN uri_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1011.360 0.000 1011.920 4.000 ;
    END
  END uri_io_in[9]
  PIN uri_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 0.000 823.760 4.000 ;
    END
  END uri_io_oeb[0]
  PIN uri_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 0.000 890.960 4.000 ;
    END
  END uri_io_oeb[10]
  PIN uri_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 0.000 897.680 4.000 ;
    END
  END uri_io_oeb[11]
  PIN uri_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 0.000 904.400 4.000 ;
    END
  END uri_io_oeb[12]
  PIN uri_io_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 910.560 0.000 911.120 4.000 ;
    END
  END uri_io_oeb[13]
  PIN uri_io_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 0.000 917.840 4.000 ;
    END
  END uri_io_oeb[14]
  PIN uri_io_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 924.000 0.000 924.560 4.000 ;
    END
  END uri_io_oeb[15]
  PIN uri_io_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 930.720 0.000 931.280 4.000 ;
    END
  END uri_io_oeb[16]
  PIN uri_io_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 0.000 938.000 4.000 ;
    END
  END uri_io_oeb[17]
  PIN uri_io_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 944.160 0.000 944.720 4.000 ;
    END
  END uri_io_oeb[18]
  PIN uri_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 0.000 830.480 4.000 ;
    END
  END uri_io_oeb[1]
  PIN uri_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 0.000 837.200 4.000 ;
    END
  END uri_io_oeb[2]
  PIN uri_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 0.000 843.920 4.000 ;
    END
  END uri_io_oeb[3]
  PIN uri_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 0.000 850.640 4.000 ;
    END
  END uri_io_oeb[4]
  PIN uri_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 0.000 857.360 4.000 ;
    END
  END uri_io_oeb[5]
  PIN uri_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 0.000 864.080 4.000 ;
    END
  END uri_io_oeb[6]
  PIN uri_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 0.000 870.800 4.000 ;
    END
  END uri_io_oeb[7]
  PIN uri_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 876.960 0.000 877.520 4.000 ;
    END
  END uri_io_oeb[8]
  PIN uri_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 0.000 884.240 4.000 ;
    END
  END uri_io_oeb[9]
  PIN uri_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 695.520 0.000 696.080 4.000 ;
    END
  END uri_io_out[0]
  PIN uri_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 0.000 763.280 4.000 ;
    END
  END uri_io_out[10]
  PIN uri_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 0.000 770.000 4.000 ;
    END
  END uri_io_out[11]
  PIN uri_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 0.000 776.720 4.000 ;
    END
  END uri_io_out[12]
  PIN uri_io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 0.000 783.440 4.000 ;
    END
  END uri_io_out[13]
  PIN uri_io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 0.000 790.160 4.000 ;
    END
  END uri_io_out[14]
  PIN uri_io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 796.320 0.000 796.880 4.000 ;
    END
  END uri_io_out[15]
  PIN uri_io_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 0.000 803.600 4.000 ;
    END
  END uri_io_out[16]
  PIN uri_io_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 809.760 0.000 810.320 4.000 ;
    END
  END uri_io_out[17]
  PIN uri_io_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 0.000 817.040 4.000 ;
    END
  END uri_io_out[18]
  PIN uri_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 702.240 0.000 702.800 4.000 ;
    END
  END uri_io_out[1]
  PIN uri_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 708.960 0.000 709.520 4.000 ;
    END
  END uri_io_out[2]
  PIN uri_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 0.000 716.240 4.000 ;
    END
  END uri_io_out[3]
  PIN uri_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 0.000 722.960 4.000 ;
    END
  END uri_io_out[4]
  PIN uri_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 0.000 729.680 4.000 ;
    END
  END uri_io_out[5]
  PIN uri_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 0.000 736.400 4.000 ;
    END
  END uri_io_out[6]
  PIN uri_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 0.000 743.120 4.000 ;
    END
  END uri_io_out[7]
  PIN uri_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 0.000 749.840 4.000 ;
    END
  END uri_io_out[8]
  PIN uri_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 0.000 756.560 4.000 ;
    END
  END uri_io_out[9]
  PIN uri_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 0.000 682.640 4.000 ;
    END
  END uri_rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 204.140 ;
    END
  END vdd
  PIN vgasp_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1401.120 216.000 1401.680 220.000 ;
    END
  END vgasp_clk
  PIN vgasp_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1414.560 216.000 1415.120 220.000 ;
    END
  END vgasp_ena
  PIN vgasp_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1831.200 216.000 1831.760 220.000 ;
    END
  END vgasp_io_in[0]
  PIN vgasp_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1764.000 216.000 1764.560 220.000 ;
    END
  END vgasp_io_in[10]
  PIN vgasp_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1757.280 216.000 1757.840 220.000 ;
    END
  END vgasp_io_in[11]
  PIN vgasp_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1750.560 216.000 1751.120 220.000 ;
    END
  END vgasp_io_in[12]
  PIN vgasp_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1743.840 216.000 1744.400 220.000 ;
    END
  END vgasp_io_in[13]
  PIN vgasp_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1737.120 216.000 1737.680 220.000 ;
    END
  END vgasp_io_in[14]
  PIN vgasp_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1730.400 216.000 1730.960 220.000 ;
    END
  END vgasp_io_in[15]
  PIN vgasp_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1723.680 216.000 1724.240 220.000 ;
    END
  END vgasp_io_in[16]
  PIN vgasp_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1716.960 216.000 1717.520 220.000 ;
    END
  END vgasp_io_in[17]
  PIN vgasp_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1710.240 216.000 1710.800 220.000 ;
    END
  END vgasp_io_in[18]
  PIN vgasp_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1703.520 216.000 1704.080 220.000 ;
    END
  END vgasp_io_in[19]
  PIN vgasp_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1824.480 216.000 1825.040 220.000 ;
    END
  END vgasp_io_in[1]
  PIN vgasp_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1696.800 216.000 1697.360 220.000 ;
    END
  END vgasp_io_in[20]
  PIN vgasp_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1690.080 216.000 1690.640 220.000 ;
    END
  END vgasp_io_in[21]
  PIN vgasp_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1683.360 216.000 1683.920 220.000 ;
    END
  END vgasp_io_in[22]
  PIN vgasp_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1676.640 216.000 1677.200 220.000 ;
    END
  END vgasp_io_in[23]
  PIN vgasp_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1669.920 216.000 1670.480 220.000 ;
    END
  END vgasp_io_in[24]
  PIN vgasp_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1663.200 216.000 1663.760 220.000 ;
    END
  END vgasp_io_in[25]
  PIN vgasp_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1656.480 216.000 1657.040 220.000 ;
    END
  END vgasp_io_in[26]
  PIN vgasp_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1649.760 216.000 1650.320 220.000 ;
    END
  END vgasp_io_in[27]
  PIN vgasp_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1643.040 216.000 1643.600 220.000 ;
    END
  END vgasp_io_in[28]
  PIN vgasp_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1636.320 216.000 1636.880 220.000 ;
    END
  END vgasp_io_in[29]
  PIN vgasp_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1817.760 216.000 1818.320 220.000 ;
    END
  END vgasp_io_in[2]
  PIN vgasp_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1629.600 216.000 1630.160 220.000 ;
    END
  END vgasp_io_in[30]
  PIN vgasp_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1622.880 216.000 1623.440 220.000 ;
    END
  END vgasp_io_in[31]
  PIN vgasp_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1616.160 216.000 1616.720 220.000 ;
    END
  END vgasp_io_in[32]
  PIN vgasp_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1609.440 216.000 1610.000 220.000 ;
    END
  END vgasp_io_in[33]
  PIN vgasp_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1602.720 216.000 1603.280 220.000 ;
    END
  END vgasp_io_in[34]
  PIN vgasp_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1596.000 216.000 1596.560 220.000 ;
    END
  END vgasp_io_in[35]
  PIN vgasp_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1589.280 216.000 1589.840 220.000 ;
    END
  END vgasp_io_in[36]
  PIN vgasp_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1582.560 216.000 1583.120 220.000 ;
    END
  END vgasp_io_in[37]
  PIN vgasp_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1811.040 216.000 1811.600 220.000 ;
    END
  END vgasp_io_in[3]
  PIN vgasp_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1804.320 216.000 1804.880 220.000 ;
    END
  END vgasp_io_in[4]
  PIN vgasp_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1797.600 216.000 1798.160 220.000 ;
    END
  END vgasp_io_in[5]
  PIN vgasp_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1790.880 216.000 1791.440 220.000 ;
    END
  END vgasp_io_in[6]
  PIN vgasp_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1784.160 216.000 1784.720 220.000 ;
    END
  END vgasp_io_in[7]
  PIN vgasp_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1777.440 216.000 1778.000 220.000 ;
    END
  END vgasp_io_in[8]
  PIN vgasp_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1770.720 216.000 1771.280 220.000 ;
    END
  END vgasp_io_in[9]
  PIN vgasp_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1407.840 216.000 1408.400 220.000 ;
    END
  END vgasp_rst
  PIN vgasp_uio_oe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1468.320 216.000 1468.880 220.000 ;
    END
  END vgasp_uio_oe[0]
  PIN vgasp_uio_oe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1461.600 216.000 1462.160 220.000 ;
    END
  END vgasp_uio_oe[1]
  PIN vgasp_uio_oe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1454.880 216.000 1455.440 220.000 ;
    END
  END vgasp_uio_oe[2]
  PIN vgasp_uio_oe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1448.160 216.000 1448.720 220.000 ;
    END
  END vgasp_uio_oe[3]
  PIN vgasp_uio_oe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1441.440 216.000 1442.000 220.000 ;
    END
  END vgasp_uio_oe[4]
  PIN vgasp_uio_oe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1434.720 216.000 1435.280 220.000 ;
    END
  END vgasp_uio_oe[5]
  PIN vgasp_uio_oe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1428.000 216.000 1428.560 220.000 ;
    END
  END vgasp_uio_oe[6]
  PIN vgasp_uio_oe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1421.280 216.000 1421.840 220.000 ;
    END
  END vgasp_uio_oe[7]
  PIN vgasp_uio_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1522.080 216.000 1522.640 220.000 ;
    END
  END vgasp_uio_out[0]
  PIN vgasp_uio_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1515.360 216.000 1515.920 220.000 ;
    END
  END vgasp_uio_out[1]
  PIN vgasp_uio_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1508.640 216.000 1509.200 220.000 ;
    END
  END vgasp_uio_out[2]
  PIN vgasp_uio_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1501.920 216.000 1502.480 220.000 ;
    END
  END vgasp_uio_out[3]
  PIN vgasp_uio_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1495.200 216.000 1495.760 220.000 ;
    END
  END vgasp_uio_out[4]
  PIN vgasp_uio_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1488.480 216.000 1489.040 220.000 ;
    END
  END vgasp_uio_out[5]
  PIN vgasp_uio_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1481.760 216.000 1482.320 220.000 ;
    END
  END vgasp_uio_out[6]
  PIN vgasp_uio_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1475.040 216.000 1475.600 220.000 ;
    END
  END vgasp_uio_out[7]
  PIN vgasp_uo_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1575.840 216.000 1576.400 220.000 ;
    END
  END vgasp_uo_out[0]
  PIN vgasp_uo_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1569.120 216.000 1569.680 220.000 ;
    END
  END vgasp_uo_out[1]
  PIN vgasp_uo_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1562.400 216.000 1562.960 220.000 ;
    END
  END vgasp_uo_out[2]
  PIN vgasp_uo_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1555.680 216.000 1556.240 220.000 ;
    END
  END vgasp_uo_out[3]
  PIN vgasp_uo_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1548.960 216.000 1549.520 220.000 ;
    END
  END vgasp_uo_out[4]
  PIN vgasp_uo_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1542.240 216.000 1542.800 220.000 ;
    END
  END vgasp_uo_out[5]
  PIN vgasp_uo_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1535.520 216.000 1536.080 220.000 ;
    END
  END vgasp_uo_out[6]
  PIN vgasp_uo_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1528.800 216.000 1529.360 220.000 ;
    END
  END vgasp_uo_out[7]
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 204.140 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.200 4.000 11.760 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.720 4.000 7.280 ;
    END
  END wb_rst_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 2392.880 208.730 ;
      LAYER Metal2 ;
        RECT 8.540 215.700 63.540 216.580 ;
        RECT 64.700 215.700 70.260 216.580 ;
        RECT 71.420 215.700 76.980 216.580 ;
        RECT 78.140 215.700 83.700 216.580 ;
        RECT 84.860 215.700 90.420 216.580 ;
        RECT 91.580 215.700 97.140 216.580 ;
        RECT 98.300 215.700 103.860 216.580 ;
        RECT 105.020 215.700 110.580 216.580 ;
        RECT 111.740 215.700 117.300 216.580 ;
        RECT 118.460 215.700 124.020 216.580 ;
        RECT 125.180 215.700 130.740 216.580 ;
        RECT 131.900 215.700 137.460 216.580 ;
        RECT 138.620 215.700 144.180 216.580 ;
        RECT 145.340 215.700 150.900 216.580 ;
        RECT 152.060 215.700 157.620 216.580 ;
        RECT 158.780 215.700 164.340 216.580 ;
        RECT 165.500 215.700 171.060 216.580 ;
        RECT 172.220 215.700 177.780 216.580 ;
        RECT 178.940 215.700 184.500 216.580 ;
        RECT 185.660 215.700 191.220 216.580 ;
        RECT 192.380 215.700 197.940 216.580 ;
        RECT 199.100 215.700 204.660 216.580 ;
        RECT 205.820 215.700 211.380 216.580 ;
        RECT 212.540 215.700 218.100 216.580 ;
        RECT 219.260 215.700 224.820 216.580 ;
        RECT 225.980 215.700 231.540 216.580 ;
        RECT 232.700 215.700 238.260 216.580 ;
        RECT 239.420 215.700 244.980 216.580 ;
        RECT 246.140 215.700 251.700 216.580 ;
        RECT 252.860 215.700 258.420 216.580 ;
        RECT 259.580 215.700 265.140 216.580 ;
        RECT 266.300 215.700 271.860 216.580 ;
        RECT 273.020 215.700 278.580 216.580 ;
        RECT 279.740 215.700 285.300 216.580 ;
        RECT 286.460 215.700 292.020 216.580 ;
        RECT 293.180 215.700 298.740 216.580 ;
        RECT 299.900 215.700 305.460 216.580 ;
        RECT 306.620 215.700 312.180 216.580 ;
        RECT 313.340 215.700 318.900 216.580 ;
        RECT 320.060 215.700 325.620 216.580 ;
        RECT 326.780 215.700 332.340 216.580 ;
        RECT 333.500 215.700 339.060 216.580 ;
        RECT 340.220 215.700 345.780 216.580 ;
        RECT 346.940 215.700 352.500 216.580 ;
        RECT 353.660 215.700 359.220 216.580 ;
        RECT 360.380 215.700 365.940 216.580 ;
        RECT 367.100 215.700 372.660 216.580 ;
        RECT 373.820 215.700 379.380 216.580 ;
        RECT 380.540 215.700 386.100 216.580 ;
        RECT 387.260 215.700 392.820 216.580 ;
        RECT 393.980 215.700 399.540 216.580 ;
        RECT 400.700 215.700 406.260 216.580 ;
        RECT 407.420 215.700 412.980 216.580 ;
        RECT 414.140 215.700 419.700 216.580 ;
        RECT 420.860 215.700 426.420 216.580 ;
        RECT 427.580 215.700 433.140 216.580 ;
        RECT 434.300 215.700 439.860 216.580 ;
        RECT 441.020 215.700 446.580 216.580 ;
        RECT 447.740 215.700 453.300 216.580 ;
        RECT 454.460 215.700 460.020 216.580 ;
        RECT 461.180 215.700 466.740 216.580 ;
        RECT 467.900 215.700 473.460 216.580 ;
        RECT 474.620 215.700 480.180 216.580 ;
        RECT 481.340 215.700 486.900 216.580 ;
        RECT 488.060 215.700 493.620 216.580 ;
        RECT 494.780 215.700 500.340 216.580 ;
        RECT 501.500 215.700 507.060 216.580 ;
        RECT 508.220 215.700 513.780 216.580 ;
        RECT 514.940 215.700 520.500 216.580 ;
        RECT 521.660 215.700 594.420 216.580 ;
        RECT 595.580 215.700 601.140 216.580 ;
        RECT 602.300 215.700 607.860 216.580 ;
        RECT 609.020 215.700 614.580 216.580 ;
        RECT 615.740 215.700 621.300 216.580 ;
        RECT 622.460 215.700 628.020 216.580 ;
        RECT 629.180 215.700 634.740 216.580 ;
        RECT 635.900 215.700 641.460 216.580 ;
        RECT 642.620 215.700 648.180 216.580 ;
        RECT 649.340 215.700 654.900 216.580 ;
        RECT 656.060 215.700 661.620 216.580 ;
        RECT 662.780 215.700 668.340 216.580 ;
        RECT 669.500 215.700 742.260 216.580 ;
        RECT 743.420 215.700 748.980 216.580 ;
        RECT 750.140 215.700 755.700 216.580 ;
        RECT 756.860 215.700 762.420 216.580 ;
        RECT 763.580 215.700 769.140 216.580 ;
        RECT 770.300 215.700 775.860 216.580 ;
        RECT 777.020 215.700 782.580 216.580 ;
        RECT 783.740 215.700 789.300 216.580 ;
        RECT 790.460 215.700 796.020 216.580 ;
        RECT 797.180 215.700 802.740 216.580 ;
        RECT 803.900 215.700 809.460 216.580 ;
        RECT 810.620 215.700 816.180 216.580 ;
        RECT 817.340 215.700 822.900 216.580 ;
        RECT 824.060 215.700 829.620 216.580 ;
        RECT 830.780 215.700 836.340 216.580 ;
        RECT 837.500 215.700 843.060 216.580 ;
        RECT 844.220 215.700 849.780 216.580 ;
        RECT 850.940 215.700 856.500 216.580 ;
        RECT 857.660 215.700 863.220 216.580 ;
        RECT 864.380 215.700 869.940 216.580 ;
        RECT 871.100 215.700 876.660 216.580 ;
        RECT 877.820 215.700 883.380 216.580 ;
        RECT 884.540 215.700 890.100 216.580 ;
        RECT 891.260 215.700 896.820 216.580 ;
        RECT 897.980 215.700 903.540 216.580 ;
        RECT 904.700 215.700 910.260 216.580 ;
        RECT 911.420 215.700 916.980 216.580 ;
        RECT 918.140 215.700 923.700 216.580 ;
        RECT 924.860 215.700 930.420 216.580 ;
        RECT 931.580 215.700 937.140 216.580 ;
        RECT 938.300 215.700 943.860 216.580 ;
        RECT 945.020 215.700 950.580 216.580 ;
        RECT 951.740 215.700 957.300 216.580 ;
        RECT 958.460 215.700 964.020 216.580 ;
        RECT 965.180 215.700 970.740 216.580 ;
        RECT 971.900 215.700 977.460 216.580 ;
        RECT 978.620 215.700 984.180 216.580 ;
        RECT 985.340 215.700 990.900 216.580 ;
        RECT 992.060 215.700 997.620 216.580 ;
        RECT 998.780 215.700 1004.340 216.580 ;
        RECT 1005.500 215.700 1011.060 216.580 ;
        RECT 1012.220 215.700 1017.780 216.580 ;
        RECT 1018.940 215.700 1024.500 216.580 ;
        RECT 1025.660 215.700 1031.220 216.580 ;
        RECT 1032.380 215.700 1037.940 216.580 ;
        RECT 1039.100 215.700 1044.660 216.580 ;
        RECT 1045.820 215.700 1051.380 216.580 ;
        RECT 1052.540 215.700 1058.100 216.580 ;
        RECT 1059.260 215.700 1064.820 216.580 ;
        RECT 1065.980 215.700 1071.540 216.580 ;
        RECT 1072.700 215.700 1078.260 216.580 ;
        RECT 1079.420 215.700 1084.980 216.580 ;
        RECT 1086.140 215.700 1091.700 216.580 ;
        RECT 1092.860 215.700 1098.420 216.580 ;
        RECT 1099.580 215.700 1105.140 216.580 ;
        RECT 1106.300 215.700 1111.860 216.580 ;
        RECT 1113.020 215.700 1118.580 216.580 ;
        RECT 1119.740 215.700 1125.300 216.580 ;
        RECT 1126.460 215.700 1132.020 216.580 ;
        RECT 1133.180 215.700 1138.740 216.580 ;
        RECT 1139.900 215.700 1145.460 216.580 ;
        RECT 1146.620 215.700 1152.180 216.580 ;
        RECT 1153.340 215.700 1158.900 216.580 ;
        RECT 1160.060 215.700 1165.620 216.580 ;
        RECT 1166.780 215.700 1172.340 216.580 ;
        RECT 1173.500 215.700 1179.060 216.580 ;
        RECT 1180.220 215.700 1185.780 216.580 ;
        RECT 1186.940 215.700 1192.500 216.580 ;
        RECT 1193.660 215.700 1199.220 216.580 ;
        RECT 1200.380 215.700 1273.140 216.580 ;
        RECT 1274.300 215.700 1279.860 216.580 ;
        RECT 1281.020 215.700 1286.580 216.580 ;
        RECT 1287.740 215.700 1293.300 216.580 ;
        RECT 1294.460 215.700 1300.020 216.580 ;
        RECT 1301.180 215.700 1306.740 216.580 ;
        RECT 1307.900 215.700 1313.460 216.580 ;
        RECT 1314.620 215.700 1320.180 216.580 ;
        RECT 1321.340 215.700 1326.900 216.580 ;
        RECT 1328.060 215.700 1400.820 216.580 ;
        RECT 1401.980 215.700 1407.540 216.580 ;
        RECT 1408.700 215.700 1414.260 216.580 ;
        RECT 1415.420 215.700 1420.980 216.580 ;
        RECT 1422.140 215.700 1427.700 216.580 ;
        RECT 1428.860 215.700 1434.420 216.580 ;
        RECT 1435.580 215.700 1441.140 216.580 ;
        RECT 1442.300 215.700 1447.860 216.580 ;
        RECT 1449.020 215.700 1454.580 216.580 ;
        RECT 1455.740 215.700 1461.300 216.580 ;
        RECT 1462.460 215.700 1468.020 216.580 ;
        RECT 1469.180 215.700 1474.740 216.580 ;
        RECT 1475.900 215.700 1481.460 216.580 ;
        RECT 1482.620 215.700 1488.180 216.580 ;
        RECT 1489.340 215.700 1494.900 216.580 ;
        RECT 1496.060 215.700 1501.620 216.580 ;
        RECT 1502.780 215.700 1508.340 216.580 ;
        RECT 1509.500 215.700 1515.060 216.580 ;
        RECT 1516.220 215.700 1521.780 216.580 ;
        RECT 1522.940 215.700 1528.500 216.580 ;
        RECT 1529.660 215.700 1535.220 216.580 ;
        RECT 1536.380 215.700 1541.940 216.580 ;
        RECT 1543.100 215.700 1548.660 216.580 ;
        RECT 1549.820 215.700 1555.380 216.580 ;
        RECT 1556.540 215.700 1562.100 216.580 ;
        RECT 1563.260 215.700 1568.820 216.580 ;
        RECT 1569.980 215.700 1575.540 216.580 ;
        RECT 1576.700 215.700 1582.260 216.580 ;
        RECT 1583.420 215.700 1588.980 216.580 ;
        RECT 1590.140 215.700 1595.700 216.580 ;
        RECT 1596.860 215.700 1602.420 216.580 ;
        RECT 1603.580 215.700 1609.140 216.580 ;
        RECT 1610.300 215.700 1615.860 216.580 ;
        RECT 1617.020 215.700 1622.580 216.580 ;
        RECT 1623.740 215.700 1629.300 216.580 ;
        RECT 1630.460 215.700 1636.020 216.580 ;
        RECT 1637.180 215.700 1642.740 216.580 ;
        RECT 1643.900 215.700 1649.460 216.580 ;
        RECT 1650.620 215.700 1656.180 216.580 ;
        RECT 1657.340 215.700 1662.900 216.580 ;
        RECT 1664.060 215.700 1669.620 216.580 ;
        RECT 1670.780 215.700 1676.340 216.580 ;
        RECT 1677.500 215.700 1683.060 216.580 ;
        RECT 1684.220 215.700 1689.780 216.580 ;
        RECT 1690.940 215.700 1696.500 216.580 ;
        RECT 1697.660 215.700 1703.220 216.580 ;
        RECT 1704.380 215.700 1709.940 216.580 ;
        RECT 1711.100 215.700 1716.660 216.580 ;
        RECT 1717.820 215.700 1723.380 216.580 ;
        RECT 1724.540 215.700 1730.100 216.580 ;
        RECT 1731.260 215.700 1736.820 216.580 ;
        RECT 1737.980 215.700 1743.540 216.580 ;
        RECT 1744.700 215.700 1750.260 216.580 ;
        RECT 1751.420 215.700 1756.980 216.580 ;
        RECT 1758.140 215.700 1763.700 216.580 ;
        RECT 1764.860 215.700 1770.420 216.580 ;
        RECT 1771.580 215.700 1777.140 216.580 ;
        RECT 1778.300 215.700 1783.860 216.580 ;
        RECT 1785.020 215.700 1790.580 216.580 ;
        RECT 1791.740 215.700 1797.300 216.580 ;
        RECT 1798.460 215.700 1804.020 216.580 ;
        RECT 1805.180 215.700 1810.740 216.580 ;
        RECT 1811.900 215.700 1817.460 216.580 ;
        RECT 1818.620 215.700 1824.180 216.580 ;
        RECT 1825.340 215.700 1830.900 216.580 ;
        RECT 1832.060 215.700 1904.820 216.580 ;
        RECT 1905.980 215.700 1911.540 216.580 ;
        RECT 1912.700 215.700 1918.260 216.580 ;
        RECT 1919.420 215.700 1924.980 216.580 ;
        RECT 1926.140 215.700 1931.700 216.580 ;
        RECT 1932.860 215.700 1938.420 216.580 ;
        RECT 1939.580 215.700 1945.140 216.580 ;
        RECT 1946.300 215.700 1951.860 216.580 ;
        RECT 1953.020 215.700 1958.580 216.580 ;
        RECT 1959.740 215.700 1965.300 216.580 ;
        RECT 1966.460 215.700 1972.020 216.580 ;
        RECT 1973.180 215.700 1978.740 216.580 ;
        RECT 1979.900 215.700 1985.460 216.580 ;
        RECT 1986.620 215.700 1992.180 216.580 ;
        RECT 1993.340 215.700 1998.900 216.580 ;
        RECT 2000.060 215.700 2005.620 216.580 ;
        RECT 2006.780 215.700 2012.340 216.580 ;
        RECT 2013.500 215.700 2019.060 216.580 ;
        RECT 2020.220 215.700 2025.780 216.580 ;
        RECT 2026.940 215.700 2032.500 216.580 ;
        RECT 2033.660 215.700 2039.220 216.580 ;
        RECT 2040.380 215.700 2045.940 216.580 ;
        RECT 2047.100 215.700 2052.660 216.580 ;
        RECT 2053.820 215.700 2059.380 216.580 ;
        RECT 2060.540 215.700 2066.100 216.580 ;
        RECT 2067.260 215.700 2072.820 216.580 ;
        RECT 2073.980 215.700 2079.540 216.580 ;
        RECT 2080.700 215.700 2086.260 216.580 ;
        RECT 2087.420 215.700 2092.980 216.580 ;
        RECT 2094.140 215.700 2099.700 216.580 ;
        RECT 2100.860 215.700 2106.420 216.580 ;
        RECT 2107.580 215.700 2113.140 216.580 ;
        RECT 2114.300 215.700 2119.860 216.580 ;
        RECT 2121.020 215.700 2126.580 216.580 ;
        RECT 2127.740 215.700 2133.300 216.580 ;
        RECT 2134.460 215.700 2140.020 216.580 ;
        RECT 2141.180 215.700 2146.740 216.580 ;
        RECT 2147.900 215.700 2153.460 216.580 ;
        RECT 2154.620 215.700 2160.180 216.580 ;
        RECT 2161.340 215.700 2166.900 216.580 ;
        RECT 2168.060 215.700 2173.620 216.580 ;
        RECT 2174.780 215.700 2180.340 216.580 ;
        RECT 2181.500 215.700 2187.060 216.580 ;
        RECT 2188.220 215.700 2193.780 216.580 ;
        RECT 2194.940 215.700 2200.500 216.580 ;
        RECT 2201.660 215.700 2207.220 216.580 ;
        RECT 2208.380 215.700 2213.940 216.580 ;
        RECT 2215.100 215.700 2220.660 216.580 ;
        RECT 2221.820 215.700 2227.380 216.580 ;
        RECT 2228.540 215.700 2234.100 216.580 ;
        RECT 2235.260 215.700 2240.820 216.580 ;
        RECT 2241.980 215.700 2247.540 216.580 ;
        RECT 2248.700 215.700 2254.260 216.580 ;
        RECT 2255.420 215.700 2260.980 216.580 ;
        RECT 2262.140 215.700 2267.700 216.580 ;
        RECT 2268.860 215.700 2391.620 216.580 ;
        RECT 8.540 4.300 2391.620 215.700 ;
        RECT 8.540 1.770 50.100 4.300 ;
        RECT 51.260 1.770 56.820 4.300 ;
        RECT 57.980 1.770 63.540 4.300 ;
        RECT 64.700 1.770 70.260 4.300 ;
        RECT 71.420 1.770 76.980 4.300 ;
        RECT 78.140 1.770 83.700 4.300 ;
        RECT 84.860 1.770 90.420 4.300 ;
        RECT 91.580 1.770 97.140 4.300 ;
        RECT 98.300 1.770 103.860 4.300 ;
        RECT 105.020 1.770 110.580 4.300 ;
        RECT 111.740 1.770 117.300 4.300 ;
        RECT 118.460 1.770 124.020 4.300 ;
        RECT 125.180 1.770 130.740 4.300 ;
        RECT 131.900 1.770 137.460 4.300 ;
        RECT 138.620 1.770 144.180 4.300 ;
        RECT 145.340 1.770 150.900 4.300 ;
        RECT 152.060 1.770 157.620 4.300 ;
        RECT 158.780 1.770 164.340 4.300 ;
        RECT 165.500 1.770 171.060 4.300 ;
        RECT 172.220 1.770 177.780 4.300 ;
        RECT 178.940 1.770 184.500 4.300 ;
        RECT 185.660 1.770 191.220 4.300 ;
        RECT 192.380 1.770 197.940 4.300 ;
        RECT 199.100 1.770 204.660 4.300 ;
        RECT 205.820 1.770 211.380 4.300 ;
        RECT 212.540 1.770 218.100 4.300 ;
        RECT 219.260 1.770 224.820 4.300 ;
        RECT 225.980 1.770 231.540 4.300 ;
        RECT 232.700 1.770 238.260 4.300 ;
        RECT 239.420 1.770 244.980 4.300 ;
        RECT 246.140 1.770 251.700 4.300 ;
        RECT 252.860 1.770 258.420 4.300 ;
        RECT 259.580 1.770 265.140 4.300 ;
        RECT 266.300 1.770 271.860 4.300 ;
        RECT 273.020 1.770 278.580 4.300 ;
        RECT 279.740 1.770 285.300 4.300 ;
        RECT 286.460 1.770 292.020 4.300 ;
        RECT 293.180 1.770 298.740 4.300 ;
        RECT 299.900 1.770 305.460 4.300 ;
        RECT 306.620 1.770 312.180 4.300 ;
        RECT 313.340 1.770 318.900 4.300 ;
        RECT 320.060 1.770 325.620 4.300 ;
        RECT 326.780 1.770 332.340 4.300 ;
        RECT 333.500 1.770 339.060 4.300 ;
        RECT 340.220 1.770 345.780 4.300 ;
        RECT 346.940 1.770 352.500 4.300 ;
        RECT 353.660 1.770 359.220 4.300 ;
        RECT 360.380 1.770 365.940 4.300 ;
        RECT 367.100 1.770 372.660 4.300 ;
        RECT 373.820 1.770 379.380 4.300 ;
        RECT 380.540 1.770 386.100 4.300 ;
        RECT 387.260 1.770 392.820 4.300 ;
        RECT 393.980 1.770 399.540 4.300 ;
        RECT 400.700 1.770 406.260 4.300 ;
        RECT 407.420 1.770 412.980 4.300 ;
        RECT 414.140 1.770 419.700 4.300 ;
        RECT 420.860 1.770 426.420 4.300 ;
        RECT 427.580 1.770 433.140 4.300 ;
        RECT 434.300 1.770 439.860 4.300 ;
        RECT 441.020 1.770 446.580 4.300 ;
        RECT 447.740 1.770 453.300 4.300 ;
        RECT 454.460 1.770 460.020 4.300 ;
        RECT 461.180 1.770 466.740 4.300 ;
        RECT 467.900 1.770 473.460 4.300 ;
        RECT 474.620 1.770 480.180 4.300 ;
        RECT 481.340 1.770 486.900 4.300 ;
        RECT 488.060 1.770 493.620 4.300 ;
        RECT 494.780 1.770 500.340 4.300 ;
        RECT 501.500 1.770 507.060 4.300 ;
        RECT 508.220 1.770 513.780 4.300 ;
        RECT 514.940 1.770 520.500 4.300 ;
        RECT 521.660 1.770 527.220 4.300 ;
        RECT 528.380 1.770 533.940 4.300 ;
        RECT 535.100 1.770 540.660 4.300 ;
        RECT 541.820 1.770 547.380 4.300 ;
        RECT 548.540 1.770 554.100 4.300 ;
        RECT 555.260 1.770 560.820 4.300 ;
        RECT 561.980 1.770 567.540 4.300 ;
        RECT 568.700 1.770 574.260 4.300 ;
        RECT 575.420 1.770 580.980 4.300 ;
        RECT 582.140 1.770 587.700 4.300 ;
        RECT 588.860 1.770 594.420 4.300 ;
        RECT 595.580 1.770 601.140 4.300 ;
        RECT 602.300 1.770 675.060 4.300 ;
        RECT 676.220 1.770 681.780 4.300 ;
        RECT 682.940 1.770 688.500 4.300 ;
        RECT 689.660 1.770 695.220 4.300 ;
        RECT 696.380 1.770 701.940 4.300 ;
        RECT 703.100 1.770 708.660 4.300 ;
        RECT 709.820 1.770 715.380 4.300 ;
        RECT 716.540 1.770 722.100 4.300 ;
        RECT 723.260 1.770 728.820 4.300 ;
        RECT 729.980 1.770 735.540 4.300 ;
        RECT 736.700 1.770 742.260 4.300 ;
        RECT 743.420 1.770 748.980 4.300 ;
        RECT 750.140 1.770 755.700 4.300 ;
        RECT 756.860 1.770 762.420 4.300 ;
        RECT 763.580 1.770 769.140 4.300 ;
        RECT 770.300 1.770 775.860 4.300 ;
        RECT 777.020 1.770 782.580 4.300 ;
        RECT 783.740 1.770 789.300 4.300 ;
        RECT 790.460 1.770 796.020 4.300 ;
        RECT 797.180 1.770 802.740 4.300 ;
        RECT 803.900 1.770 809.460 4.300 ;
        RECT 810.620 1.770 816.180 4.300 ;
        RECT 817.340 1.770 822.900 4.300 ;
        RECT 824.060 1.770 829.620 4.300 ;
        RECT 830.780 1.770 836.340 4.300 ;
        RECT 837.500 1.770 843.060 4.300 ;
        RECT 844.220 1.770 849.780 4.300 ;
        RECT 850.940 1.770 856.500 4.300 ;
        RECT 857.660 1.770 863.220 4.300 ;
        RECT 864.380 1.770 869.940 4.300 ;
        RECT 871.100 1.770 876.660 4.300 ;
        RECT 877.820 1.770 883.380 4.300 ;
        RECT 884.540 1.770 890.100 4.300 ;
        RECT 891.260 1.770 896.820 4.300 ;
        RECT 897.980 1.770 903.540 4.300 ;
        RECT 904.700 1.770 910.260 4.300 ;
        RECT 911.420 1.770 916.980 4.300 ;
        RECT 918.140 1.770 923.700 4.300 ;
        RECT 924.860 1.770 930.420 4.300 ;
        RECT 931.580 1.770 937.140 4.300 ;
        RECT 938.300 1.770 943.860 4.300 ;
        RECT 945.020 1.770 950.580 4.300 ;
        RECT 951.740 1.770 957.300 4.300 ;
        RECT 958.460 1.770 964.020 4.300 ;
        RECT 965.180 1.770 970.740 4.300 ;
        RECT 971.900 1.770 977.460 4.300 ;
        RECT 978.620 1.770 984.180 4.300 ;
        RECT 985.340 1.770 990.900 4.300 ;
        RECT 992.060 1.770 997.620 4.300 ;
        RECT 998.780 1.770 1004.340 4.300 ;
        RECT 1005.500 1.770 1011.060 4.300 ;
        RECT 1012.220 1.770 1017.780 4.300 ;
        RECT 1018.940 1.770 1024.500 4.300 ;
        RECT 1025.660 1.770 1031.220 4.300 ;
        RECT 1032.380 1.770 1037.940 4.300 ;
        RECT 1039.100 1.770 1044.660 4.300 ;
        RECT 1045.820 1.770 1051.380 4.300 ;
        RECT 1052.540 1.770 1058.100 4.300 ;
        RECT 1059.260 1.770 1064.820 4.300 ;
        RECT 1065.980 1.770 1071.540 4.300 ;
        RECT 1072.700 1.770 1078.260 4.300 ;
        RECT 1079.420 1.770 1084.980 4.300 ;
        RECT 1086.140 1.770 1091.700 4.300 ;
        RECT 1092.860 1.770 1098.420 4.300 ;
        RECT 1099.580 1.770 1105.140 4.300 ;
        RECT 1106.300 1.770 1111.860 4.300 ;
        RECT 1113.020 1.770 1118.580 4.300 ;
        RECT 1119.740 1.770 1125.300 4.300 ;
        RECT 1126.460 1.770 1132.020 4.300 ;
        RECT 1133.180 1.770 1138.740 4.300 ;
        RECT 1139.900 1.770 1145.460 4.300 ;
        RECT 1146.620 1.770 1152.180 4.300 ;
        RECT 1153.340 1.770 1158.900 4.300 ;
        RECT 1160.060 1.770 1165.620 4.300 ;
        RECT 1166.780 1.770 1172.340 4.300 ;
        RECT 1173.500 1.770 1179.060 4.300 ;
        RECT 1180.220 1.770 1185.780 4.300 ;
        RECT 1186.940 1.770 1192.500 4.300 ;
        RECT 1193.660 1.770 1199.220 4.300 ;
        RECT 1200.380 1.770 1273.140 4.300 ;
        RECT 1274.300 1.770 1279.860 4.300 ;
        RECT 1281.020 1.770 1286.580 4.300 ;
        RECT 1287.740 1.770 1293.300 4.300 ;
        RECT 1294.460 1.770 1300.020 4.300 ;
        RECT 1301.180 1.770 1306.740 4.300 ;
        RECT 1307.900 1.770 1313.460 4.300 ;
        RECT 1314.620 1.770 1320.180 4.300 ;
        RECT 1321.340 1.770 1326.900 4.300 ;
        RECT 1328.060 1.770 1333.620 4.300 ;
        RECT 1334.780 1.770 1340.340 4.300 ;
        RECT 1341.500 1.770 1347.060 4.300 ;
        RECT 1348.220 1.770 1353.780 4.300 ;
        RECT 1354.940 1.770 1360.500 4.300 ;
        RECT 1361.660 1.770 1367.220 4.300 ;
        RECT 1368.380 1.770 1373.940 4.300 ;
        RECT 1375.100 1.770 1515.060 4.300 ;
        RECT 1516.220 1.770 1521.780 4.300 ;
        RECT 1522.940 1.770 1528.500 4.300 ;
        RECT 1529.660 1.770 1535.220 4.300 ;
        RECT 1536.380 1.770 1541.940 4.300 ;
        RECT 1543.100 1.770 1548.660 4.300 ;
        RECT 1549.820 1.770 1555.380 4.300 ;
        RECT 1556.540 1.770 1562.100 4.300 ;
        RECT 1563.260 1.770 1568.820 4.300 ;
        RECT 1569.980 1.770 1575.540 4.300 ;
        RECT 1576.700 1.770 1582.260 4.300 ;
        RECT 1583.420 1.770 1588.980 4.300 ;
        RECT 1590.140 1.770 1595.700 4.300 ;
        RECT 1596.860 1.770 1602.420 4.300 ;
        RECT 1603.580 1.770 1609.140 4.300 ;
        RECT 1610.300 1.770 1615.860 4.300 ;
        RECT 1617.020 1.770 1622.580 4.300 ;
        RECT 1623.740 1.770 1629.300 4.300 ;
        RECT 1630.460 1.770 1636.020 4.300 ;
        RECT 1637.180 1.770 1642.740 4.300 ;
        RECT 1643.900 1.770 1649.460 4.300 ;
        RECT 1650.620 1.770 1656.180 4.300 ;
        RECT 1657.340 1.770 1662.900 4.300 ;
        RECT 1664.060 1.770 1669.620 4.300 ;
        RECT 1670.780 1.770 1676.340 4.300 ;
        RECT 1677.500 1.770 1683.060 4.300 ;
        RECT 1684.220 1.770 1689.780 4.300 ;
        RECT 1690.940 1.770 1696.500 4.300 ;
        RECT 1697.660 1.770 1703.220 4.300 ;
        RECT 1704.380 1.770 1709.940 4.300 ;
        RECT 1711.100 1.770 1716.660 4.300 ;
        RECT 1717.820 1.770 1723.380 4.300 ;
        RECT 1724.540 1.770 1730.100 4.300 ;
        RECT 1731.260 1.770 1736.820 4.300 ;
        RECT 1737.980 1.770 1743.540 4.300 ;
        RECT 1744.700 1.770 1750.260 4.300 ;
        RECT 1751.420 1.770 1756.980 4.300 ;
        RECT 1758.140 1.770 1763.700 4.300 ;
        RECT 1764.860 1.770 1770.420 4.300 ;
        RECT 1771.580 1.770 1777.140 4.300 ;
        RECT 1778.300 1.770 1783.860 4.300 ;
        RECT 1785.020 1.770 1790.580 4.300 ;
        RECT 1791.740 1.770 1797.300 4.300 ;
        RECT 1798.460 1.770 1804.020 4.300 ;
        RECT 1805.180 1.770 1810.740 4.300 ;
        RECT 1811.900 1.770 1817.460 4.300 ;
        RECT 1818.620 1.770 1824.180 4.300 ;
        RECT 1825.340 1.770 1830.900 4.300 ;
        RECT 1832.060 1.770 1837.620 4.300 ;
        RECT 1838.780 1.770 1844.340 4.300 ;
        RECT 1845.500 1.770 1851.060 4.300 ;
        RECT 1852.220 1.770 1857.780 4.300 ;
        RECT 1858.940 1.770 1864.500 4.300 ;
        RECT 1865.660 1.770 1871.220 4.300 ;
        RECT 1872.380 1.770 1877.940 4.300 ;
        RECT 1879.100 1.770 1884.660 4.300 ;
        RECT 1885.820 1.770 1891.380 4.300 ;
        RECT 1892.540 1.770 1898.100 4.300 ;
        RECT 1899.260 1.770 1904.820 4.300 ;
        RECT 1905.980 1.770 1911.540 4.300 ;
        RECT 1912.700 1.770 1918.260 4.300 ;
        RECT 1919.420 1.770 1924.980 4.300 ;
        RECT 1926.140 1.770 1931.700 4.300 ;
        RECT 1932.860 1.770 1938.420 4.300 ;
        RECT 1939.580 1.770 1945.140 4.300 ;
        RECT 1946.300 1.770 1951.860 4.300 ;
        RECT 1953.020 1.770 1958.580 4.300 ;
        RECT 1959.740 1.770 1965.300 4.300 ;
        RECT 1966.460 1.770 1972.020 4.300 ;
        RECT 1973.180 1.770 1978.740 4.300 ;
        RECT 1979.900 1.770 1985.460 4.300 ;
        RECT 1986.620 1.770 1992.180 4.300 ;
        RECT 1993.340 1.770 1998.900 4.300 ;
        RECT 2000.060 1.770 2005.620 4.300 ;
        RECT 2006.780 1.770 2012.340 4.300 ;
        RECT 2013.500 1.770 2019.060 4.300 ;
        RECT 2020.220 1.770 2025.780 4.300 ;
        RECT 2026.940 1.770 2032.500 4.300 ;
        RECT 2033.660 1.770 2039.220 4.300 ;
        RECT 2040.380 1.770 2045.940 4.300 ;
        RECT 2047.100 1.770 2052.660 4.300 ;
        RECT 2053.820 1.770 2059.380 4.300 ;
        RECT 2060.540 1.770 2066.100 4.300 ;
        RECT 2067.260 1.770 2072.820 4.300 ;
        RECT 2073.980 1.770 2079.540 4.300 ;
        RECT 2080.700 1.770 2086.260 4.300 ;
        RECT 2087.420 1.770 2092.980 4.300 ;
        RECT 2094.140 1.770 2099.700 4.300 ;
        RECT 2100.860 1.770 2106.420 4.300 ;
        RECT 2107.580 1.770 2113.140 4.300 ;
        RECT 2114.300 1.770 2119.860 4.300 ;
        RECT 2121.020 1.770 2126.580 4.300 ;
        RECT 2127.740 1.770 2133.300 4.300 ;
        RECT 2134.460 1.770 2140.020 4.300 ;
        RECT 2141.180 1.770 2146.740 4.300 ;
        RECT 2147.900 1.770 2153.460 4.300 ;
        RECT 2154.620 1.770 2160.180 4.300 ;
        RECT 2161.340 1.770 2166.900 4.300 ;
        RECT 2168.060 1.770 2173.620 4.300 ;
        RECT 2174.780 1.770 2180.340 4.300 ;
        RECT 2181.500 1.770 2187.060 4.300 ;
        RECT 2188.220 1.770 2193.780 4.300 ;
        RECT 2194.940 1.770 2200.500 4.300 ;
        RECT 2201.660 1.770 2207.220 4.300 ;
        RECT 2208.380 1.770 2213.940 4.300 ;
        RECT 2215.100 1.770 2391.620 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 214.740 2395.700 215.460 ;
        RECT 4.000 213.660 2396.000 214.740 ;
        RECT 4.300 212.540 2396.000 213.660 ;
        RECT 4.300 212.500 2395.700 212.540 ;
        RECT 4.000 211.380 2395.700 212.500 ;
        RECT 4.000 209.180 2396.000 211.380 ;
        RECT 4.300 208.020 2395.700 209.180 ;
        RECT 4.000 205.820 2396.000 208.020 ;
        RECT 4.000 204.700 2395.700 205.820 ;
        RECT 4.300 204.660 2395.700 204.700 ;
        RECT 4.300 203.540 2396.000 204.660 ;
        RECT 4.000 202.460 2396.000 203.540 ;
        RECT 4.000 201.300 2395.700 202.460 ;
        RECT 4.000 200.220 2396.000 201.300 ;
        RECT 4.300 199.100 2396.000 200.220 ;
        RECT 4.300 199.060 2395.700 199.100 ;
        RECT 4.000 197.940 2395.700 199.060 ;
        RECT 4.000 195.740 2396.000 197.940 ;
        RECT 4.300 194.580 2395.700 195.740 ;
        RECT 4.000 192.380 2396.000 194.580 ;
        RECT 4.000 191.260 2395.700 192.380 ;
        RECT 4.300 191.220 2395.700 191.260 ;
        RECT 4.300 190.100 2396.000 191.220 ;
        RECT 4.000 189.020 2396.000 190.100 ;
        RECT 4.000 187.860 2395.700 189.020 ;
        RECT 4.000 186.780 2396.000 187.860 ;
        RECT 4.300 185.660 2396.000 186.780 ;
        RECT 4.300 185.620 2395.700 185.660 ;
        RECT 4.000 184.500 2395.700 185.620 ;
        RECT 4.000 182.300 2396.000 184.500 ;
        RECT 4.300 181.140 2395.700 182.300 ;
        RECT 4.000 178.940 2396.000 181.140 ;
        RECT 4.000 177.820 2395.700 178.940 ;
        RECT 4.300 177.780 2395.700 177.820 ;
        RECT 4.300 176.660 2396.000 177.780 ;
        RECT 4.000 175.580 2396.000 176.660 ;
        RECT 4.000 174.420 2395.700 175.580 ;
        RECT 4.000 173.340 2396.000 174.420 ;
        RECT 4.300 172.220 2396.000 173.340 ;
        RECT 4.300 172.180 2395.700 172.220 ;
        RECT 4.000 171.060 2395.700 172.180 ;
        RECT 4.000 168.860 2396.000 171.060 ;
        RECT 4.300 167.700 2395.700 168.860 ;
        RECT 4.000 165.500 2396.000 167.700 ;
        RECT 4.000 164.380 2395.700 165.500 ;
        RECT 4.300 164.340 2395.700 164.380 ;
        RECT 4.300 163.220 2396.000 164.340 ;
        RECT 4.000 162.140 2396.000 163.220 ;
        RECT 4.000 160.980 2395.700 162.140 ;
        RECT 4.000 159.900 2396.000 160.980 ;
        RECT 4.300 158.780 2396.000 159.900 ;
        RECT 4.300 158.740 2395.700 158.780 ;
        RECT 4.000 157.620 2395.700 158.740 ;
        RECT 4.000 155.420 2396.000 157.620 ;
        RECT 4.300 154.260 2395.700 155.420 ;
        RECT 4.000 152.060 2396.000 154.260 ;
        RECT 4.000 150.940 2395.700 152.060 ;
        RECT 4.300 150.900 2395.700 150.940 ;
        RECT 4.300 149.780 2396.000 150.900 ;
        RECT 4.000 148.700 2396.000 149.780 ;
        RECT 4.000 147.540 2395.700 148.700 ;
        RECT 4.000 146.460 2396.000 147.540 ;
        RECT 4.300 145.340 2396.000 146.460 ;
        RECT 4.300 145.300 2395.700 145.340 ;
        RECT 4.000 144.180 2395.700 145.300 ;
        RECT 4.000 141.980 2396.000 144.180 ;
        RECT 4.300 140.820 2395.700 141.980 ;
        RECT 4.000 138.620 2396.000 140.820 ;
        RECT 4.000 137.500 2395.700 138.620 ;
        RECT 4.300 137.460 2395.700 137.500 ;
        RECT 4.300 136.340 2396.000 137.460 ;
        RECT 4.000 135.260 2396.000 136.340 ;
        RECT 4.000 134.100 2395.700 135.260 ;
        RECT 4.000 133.020 2396.000 134.100 ;
        RECT 4.300 131.900 2396.000 133.020 ;
        RECT 4.300 131.860 2395.700 131.900 ;
        RECT 4.000 130.740 2395.700 131.860 ;
        RECT 4.000 128.540 2396.000 130.740 ;
        RECT 4.300 127.380 2395.700 128.540 ;
        RECT 4.000 125.180 2396.000 127.380 ;
        RECT 4.000 124.060 2395.700 125.180 ;
        RECT 4.300 124.020 2395.700 124.060 ;
        RECT 4.300 122.900 2396.000 124.020 ;
        RECT 4.000 121.820 2396.000 122.900 ;
        RECT 4.000 120.660 2395.700 121.820 ;
        RECT 4.000 119.580 2396.000 120.660 ;
        RECT 4.300 118.460 2396.000 119.580 ;
        RECT 4.300 118.420 2395.700 118.460 ;
        RECT 4.000 117.300 2395.700 118.420 ;
        RECT 4.000 115.100 2396.000 117.300 ;
        RECT 4.300 113.940 2395.700 115.100 ;
        RECT 4.000 111.740 2396.000 113.940 ;
        RECT 4.000 110.620 2395.700 111.740 ;
        RECT 4.300 110.580 2395.700 110.620 ;
        RECT 4.300 109.460 2396.000 110.580 ;
        RECT 4.000 108.380 2396.000 109.460 ;
        RECT 4.000 107.220 2395.700 108.380 ;
        RECT 4.000 106.140 2396.000 107.220 ;
        RECT 4.300 105.020 2396.000 106.140 ;
        RECT 4.300 104.980 2395.700 105.020 ;
        RECT 4.000 103.860 2395.700 104.980 ;
        RECT 4.000 101.660 2396.000 103.860 ;
        RECT 4.300 100.500 2395.700 101.660 ;
        RECT 4.000 98.300 2396.000 100.500 ;
        RECT 4.000 97.180 2395.700 98.300 ;
        RECT 4.300 97.140 2395.700 97.180 ;
        RECT 4.300 96.020 2396.000 97.140 ;
        RECT 4.000 94.940 2396.000 96.020 ;
        RECT 4.000 93.780 2395.700 94.940 ;
        RECT 4.000 92.700 2396.000 93.780 ;
        RECT 4.300 91.580 2396.000 92.700 ;
        RECT 4.300 91.540 2395.700 91.580 ;
        RECT 4.000 90.420 2395.700 91.540 ;
        RECT 4.000 88.220 2396.000 90.420 ;
        RECT 4.300 87.060 2395.700 88.220 ;
        RECT 4.000 84.860 2396.000 87.060 ;
        RECT 4.000 83.740 2395.700 84.860 ;
        RECT 4.300 83.700 2395.700 83.740 ;
        RECT 4.300 82.580 2396.000 83.700 ;
        RECT 4.000 81.500 2396.000 82.580 ;
        RECT 4.000 80.340 2395.700 81.500 ;
        RECT 4.000 79.260 2396.000 80.340 ;
        RECT 4.300 78.140 2396.000 79.260 ;
        RECT 4.300 78.100 2395.700 78.140 ;
        RECT 4.000 76.980 2395.700 78.100 ;
        RECT 4.000 74.780 2396.000 76.980 ;
        RECT 4.300 73.620 2395.700 74.780 ;
        RECT 4.000 71.420 2396.000 73.620 ;
        RECT 4.000 70.300 2395.700 71.420 ;
        RECT 4.300 70.260 2395.700 70.300 ;
        RECT 4.300 69.140 2396.000 70.260 ;
        RECT 4.000 68.060 2396.000 69.140 ;
        RECT 4.000 66.900 2395.700 68.060 ;
        RECT 4.000 65.820 2396.000 66.900 ;
        RECT 4.300 64.700 2396.000 65.820 ;
        RECT 4.300 64.660 2395.700 64.700 ;
        RECT 4.000 63.540 2395.700 64.660 ;
        RECT 4.000 61.340 2396.000 63.540 ;
        RECT 4.300 60.180 2395.700 61.340 ;
        RECT 4.000 57.980 2396.000 60.180 ;
        RECT 4.000 56.860 2395.700 57.980 ;
        RECT 4.300 56.820 2395.700 56.860 ;
        RECT 4.300 55.700 2396.000 56.820 ;
        RECT 4.000 54.620 2396.000 55.700 ;
        RECT 4.000 53.460 2395.700 54.620 ;
        RECT 4.000 52.380 2396.000 53.460 ;
        RECT 4.300 51.260 2396.000 52.380 ;
        RECT 4.300 51.220 2395.700 51.260 ;
        RECT 4.000 50.100 2395.700 51.220 ;
        RECT 4.000 47.900 2396.000 50.100 ;
        RECT 4.300 46.740 2395.700 47.900 ;
        RECT 4.000 44.540 2396.000 46.740 ;
        RECT 4.000 43.420 2395.700 44.540 ;
        RECT 4.300 43.380 2395.700 43.420 ;
        RECT 4.300 42.260 2396.000 43.380 ;
        RECT 4.000 41.180 2396.000 42.260 ;
        RECT 4.000 40.020 2395.700 41.180 ;
        RECT 4.000 38.940 2396.000 40.020 ;
        RECT 4.300 37.820 2396.000 38.940 ;
        RECT 4.300 37.780 2395.700 37.820 ;
        RECT 4.000 36.660 2395.700 37.780 ;
        RECT 4.000 34.460 2396.000 36.660 ;
        RECT 4.300 33.300 2395.700 34.460 ;
        RECT 4.000 31.100 2396.000 33.300 ;
        RECT 4.000 29.980 2395.700 31.100 ;
        RECT 4.300 29.940 2395.700 29.980 ;
        RECT 4.300 28.820 2396.000 29.940 ;
        RECT 4.000 27.740 2396.000 28.820 ;
        RECT 4.000 26.580 2395.700 27.740 ;
        RECT 4.000 25.500 2396.000 26.580 ;
        RECT 4.300 24.380 2396.000 25.500 ;
        RECT 4.300 24.340 2395.700 24.380 ;
        RECT 4.000 23.220 2395.700 24.340 ;
        RECT 4.000 21.020 2396.000 23.220 ;
        RECT 4.300 19.860 2395.700 21.020 ;
        RECT 4.000 17.660 2396.000 19.860 ;
        RECT 4.000 16.540 2395.700 17.660 ;
        RECT 4.300 16.500 2395.700 16.540 ;
        RECT 4.300 15.380 2396.000 16.500 ;
        RECT 4.000 14.300 2396.000 15.380 ;
        RECT 4.000 13.140 2395.700 14.300 ;
        RECT 4.000 12.060 2396.000 13.140 ;
        RECT 4.300 10.940 2396.000 12.060 ;
        RECT 4.300 10.900 2395.700 10.940 ;
        RECT 4.000 9.780 2395.700 10.900 ;
        RECT 4.000 7.580 2396.000 9.780 ;
        RECT 4.300 6.420 2395.700 7.580 ;
        RECT 4.000 4.220 2396.000 6.420 ;
        RECT 4.000 3.060 2395.700 4.220 ;
        RECT 4.000 1.820 2396.000 3.060 ;
      LAYER Metal4 ;
        RECT 409.500 18.010 482.740 201.510 ;
        RECT 484.940 18.010 559.540 201.510 ;
        RECT 561.740 18.010 636.340 201.510 ;
        RECT 638.540 18.010 713.140 201.510 ;
        RECT 715.340 18.010 789.940 201.510 ;
        RECT 792.140 18.010 866.740 201.510 ;
        RECT 868.940 18.010 943.540 201.510 ;
        RECT 945.740 18.010 1020.340 201.510 ;
        RECT 1022.540 18.010 1097.140 201.510 ;
        RECT 1099.340 18.010 1173.940 201.510 ;
        RECT 1176.140 18.010 1250.740 201.510 ;
        RECT 1252.940 18.010 1327.540 201.510 ;
        RECT 1329.740 18.010 1404.340 201.510 ;
        RECT 1406.540 18.010 1481.140 201.510 ;
        RECT 1483.340 18.010 1557.940 201.510 ;
        RECT 1560.140 18.010 1600.340 201.510 ;
  END
END top_design_mux
END LIBRARY

