* NGSPICE file created from top_vga_spi_rom.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

.subckt top_vga_spi_rom clk rst ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5]
+ ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6]
+ uio_in[7] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] vdd vss uio_oe[0]
+ uio_out[6]
XANTENNA__1343__B _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2037_ net39 clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.r_rgb\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_52_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1270_ _0380_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[18\] _0671_ _0457_
+ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_46_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1606_ _0579_ _0905_ _0181_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1295__S0 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0985_ _0390_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1537_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[9\] _0907_ _0912_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1399_ _0800_ net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1468_ _0856_ _0837_ _0858_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_49_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__A1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[64\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1672__I _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1322_ _0722_ _0723_ _0496_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1253_ _0363_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1184_ _0492_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1340__C _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0968_ _0376_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1940_ _0057_ clknet_4_6_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[45\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1871_ _0332_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_24_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1236_ _0613_ _0619_ _0636_ _0637_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1305_ _0405_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_19_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1167_ _0568_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[47\] _0569_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1098_ _0494_ _0502_ _0505_ net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_42_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1030__A2 _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_44_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1021_ _0425_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1923_ _0040_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1854_ _0329_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1785_ _0284_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1219_ _0427_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1251__A2 _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1570_ _0930_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1004_ _0347_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1906_ _0023_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1768_ _0275_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1837_ _0536_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1699_ _0235_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_11_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput20 net20 uo_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1942__CLKN clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1622_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[45\] _0184_ _0192_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1957__CLKN clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1553_ _0920_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1484_ _0549_ _0822_ _0868_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_52_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2036_ _0153_ clknet_4_8_0_clk tt_um_algofoogle_vga_spi_rom.r_rgb\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1896__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0984_ _0387_ _0392_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1605_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[39\] _0907_ _0181_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1536_ _0651_ _0909_ _0911_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1295__S1 _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1354__B _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1467_ _0857_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1398_ _0799_ tt_um_algofoogle_vga_spi_rom.r_rgb\[2\] _0553_ _0800_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2019_ _0136_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[124\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1363__A1 _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1252_ _0560_ _0646_ _0653_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1321_ _0494_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[106\] _0723_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1183_ _0379_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0967_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.quad _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_58_Left_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1519_ _0899_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_25_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1336__A1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1870_ _0375_ _0335_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1327__A1 _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1887__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1166_ _0431_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1304_ _0364_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[114\] _0704_
+ _0705_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1235_ _0418_ _0453_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1097_ _0401_ _0502_ _0504_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1999_ _0116_ clknet_4_4_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[104\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_30_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2042__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output12_I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1020_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[3\] _0426_ _0428_
+ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1922_ _0039_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1853_ _0326_ _0799_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1784_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[116\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[115\]
+ _0281_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1149_ _0549_ _0551_ _0543_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1218_ _0426_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_7_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1003_ _0352_ _0405_ _0409_ _0411_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_44_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1905_ _0022_ clknet_4_6_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_32_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1698_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[79\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[78\]
+ _0231_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1767_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[108\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[107\]
+ _0274_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1836_ _0696_ _0817_ _0443_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1871__I _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1267__B _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 net21 uo_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1552_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[17\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[16\]
+ _0918_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1621_ _0191_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1691__I _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1483_ _0859_ _0870_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input3_I ui_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2035_ _0152_ clknet_4_8_0_clk tt_um_algofoogle_vga_spi_rom.r_rgb\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1819_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[131\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[130\]
+ _0302_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0983_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.quad _0388_ _0390_ _0391_ _0392_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_13_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1604_ _0180_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1535_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[9\] _0910_ _0911_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1372__A2 _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1466_ net1 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1397_ _0794_ _0797_ _0798_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2018_ _0135_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[123\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1956__CLKN clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1909__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1354__A2 _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1320_ _0364_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[107\] _0722_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1251_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[9\] _0574_ _0650_ _0652_
+ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1182_ _0583_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_19_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0966_ _0369_ _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1518_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[4\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[3\]
+ _0896_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1365__B _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1449_ _0840_ _0842_ _0843_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1281__A1 _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1336__A2 _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2009__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1024__A1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1303_ _0629_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1234_ _0623_ _0627_ _0630_ _0634_ _0635_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1165_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[46\] _0567_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1096_ _0503_ _0387_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1998_ _0115_ clknet_4_4_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[103\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0949_ _0354_ _0357_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1309__A2 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1921_ _0038_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1852_ _0328_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1783_ _0283_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1217_ _0615_ _0618_ _0466_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_35_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1079_ _0411_ _0465_ _0483_ _0487_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_1_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1148_ _0550_ net37 _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1109__I _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold10 _0810_ net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_41_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1779__I _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1002_ _0410_ _0383_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1904_ _0021_ clknet_4_6_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_32_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1769__A2 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1835_ _0813_ _0311_ _0314_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1697_ _0234_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1766_ _0261_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2032__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xoutput22 net22 uo_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1551_ _0919_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1620_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[45\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[44\]
+ _0189_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1482_ _0549_ _0869_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2034_ _0151_ clknet_4_2_0_clk tt_um_algofoogle_vga_spi_rom.r_rgb\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1818_ _0303_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1749_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[100\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[99\]
+ _0262_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtop_vga_spi_rom_30 uio_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_7_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1278__B _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0982_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[8\] _0391_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1603_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[39\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[38\]
+ _0176_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1534_ _0890_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1465_ _0821_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1396_ _0541_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2017_ _0134_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[122\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_13_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1117__I tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1250_ _0651_ _0441_ _0626_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1181_ _0404_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_19_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0965_ _0373_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1517_ _0898_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1448_ _0841_ _0815_ _0824_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1379_ _0620_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[74\] _0780_ _0629_
+ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_45_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1033__A2 _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1233_ _0352_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1302_ _0703_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[115\] _0704_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_59_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1164_ _0565_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1095_ _0464_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1940__CLKN clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1997_ _0114_ clknet_4_4_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[102\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_0948_ _0355_ _0356_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1376__B _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1955__CLKN clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1908__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1920_ _0037_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1851_ _0326_ net45 _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1782_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[115\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[114\]
+ _0281_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1556__I0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1216_ _0616_ _0617_ _0459_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_35_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1078_ _0484_ _0421_ _0407_ _0486_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1147_ net11 _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2008__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold11 net49 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_11_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1463__C _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1001_ _0370_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1903_ _0020_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_32_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1765_ _0273_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1834_ _0444_ _0312_ _0386_ _0313_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_1696_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[78\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[77\]
+ _0231_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1209__A2 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput12 net12 uio_oe[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput23 net23 uo_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1550_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[16\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[15\]
+ _0918_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1481_ _0822_ _0868_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2033_ net43 clknet_4_2_0_clk tt_um_algofoogle_vga_spi_rom.r_rgb\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1748_ _0264_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1817_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[130\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[129\]
+ _0302_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_15_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1679_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[71\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[70\]
+ _0220_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtop_vga_spi_rom_31 uio_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0981_ _0389_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[7\] _0390_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1602_ _0179_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1357__A1 _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1533_ _0904_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1395_ _0491_ _0796_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1464_ _0829_ _0822_ _0854_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2016_ _0133_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[121\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_57_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2045__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1180_ _0560_ _0572_ _0581_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1043__I _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1199__B _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0964_ _0370_ _0371_ _0372_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1516_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[3\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[2\]
+ _0896_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1447_ _0815_ _0823_ _0841_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1378_ _0621_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[75\] _0780_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1128__I tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1798__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Left_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_24_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_6_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1232_ _0631_ _0633_ _0583_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1301_ _0492_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1163_ _0355_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1094_ _0393_ _0399_ _0501_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_19_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1996_ _0113_ clknet_4_4_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[101\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_0947_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[1\] _0356_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_30_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1286__C _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_3_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1850_ _0840_ _0805_ net42 _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1781_ _0282_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1215_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[53\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[52\]
+ _0598_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1146_ _0548_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1077_ _0485_ _0415_ _0480_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1979_ _0096_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[84\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
Xhold12 net48 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_58_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1000_ _0408_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1954__CLKN clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1902_ _0019_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1710__I1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[83\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1969__CLKN clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1764_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[107\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[106\]
+ _0267_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1833_ _0560_ _0384_ _0503_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1907__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1695_ _0233_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1162__S _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1129_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[0\] _0533_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_14_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput24 net24 uo_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput13 net13 uio_oe[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_hold5_I uio_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2007__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1480_ _0864_ _0865_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2032_ _0149_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.r_hsync vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1747_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[99\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[98\]
+ _0262_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1678_ _0223_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1816_ _0286_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xtop_vga_spi_rom_32 uio_oe[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1054__A1 _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0980_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[6\] _0389_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1601_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[38\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[37\]
+ _0176_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1532_ _0651_ _0905_ _0908_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input1_I rst vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1394_ _0550_ net9 _0795_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1463_ _0851_ _0853_ _0854_ _0823_ _0813_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_49_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2015_ _0132_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[120\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1379__C _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1348__A2 _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1289__C _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_2_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0963_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[5\] _0372_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1027__A1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1515_ _0897_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1377_ _0776_ _0778_ _0466_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1446_ _0532_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1231_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[57\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[56\]
+ _0632_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1162_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[45\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[44\]
+ _0563_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1300_ _0695_ _0701_ _0384_ _0506_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1248__A1 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1093_ _0496_ _0498_ _0400_ _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_1995_ _0112_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[100\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_42_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0946_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[0\] _0355_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2035__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1420__A1 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1392__C _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1429_ _0530_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1780_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[114\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[113\]
+ _0281_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1512__I _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1214_ _0414_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1145_ _0462_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1076_ _0413_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1387__C _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1978_ _0095_ clknet_4_13_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[83\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_30_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_10_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold13 uio_in[2] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1901_ _0018_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1832_ _0402_ _0450_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1763_ _0725_ _0251_ _0272_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1694_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[77\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[76\]
+ _0231_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1862__A1 _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1059_ _0465_ _0467_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1128_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[1\] _0532_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput14 net14 uio_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput25 net25 uo_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1417__I _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1853__A1 _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1890__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2031_ _0148_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.hsync vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1844__A1 _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1815_ _0301_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1746_ _0263_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1677_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[70\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[69\]
+ _0220_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtop_vga_spi_rom_33 uio_oe[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_0_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1700__I _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1835__A1 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1953__CLKN clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1968__CLKN clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1610__I _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1906__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1600_ _0178_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1531_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[7\] _0907_ _0908_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1462_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[4\] _0833_ _0852_
+ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_38_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1393_ _0548_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2014_ _0131_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[119\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_5_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1729_ _0752_ _0251_ _0253_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_5_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2006__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0962_ _0361_ _0347_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_index\[3\] _0348_
+ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_6_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1496__B _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1514_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[2\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[1\]
+ _0896_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1445_ _0815_ _0823_ _0839_ _0840_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1376_ _0616_ _0777_ _0626_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_2_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1193__A1 _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1230_ _0431_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1161_ _0562_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1092_ _0450_ _0499_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_19_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1994_ _0111_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[99\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_19_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0945_ _0348_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1428_ _0821_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1359_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[84\] _0674_ _0761_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1175__A1 _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1213_ _0484_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[54\] _0614_ _0608_
+ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1075_ _0379_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1144_ _0547_ net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1977_ _0094_ clknet_4_14_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[82\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_7_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold14 ui_in[0] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_11_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1814__S _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1320__A1 _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1900_ _0017_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_32_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1831_ _0498_ _0500_ _0726_ _0310_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1762_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[106\] _0252_ _0272_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1693_ _0232_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1862__A2 _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1058_ _0466_ _0444_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1127_ _0522_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput15 net15 uio_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2048__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1369__A1 _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2030_ _0147_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[135\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1745_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[98\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[97\]
+ _0262_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1814_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[129\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[128\]
+ _0297_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1676_ _0222_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtop_vga_spi_rom_34 uio_oe[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1530_ _0906_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1461_ _0848_ _0823_ _0852_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1392_ _0555_ net9 _0793_ _0378_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2013_ _0130_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[118\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XPHY_EDGE_ROW_19_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1728_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[91\] _0252_ _0253_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1659_ _0207_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_5_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1158__I _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0961_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[4\] _0370_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1513_ _0895_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1375_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[69\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[68\]
+ _0632_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1444_ _0812_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1952__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1967__CLKN clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1905__CLKN clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1160_ _0346_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1091_ _0417_ _0365_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_51_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1993_ _0110_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[98\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XPHY_EDGE_ROW_41_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0944_ _0352_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_Left_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1358_ _0585_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[86\] _0759_ _0457_
+ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2005__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1427_ _0822_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1289_ _0684_ _0686_ _0688_ _0690_ _0635_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_33_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1212_ _0576_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[55\] _0614_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_47_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1074_ _0480_ _0481_ _0482_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1143_ _0546_ tt_um_algofoogle_vga_spi_rom.r_rgb\[4\] _0511_ _0547_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1976_ _0093_ clknet_4_14_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[81\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold15 uio_in[7] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_38_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_7_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1093__A1 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1166__I _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1761_ _0725_ _0248_ _0271_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1830_ _0536_ _0506_ _0309_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1692_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[76\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[75\]
+ _0231_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1126_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[9\] _0530_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1057_ _0417_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1959_ _0076_ clknet_4_11_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[64\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_28_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput16 net36 uio_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1825__S _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1744_ _0261_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1813_ _0300_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1675_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[69\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[68\]
+ _0220_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtop_vga_spi_rom_35 uio_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_7_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1109_ _0513_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1296__A1 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1709__I _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1444__I _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1380__S _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1211__A1 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1460_ _0388_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[1\] _0533_
+ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1391_ _0694_ _0702_ _0792_ _0555_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1278__A1 _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2012_ _0129_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[117\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_45_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2038__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1727_ _0890_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1658_ _0212_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1589_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[33\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[32\]
+ _0170_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0960_ _0368_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1512_ _0894_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1374_ _0484_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[70\] _0775_ _0608_
+ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_4_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1443_ _0815_ _0838_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1499__A1 _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1423__A1 _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1090_ _0497_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1992_ _0109_ clknet_4_4_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[97\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_27_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0943_ _0351_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1807__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1357_ _0586_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[87\] _0759_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1288_ _0608_ _0689_ _0626_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1426_ _0821_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1951__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1211_ _0497_ _0609_ _0611_ _0612_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1142_ _0543_ _0545_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1073_ _0376_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_23_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1904__CLKN clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1975_ _0092_ clknet_4_14_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[80\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_15_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1919__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1409_ _0808_ net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1093__A2 _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_40_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1760_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[104\] _0249_ _0271_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1691_ _0230_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2004__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2019__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1125_ _0513_ _0528_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1056_ _0464_ _0393_ _0399_ _0400_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_43_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1958_ _0075_ clknet_4_11_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[63\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_3_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput17 net17 uio_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1889_ _0006_ clknet_4_2_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1216__B _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1838__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1730__I _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1674_ _0221_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1743_ _0206_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1812_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[128\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[127\]
+ _0297_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1108_ net2 _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1039_ _0360_ _0382_ _0423_ _0447_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_48_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_10_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1390_ _0721_ _0747_ _0790_ _0791_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_57_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2011_ _0128_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[116\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1588_ _0171_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1726_ _0891_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1657_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[61\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[60\]
+ _0208_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1269__A2 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1511_ _0889_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1442_ _0824_ _0837_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1373_ _0568_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[71\] _0775_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1499__A2 _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1709_ _0230_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_51_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0973__B _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1991_ _0108_ clknet_4_4_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[96\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1169__A1 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1405__A2 _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0942_ _0350_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1425_ _0816_ _0819_ _0820_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1287_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[31\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[30\]
+ _0632_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1356_ _0635_ _0751_ _0757_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_33_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1707__I0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[83\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1210_ _0585_ _0597_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[49\] _0612_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1072_ _0415_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1141_ net37 _0544_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1974_ _0091_ clknet_4_14_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[79\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_28_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1311__C _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1408_ _0807_ tt_um_algofoogle_vga_spi_rom.r_rgb\[0\] _0553_ _0808_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1339_ _0493_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[101\] _0741_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1865__A2 _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1221__C _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1690_ _0206_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1306__C _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1322__B _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1055_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[9\] _0464_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1124_ _0462_ _0521_ _0527_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1957_ _0074_ clknet_4_11_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[62\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_43_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput18 net18 uo_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1888_ _0005_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1883__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1838__A2 _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1950__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1918__CLKN clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1903__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1811_ _0299_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1742_ _0260_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1673_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[68\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[67\]
+ _0220_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtop_vga_spi_rom_26 uio_oe[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_7_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1038_ _0360_ _0446_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1107_ _0512_ net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2003__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2018__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2010_ _0127_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[115\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_54_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1725_ _0752_ _0248_ _0250_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1587_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[32\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[31\]
+ _0170_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1656_ _0211_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1510_ _0893_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_10_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1441_ _0825_ _0827_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1372_ _0770_ _0726_ _0772_ _0773_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1314__C _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1708_ _0240_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1639_ _0175_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_36_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1178__A2 _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1990_ _0107_ clknet_4_4_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[95\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_0941_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_index\[3\] _0350_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_15_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1309__C _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1355_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[89\] _0574_ _0754_ _0756_
+ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1424_ _0712_ _0536_ _0590_ _0411_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_38_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1286_ _0682_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[28\] _0687_ _0485_
+ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_46_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1332__A2 _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1196__I _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1020__A1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1071_ _0350_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1140_ _0378_ net11 _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_55_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ _0090_ clknet_4_11_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[78\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_23_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1338_ _0452_ _0737_ _0738_ _0739_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1407_ _0805_ _0806_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1314__A2 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1269_ _0648_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[19\] _0671_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1744__I _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1054_ _0452_ _0458_ _0461_ _0462_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1123_ _0523_ _0526_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1887_ _0004_ clknet_4_2_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1956_ _0073_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[61\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 uo_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1741_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[97\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[96\]
+ _0254_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1810_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[127\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[126\]
+ _0297_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1672_ _0207_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xtop_vga_spi_rom_27 uio_oe[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1317__C _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1106_ tt_um_algofoogle_vga_spi_rom.hsync tt_um_algofoogle_vga_spi_rom.r_hsync _0511_
+ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1037_ _0430_ _0434_ _0437_ _0440_ _0442_ _0445_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__1205__A1 _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1939_ _0056_ clknet_4_6_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[44\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_16_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_48_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_57_Left_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1724_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[89\] _0249_ _0250_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1586_ _0923_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_0_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1655_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[60\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[59\]
+ _0208_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1902__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1979__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1917__CLKN clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold1_I uio_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1371_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[64\] _0460_ _0600_ _0773_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1440_ _0830_ _0831_ _0832_ _0835_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2002__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1638_ _0200_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1707_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[83\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[82\]
+ _0236_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2017__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1569_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[24\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[23\]
+ _0929_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1670__I1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[66\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0940_ _0346_ _0347_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_index\[3\] _0348_
+ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1285_ _0621_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[29\] _0687_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1354_ _0755_ _0441_ _0451_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1423_ _0452_ _0817_ _0503_ _0818_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_46_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1317__B1 _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output17_I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1070_ _0470_ _0478_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_55_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1972_ _0089_ clknet_4_11_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[77\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1337_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[96\] _0590_ _0739_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1406_ net41 _0544_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1268_ _0449_ _0499_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1199_ _0597_ _0599_ _0600_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1250__A2 _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1122_ _0524_ _0525_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[4\]
+ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_20_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1053_ _0376_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1886_ _0003_ clknet_4_2_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1955_ _0072_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[60\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1671_ _0219_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1740_ _0259_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtop_vga_spi_rom_28 uio_oe[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_7_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1333__C _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1105_ net4 _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1036_ _0358_ _0444_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1938_ _0055_ clknet_4_6_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[43\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1869_ _0334_ _0335_ _0336_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_39_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1723_ _0895_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1199__A1 _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1654_ _0210_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1585_ _0169_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1344__B _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1371__A1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[64\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1019_ _0388_ _0427_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_4_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1370_ _0682_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[66\] _0771_ _0624_
+ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_26_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1637_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[53\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[52\]
+ _0196_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1706_ _0239_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1568_ _0923_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_1_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1499_ _0513_ _0812_ _0877_ _0884_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_36_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1422_ net2 _0395_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1901__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1978__CLKN clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1284_ _0631_ _0685_ _0583_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1353_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[88\] _0755_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1916__CLKN clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0999_ _0346_ _0347_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1317__B2 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[121\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1317__A1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[120\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1886__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1308__A1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2041__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2016__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1971_ _0088_ clknet_4_11_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[76\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_11_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1405_ _0795_ _0560_ _0490_ _0541_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1267_ _0662_ _0668_ _0604_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1336_ _0659_ _0561_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[97\] _0738_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1198_ _0404_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput1 rst net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_4_9_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1121_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[5\] _0525_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1052_ _0459_ _0443_ _0460_ _0454_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_31_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1954_ _0071_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[59\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_3_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1885_ _0002_ clknet_4_2_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1861__I _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1319_ _0637_ _0713_ _0720_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_19_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1231__I0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[57\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[67\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[66\]
+ _0213_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0973__A2 _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtop_vga_spi_rom_29 uio_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1681__I _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1035_ _0404_ _0443_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1104_ _0506_ _0387_ _0392_ _0510_ net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1937_ _0054_ clknet_4_3_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[42\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_16_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1799_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[122\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[121\]
+ _0292_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1868_ _0410_ _0371_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1295__I3 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[128\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1766__I _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1507__I1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1584_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[31\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[30\]
+ _0934_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1722_ _0904_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1653_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[59\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[58\]
+ _0208_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1371__A2 _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1018_ _0361_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1362__A2 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[83\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_31_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1705_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[82\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[81\]
+ _0236_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1664__I0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[64\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1567_ _0928_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1636_ _0199_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1498_ _0530_ _0826_ _0538_ _0883_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_24_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1265__B _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1271__A1 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1646__I0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[57\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1326__A2 _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1421_ _0398_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1283_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[25\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[24\]
+ _0632_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1352_ _0566_ _0752_ _0753_ _0495_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_46_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1262__A1 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0998_ _0402_ _0406_ _0383_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1619_ _0190_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1317__A2 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_5_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1244__A1 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1970_ _0087_ clknet_4_9_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[75\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_15_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1335_ _0592_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[98\] _0736_ _0657_
+ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1404_ _0804_ net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1197_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[33\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[32\]
+ _0598_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1266_ _0664_ _0667_ _0602_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 net46 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1262__C _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1900__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1915__CLKN clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1051_ _0408_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1120_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[6\] _0524_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_31_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1884_ _0001_ clknet_4_2_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1953_ _0070_ clknet_4_9_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[58\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_43_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1318_ _0715_ _0716_ _0718_ _0719_ _0635_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_54_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1249_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[8\] _0651_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2015__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2031__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1034_ _0355_ _0356_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__1438__A1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1103_ _0400_ _0509_ _0399_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1936_ _0053_ clknet_4_6_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[41\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1297__S0 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1867_ _0332_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1798_ _0286_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_4_13_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1668__A1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[66\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1223__S _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1178__B _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1721_ _0755_ _0186_ _0247_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1583_ _0168_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1652_ _0209_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_53_Left_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1831__A1 _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1867__I _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1682__I1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[71\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1017_ _0362_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1919_ _0036_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_8_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1270__C _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1017__I _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1704_ _0238_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1566_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[23\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[22\]
+ _0924_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1635_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[52\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[51\]
+ _0196_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1497_ _0532_ _0879_ _0873_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_55_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1371__B _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1271__A2 _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1023__A2 _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1351_ _0568_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[91\] _0753_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1420_ _0584_ _0535_ _0420_ _0394_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA_clkbuf_4_1_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1282_ _0682_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[26\] _0683_ _0624_
+ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_46_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1366__B _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1618_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[44\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[43\]
+ _0189_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0997_ _0352_ _0405_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1573__I0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1549_ _0895_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_5_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1120__I tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1334_ _0493_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[99\] _0736_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1265_ _0665_ _0666_ _0600_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1180__A1 _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1403_ _0803_ tt_um_algofoogle_vga_spi_rom.r_rgb\[3\] _0553_ _0804_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1196_ _0427_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 ui_in[1] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1794__I0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[120\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1171__A1 _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0954__I _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1050_ _0354_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1952_ _0069_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[57\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_43_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1883_ _0000_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.r_vsync vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1363__C _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1248_ _0642_ _0647_ _0649_ _0570_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1317_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[120\] _0674_ _0574_
+ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[121\] _0707_ _0719_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_54_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1179_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[41\] _0574_ _0578_ _0580_
+ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_2_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1102_ _0508_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_51_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1033_ _0357_ _0441_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_17_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1935_ _0052_ clknet_4_6_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[40\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1358__C _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1961__CLKN clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1797_ _0291_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1297__S1 _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1866_ _0410_ _0371_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1914__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1929__CLKN clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1303__I _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1720_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[89\] _0187_ _0247_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_13_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1651_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[58\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[57\]
+ _0208_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1582_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[30\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[29\]
+ _0934_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1356__A1 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I ui_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1016_ _0424_ _0366_ _0349_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2014__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1918_ _0035_ clknet_4_13_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1849_ _0327_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2029__CLKN clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1889__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1338__A1 _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2044__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1634_ _0198_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1703_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[81\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[80\]
+ _0236_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1565_ _0927_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1496_ _0875_ _0881_ _0514_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_18_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2048_ _0165_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1281_ _0563_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[27\] _0683_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1350_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[90\] _0752_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0996_ _0404_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1617_ _0175_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1548_ _0643_ _0909_ _0917_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1479_ _0840_ _0867_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_37_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1402_ _0794_ _0802_ _0798_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1264_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[1\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[0\]
+ _0641_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1333_ _0724_ _0728_ _0731_ _0734_ _0712_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
Xinput4 ui_in[2] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1195_ _0414_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0979_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[2\] _0388_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1171__A2 _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0970__I _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1131__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1951_ _0068_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[56\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_22_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1882_ _0335_ _0344_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1247_ _0648_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[11\] _0649_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1178_ _0579_ _0441_ _0451_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1316_ _0659_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[122\] _0717_
+ _0705_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_54_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1392__A2 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1032_ _0355_ _0356_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_17_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1101_ _0449_ _0507_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1934_ _0051_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[39\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1865_ _0471_ _0333_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1796_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[121\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[120\]
+ _0287_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1581_ _0167_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_13_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1650_ _0207_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1194__C _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1015_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[4\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[5\]
+ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1917_ _0034_ clknet_4_13_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_48_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1831__A3 _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1385__B _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1848_ _0326_ tt_um_algofoogle_vga_spi_rom.hsync _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1779_ _0261_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold15_I uio_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1274__A1 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1026__A1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1564_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[22\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[21\]
+ _0924_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1633_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[51\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[50\]
+ _0196_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1702_ _0237_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1913__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1495_ _0825_ _0795_ _0880_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1928__CLKN clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1265__A1 _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2047_ _0164_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1812__I0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[128\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1256__A1 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1280_ _0379_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2013__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2028__CLKN clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0995_ _0403_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[15\] _0910_ _0917_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1219__I _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1616_ _0575_ _0186_ _0188_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1478_ _0828_ _0856_ _0838_ _0866_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2034__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1401_ _0491_ _0801_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1194_ _0585_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[34\] _0595_ _0588_
+ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1263_ _0495_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1332_ _0732_ _0726_ _0733_ _0707_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xinput5 ui_in[5] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0978_ _0384_ _0385_ _0386_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_52_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1950_ _0067_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[55\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1870__A1 _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1881_ _0503_ _0343_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_22_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1315_ _0703_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[123\] _0717_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1177_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[40\] _0579_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1246_ _0562_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1100_ _0482_ _0353_ _0410_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1031_ _0368_ _0373_ _0439_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1933_ _0050_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[38\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1843__A1 _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1864_ _0472_ _0333_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1227__I _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1795_ _0290_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1229_ _0414_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1580_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[29\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[28\]
+ _0934_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1047__I _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1014_ _0401_ _0422_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1916_ _0033_ clknet_4_12_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_29_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1847_ _0858_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1778_ _0280_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_40_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1035__A2 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1701_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[80\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[79\]
+ _0236_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1026__A2 _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1563_ _0926_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1632_ _0197_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1494_ _0848_ _0555_ _0841_ _0879_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__1240__I _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2046_ _0163_ clknet_4_9_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1192__A1 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0994_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[2\] _0403_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1546_ _0643_ _0905_ _0916_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1615_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[43\] _0187_ _0188_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1477_ _0864_ _0865_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_37_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2029_ _0146_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[134\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_17_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1346__S _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1989__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1912__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1927__CLKN clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1331_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[108\] _0460_ _0733_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1400_ _0795_ _0550_ net9 _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1193_ _0586_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[35\] _0595_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1262_ _0655_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[2\] _0663_ _0588_
+ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_36_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 ui_in[6] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0977_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[6\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[7\]
+ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_14_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1529_ _0889_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2012__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2027__CLKN clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ _0317_ _0341_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1138__A1 _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1314_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[124\] _0610_ _0573_
+ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[125\] _0459_ _0716_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1245_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[10\] _0647_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1176_ _0566_ _0575_ _0577_ _0570_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_42_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2047__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1030_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[5\] _0362_ _0438_
+ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1932_ _0049_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[37\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1863_ _0442_ _0333_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1794_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[120\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[119\]
+ _0287_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1228_ _0620_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[58\] _0628_ _0629_
+ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_59_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1159_ _0495_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1264__S _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1013_ _0407_ _0412_ _0419_ _0421_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1915_ _0032_ clknet_4_13_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_29_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1777_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[113\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[112\]
+ _0274_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1846_ _0325_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__1812__S _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1631_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[50\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[49\]
+ _0196_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1700_ _0230_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1562_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[21\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[20\]
+ _0924_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1493_ _0533_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_49_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I ui_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2045_ _0162_ clknet_4_9_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1829_ _0696_ _0817_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_23_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0993_ _0365_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1614_ _0890_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1545_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[13\] _0907_ _0916_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1476_ _0524_ _0829_ _0854_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_37_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2028_ _0145_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[133\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_17_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1261_ _0586_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[3\] _0663_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_31_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1330_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[109\] _0732_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1192_ _0584_ _0589_ _0591_ _0593_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_36_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 ui_in[7] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0976_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.quad tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[2\]
+ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1528_ _0904_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1459_ _0826_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1138__A2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1244_ _0496_ _0640_ _0645_ _0497_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_2_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1313_ _0364_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[126\] _0714_
+ _0705_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1175_ _0576_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[43\] _0577_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1973__CLKN clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0959_ _0350_ _0365_ _0366_ _0367_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_6_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1911__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1926__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1065__A1 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1679__I0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[71\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1931_ _0048_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[36\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1359__A2 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1862_ _0494_ _0333_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1793_ _0289_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput10 net16 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1158_ _0353_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1227_ _0455_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2011__CLKN clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1089_ _0415_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2026__CLKN clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1012_ _0420_ _0387_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1914_ _0031_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1776_ _0279_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1845_ _0315_ tt_um_algofoogle_vga_spi_rom.hsync _0324_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_4_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1203__B _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2037__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1164__I _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1630_ _0175_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_38_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1561_ _0925_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1492_ _0876_ _0877_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_49_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2044_ _0161_ clknet_4_9_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1422__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1759_ _0270_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1828_ _0308_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_15_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold13_I uio_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0992_ _0383_ _0393_ _0399_ _0400_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1544_ _0915_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1613_ _0891_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1475_ _0828_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_37_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2027_ _0144_ clknet_4_9_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[132\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_45_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1260_ _0584_ _0658_ _0660_ _0661_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1191_ _0592_ _0561_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[37\] _0593_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_36_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 net40 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1892__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0975_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[8\] _0384_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_6_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1527__I _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1527_ _0894_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1458_ _0814_ _0850_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1389_ _0517_ _0557_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1437__I tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1855__A1 _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1243_ _0642_ _0643_ _0644_ _0570_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1174_ _0562_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1082__I _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1312_ _0566_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[127\] _0714_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_59_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1074__A2 _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1031__B _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0958_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[0\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[1\]
+ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[2\] _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_6_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1930_ _0047_ clknet_4_12_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[35\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XPHY_EDGE_ROW_26_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 net44 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1792_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[119\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[118\]
+ _0287_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1861_ _0332_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1157_ _0518_ _0558_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1226_ _0621_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[59\] _0628_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_59_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1088_ _0495_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1210__A2 _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1972__CLKN clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1011_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[9\] _0420_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1913_ _0030_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_29_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1029__A2 _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1925__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1910__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1775_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[112\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[111\]
+ _0274_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1844_ _0514_ _0320_ _0323_ _0812_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_8_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1209_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[48\] _0610_ _0611_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1259__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1560_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[20\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[19\]
+ _0924_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2025__CLKN clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2010__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1491_ _0530_ _0826_ _0538_ _0835_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_55_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1090__I _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2043_ _0160_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[135\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[134\]
+ _0906_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1758_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[104\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[103\]
+ _0267_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1689_ _0229_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_13_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1110__A1 _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0991_ _0389_ _0385_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1543_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[13\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[12\]
+ _0901_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1085__I _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1612_ _0575_ _0183_ _0185_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1474_ _0814_ _0863_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2026_ _0143_ clknet_4_9_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[131\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_9_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1190_ _0363_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput9 net47 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_52_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0974_ _0366_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1526_ _0903_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1457_ _0848_ _0846_ _0849_ _0838_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1388_ _0758_ _0769_ _0670_ _0789_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1864__A2 _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1313__A1 _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2009_ _0126_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[114\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1304__A1 _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_36_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1311_ _0706_ _0708_ _0710_ _0711_ _0712_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_EDGE_ROW_56_Left_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1242_ _0576_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[15\] _0644_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1173_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[42\] _0575_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0957_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[5\] _0366_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1509_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[1\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[0\]
+ _0891_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_53_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1384__S _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_1_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1860_ _0858_ _0856_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1791_ _0288_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1087_ _0413_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1225_ _0624_ _0625_ _0626_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1156_ _0397_ _0557_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1989_ _0106_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[94\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_30_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1010_ _0416_ _0418_ _0376_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1912_ _0029_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1843_ _0514_ _0444_ _0313_ _0322_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1774_ _0278_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1816__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1208_ _0409_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1139_ _0491_ _0541_ _0542_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1490_ _0874_ _0875_ _0857_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2042_ _0159_ clknet_4_11_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_index\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold1 uio_in[6] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_49_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ _0307_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1757_ _0269_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1688_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[75\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[74\]
+ _0225_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1971__CLKN clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1405__B _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1924__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__CLKN clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1611_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[41\] _0184_ _0185_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0990_ _0385_ _0394_ _0396_ _0398_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_14_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1542_ _0914_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1473_ _0524_ _0855_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_49_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2025_ _0142_ clknet_4_8_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[130\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_49_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1809_ _0298_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1225__B _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1331__A2 _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__CLKN clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1186__I _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0973_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[9\] _0364_ _0375_
+ _0381_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1525_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[7\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[6\]
+ _0901_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1387_ _0774_ _0779_ _0788_ _0604_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1456_ _0848_ _0844_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1077__A1 _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2008_ _0125_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[113\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_45_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1845__S _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1241_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[14\] _0643_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1310_ _0480_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1172_ _0573_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0956_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[4\] _0365_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1508_ _0892_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1298__A1 _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1439_ _0833_ _0531_ _0834_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1790_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[118\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[117\]
+ _0287_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_4_8_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1224_ _0354_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1086_ _0493_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1155_ _0372_ _0499_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0939_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[2\] _0348_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1988_ _0105_ clknet_4_3_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[93\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_15_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_38_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1911_ _0028_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_29_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1773_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[111\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[110\]
+ _0274_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1842_ _0321_ _0394_ _0411_ _0309_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_12_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1207_ _0484_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[50\] _0607_ _0608_
+ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1069_ _0472_ _0473_ _0475_ _0476_ _0477_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1138_ _0378_ net14 _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2041_ _0158_ clknet_4_11_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold2 net10 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_57_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1756_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[103\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[102\]
+ _0267_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1825_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[134\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[133\]
+ _0906_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1687_ _0228_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1610_ _0906_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1541_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[12\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[11\]
+ _0901_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1472_ _0862_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2024_ _0141_ clknet_4_8_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[129\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1651__I1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[57\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1739_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[96\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[95\]
+ _0254_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1808_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[126\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[125\]
+ _0297_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_42_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0972_ _0378_ _0380_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1524_ _0902_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1386_ _0781_ _0783_ _0785_ _0787_ _0353_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1455_ _0833_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2007_ _0124_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[112\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1970__CLKN clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1923__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1236__B _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1938__CLKN clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1240_ _0641_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_4_4_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1171_ _0492_ _0455_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_2_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0955_ _0363_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_6_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1507_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[0\] net9 _0891_ _0892_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2023__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1369_ _0563_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[67\] _0771_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1438_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[1\] _0533_ _0834_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0972__A1 _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1223_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[63\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[62\]
+ _0565_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1154_ _0395_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1085_ _0492_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0938_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[1\] _0347_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1987_ _0104_ clknet_4_4_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[92\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_30_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1140__A1 _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1910_ _0027_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1772_ _0732_ _0251_ _0277_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1841_ _0312_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1318__C _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1206_ _0456_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1137_ _0513_ _0520_ _0529_ _0530_ _0540_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_18_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1068_ _0474_ _0425_ _0436_ _0472_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_50_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_12_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1228__C _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1361__A1 _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1352__A1 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2040_ _0157_ clknet_4_11_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold3 _0545_ net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1755_ _0268_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1329__B _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1824_ _0306_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1686_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[74\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[73\]
+ _0225_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1753__I _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1540_ _0647_ _0909_ _0913_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1471_ _0855_ _0861_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2023_ _0140_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[128\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1807_ _0286_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_17_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_20_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1738_ _0258_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1669_ _0770_ _0186_ _0218_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1316__A1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1885__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0971_ _0379_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_0_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1523_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[6\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[5\]
+ _0901_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1326__C _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1454_ _0814_ _0847_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1342__B _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1385_ _0624_ _0786_ _0451_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2040__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2006_ _0123_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[111\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1236__C _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1560__I1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1170_ _0561_ _0564_ _0571_ _0481_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_42_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0954_ _0362_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1506_ _0890_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1437_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[3\] _0833_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_43_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1368_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[65\] _0770_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1299_ _0696_ _0500_ _0698_ _0700_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XPHY_EDGE_ROW_52_Left_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0972__A2 _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1222_ _0455_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1084_ _0346_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1153_ _0522_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_50_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1922__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1986_ _0103_ clknet_4_3_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[91\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_0937_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[0\] _0346_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1067__B _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2022__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1840_ _0319_ _0311_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_52_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1771_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[110\] _0252_ _0277_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1370__A2 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[66\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1205_ _0576_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[51\] _0607_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1136_ _0531_ _0532_ _0534_ _0535_ _0539_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_1067_ _0369_ _0374_ _0439_ _0442_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_47_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1189__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ _0086_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[74\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1244__C _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold4 _0154_ net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_17_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1823_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[133\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[132\]
+ _0302_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1754_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[102\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[101\]
+ _0267_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1345__B _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1685_ _0227_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1119_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[3\] _0522_ _0523_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1098__A1 _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1270__A1 _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1470_ _0859_ _0860_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1325__A2 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2022_ _0139_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[127\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_9_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1261__A1 _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1806_ _0296_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1599_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[37\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[36\]
+ _0176_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1737_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[95\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[94\]
+ _0254_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1668_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[66\] _0187_ _0218_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1252__A1 _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_34_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1243__A1 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0970_ _0362_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1522_ _0895_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1453_ _0531_ _0843_ _0846_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1384_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[79\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[78\]
+ _0565_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2005_ _0122_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[110\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0953_ _0361_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1367_ _0763_ _0768_ _0637_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1505_ _0889_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1436_ _0462_ _0521_ _0525_ _0535_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_1298_ _0498_ _0699_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1221_ _0620_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[60\] _0622_ _0485_
+ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_20_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1083_ _0491_ net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1152_ _0554_ net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1985_ _0102_ clknet_4_3_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[90\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_0936_ _0345_ net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1419_ _0534_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1770_ _0732_ _0248_ _0276_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1204_ _0372_ _0499_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1066_ _0474_ _0425_ _0429_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1135_ _0537_ _0538_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1899_ _0016_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_47_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1968_ _0085_ clknet_4_10_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[73\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_3_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1921__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold5 uio_in[1] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1936__CLKN clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1170__C _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1753_ _0261_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1822_ _0305_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1684_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[73\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[72\]
+ _0225_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1049_ _0377_ _0357_ _0454_ _0457_ _0402_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1118_ _0388_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2021__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2021_ _0138_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[126\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_57_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1736_ _0749_ _0251_ _0257_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1805_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[125\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[124\]
+ _0292_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1598_ _0177_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1667_ _0770_ _0183_ _0217_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1266__B _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1521_ _0900_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1383_ _0620_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[76\] _0784_ _0485_
+ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1452_ _0824_ _0845_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2004_ _0121_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[109\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_45_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1414__1_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1719_ _0755_ _0183_ _0246_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1170__A1 _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0952_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[0\] _0361_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1504_ _0482_ _0522_ _0520_ _0888_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1366_ _0765_ _0767_ _0602_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1435_ _0532_ _0534_ _0523_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1297_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[135\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[134\]
+ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[133\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[132\]
+ _0642_ _0665_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__1595__I _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_41_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1382__A1 _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1220_ _0621_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[61\] _0622_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1151_ _0552_ tt_um_algofoogle_vga_spi_rom.r_rgb\[5\] _0553_ _0554_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1082_ _0490_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1984_ _0101_ clknet_4_3_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[89\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_23_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0935_ net6 net5 net7 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_15_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1373__A1 _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1349_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[92\] _0610_ _0748_ _0657_
+ _0750_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1418_ _0814_ _0515_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1125__A1 _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1203_ _0594_ _0603_ _0604_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1134_ _0482_ _0521_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[6\]
+ _0525_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_34_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1065_ _0443_ _0408_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1898_ _0015_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_28_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1967_ _0084_ clknet_4_9_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[72\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_59_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold6 net8 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1888__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1752_ _0266_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1821_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[132\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[131\]
+ _0302_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1683_ _0226_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1328__A1 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2043__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1117_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[7\] _0521_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1048_ _0456_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1319__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1108__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ _0137_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[125\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_15_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1666_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[64\] _0184_ _0217_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1735_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[94\] _0252_ _0257_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1804_ _0295_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1597_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[36\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[35\]
+ _0176_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1982__CLKN clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1920__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1935__CLKN clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1301__I _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1520_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[5\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[4\]
+ _0896_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1382_ _0641_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[77\] _0784_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1451_ _0837_ _0844_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2003_ _0120_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[108\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_26_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1367__B _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2020__CLKN clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1718_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[87\] _0184_ _0246_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1649_ _0206_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_56_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0951_ _0349_ _0359_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1503_ _0449_ _0394_ _0464_ _0391_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__1206__I _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1365_ _0616_ _0766_ _0600_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1296_ _0584_ _0697_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1434_ _0548_ _0828_ _0829_ _0535_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1150_ net4 _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1081_ _0448_ _0469_ _0489_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1983_ _0100_ clknet_4_3_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[88\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_48_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1373__A2 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[71\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1417_ _0813_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1279_ _0678_ _0680_ _0466_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1348_ _0703_ _0629_ _0749_ _0405_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_6_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1052__A1 _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1355__A2 _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1202_ _0454_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1133_ _0397_ _0536_ _0464_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1064_ _0368_ _0374_ _0433_ _0442_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1966_ _0083_ clknet_4_14_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[71\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_34_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1897_ _0014_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1337__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold7 _0806_ net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ _0304_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1751_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[101\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[100\]
+ _0262_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1682_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[72\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[71\]
+ _0225_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1047_ _0455_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1116_ _0420_ _0519_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1949_ _0066_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[54\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_16_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1803_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[124\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[123\]
+ _0292_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1596_ _0175_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1665_ _0216_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1734_ _0749_ _0248_ _0256_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1789__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2033__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1450_ _0531_ _0841_ _0534_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1381_ _0631_ _0782_ _0583_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2002_ _0119_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[107\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_26_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1579_ _0166_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1717_ _0245_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1648_ _0889_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1981__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1187__C _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0950_ _0353_ _0358_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1502_ _0887_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1433_ _0525_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1364_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[81\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[80\]
+ _0598_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1295_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[131\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[130\]
+ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[129\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[128\]
+ _0642_ _0665_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_58_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1934__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1222__I _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1949__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1851__A1 _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1288__B _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1080_ _0382_ _0471_ _0479_ _0488_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__1134__A3 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1982_ _0099_ clknet_4_6_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[87\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_30_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1347_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[93\] _0749_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1416_ _0812_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1278_ _0588_ _0679_ _0459_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1833__A1 _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1290__C _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1238__S _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1052__A2 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1201_ _0596_ _0601_ _0602_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1063_ _0403_ _0408_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_25_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1132_ _0391_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1965_ _0082_ clknet_4_14_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[70\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1896_ _0013_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_11_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1282__A2 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold8 _0150_ net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1273__A2 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1750_ _0265_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _0207_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_20_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1230__I _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1046_ _0356_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_0_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1115_ _0391_ _0518_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1948_ _0065_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[53\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1879_ _0317_ _0341_ _0342_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1341__S _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_57_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1733_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[92\] _0249_ _0256_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1802_ _0294_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1595_ _0894_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1664_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[64\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[63\]
+ _0213_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1029_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[4\] _0431_ _0438_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1796__I0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[121\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1380_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[73\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[72\]
+ _0565_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2001_ _0118_ clknet_4_1_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[106\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_42_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1716_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[87\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[86\]
+ _0241_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1578_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[28\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[27\]
+ _0934_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1647_ _0205_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1383__C _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1363_ _0380_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[82\] _0764_ _0457_
+ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1501_ _0878_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.vsync _0886_ _0887_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1137__A1 _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1432_ _0521_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_53_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1294_ _0395_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1119__A1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1981_ _0098_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[86\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_48_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1346_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[95\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[94\]
+ _0563_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1415_ net1 _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1414__1 clknet_4_8_0_clk net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2046__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1277_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[23\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[22\]
+ _0598_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1980__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1995__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1052__A3 _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1933__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1200_ _0480_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_0_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1948__CLKN clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1062_ _0470_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1131_ net2 _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1895_ _0012_ clknet_4_4_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1964_ _0081_ clknet_4_14_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[69\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1329_ _0729_ _0730_ _0496_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2059__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold9 net50 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_57_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1048__I _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1680_ _0224_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1114_ _0398_ _0517_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1045_ _0418_ _0453_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1947_ _0064_ clknet_4_13_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[52\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_31_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1386__C _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1878_ _0317_ _0341_ _0337_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1575__I1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1191__A2 _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1732_ _0255_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1663_ _0215_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1801_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[123\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[122\]
+ _0292_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1594_ _0174_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1028_ _0425_ _0436_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1796__I1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[120\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1844__C _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1416__I _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1400__A3 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2000_ _0117_ clknet_4_4_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[105\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_26_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1715_ _0244_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1646_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[57\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[56\]
+ _0201_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1577_ _0923_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_6_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1394__A2 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1810__S _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1500_ _0876_ _0882_ _0885_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1362_ _0648_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[83\] _0764_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_37_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1431_ _0524_ _0826_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1293_ _0397_ _0557_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1629_ _0195_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1980_ _0097_ clknet_4_7_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[85\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1276_ _0380_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[20\] _0677_ _0616_
+ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1345_ _0735_ _0746_ _0606_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1349__A2 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1760__A2 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1130_ _0533_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1276__A1 _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1061_ _0417_ _0367_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1963_ _0080_ clknet_4_14_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[68\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_7_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1894_ _0011_ clknet_4_0_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.vsync
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_11_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1259_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[4\] _0590_ _0661_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1328_ _0655_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[111\] _0730_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1258__A1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2036__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1733__A2 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1113_ _0366_ _0389_ _0453_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1044_ _0351_ _0370_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1946_ _0063_ clknet_4_13_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[51\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_43_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1877_ _0817_ _0339_ _0341_ _0335_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_16_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1994__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1724__A2 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1932__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1947__CLKN clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1800_ _0293_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1731_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[92\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[91\]
+ _0254_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1662_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[63\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[62\]
+ _0213_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1593_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[35\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[34\]
+ _0170_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1027_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[7\] _0426_ _0435_
+ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1929_ _0046_ clknet_4_13_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[34\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Left_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1808__S _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1714_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[86\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[85\]
+ _0241_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1576_ _0933_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1645_ _0204_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1201__B _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2059_ net3 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1891__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1430_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[4\] _0826_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1361_ _0707_ _0760_ _0761_ _0762_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1292_ _0559_ _0639_ _0693_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_53_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1559_ _0923_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1628_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[49\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[48\]
+ _0189_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1413_ _0811_ net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1275_ _0648_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[21\] _0677_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1344_ _0740_ _0745_ _0604_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1530__I _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_4_7_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1060_ _0402_ _0450_ _0463_ _0468_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1962_ _0079_ clknet_4_14_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[67\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_34_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ _0010_ clknet_4_3_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1189_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[36\] _0590_ _0591_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1258_ _0659_ _0561_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[5\] _0660_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1327_ _0494_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[110\] _0729_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1814__I1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[128\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1019__A2 _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0950__A1 _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1258__A2 _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1043_ _0451_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1112_ _0511_ _0515_ _0516_ net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1945_ _0062_ clknet_4_12_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[50\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_0_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1185__A1 _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1255__I _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1876_ _0369_ _0386_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_39_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1176__A1 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1592_ _0173_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1730_ _0230_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1167__A1 _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1661_ _0214_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input7_I ui_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1026_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[6\] _0427_ _0435_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1928_ _0045_ clknet_4_13_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[33\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1859_ _0331_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_15_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1321__A1 _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1713_ _0243_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1993__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1931__CLKN clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1575_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[27\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[26\]
+ _0929_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1644_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[56\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[55\]
+ _0201_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1946__CLKN clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1863__A2 _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1312__A1 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1009_ _0417_ _0365_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1360_ _0592_ _0665_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[85\] _0762_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_2_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1291_ _0654_ _0669_ _0670_ _0692_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_37_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1558_ _0894_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1627_ _0194_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1489_ _0828_ _0526_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1049__B1 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_3_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1343_ _0742_ _0744_ _0602_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1412_ _0810_ tt_um_algofoogle_vga_spi_rom.r_rgb\[1\] net4 _0811_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1274_ _0497_ _0672_ _0673_ _0675_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_13_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0989_ _0397_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_52_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1961_ _0078_ clknet_4_12_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[66\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_28_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1892_ _0009_ clknet_4_2_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.quad vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_7_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1326_ _0725_ _0726_ _0727_ _0452_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1188_ _0409_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1257_ _0363_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1827__S _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1042_ _0354_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1111_ _0511_ tt_um_algofoogle_vga_spi_rom.r_vsync _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1944_ _0061_ clknet_4_12_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[49\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_31_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1875_ _0340_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_39_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1309_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[116\] _0610_ _0573_
+ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[117\] _0481_ _0711_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_19_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_11_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1799__I1 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[121\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1100__A2 _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1591_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[34\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[33\]
+ _0170_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[62\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[61\]
+ _0213_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1025_ _0368_ _0374_ _0433_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1927_ _0044_ clknet_4_13_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[32\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1858_ _0858_ _0552_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1789_ _0286_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_30_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1712_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[85\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[84\]
+ _0241_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1643_ _0203_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1574_ _0932_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1008_ _0350_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1290_ _0676_ _0681_ _0691_ _0637_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_41_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1626_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[48\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[47\]
+ _0189_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1557_ _0922_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1488_ _0825_ _0548_ _0834_ _0873_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_52_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1836__A3 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1930__CLKN clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2039__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1945__CLKN clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1212__A1 _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1273_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[16\] _0674_ _0675_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1342_ _0657_ _0743_ _0481_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1411_ _0549_ _0809_ _0805_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0988_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[7\] _0397_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1609_ _0904_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2030__CLKN clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1184__I _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1960_ _0077_ clknet_4_3_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[65\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1891_ _0008_ clknet_4_8_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1899__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1256_ _0655_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[6\] _0656_ _0657_
+ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1325_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[104\] _0674_ _0727_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1187_ _0585_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[38\] _0587_ _0588_
+ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_24_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1424__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1110_ _0514_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.vsync _0515_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1041_ _0449_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1943_ _0060_ clknet_4_12_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[48\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_24_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1874_ _0337_ _0338_ _0339_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_51_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1239_ _0562_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1308_ _0659_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[118\] _0709_
+ _0705_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_47_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1894__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1590_ _0172_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1024_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[1\] _0426_ _0432_
+ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_44_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1926_ _0043_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1788_ _0206_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1857_ _0813_ _0543_ net38 _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_39_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1857__A1 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Left_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1711_ _0242_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1642_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[55\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[54\]
+ _0201_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_5_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1573_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[26\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[25\]
+ _0929_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1848__A1 _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1007_ _0414_ _0415_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1909_ _0026_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_36_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1650__I _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1556_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[19\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[18\]
+ _0918_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1625_ _0567_ _0186_ _0193_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1487_ _0833_ _0555_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_52_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2039_ _0156_ clknet_4_12_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1460__A2 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1410_ net41 _0550_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1341_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[103\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[102\]
+ _0641_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1272_ _0409_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0987_ _0395_ _0385_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1539_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[11\] _0910_ _0913_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1608_ _0579_ _0909_ _0182_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1890_ _0007_ clknet_4_2_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1186_ _0456_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1255_ _0456_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1324_ _0682_ _0631_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_46_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1944__CLKN clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1959__CLKN clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output14_I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1351__A1 _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1040_ _0383_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1942_ _0059_ clknet_4_6_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[47\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_28_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1873_ _0450_ _0696_ _0334_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1238_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[13\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[12\]
+ _0568_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1169_ _0566_ _0567_ _0569_ _0570_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1307_ _0703_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[119\] _0709_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_51_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1898__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1023_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[0\] _0431_ _0432_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1925_ _0042_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_44_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1856_ _0330_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1787_ _0285_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1572_ _0931_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1710_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[84\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[83\]
+ _0241_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1641_ _0202_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input5_I ui_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1884__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1006_ _0348_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1908_ _0025_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__1558__I _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1839_ _0312_ _0316_ _0318_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_4_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1555_ _0921_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1624_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[47\] _0187_ _0193_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1486_ _0859_ _0872_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2038_ _0155_ clknet_4_2_0_clk tt_um_algofoogle_vga_spi_rom.r_rgb\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__1237__B _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1340_ _0592_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[100\] _0741_
+ _0597_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1271_ _0655_ _0597_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[17\] _0673_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0986_ _0389_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1538_ _0647_ _0905_ _0912_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1607_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[41\] _0910_ _0182_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1469_ _0824_ _0854_ _0829_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1323_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[105\] _0725_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1185_ _0586_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[39\] _0587_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1254_ _0493_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[7\] _0656_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_46_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1424__A3 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0969_ _0377_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1360__A2 _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1234__C _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1250__B _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1179__A2 _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1941_ _0058_ clknet_4_3_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[46\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_28_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1872_ _0556_ _0369_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1306_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[112\] _0460_ _0573_
+ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[113\] _0707_ _0708_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1237_ _0582_ _0605_ _0606_ _0638_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1168_ _0413_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1099_ _0420_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_34_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1022_ _0361_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1924_ _0041_ clknet_4_15_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_44_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1260__A1 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1855_ _0326_ _0803_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1943__CLKN clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1786_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[117\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[116\]
+ _0281_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1958__CLKN clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1306__A2 _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1242__A1 _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1571_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[25\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[24\]
+ _0929_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1640_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[54\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[53\]
+ _0201_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1332__C _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1005_ _0413_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1907_ _0024_ clknet_4_5_0_clk tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1838_ _0712_ _0498_ _0317_ _0506_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__1897__CLKN clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1769_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[108\] _0249_ _0276_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_hold14_I ui_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1659__I _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1554_ tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[18\] tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[17\]
+ _0918_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1623_ _0567_ _0183_ _0192_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1485_ _0825_ _0871_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
.ends

