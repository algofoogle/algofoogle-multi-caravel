// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * Our main top design macro (top_raybox_zero_fsm) is
 * instantiated in this UPW.
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper (
`ifdef USE_POWER_PINS
    inout vdd,      // User area 5.0V supply
    inout vss,      // User area ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [63:0] la_data_in,
    output [63:0] la_data_out,
    input  [63:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

/*--------------------------------------*/
/* User project is instantiated  here   */
/*--------------------------------------*/

    //// BEGIN: INSTANTIATION OF ANTON'S DESIGN (top_raybox_zero_fsm) (GFMPW1_SNIPPET_top_raybox_zero_fsm) ---------------------

    // This snippet comes from here:
    // https://github.com/algofoogle/raybox-zero/blob/gf180/src/rtl/gfmpw1_snippets/GFMPW1_SNIPPET_top_raybox_zero_fsm.v

    wire rbz_fsm_clock_in = wb_clk_i;
    wire rbz_fsm_reset = wb_rst_i;
    wire rbz_fsm_reset_alt = rbz_fsm_la_in[0]; // Reset by SoC reset OR LA.
    wire [12:0] rbz_fsm_la_in = la_data_in[12:0]; // Can be reassigned, if desired.
    wire [15:0] a0s, a1s;                   // Low and high signals from our design that we can use to mix constants.
    assign io_out[34:19] = a0s[15:0]; // Irrelevant.
    assign io_out[7:0] = a0s[15:8];  // Irrelevant.

    wire rbz_fsm_tex_oeb0;
    assign io_oeb = {
        a0s[15:13],         // 37:35 are OUT
        a1s[15:0],          // 34:19 are IN
        rbz_fsm_tex_oeb0,   // 18 is bidir (tex_io0)
        a0s[12:3],          // 17:8 are OUT
        a1s[15:8],          // 7:0 are IN or not otherwise used (i.e. under SoC control).
    }; // 0001111111111111111*000000000011111111 where *=tex_io0 dir.

    top_raybox_zero_fsm top_raybox_zero_fsm(
    `ifdef USE_POWER_PINS
        .vdd(vdd),        // User area 1 1.8V power
        .vss(vss),        // User area 1 digital ground
    `endif

        .i_clk                  (rbz_fsm_clock_in),
        .i_reset                (rbz_fsm_reset),
        .i_reset_alt            (rbz_fsm_reset_alt),

        .zeros                  (a0s),  // A source of 16 constant '0' signals.
        .ones                   (a1s),  // A source of 16 constant '1' signals.

        .o_hsync                (io_out[8]),
        .o_vsync                (io_out[9]),
        .o_rgb                  (io_out[15:10]),

        .o_tex_csb              (io_out[16]),
        .o_tex_sclk             (io_out[17]),
        .o_tex_oeb0             (rbz_fsm_tex_oeb0), // My only bidirectional pad.
        .o_tex_out0             (io_out[18]),
        .i_tex_in               (io_in[21:18]),

        .i_vec_csb              (io_in[22]),
        .i_vec_sclk             (io_in[23]),
        .i_vec_mosi             (io_in[24]),

        .i_reg_csb              (io_in[25]),
        .i_reg_sclk             (io_in[26]),
        .i_reg_mosi             (io_in[27]),

        .i_debug_vec_overlay    (io_in[28]),
        .i_debug_map_overlay    (io_in[29]),
        .i_debug_trace_overlay  (io_in[30]),
        .i_reg_outs_enb         (io_in[31]),
        .i_mode                 (io_in[34:32]),

        .o_gpout                (io_out[37:35]),
        .i_gpout0_sel           (rbz_fsm_la_in[4:1]),
        .i_gpout1_sel           (rbz_fsm_la_in[8:5]),
        .i_gpout2_sel           (rbz_fsm_la_in[12:9])
    );

    //// END: INSTANTIATION OF ANTON'S DESIGN (top_raybox_zero_fsm) (GFMPW1_SNIPPET_top_raybox_zero_fsm) ---------------------

endmodule	// user_project_wrapper

`default_nettype wire
