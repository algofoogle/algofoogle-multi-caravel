* NGSPICE file created from urish_simon_says.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

.subckt urish_simon_says io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[2] io_oeb[30]
+ io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4]
+ io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[3] io_out[4] io_out[7] io_out[8] io_out[9] vdd vss wb_clk_i wb_rst_i
+ io_oeb[20] io_out[37] io_out[11] io_out[0] io_out[36] io_oeb[25] io_out[35] io_out[10]
+ io_oeb[24] io_out[34] io_out[33] io_oeb[23] io_oeb[22] io_out[32] io_out[31] io_oeb[21]
+ io_out[6] io_oeb[29] io_oeb[28] io_out[30] io_out[5] io_oeb[27] io_oeb[26] io_oeb[1]
+ io_oeb[11] io_oeb[35]
X_2037_ _0291_ _0294_ _0300_ _0301_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_2106_ _0351_ _0359_ _0365_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2182__A2 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1996__A2 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1920__A2 _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1606_ _0729_ _0745_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2724_ _0153_ clknet_4_8_0_wb_clk_i simon1.seq\[19\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2655_ _0084_ clknet_4_8_0_wb_clk_i simon1.play1.tick_counter\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1399_ _0836_ simon1.seq_length\[0\] _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2586_ _0032_ clknet_4_4_0_wb_clk_i simon1.seq\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1468_ _0889_ _0900_ _0904_ _0905_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1537_ _0004_ _0963_ _0974_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_22_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2672__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2440_ _0637_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1322_ _0748_ _0742_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2371_ simon1.tick_counter\[3\] simon1.tick_counter\[4\] _0588_ _0591_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_61_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2707_ _0136_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2638_ _0067_ clknet_4_14_0_wb_clk_i simon1.play1.tick_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2569_ _0015_ clknet_4_4_0_wb_clk_i simon1.seq\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2695__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1940_ _0211_ _0217_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1871_ _1243_ _1244_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2423_ _0622_ _0627_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2119__A2 _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2354_ _0577_ _0578_ _0579_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1305_ _0746_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2285_ _0991_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2357__B _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2710__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_21_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2070_ _0320_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1854_ _1223_ _1227_ _1228_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1785_ _1173_ _1174_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1923_ _0201_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2406_ simon1.tick_counter\[14\] _0613_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2199_ _0416_ _0984_ _0442_ _0419_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2268_ _0506_ _0507_ _0998_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2337_ _0566_ _0557_ _0522_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2733__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2028__A1 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xurish_simon_says_52 io_out[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_74 io_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_30 io_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_41 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_63 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_53_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1945__I _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _0999_ _1004_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2606__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2053_ simon1.play1.tick_counter\[16\] _0277_ _0292_ _0319_ _0320_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2756__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2122_ _0379_ _0374_ _0380_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_29_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1906_ _1221_ _1223_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1837_ _1212_ _1213_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1768_ _1161_ _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2430__A1 _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1699_ _1080_ simon1.seq\[16\]\[0\] _1113_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2629__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput20 net20 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput7 net7 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_46_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1622_ _0772_ _0777_ _1038_ _0783_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2671_ _0100_ clknet_4_13_0_wb_clk_i simon1.tone_sequence_counter\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2740_ _0169_ clknet_4_3_0_wb_clk_i simon1.seq\[24\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1553_ _0787_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1484_ _0004_ _0907_ _0921_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_37_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2036_ _1267_ _0300_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2105_ _0353_ _0359_ _0365_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_15_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2723_ _0152_ clknet_4_8_0_wb_clk_i simon1.seq\[19\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1605_ _1032_ _1036_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2654_ _0083_ clknet_4_10_0_wb_clk_i simon1.play1.tick_counter\[23\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2585_ _0031_ clknet_4_4_0_wb_clk_i simon1.seq\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1536_ _0886_ _0968_ _0973_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1398_ simon1.seq_counter\[0\] _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1467_ _0871_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2019_ _0279_ _0283_ _0289_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ _0585_ _0590_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1321_ _0747_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_59_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2706_ _0135_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2637_ _0066_ clknet_4_11_0_wb_clk_i simon1.play1.tick_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2568_ _0728_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2499_ _0670_ simon1.seq\[27\]\[0\] _0684_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1519_ _0889_ _0952_ _0956_ _0898_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_45_Left_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_54_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1870_ simon1.play1.tick_counter\[20\] _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2353_ _0421_ _0576_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2422_ _1110_ _0626_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1304_ simon1.score1.ones\[0\] simon1.score1.tens\[0\] _0745_ _0746_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2447__C _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2284_ _0461_ _0464_ _0520_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1999_ _0261_ _0262_ _0267_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2662__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1557__A1 _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1922_ _0200_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1853_ _1223_ _1227_ _1199_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2685__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1784_ simon1.seq_counter\[4\] _1167_ _1168_ _0834_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2405_ simon1.tick_counter\[14\] _0613_ _0614_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2336_ _0534_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2198_ simon1.state\[7\] _0811_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2267_ _1224_ _0487_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1711__A1 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xurish_simon_says_53 io_out[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_75 io_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_31 io_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_42 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_64 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_53_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2278__B _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2052_ _1258_ _1242_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2121_ _0379_ _0372_ _0350_ _0364_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1905_ simon1.play1.freq\[6\] simon1.play1.tick_counter\[6\] _1279_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1836_ _1205_ _1206_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1767_ _0828_ _1004_ _1158_ _1160_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1698_ _1109_ _1112_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2700__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2319_ _0522_ _0794_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1820__B _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput10 net10 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput8 net8 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__1932__A1 _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2098__B _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_46_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1621_ _1047_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2670_ _0099_ clknet_4_13_0_wb_clk_i simon1.tone_sequence_counter\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1552_ _0829_ _0987_ _0989_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2723__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I io_in[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2104_ _0362_ _0363_ _0364_ _0350_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__2479__A2 _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1483_ _0886_ _0912_ _0920_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_37_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2035_ _0299_ _1241_ _0303_ _0304_ _0246_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_27_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1819_ _1104_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2746__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2722_ _0151_ clknet_4_13_0_wb_clk_i net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2149__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1604_ simon1.state\[1\] _1033_ _1034_ _0985_ _1035_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2653_ _0082_ clknet_4_10_0_wb_clk_i simon1.play1.tick_counter\[22\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2584_ _0030_ clknet_4_0_0_wb_clk_i simon1.seq\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1535_ _0913_ _0969_ _0972_ _0898_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2619__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2321__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1397_ simon1.seq_counter\[1\] simon1.seq_counter\[0\] _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_1466_ _0892_ _0901_ _0903_ _0896_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_64_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2018_ _0193_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_45_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2220__I _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1320_ _0743_ _0751_ _0756_ _0761_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_51_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2286__B _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_19_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2636_ _0065_ clknet_4_14_0_wb_clk_i simon1.play1.tick_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2705_ _0134_ clknet_4_4_0_wb_clk_i simon1.tick_counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2567_ _1077_ simon1.seq\[9\]\[1\] _0726_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1449_ _0880_ _0885_ _0886_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2498_ _1131_ _0683_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1518_ _0953_ _0892_ _0896_ _0955_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2591__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1303_ _0731_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2352_ _0496_ _1004_ _0474_ _0561_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2283_ _0460_ _0517_ _0518_ _0519_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2421_ _0623_ _1130_ _0618_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_67_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2619_ _0192_ clknet_4_13_0_wb_clk_i net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1998_ _0259_ _1255_ _0251_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_30_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1852_ _1220_ _1225_ _1226_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1921_ _1231_ _1238_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1783_ _1031_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2335_ _0563_ _0564_ _0565_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2404_ simon1.tick_counter\[14\] _0613_ _0602_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2266_ _0503_ _0505_ _0484_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2197_ _0439_ _0429_ _0441_ _0428_ _0417_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_47_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1539__A2 _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1711__A2 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xurish_simon_says_21 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xurish_simon_says_54 io_out[33] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_76 io_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_32 io_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_43 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_65 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2120_ simon1.play1.tick_counter\[27\] _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_49_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2051_ simon1.play1.tick_counter\[18\] _1267_ _0300_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2652__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1835_ simon1.play1.freq\[2\] simon1.play1.tick_counter\[2\] _1212_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1904_ _1277_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1766_ _1000_ _0791_ _1159_ _1021_ _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1697_ _1110_ _1089_ _1111_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_12_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2318_ _0534_ _0539_ _0550_ _0551_ _0390_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2249_ _0463_ _0460_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1599__I _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1457__A1 _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput9 net9 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput11 net11 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2675__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1620_ _0782_ _1041_ _1046_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1551_ _0988_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1482_ _0913_ _0914_ _0919_ _0898_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2103_ _0362_ _1273_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2034_ _0296_ _0302_ _0198_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2100__A2 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1818_ simon1.play1.freq\[0\] _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2698__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1749_ _1147_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2158__A2 _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2094__A1 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2721_ _0150_ clknet_4_13_0_wb_clk_i net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2149__A2 _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2652_ _0081_ clknet_4_10_0_wb_clk_i simon1.play1.tick_counter\[21\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1603_ _1025_ _1028_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2583_ _0029_ clknet_4_0_0_wb_clk_i simon1.seq\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1465_ _0902_ simon1.seq\[4\]\[1\] _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1534_ _0915_ _0970_ _0971_ _0918_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2321__A2 _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1396_ simon1.seq_counter\[4\] _0833_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2017_ _0200_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_65_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1363__A3 _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1787__I _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2713__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2635_ _0064_ clknet_4_14_0_wb_clk_i simon1.play1.tick_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2704_ _0133_ clknet_4_4_0_wb_clk_i simon1.tick_counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2566_ _0727_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2736__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1448_ _0003_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1517_ simon1.seq\[0\]\[0\] _0954_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2497_ _0623_ _0682_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1379_ simon1.millis_counter\[6\] _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_2_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2297__B2 _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2609__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2420_ _0622_ _0625_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2351_ _0421_ _0576_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1302_ _0737_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2282_ _0496_ _0434_ _0441_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_59_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1997_ simon1.play1.tick_counter\[13\] _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2618_ _0191_ clknet_4_13_0_wb_clk_i net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2549_ simon1.seq\[25\]\[0\] _0705_ _0716_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1851_ _1224_ simon1.play1.tick_counter\[4\] _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1920_ _1230_ _1241_ _1286_ _0199_ _0790_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2403_ _0597_ _0612_ _0613_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1782_ _1032_ _1172_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2581__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2196_ _0825_ _0431_ _0440_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2334_ _0798_ _0559_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2265_ _0995_ _0454_ _0504_ _0495_ _0450_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xurish_simon_says_55 io_out[34] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_33 io_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_44 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_22 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xurish_simon_says_77 io_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_66 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_21_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ _0289_ _0308_ _0312_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_52_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1834_ _1208_ _1210_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1765_ simon1.state\[5\] _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1903_ _1263_ _1270_ _1276_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_TAPCELL_ROW_32_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1696_ simon1.seq_length\[4\] _1065_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2179_ _0815_ _0824_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2317_ _0821_ _0549_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2248_ _1006_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput12 net12 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_50_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1550_ _0788_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1481_ _0915_ _0916_ _0917_ _0918_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2033_ _0296_ _0302_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_27_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2102_ _1273_ _0335_ _0347_ _0349_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_57_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1817_ _1189_ _1195_ _1197_ _1175_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1375__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1748_ _1139_ simon1.seq\[4\]\[1\] _1145_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1679_ simon1.seq_length\[0\] _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2642__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2409__I _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2720_ _0149_ clknet_4_7_0_wb_clk_i net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1602_ _0849_ _0978_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2582_ _0028_ clknet_4_0_0_wb_clk_i simon1.seq\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2651_ _0080_ clknet_4_10_0_wb_clk_i simon1.play1.tick_counter\[20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1395_ _0831_ _0832_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1533_ _0954_ simon1.seq\[8\]\[0\] _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1464_ _0000_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_65_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2016_ _1252_ _0276_ _0286_ _0287_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_19_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2665__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2076__A2 _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2688__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2703_ _0132_ clknet_4_4_0_wb_clk_i simon1.tick_counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2634_ _0063_ clknet_4_11_0_wb_clk_i simon1.play1.tick_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2565_ _1061_ simon1.seq\[9\]\[0\] _0726_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1516_ _0855_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1378_ simon1.millis_counter\[5\] _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_49_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2496_ simon1.seq_length\[4\] _1068_ _1092_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1447_ _0851_ _0881_ _0884_ _0872_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_53_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2058__A2 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1301_ _0729_ _0734_ _0742_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2350_ _0567_ _0575_ _0576_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2281_ _0468_ _0436_ _0508_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_32_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1996_ _0259_ _0249_ _0269_ _1166_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_15_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2617_ _0190_ clknet_4_13_0_wb_clk_i net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2703__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2548_ _1067_ _0687_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2479_ _1082_ _1153_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_65_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_21_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1850_ _1224_ simon1.play1.tick_counter\[4\] _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1781_ simon1.seq_counter\[3\] _1167_ _1168_ _0844_ _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2726__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2333_ _0798_ _0559_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2402_ simon1.tick_counter\[13\] _0610_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2195_ _0416_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2264_ _0801_ _0492_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ _0247_ _0253_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xurish_simon_says_56 io_out[35] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_78 io_oeb[33] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_45 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_67 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_34 io_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_23 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_7_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2749__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2360__A1 _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1902_ _1271_ _1272_ _1274_ _1275_ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_32_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1764_ _1053_ _1034_ _1157_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1833_ _1209_ simon1.play1.tick_counter\[3\] _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2316_ _0821_ _0549_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1695_ simon1.seq_length\[3\] _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2178_ _0791_ _0808_ _1021_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_48_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2247_ _0485_ _0488_ _0998_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput13 net13 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_50_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2571__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1480_ _0861_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_37_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2032_ _0300_ _0301_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2101_ simon1.play1.tick_counter\[25\] _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_27_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1816_ simon1.score1.tens\[3\] _1196_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1375__A2 _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1678_ _1097_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1747_ _1146_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2594__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_42_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1601_ _1016_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1532_ simon1.seq\[9\]\[0\] _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2650_ _0079_ clknet_4_10_0_wb_clk_i simon1.play1.tick_counter\[19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2581_ _0027_ clknet_4_0_0_wb_clk_i simon1.seq\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input1_I io_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1394_ simon1.seq_counter\[2\] simon1.seq_counter\[1\] simon1.seq_counter\[0\] _0832_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_1_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1463_ simon1.seq\[5\]\[1\] _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2015_ _0988_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1414__I _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2702_ _0131_ clknet_4_4_0_wb_clk_i simon1.tick_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2633_ _0062_ clknet_4_11_0_wb_clk_i simon1.play1.tick_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2564_ _1141_ _1091_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2495_ _0681_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1515_ simon1.seq\[1\]\[0\] _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1377_ simon1.state\[3\] _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1446_ _0857_ _0882_ _0883_ _0862_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2632__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1853__B _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2509__A1 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1300_ _0734_ _0737_ _0741_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2280_ _0502_ _0497_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2655__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2616_ _0189_ clknet_4_13_0_wb_clk_i net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1995_ _0260_ _0268_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1971__A2 _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1429_ simon1.seq\[29\]\[1\] _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2547_ _0715_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2478_ _1079_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2523__I _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2678__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1780_ _1032_ _1171_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_12_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2332_ _0522_ _0562_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2401_ simon1.tick_counter\[13\] _0610_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2194_ _0826_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2263_ _0501_ _0502_ _1011_ _0460_ _0466_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_46_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_23_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1978_ _0234_ _0240_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_15_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xurish_simon_says_57 io_out[36] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_79 io_oeb[34] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_46 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_68 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_35 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_24 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_21_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1832_ simon1.play1.freq\[3\] _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1901_ simon1.play1.tick_counter\[29\] simon1.play1.tick_counter\[28\] simon1.play1.tick_counter\[27\]
+ simon1.play1.tick_counter\[26\] _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1763_ _0979_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1694_ _1081_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2315_ _0548_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2246_ simon1.play1.freq\[2\] _0487_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2177_ _0416_ _1010_ _0419_ _0423_ _0808_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_48_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput14 net14 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_31_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1417__I _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2716__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2100_ _0357_ _0276_ _0361_ _0287_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2031_ _0280_ _0293_ _1259_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_27_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1815_ simon1.score1.tens\[2\] simon1.score1.tens\[1\] _1188_ _1196_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_40_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1677_ simon1.seq\[11\]\[1\] _1077_ _1095_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1746_ _1136_ simon1.seq\[4\]\[0\] _1145_ _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2229_ _0436_ _0471_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2739__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2531__I _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1600_ _1031_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1531_ simon1.seq\[10\]\[0\] simon1.seq\[11\]\[0\] _0902_ _0969_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1462_ simon1.seq\[6\]\[1\] simon1.seq\[7\]\[1\] _0890_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2580_ _0026_ clknet_4_3_0_wb_clk_i simon1.seq\[16\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1393_ simon1.seq_counter\[3\] _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2014_ _0279_ _0284_ _0285_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1729_ _1134_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1586__B _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2472__A1 _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2701_ _0130_ clknet_4_4_0_wb_clk_i simon1.tick_counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2632_ _0061_ clknet_4_9_0_wb_clk_i simon1.play1.tick_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2584__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2494_ simon1.seq\[28\]\[1\] _0668_ _0679_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1445_ _0868_ simon1.seq\[20\]\[1\] _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1514_ simon1.seq\[2\]\[0\] simon1.seq\[3\]\[0\] _0890_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2563_ _0725_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1376_ _0790_ _0792_ _0806_ _0814_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_4_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ _0263_ _0267_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_15_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2615_ _0188_ clknet_4_13_0_wb_clk_i net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2546_ simon1.seq\[23\]\[1\] _0708_ _0713_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1428_ simon1.seq\[30\]\[1\] simon1.seq\[31\]\[1\] _0853_ _0866_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2477_ _0669_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1359_ _0797_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _0610_ _0611_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_12_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2331_ _1026_ _1022_ _0536_ _0561_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2262_ _0410_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2622__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2193_ _0429_ _0437_ _0438_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ _1255_ _0251_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2529_ _0700_ simon1.seq\[18\]\[1\] _0702_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1703__I _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xurish_simon_says_58 io_out[37] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_69 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_36 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_47 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_25 io_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2645__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1831_ simon1.play1.freq\[3\] simon1.play1.tick_counter\[3\] _1208_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_32_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1900_ simon1.play1.tick_counter\[25\] _1273_ simon1.play1.tick_counter\[23\] _1274_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_40_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1693_ _1108_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1762_ _1156_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2176_ _0981_ _1001_ _0420_ _0422_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_2314_ _0541_ _0543_ _0545_ _0547_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2245_ _0486_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2668__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput15 net15 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2030_ simon1.play1.tick_counter\[16\] _0278_ _0293_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_27_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1814_ _1190_ _1191_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1745_ _1109_ _1132_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1676_ _1096_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2159_ _1015_ _1019_ _0409_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2228_ _0423_ _0470_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1392_ simon1.seq_length\[4\] _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_1461_ _0889_ _0891_ _0897_ _0898_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1530_ _0913_ _0964_ _0967_ _0905_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2013_ _0279_ _0284_ _0208_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2706__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1728_ simon1.seq\[7\]\[0\] _1116_ _1133_ _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1659_ _1081_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_56_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_64_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2700_ _0129_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2631_ _0060_ clknet_4_9_0_wb_clk_i simon1.play1.tick_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2729__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2562_ _0700_ simon1.seq\[31\]\[1\] _0723_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1375_ _0807_ _0809_ _0813_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1444_ simon1.seq\[21\]\[1\] _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2493_ _0680_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1513_ _0939_ _0950_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1993_ _0248_ _0264_ _0265_ _0266_ _1277_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_27_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2614_ _0187_ clknet_4_13_0_wb_clk_i net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2545_ _0714_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1358_ simon1.millis_counter\[3\] _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2476_ simon1.seq\[19\]\[1\] _0668_ _0666_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1427_ _0851_ _0854_ _0863_ _0864_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1289_ simon1.score1.active_digit _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1947__A1 _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2574__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2192_ _0432_ _0427_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2330_ _0993_ _1105_ _0537_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2261_ simon1.user_input\[0\] _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1976_ _0239_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2597__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2528_ _0703_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2459_ _0646_ _0643_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xurish_simon_says_37 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_26 io_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_53_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xurish_simon_says_48 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_59 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1830_ _1173_ _1207_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1761_ simon1.seq\[21\]\[1\] _1119_ _1154_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2313_ simon1.tick_counter\[12\] _0546_ simon1.tick_counter\[14\] simon1.tick_counter\[15\]
+ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_52_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1692_ simon1.seq\[0\]\[1\] _1077_ _1106_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2175_ simon1.millis_counter\[9\] _0421_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2244_ _0443_ _0445_ _0446_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1959_ _0218_ _0220_ _0231_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_31_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput16 net16 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2612__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1813_ _1129_ _1194_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1744_ _1144_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1675_ simon1.seq\[11\]\[0\] _1061_ _1095_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2158_ _0408_ _1019_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2635__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2227_ _0794_ _0469_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2089_ _0351_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_39_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2548__A1 _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_57_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1391_ _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2658__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1460_ _0002_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_66_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2012_ _0219_ _0283_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1727_ _1131_ _1132_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1658_ _1062_ _1064_ _1065_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1589_ _1021_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_64_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2630_ _0059_ clknet_4_15_0_wb_clk_i simon1.score1.tens\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1349__I _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1983__A2 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2492_ simon1.seq\[28\]\[0\] _0665_ _0679_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1512_ _0944_ _0949_ _0886_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2561_ _0724_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1374_ _0787_ _0812_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1443_ simon1.seq\[22\]\[1\] simon1.seq\[23\]\[1\] _0853_ _0881_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1722__I _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1956__A2 _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1992_ _0196_ _0206_ _0218_ _0231_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_15_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2613_ _0186_ clknet_4_13_0_wb_clk_i net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2544_ simon1.seq\[23\]\[0\] _0705_ _0713_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2475_ _1076_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1357_ _0795_ simon1.millis_counter\[8\] _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1288_ simon1.score1.ones\[3\] _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2133__A2 _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1426_ _0002_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2719__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2041__C _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2191_ _0433_ _0434_ _0436_ _0809_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2260_ _0489_ _0500_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1975_ _0235_ _0241_ _1278_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2458_ _0630_ _0654_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1981__B _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1409_ _0843_ _0844_ _0846_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2527_ _0697_ simon1.seq\[18\]\[0\] _0702_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2389_ simon1.tick_counter\[9\] _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_26_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xurish_simon_says_49 io_out[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_38 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_27 io_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2290__A1 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2345__A2 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2691__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1691_ _1107_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1760_ _1155_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2312_ simon1.tick_counter\[13\] _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_27_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2174_ simon1.millis_counter\[8\] _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1847__A1 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2243_ _0482_ _0483_ _0484_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_11_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput17 net17 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_43_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1958_ simon1.play1.tick_counter\[10\] _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1889_ _1242_ _1245_ _1257_ _1261_ _1262_ _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_31_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2587__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2471__I _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1812_ simon1.score1.tens\[2\] _1193_ _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1674_ _1091_ _1094_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1743_ _1139_ simon1.seq\[5\]\[1\] _1142_ _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2226_ simon1.millis_counter\[0\] simon1.millis_counter\[1\] _0469_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2157_ simon1.user_input\[0\] _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2088_ simon1.play1.tick_counter\[23\] _0348_ _0350_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_48_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1390_ _0815_ _0827_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_54_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2011_ _0266_ _0265_ _0280_ _0281_ _0282_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2415__B _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1588_ _0815_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1657_ _1079_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1726_ _0830_ _1069_ _1070_ _1090_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_56_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2209_ _0440_ _0452_ _0431_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2752__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2602__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2625__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2491_ _1082_ _0678_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1511_ _0925_ _0945_ _0948_ _0872_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1442_ _0851_ _0876_ _0879_ _0864_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2560_ _0697_ simon1.seq\[31\]\[0\] _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1373_ _0811_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1476__S _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2689_ _0118_ clknet_4_5_0_wb_clk_i simon1.millis_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1709_ _1120_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2648__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1991_ _1255_ _0251_ _0253_ _0247_ _0264_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_2612_ _0050_ clknet_4_6_0_wb_clk_i _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_27_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2543_ _1093_ _1153_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1425_ _0857_ _0858_ _0860_ _0862_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2474_ _0667_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_66_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1287_ net3 _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1356_ simon1.millis_counter\[9\] _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_46_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1571__A1 _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2190_ _0435_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1974_ _0198_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2457_ net8 _0633_ _0653_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1553__I _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2388_ _0601_ _0603_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1562__A1 _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1408_ _0843_ _0844_ _0845_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2526_ _1100_ _1112_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_66_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1339_ _0757_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_26_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xurish_simon_says_39 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_28 io_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1690_ simon1.seq\[0\]\[0\] _1061_ _1106_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2242_ _0447_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2311_ simon1.tick_counter\[11\] _0544_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2173_ _0797_ simon1.millis_counter\[7\] _0804_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_48_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1957_ _0202_ _0232_ _0233_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_31_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2709__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_23_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput18 net18 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1888_ simon1.play1.tick_counter\[22\] _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2509_ _1121_ _0678_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_66_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2063__B _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1811_ _1190_ _1188_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1742_ _1143_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1673_ _1093_ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2225_ _0442_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2156_ _0407_ _0987_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2087_ _0335_ _0347_ _0349_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2681__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1995__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ _0247_ _0241_ _0261_ _0262_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__2482__I _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1725_ _1130_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1587_ _0791_ _0806_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1656_ _1059_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2208_ _0451_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2139_ _0387_ _0395_ _0275_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1736__I _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2154__A1 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2577__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2490_ _1088_ _1068_ _1069_ _1092_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_10_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1510_ _0927_ _0946_ _0947_ _0931_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1441_ _0857_ _0877_ _0878_ _0862_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1372_ net4 net1 _0810_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_65_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_61_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2145__C _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2688_ _0117_ clknet_4_5_0_wb_clk_i simon1.millis_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1708_ simon1.seq\[15\]\[1\] _1119_ _1117_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1639_ simon1.seq_length\[0\] _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_1_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1990_ simon1.play1.tick_counter\[10\] _0240_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_7_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2611_ _0049_ clknet_4_6_0_wb_clk_i _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2542_ _0712_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2742__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1355_ _0793_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__2118__A1 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2473_ simon1.seq\[19\]\[0\] _0665_ _0666_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1424_ _0861_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2109__A1 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2615__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2520__A1 _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1973_ _0247_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_15_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2525_ _0701_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1338_ _0744_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2456_ _0645_ _0651_ _0652_ _0634_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2638__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2387_ simon1.tick_counter\[8\] _0599_ _0602_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1407_ simon1.seq_counter\[4\] _0833_ _0830_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_26_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xurish_simon_says_29 io_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_61_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2172_ _0417_ _0418_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_2241_ _0462_ _0461_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2310_ simon1.tick_counter\[8\] simon1.tick_counter\[9\] simon1.tick_counter\[10\]
+ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_20_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1956_ simon1.play1.tick_counter\[9\] _0209_ _0223_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1887_ simon1.play1.tick_counter\[22\] _1258_ _1260_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_31_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2508_ _0690_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2439_ _0635_ _1054_ _0636_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_39_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1810_ _1190_ _1189_ _1192_ _1129_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_57_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1741_ _1136_ simon1.seq\[5\]\[0\] _1142_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1672_ _1063_ _1064_ _1092_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_2224_ _0465_ _0466_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2155_ _1006_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_36_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2086_ simon1.play1.tick_counter\[23\] simon1.play1.tick_counter\[22\] _0349_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1939_ _1283_ _0212_ _0213_ _1220_ _0216_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2058__C _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_35_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_44_Left_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1724_ _1062_ simon1.seq_length\[0\] _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1586_ _1007_ _1011_ _1019_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1655_ _1078_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2207_ _0825_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_53_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2138_ _0391_ _0392_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2069_ _0332_ _0333_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_64_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_62_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1371_ net5 net2 _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_50_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2145__A2 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1440_ _0859_ simon1.seq\[16\]\[1\] _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2671__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2687_ _0116_ clknet_4_5_0_wb_clk_i simon1.millis_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2756_ _0185_ clknet_4_4_0_wb_clk_i simon1.seq\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1638_ _1062_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1707_ _1076_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1569_ _1000_ _1003_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_52_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1647__A1 _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_9_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2694__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2610_ _0048_ clknet_4_6_0_wb_clk_i _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1657__I _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2541_ simon1.seq\[29\]\[1\] _0708_ _0710_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2472_ _1094_ _1112_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1354_ simon1.millis_counter\[0\] simon1.millis_counter\[1\] _0793_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1423_ _0001_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2739_ _0168_ clknet_4_3_0_wb_clk_i simon1.seq\[24\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2045__A1 _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2066__C _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1859__A1 simon1.play1.freq\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1972_ simon1.play1.tick_counter\[11\] _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2455_ _0404_ _0796_ _0638_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2524_ _0700_ simon1.seq\[24\]\[1\] _0698_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1337_ _0748_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2386_ _0584_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1406_ _0831_ _0832_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2167__B _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2732__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2171_ simon1.tone_sequence_counter\[0\] simon1.tone_sequence_counter\[1\] _0418_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2240_ _0994_ _0434_ _0481_ _1011_ _0411_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1955_ _0225_ _0231_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_31_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1886_ simon1.play1.tick_counter\[21\] simon1.play1.tick_counter\[20\] _1259_ _1242_
+ _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_7_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2438_ _1159_ _0999_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2605__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2507_ simon1.seq\[26\]\[1\] _0668_ _0688_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2369_ simon1.tick_counter\[3\] _0588_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2755__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2628__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1671_ _1057_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1740_ _1141_ _1132_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2154_ _1216_ _0406_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2223_ _0462_ _0463_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2085_ _0345_ _0335_ _0347_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1938_ _1234_ _1248_ _0215_ _1235_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_31_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1869_ simon1.play1.tick_counter\[21\] _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1723_ _0745_ _1129_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1654_ simon1.seq\[13\]\[1\] _1077_ _1072_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2163__A3 _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2206_ _1022_ _0449_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1585_ _1018_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2137_ _0368_ _0382_ _0386_ _0393_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_2068_ _1243_ _1244_ _0321_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1674__A2 _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1370_ _0808_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2686_ _0115_ clknet_4_5_0_wb_clk_i simon1.millis_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2755_ _0184_ clknet_4_4_0_wb_clk_i simon1.seq\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1637_ simon1.seq_length\[1\] _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1706_ _1118_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_18_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1568_ _1002_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1647__A2 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1499_ _0927_ _0935_ _0936_ _0931_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_52_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2540_ _0711_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2471_ _1060_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1422_ _0859_ simon1.seq\[24\]\[1\] _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1673__I _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1353_ _0791_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_46_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2738_ _0167_ clknet_4_1_0_wb_clk_i simon1.seq\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2669_ _0098_ clknet_4_9_0_wb_clk_i simon1.next_random\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_29_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1556__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2661__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1971_ _0234_ _1241_ _0242_ _0245_ _0246_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_15_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2454_ _0646_ _0648_ _0650_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2385_ _0600_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1405_ simon1.seq_length\[3\] _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2523_ _1085_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput1 io_in[10] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1336_ _0762_ _0776_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1786__A1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2027__A2 _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2684__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2170_ simon1.tone_sequence_counter\[2\] _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2268__B _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1954_ _0227_ _0230_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_48_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1885_ simon1.play1.tick_counter\[16\] _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_31_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2368_ _0587_ _0588_ _0589_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2437_ _1021_ simon1.state\[1\] _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2506_ _0689_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1319_ _0729_ _0758_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2299_ _0489_ _0533_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_6_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ _1088_ _1089_ _1090_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2222_ _0464_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2153_ _0807_ _0405_ simon1.score1.ena _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2084_ _0346_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_63_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1937_ _0214_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2722__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1799_ simon1.score1.inc simon1.score1.ones\[0\] _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1868_ simon1.play1.tick_counter\[19\] simon1.play1.tick_counter\[18\] _1242_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_58_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1722_ _1128_ _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1584_ _1017_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2148__A1 _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1653_ _1076_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2745__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2205_ _0416_ simon1.tone_sequence_counter\[1\] _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2136_ simon1.play1.tick_counter\[29\] _0392_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2067_ _1244_ _0321_ _1243_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_63_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2618__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1705_ simon1.seq\[15\]\[0\] _1116_ _1117_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2754_ _0183_ clknet_4_8_0_wb_clk_i simon1.seq\[31\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1567_ _0797_ _0796_ _0818_ _1001_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2685_ _0114_ clknet_4_5_0_wb_clk_i simon1.millis_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1636_ _1060_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_1_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1498_ _0929_ simon1.seq\[28\]\[0\] _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2119_ _0372_ _0326_ _0376_ _0378_ _0246_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_52_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2532__A1 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2590__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2470_ _0630_ _0664_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1421_ _0852_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1352_ simon1.state\[4\] _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2668_ _0097_ clknet_4_9_0_wb_clk_i simon1.next_random\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2737_ _0166_ clknet_4_1_0_wb_clk_i simon1.seq\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1619_ _0763_ _0770_ _0767_ _1044_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2599_ _0037_ clknet_4_0_0_wb_clk_i simon1.seq\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2514__A1 _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ _0789_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2522_ _0699_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1335_ _0765_ _0775_ _0764_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2453_ _0501_ _1009_ _0649_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2384_ simon1.tick_counter\[8\] _0599_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1404_ simon1.seq_length\[1\] _0835_ _0838_ _0841_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_23_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 io_in[11] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_25_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ _0228_ _0229_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1884_ simon1.play1.tick_counter\[17\] _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2505_ simon1.seq\[26\]\[0\] _0665_ _0688_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2367_ simon1.tick_counter\[1\] _0542_ simon1.tick_counter\[2\] _0589_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2436_ _0632_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1318_ _0744_ _0759_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2298_ simon1.play1.freq\[9\] _0515_ _0503_ _0532_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_22_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2651__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1931__A2 _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2152_ _0404_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2221_ _0462_ _0463_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2674__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2083_ simon1.play1.tick_counter\[21\] simon1.play1.tick_counter\[20\] _0346_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1936_ _1234_ simon1.play1.tick_counter\[7\] _1229_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1867_ _1240_ _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1798_ _1175_ _1182_ _1183_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2419_ _0623_ _0624_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2697__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1721_ simon1.score_rst _0788_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_38_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1583_ simon1.state\[1\] _0813_ _1016_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1652_ _1075_ _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2204_ _0447_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2135_ simon1.play1.tick_counter\[28\] _0380_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2066_ _0325_ _0326_ _0330_ _0331_ _0246_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1919_ _0195_ _0196_ _0198_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_55_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2712__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2684_ _0113_ clknet_4_5_0_wb_clk_i simon1.millis_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1704_ _1071_ _1093_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2753_ _0182_ clknet_4_3_0_wb_clk_i simon1.seq\[31\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1566_ simon1.millis_counter\[2\] _0793_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1635_ _1059_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1497_ simon1.seq\[29\]\[0\] _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2118_ _0243_ _0377_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2057__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2049_ simon1.play1.tick_counter\[19\] _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2532__A2 _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2735__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2048__A1 _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1351_ _0789_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1420_ simon1.seq\[25\]\[1\] _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2667_ _0096_ clknet_4_7_0_wb_clk_i simon1.user_input\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1618_ _0778_ _0775_ _1043_ _1045_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2211__A1 _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2608__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2736_ _0165_ clknet_4_8_0_wb_clk_i simon1.seq\[30\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1549_ _0849_ _0986_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_5_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2598_ _0036_ clknet_4_0_0_wb_clk_i simon1.seq\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2269__A1 _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2521_ _0697_ simon1.seq\[24\]\[0\] _0698_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1334_ _0758_ _0767_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2383_ _0597_ _0598_ _0599_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2452_ _1008_ _0463_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1403_ simon1.seq_length\[2\] _0840_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 io_in[26] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2432__A1 _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2719_ _0148_ clknet_4_13_0_wb_clk_i net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1824__B _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2580__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1952_ simon1.play1.freq\[9\] simon1.play1.tick_counter\[9\] _0229_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1883_ _1246_ _1247_ _1256_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2435_ _0632_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2504_ _1121_ _0687_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_24_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2366_ simon1.tick_counter\[1\] simon1.tick_counter\[0\] simon1.tick_counter\[2\]
+ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1317_ _0746_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2297_ _0450_ _0529_ _0531_ _0995_ _0457_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2151_ _0812_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2220_ _0976_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2082_ simon1.play1.tick_counter\[22\] _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_17_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1797_ simon1.score1.ones\[2\] _1179_ _1177_ _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1935_ _1280_ _0212_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1866_ _1239_ _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1374__A1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2418_ _1130_ _0619_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2349_ _0803_ _0804_ _0571_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_62_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2093__A2 _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1651_ _1074_ _1058_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1720_ _1127_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1582_ _0810_ _1012_ _1013_ _1015_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2641__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input6_I wb_rst_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2203_ _0443_ _0445_ _0446_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2134_ simon1.play1.tick_counter\[29\] _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2065_ _0327_ _0329_ _0198_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1849_ simon1.play1.freq\[4\] _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1918_ _0197_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2219__I _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2664__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1586__A1 _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2066__A2 _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2683_ _0112_ clknet_4_4_0_wb_clk_i simon1.millis_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1634_ _1048_ _1058_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2752_ _0181_ clknet_4_3_0_wb_clk_i simon1.seq\[17\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1703_ _1060_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1565_ simon1.state\[6\] _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1496_ simon1.seq\[30\]\[0\] simon1.seq\[31\]\[0\] _0868_ _0934_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2048_ _0202_ _0314_ _0315_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2117_ _0369_ _0375_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2687__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1562__B _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1740__A1 _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_Left_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1350_ _0788_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_66_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1617_ _0743_ _1044_ _0764_ _0766_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2666_ _0095_ clknet_4_7_0_wb_clk_i simon1.user_input\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2597_ _0035_ clknet_4_0_0_wb_clk_i simon1.seq\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2735_ _0164_ clknet_4_8_0_wb_clk_i simon1.seq\[30\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1548_ _0978_ _0985_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1479_ _0902_ simon1.seq\[8\]\[1\] _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2702__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2451_ _0555_ _0467_ _0647_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1952__A1 simon1.play1.freq\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1402_ simon1.seq_counter\[2\] _0839_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2520_ _1109_ _0683_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[8] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1333_ _0774_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2382_ simon1.tick_counter\[7\] _0596_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1704__A1 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2718_ _0147_ clknet_4_6_0_wb_clk_i simon1.seq_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2725__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2649_ _0078_ clknet_4_10_0_wb_clk_i simon1.play1.tick_counter\[18\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1951_ simon1.play1.freq\[9\] simon1.play1.tick_counter\[9\] _0228_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1882_ _1249_ _1251_ _1253_ _1255_ _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2748__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2365_ _0584_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2434_ _0792_ _0446_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2503_ _1089_ _0682_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1316_ _0757_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2296_ _0423_ _0530_ _0454_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2332__A1 _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2150_ _0790_ _0249_ _0403_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2081_ _1262_ _0343_ _0344_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1934_ _1279_ _0203_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2570__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1796_ _1179_ _1178_ simon1.score1.ones\[2\] _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1865_ _1231_ _1238_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2348_ _0804_ _0571_ _0803_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2417_ simon1.seq_length\[2\] _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2279_ _0514_ _0516_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2593__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1520__S _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1581_ _0810_ _1012_ _1014_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_41_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1650_ simon1.next_random\[1\] _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2202_ _1000_ _0984_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2553__A1 _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2133_ _0385_ _0326_ _0387_ _0389_ _0390_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_21_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2064_ _0327_ _0329_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1917_ _1239_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1848_ simon1.play1.freq\[5\] simon1.play1.tick_counter\[5\] _1223_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1779_ simon1.seq_counter\[2\] _1167_ _1168_ _0840_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2751_ _0180_ clknet_4_3_0_wb_clk_i simon1.seq\[17\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2682_ _0111_ clknet_4_12_0_wb_clk_i simon1.play1.freq\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1564_ simon1.state\[2\] _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1633_ _0990_ _1052_ _1057_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1702_ _1115_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2526__A1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1495_ _0925_ _0926_ _0932_ _0864_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2047_ simon1.play1.tick_counter\[18\] _0201_ _0223_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2116_ _0368_ _0375_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2631__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_66_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2734_ _0163_ clknet_4_8_0_wb_clk_i simon1.seq\[26\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1616_ _0741_ _0754_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2665_ _0094_ clknet_4_12_0_wb_clk_i simon1.score1.inc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1547_ _0979_ _0984_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2596_ _0034_ clknet_4_0_0_wb_clk_i simon1.seq\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1478_ simon1.seq\[9\]\[1\] _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2654__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2381_ simon1.tick_counter\[7\] _0596_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2450_ _1008_ _0473_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1401_ simon1.seq_counter\[1\] simon1.seq_counter\[0\] _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1704__A2 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 io_in[9] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1332_ _0762_ _0769_ _0773_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2677__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2717_ _0146_ clknet_4_6_0_wb_clk_i simon1.seq_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2648_ _0077_ clknet_4_10_0_wb_clk_i simon1.play1.tick_counter\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2579_ _0025_ clknet_4_3_0_wb_clk_i simon1.seq\[16\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1698__A1 _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1950_ _0211_ _0217_ _0226_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1881_ _1254_ _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2502_ _0686_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2364_ _0585_ _0586_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2433_ net7 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1315_ _0733_ _0740_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1689__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2295_ _0508_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2715__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2080_ _1262_ _0343_ _0223_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1933_ simon1.play1.freq\[8\] simon1.play1.tick_counter\[8\] _0211_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_44_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1795_ _1179_ _1178_ _1181_ _1129_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1864_ _1233_ _1237_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2347_ _0573_ _0574_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2278_ _1235_ _0515_ _0992_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2416_ _1131_ _0619_ _0621_ _0622_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_10_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2738__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1600__I _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1580_ net5 net2 _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2201_ _0444_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2132_ _0789_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2063_ _0308_ _0328_ _1278_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1847_ _1216_ _1222_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1916_ _1285_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_44_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1778_ _1032_ _1170_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_63_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2681_ _0110_ clknet_4_12_0_wb_clk_i simon1.play1.freq\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2750_ _0179_ clknet_4_2_0_wb_clk_i simon1.seq\[25\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1701_ _1086_ simon1.seq\[16\]\[1\] _1113_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1563_ _0988_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1632_ _0848_ _0996_ _1056_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1494_ _0927_ _0928_ _0930_ _0931_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_55_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2110__B _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2115_ _0373_ _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2046_ _0312_ _0313_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2214__B2 _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2583__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1526__S _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2664_ _0093_ clknet_4_13_0_wb_clk_i simon1.score1.ena vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2733_ _0162_ clknet_4_8_0_wb_clk_i simon1.seq\[26\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1615_ _0753_ _0760_ _0780_ _0778_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1546_ _0983_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2595_ _0012_ clknet_4_6_0_wb_clk_i simon1.state\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1477_ _0856_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1486__A2 _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2029_ _1259_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1331_ _0759_ _0770_ _0771_ _0742_ _0772_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2380_ _0584_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1400_ simon1.seq_length\[1\] _0835_ _0837_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput6 wb_rst_i net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2716_ _0145_ clknet_4_6_0_wb_clk_i simon1.seq_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2647_ _0076_ clknet_4_10_0_wb_clk_i simon1.play1.tick_counter\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2621__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2578_ _0024_ clknet_4_6_0_wb_clk_i simon1.seq\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1529_ _0915_ _0965_ _0966_ _0918_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_25_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ simon1.play1.tick_counter\[11\] simon1.play1.tick_counter\[10\] _1254_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_38_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_47_Left_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2644__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2501_ _0673_ simon1.seq\[27\]\[1\] _0684_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2363_ simon1.tick_counter\[1\] _0542_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1314_ _0753_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2294_ _0440_ _0432_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2432_ _1007_ _1174_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_56_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_65_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2519__I _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2667__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1863_ _1234_ _1235_ _1236_ _1224_ _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1932_ _0202_ _0207_ _0210_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1794_ _1178_ _1180_ _1179_ _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2415_ _0792_ _1009_ _1104_ _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2346_ _0817_ _0571_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2277_ _0457_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2002__A2 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2200_ simon1.state\[2\] _1051_ _0426_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2062_ simon1.play1.tick_counter\[19\] _0311_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2131_ _0260_ _0388_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1846_ _1220_ _1221_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1915_ _0194_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1777_ simon1.seq_counter\[1\] _1167_ _1168_ _1169_ _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2329_ _0790_ _0559_ _0560_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_47_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2705__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2680_ _0109_ clknet_4_12_0_wb_clk_i simon1.play1.freq\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1631_ _1053_ _1049_ _1054_ _1055_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1700_ _1114_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1562_ _0995_ _0997_ _0989_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1493_ _0861_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input4_I io_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2045_ _0194_ _0308_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2114_ simon1.play1.tick_counter\[26\] _0362_ _1273_ _0358_ _0374_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_29_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1829_ _1205_ _1206_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_32_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2728__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2150__A1 _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1716__A1 _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1614_ _0772_ _1038_ _0783_ _1042_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_54_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2663_ _0092_ clknet_4_14_0_wb_clk_i net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2594_ _0011_ clknet_4_7_0_wb_clk_i simon1.state\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2732_ _0161_ clknet_4_2_0_wb_clk_i simon1.seq\[27\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1545_ simon1.millis_counter\[3\] simon1.millis_counter\[2\] _0980_ _0982_ _0983_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1476_ simon1.seq\[10\]\[1\] simon1.seq\[11\]\[1\] _0894_ _0914_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2028_ _1216_ _0298_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_20_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1330_ _0729_ _0753_ _0758_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_52_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2573__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2715_ _0144_ clknet_4_6_0_wb_clk_i simon1.seq_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2646_ _0075_ clknet_4_11_0_wb_clk_i simon1.play1.tick_counter\[15\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2577_ _0023_ clknet_4_6_0_wb_clk_i simon1.seq\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1528_ _0954_ simon1.seq\[12\]\[0\] _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1459_ _0892_ _0893_ _0895_ _0896_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_33_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2596__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2431_ _1007_ _1172_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2500_ _0685_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2362_ _0542_ _0585_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1313_ _0741_ _0754_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2293_ _0489_ _0528_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2629_ _0058_ clknet_4_15_0_wb_clk_i simon1.score1.tens\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2535__I _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2317__A1 _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1793_ _0730_ simon1.score1.ones\[2\] _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_56_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1862_ simon1.play1.freq\[5\] _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1931_ _1248_ _0209_ _1199_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2611__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2414_ _1098_ _0619_ _1063_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2345_ _1027_ _1023_ _0572_ _1104_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2276_ _0487_ _0490_ _0497_ _0513_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_30_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2634__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2538__A1 _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2061_ _1244_ _0321_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2130_ _0369_ _0382_ _0386_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1914_ _0193_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1845_ simon1.play1.freq\[4\] simon1.play1.tick_counter\[4\] _1221_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1776_ _0835_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2328_ _1027_ _0536_ _0538_ _0553_ _0800_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2657__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2259_ _1209_ _0448_ _0499_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1630_ net6 simon1.state\[4\] simon1.state\[2\] _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_41_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1561_ _0996_ _0985_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1492_ _0929_ simon1.seq\[24\]\[0\] _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2044_ _0311_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2113_ _0350_ _0364_ _0372_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_57_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ simon1.play1.freq\[2\] simon1.play1.tick_counter\[2\] _1206_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1759_ simon1.seq\[21\]\[0\] _1116_ _1154_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_9_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2150__A2 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2731_ _0160_ clknet_4_3_0_wb_clk_i simon1.seq\[27\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1613_ _1039_ _1041_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1544_ _0793_ _0796_ _0981_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2593_ _0010_ clknet_4_12_0_wb_clk_i simon1.state\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2662_ _0091_ clknet_4_9_0_wb_clk_i simon1.play1.tick_counter\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1475_ _0850_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2027_ _1246_ _0288_ _0297_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1946__A2 _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1707__I _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1598__B _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2718__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ _0143_ clknet_4_9_0_wb_clk_i simon1.seq_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2645_ _0074_ clknet_4_11_0_wb_clk_i simon1.play1.tick_counter\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1527_ simon1.seq\[13\]\[0\] _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2576_ _0022_ clknet_4_6_0_wb_clk_i simon1.seq\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1389_ _0824_ _0826_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1458_ _0861_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2361_ _0584_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2430_ _1007_ _1171_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2690__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1312_ net3 _0734_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2292_ _1232_ _0515_ _0524_ _0527_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_47_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2628_ _0057_ clknet_4_15_0_wb_clk_i simon1.score1.tens\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2559_ _1131_ _0722_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_65_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1930_ _0208_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1792_ simon1.score1.ones\[1\] _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1861_ simon1.play1.freq\[6\] _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2344_ _0554_ _0556_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2410__B _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2413_ _1098_ _0617_ _0620_ _0384_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2275_ _0509_ _0512_ _0432_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2586__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ _0275_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1913_ _1263_ _1270_ _1276_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1844_ _1205_ _1217_ _1219_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1775_ _1164_ _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2327_ _0822_ _0469_ _0548_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2258_ _0484_ _0491_ _0498_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_67_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2465__A1 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2189_ _0417_ _0418_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__2751__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1560_ _0978_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1491_ _0855_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2112_ simon1.play1.tick_counter\[26\] _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_55_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2043_ simon1.play1.tick_counter\[18\] _0310_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_17_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2119__C _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ _1201_ _1202_ _1204_ _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2624__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1689_ _1104_ _1105_ _1070_ _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1758_ _1067_ _1153_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_67_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2429__A1 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2661_ _0090_ clknet_4_9_0_wb_clk_i simon1.play1.tick_counter\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2647__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2730_ _0159_ clknet_4_2_0_wb_clk_i simon1.seq\[28\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1612_ _0765_ _0779_ _1040_ _0764_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1543_ simon1.millis_counter\[4\] _0816_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2592_ _0009_ clknet_4_4_0_wb_clk_i simon1.state\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1474_ _0889_ _0908_ _0911_ _0905_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_65_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2026_ _1231_ _1238_ _0290_ _0295_ _0296_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_17_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_17_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2644_ _0073_ clknet_4_11_0_wb_clk_i simon1.play1.tick_counter\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2713_ _0142_ clknet_4_1_0_wb_clk_i simon1.seq_length\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1971__C _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2575_ _0021_ clknet_4_1_0_wb_clk_i simon1.seq\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1526_ simon1.seq\[14\]\[0\] simon1.seq\[15\]\[0\] _0894_ _0964_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1457_ _0894_ simon1.seq\[0\]\[1\] _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1388_ simon1.tone_sequence_counter\[2\] _0825_ simon1.tone_sequence_counter\[1\]
+ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2009_ simon1.play1.tick_counter\[13\] _0271_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2041__A2 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1311_ _0752_ _0746_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2291_ _0484_ _0518_ _0525_ _0526_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2360_ _0991_ _0549_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2627_ _0056_ clknet_4_14_0_wb_clk_i simon1.score1.tens\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_34_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1509_ _0929_ simon1.seq\[20\]\[0\] _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2489_ _0677_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2558_ _0678_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_43_Left_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2708__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_52_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1860_ simon1.play1.freq\[7\] _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_44_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1791_ _1175_ _1176_ _1178_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2343_ _0563_ _0570_ _0571_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_58_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2274_ _0496_ _0452_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2412_ _1098_ _0619_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1989_ _0261_ _0262_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output11_I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2680__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1912_ _1278_ _1285_ _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1843_ _1212_ _1218_ _1210_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1774_ _1161_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2140__C _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2257_ _0468_ _0494_ _0495_ _0496_ _0411_ _0497_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_2326_ _0552_ _0553_ _0558_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2188_ _0418_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_55_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2153__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1636__I _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1490_ simon1.seq\[25\]\[0\] _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2042_ _1267_ _1259_ _0278_ _0293_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2111_ _0370_ _0371_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2576__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1826_ simon1.play1.freq\[1\] simon1.play1.tick_counter\[1\] _1204_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1688_ _1052_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_9_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1757_ _1068_ _1152_ _1111_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_2309_ simon1.tick_counter\[1\] _0542_ simon1.tick_counter\[2\] simon1.tick_counter\[3\]
+ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2599__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1611_ _0780_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ _0089_ clknet_4_3_0_wb_clk_i simon1.play1.tick_counter\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_14_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1542_ simon1.millis_counter\[7\] simon1.millis_counter\[6\] _0980_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2591_ _0008_ clknet_4_7_0_wb_clk_i simon1.state\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1473_ _0892_ _0909_ _0910_ _0896_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input2_I io_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2025_ _0290_ _0295_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1809_ _1189_ _1191_ _1190_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2741__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2614__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2338__A1 _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2643_ _0072_ clknet_4_11_0_wb_clk_i simon1.play1.tick_counter\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2712_ _0141_ clknet_4_1_0_wb_clk_i simon1.seq_length\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2574_ _0020_ clknet_4_6_0_wb_clk_i simon1.seq\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1387_ simon1.tone_sequence_counter\[0\] _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1456_ _0852_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1525_ _0874_ _0957_ _0962_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2008_ _0278_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2329__A1 _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1552__A2 _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2637__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1310_ simon1.score1.ones\[1\] simon1.score1.tens\[1\] _0745_ _0752_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2290_ _1023_ _0453_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2475__I _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1819__I _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2559__A1 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2626_ _0055_ clknet_4_14_0_wb_clk_i simon1.score1.ones\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ _0721_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2488_ _0673_ simon1.seq\[2\]\[1\] _0675_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1508_ simon1.seq\[21\]\[0\] _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1439_ simon1.seq\[17\]\[1\] _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_65_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2318__C _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1464__I _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1790_ _1177_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ _0618_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2342_ simon1.millis_counter\[5\] _0569_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2273_ _0489_ _0511_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1988_ _1254_ _0251_ _0259_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2609_ _0047_ clknet_4_6_0_wb_clk_i _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1911_ _1279_ _1284_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1842_ _1209_ simon1.play1.tick_counter\[3\] _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1773_ _0836_ _1162_ _1165_ _1166_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2187_ _0415_ _0432_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2256_ _0408_ _1157_ _1053_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2325_ simon1.millis_counter\[1\] _0550_ _0557_ _1027_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_63_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2041_ _1258_ _0276_ _0309_ _0287_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2110_ _0362_ _0288_ _0992_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_60_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1825_ _1201_ _1202_ _1203_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1756_ _1069_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2308_ simon1.tick_counter\[0\] _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1687_ _0990_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2670__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2239_ _1001_ _0480_ _0417_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2126__A2 _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1610_ _0743_ _0751_ _0756_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_54_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2590_ _0007_ clknet_4_7_0_wb_clk_i simon1.state\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1541_ simon1.state\[5\] _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2478__I _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1472_ _0902_ simon1.seq\[12\]\[1\] _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2693__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2024_ _0291_ _0294_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1808_ simon1.score1.tens\[3\] _0738_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1739_ _1063_ _1066_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2337__B _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2247__B _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1930__I _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2711_ _0140_ clknet_4_3_0_wb_clk_i simon1.seq_length\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2642_ _0071_ clknet_4_11_0_wb_clk_i simon1.play1.tick_counter\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2573_ _0019_ clknet_4_6_0_wb_clk_i simon1.seq\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1524_ _0913_ _0958_ _0961_ _0905_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1386_ simon1.millis_counter\[1\] _0819_ _0820_ _0823_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__1840__I _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1455_ simon1.seq\[1\]\[1\] _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2007_ _1247_ _0278_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_26_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2589__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2265__A1 _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2731__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2625_ _0054_ clknet_4_14_0_wb_clk_i simon1.score1.ones\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1507_ simon1.seq\[22\]\[0\] simon1.seq\[23\]\[0\] _0868_ _0945_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2487_ _0676_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2556_ _0700_ simon1.seq\[17\]\[1\] _0719_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1369_ simon1.state\[7\] _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_38_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1438_ simon1.seq\[18\]\[1\] simon1.seq\[19\]\[1\] _0853_ _0876_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2604__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2754__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2341_ simon1.millis_counter\[5\] _0569_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2410_ _0792_ _1159_ _0987_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_3_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2272_ _1236_ _0487_ _0510_ _0452_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2627__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1987_ _0259_ _1254_ _0240_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2608_ _0046_ clknet_4_3_0_wb_clk_i _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2539_ simon1.seq\[29\]\[0\] _0705_ _0710_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_58_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2345__B _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1910_ _1220_ _1280_ _1283_ _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1682__A2 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1841_ _1206_ _1208_ _1210_ _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1772_ _0988_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2324_ _0426_ _0554_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2186_ _0431_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2255_ _1022_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ _0303_ _0305_ _0308_ _0219_ _1240_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_60_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1824_ _1201_ _1202_ _1199_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1755_ _1151_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1686_ _1103_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2238_ _0800_ _0793_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2307_ _0540_ simon1.tick_counter\[5\] simon1.tick_counter\[6\] simon1.tick_counter\[7\]
+ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_2169_ simon1.tone_sequence_counter\[2\] _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1540_ _0924_ _0977_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1471_ simon1.seq\[13\]\[1\] _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_65_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2023_ _0280_ _0293_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_15_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1807_ simon1.score1.tens\[1\] _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1738_ _1140_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1669_ simon1.seq_length\[3\] _1065_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__A2 _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2710_ _0139_ clknet_4_3_0_wb_clk_i simon1.seq_length\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2641_ _0070_ clknet_4_11_0_wb_clk_i simon1.play1.tick_counter\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2660__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1454_ _0856_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1523_ _0915_ _0959_ _0960_ _0918_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2572_ _0018_ clknet_4_1_0_wb_clk_i simon1.seq\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1385_ _0821_ _0797_ _0822_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_65_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1996__C _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2006_ _0277_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1785__A1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2683__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2624_ _0053_ clknet_4_15_0_wb_clk_i simon1.score1.ones\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2555_ _0720_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2486_ _0670_ simon1.seq\[2\]\[0\] _0675_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1437_ _0865_ _0873_ _0874_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1506_ _0925_ _0940_ _0943_ _0864_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1299_ _0740_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1368_ simon1.state\[0\] _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_38_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1758__A1 _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2340_ _0567_ _0568_ _0569_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2271_ _0486_ _0509_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2579__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1986_ _0197_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2607_ _0045_ clknet_4_2_0_wb_clk_i simon1.seq\[21\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2469_ net10 _0633_ _0661_ _0663_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1912__A1 _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2538_ _1067_ _0678_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2721__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1840_ _1031_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1771_ _0836_ _1164_ _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2254_ _0440_ _0452_ _0434_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2323_ _0555_ _1052_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2185_ simon1.tone_sequence_counter\[1\] _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ _0243_ _0244_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2744__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2091__B _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2617__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1823_ simon1.play1.freq\[1\] simon1.play1.tick_counter\[1\] _1202_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1754_ _1139_ simon1.seq\[3\]\[1\] _1149_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1685_ _1086_ simon1.seq\[10\]\[1\] _1101_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2306_ simon1.tick_counter\[4\] _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2237_ _0407_ _0479_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2168_ _0825_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2099_ _0353_ _0359_ _0360_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1470_ simon1.seq\[14\]\[1\] simon1.seq\[15\]\[1\] _0890_ _0908_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_59_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2022_ _0292_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1806_ _1128_ _1187_ _1189_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1599_ _0787_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1668_ simon1.seq_length\[2\] _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1737_ _1139_ simon1.seq\[6\]\[1\] _1137_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_28_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2504__A1 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2640_ _0069_ clknet_4_11_0_wb_clk_i simon1.play1.tick_counter\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1453_ simon1.seq\[2\]\[1\] simon1.seq\[3\]\[1\] _0890_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1522_ _0954_ simon1.seq\[4\]\[0\] _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2571_ _0017_ clknet_4_1_0_wb_clk_i simon1.seq\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1384_ simon1.millis_counter\[2\] _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2005_ _0270_ _0258_ _1254_ _0239_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_26_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2623_ _0052_ clknet_4_14_0_wb_clk_i simon1.score1.ones\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2554_ _0697_ simon1.seq\[17\]\[0\] _0719_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1367_ _0794_ _0796_ _0802_ _0805_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_50_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2485_ _1100_ _1148_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1505_ _0927_ _0941_ _0942_ _0931_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1436_ _0003_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1298_ simon1.score1.ones\[2\] _0735_ _0739_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_38_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1758__A2 _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2650__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2270_ _0454_ _0508_ _0468_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1985_ _0258_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2537_ _0709_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2606_ _0044_ clknet_4_0_0_wb_clk_i simon1.seq\[21\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2468_ _0634_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2399_ simon1.tick_counter\[12\] _0609_ _0602_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2673__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1419_ _0856_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2156__A2 _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1770_ _1161_ _1163_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2696__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2184_ _0415_ _0429_ _0430_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2253_ _0436_ _0492_ _0493_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2322_ _1159_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_34_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_25_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1830__A1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1968_ _0195_ _0235_ _0241_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_31_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1899_ simon1.play1.tick_counter\[24\] _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2569__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1822_ simon1.play1.freq\[0\] simon1.play1.tick_counter\[0\] _1201_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1753_ _1150_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1684_ _1102_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2305_ _0536_ _0538_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2236_ simon1.play1.freq\[1\] _0448_ _0478_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2167_ _0413_ _0414_ _0989_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2711__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2098_ _0353_ _0359_ _0208_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2021_ simon1.play1.tick_counter\[15\] simon1.play1.tick_counter\[14\] _0292_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2734__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1805_ _1188_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1736_ _1085_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1598_ _1020_ _1030_ _0989_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1667_ simon1.seq_length\[4\] _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2219_ _0923_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2607__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2570_ _0016_ clknet_4_4_0_wb_clk_i simon1.seq\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1383_ simon1.millis_counter\[0\] _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1452_ _0855_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1521_ simon1.seq\[5\]\[0\] _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2004_ _0275_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2431__A1 _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2699_ _0128_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1719_ _1086_ simon1.seq\[8\]\[1\] _1125_ _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2498__A1 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2622_ _0051_ clknet_4_12_0_wb_clk_i simon1.score_rst vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_30_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1504_ _0929_ simon1.seq\[16\]\[0\] _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2553_ _1141_ _1112_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1366_ _0803_ _0804_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2484_ _0674_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1435_ _0851_ _0866_ _0870_ _0872_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1297_ _0738_ _0735_ simon1.score1.ena _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1984_ simon1.play1.tick_counter\[12\] _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2467_ _0404_ _0422_ _0638_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2536_ simon1.seq\[22\]\[1\] _0708_ _0706_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2605_ _0043_ clknet_4_0_0_wb_clk_i simon1.seq\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2398_ simon1.tick_counter\[12\] _0609_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1349_ _0787_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1418_ _0855_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2321_ _0807_ _0809_ _0812_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2183_ _0415_ _0427_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2252_ _0798_ _0800_ _0794_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_18_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1967_ _0197_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1898_ simon1.play1.tick_counter\[30\] _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_28_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2640__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2519_ _1079_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_54_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1783__I _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2663__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1821_ _1198_ simon1.play1.tick_counter\[0\] _1200_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1752_ _1136_ simon1.seq\[3\]\[0\] _1149_ _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1683_ _1080_ simon1.seq\[10\]\[0\] _1101_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2304_ _0993_ _1105_ _0426_ _0537_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2235_ _0461_ _0467_ _0477_ _0457_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2166_ _1074_ simon1.next_random\[0\] _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2097_ _0357_ _0358_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_51_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1552__B _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2686__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2020_ _1247_ _0280_ _1246_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1804_ simon1.score1.tens\[0\] _1185_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1735_ _1138_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1666_ _1087_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1597_ _1023_ _1024_ _1025_ _1029_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2149_ net11 _0194_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2218_ _0460_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_36_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1951__A1 simon1.play1.freq\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1520_ simon1.seq\[6\]\[0\] simon1.seq\[7\]\[0\] _0894_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1382_ simon1.millis_counter\[9\] simon1.millis_counter\[8\] _0820_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2701__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1451_ _0850_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2003_ _0197_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2698_ _0127_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1649_ _1073_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1718_ _1126_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2724__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_30_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2621_ _0014_ clknet_4_15_0_wb_clk_i net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2552_ _0718_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2483_ _0673_ simon1.seq\[20\]\[1\] _0671_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1503_ simon1.seq\[17\]\[0\] _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1365_ simon1.millis_counter\[6\] _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1296_ simon1.score1.tens\[2\] _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_38_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1434_ _0871_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2747__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1983_ _0248_ _0249_ _0257_ _1166_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_7_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2604_ _0042_ clknet_4_0_0_wb_clk_i simon1.seq\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2466_ _0648_ _0655_ _0645_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2535_ _1076_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1417_ _0000_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2397_ _0597_ _0608_ _0609_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1348_ net6 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2251_ _0799_ _0480_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2320_ _0469_ _0549_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2182_ _0809_ _1023_ _0428_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2592__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1966_ _0195_ _0235_ _0241_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1897_ simon1.play1.tick_counter\[31\] _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2449_ _0555_ _0999_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2543__A1 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ _0696_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_54_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1820_ _1198_ simon1.play1.tick_counter\[0\] _1199_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1682_ _1091_ _1100_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1751_ _1094_ _1148_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2303_ _1010_ _0435_ _0442_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2234_ _0468_ _0472_ _0473_ _0474_ _0476_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_29_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_51_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2165_ simon1.next_random\[1\] _1048_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2096_ _0320_ _0347_ _0349_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_63_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1949_ _1232_ _1250_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2630__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1803_ simon1.score1.tens\[0\] _1185_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1596_ _1028_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1734_ _1136_ simon1.seq\[6\]\[0\] _1137_ _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1665_ _1086_ simon1.seq\[12\]\[1\] _1083_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2217_ _1051_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_37_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_46_Left_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2148_ _0288_ _0402_ _1271_ _0384_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_36_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2079_ _1240_ _0342_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_55_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2653__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1450_ _0875_ _0887_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1381_ _0818_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1920__C _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2002_ _0270_ _0249_ _0274_ _1166_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_33_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1579_ net4 net1 _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2697_ _0126_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1648_ simon1.seq\[13\]\[0\] _1061_ _1072_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1717_ _1080_ simon1.seq\[8\]\[0\] _1125_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2676__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1630__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2110__A2 _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2620_ _0013_ clknet_4_15_0_wb_clk_i net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2699__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2551_ simon1.seq\[25\]\[1\] _0708_ _0716_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2482_ _1085_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1433_ _0002_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1502_ simon1.seq\[18\]\[0\] simon1.seq\[19\]\[0\] _0859_ _0940_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1364_ simon1.millis_counter\[7\] _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1295_ simon1.score1.ones\[1\] _0735_ _0736_ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1931__B _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2749_ _0178_ clknet_4_2_0_wb_clk_i simon1.seq\[25\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2159__A2 _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1982_ _0250_ _0255_ _0256_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2534_ _0707_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2603_ _0041_ clknet_4_1_0_wb_clk_i simon1.seq\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1347_ _0786_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2465_ _0630_ _0660_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2396_ simon1.tick_counter\[11\] _0606_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1416_ simon1.seq\[26\]\[1\] simon1.seq\[27\]\[1\] _0853_ _0854_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2714__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2250_ _0462_ _0490_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2001__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2181_ _0427_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2737__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1965_ _0234_ _0240_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1896_ _1265_ _1269_ _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2543__A2 _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2517_ _0673_ simon1.seq\[1\]\[1\] _0694_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2448_ _0639_ _0637_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2379_ _0587_ _0595_ _0596_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1806__A1 _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2298__A1 simon1.play1.freq\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2470__A1 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1750_ _1088_ _1110_ _1089_ _1070_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XPHY_EDGE_ROW_29_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1681_ _1098_ _1099_ _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2233_ _0450_ _0475_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2302_ _1157_ _0535_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2164_ _0407_ simon1.next_random\[0\] _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_51_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2095_ simon1.play1.tick_counter\[24\] _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1948_ _1278_ _0218_ _0220_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1879_ _1246_ _1252_ simon1.play1.tick_counter\[13\] simon1.play1.tick_counter\[12\]
+ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_8_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2582__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1802_ _1175_ _1185_ _1186_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1733_ _1100_ _1132_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1595_ _1027_ _1002_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1664_ _1085_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2216_ _0407_ _0459_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2147_ _0394_ _0401_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2078_ _0219_ _0338_ _0333_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1380_ simon1.millis_counter\[4\] _0816_ simon1.millis_counter\[7\] _0817_ _0818_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2001_ _0260_ _0273_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2416__A1 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2696_ _0125_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1716_ _1109_ _1091_ _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1578_ net4 net1 _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1647_ _1067_ _1071_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_49_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_24_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2620__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1385__A1 _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2550_ _0717_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1363_ _0799_ _0800_ _0801_ simon1.millis_counter\[5\] _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2481_ _0672_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1432_ _0857_ _0867_ _0869_ _0862_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1501_ _0933_ _0938_ _0874_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1294_ simon1.score1.tens\[1\] _0731_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_58_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1376__A1 _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2679_ _0108_ clknet_4_12_0_wb_clk_i simon1.play1.freq\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2643__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2748_ _0177_ clknet_4_2_0_wb_clk_i simon1.seq\[23\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2002__C _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2666__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1981_ _0250_ _0255_ _0208_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2533_ simon1.seq\[22\]\[0\] _0705_ _0706_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2602_ _0040_ clknet_4_1_0_wb_clk_i simon1.seq\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1346_ _0776_ _0782_ _0785_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2464_ net9 _0633_ _0656_ _0659_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2395_ simon1.tick_counter\[11\] _0606_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1415_ _0852_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_65_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1597__A1 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2013__B _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2689__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2180_ _0990_ _0424_ _0425_ _0426_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_20_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ _0239_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1895_ _1260_ _1266_ _1268_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_31_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2447_ _0631_ _0633_ _0641_ _0644_ _1031_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_11_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2516_ _0695_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1751__A1 _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1329_ _0765_ _0763_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2378_ simon1.tick_counter\[6\] _0593_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_3_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2301_ _1010_ _1034_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2704__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1680_ _1062_ _1092_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1733__A1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2163_ net4 net5 _1019_ _0412_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2232_ _0451_ _0431_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2100__C _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2094_ _1216_ _0356_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1947_ _0202_ _0222_ _0224_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1878_ _1247_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_28_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2727__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1801_ _0730_ _1183_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1663_ _1075_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1732_ _1079_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1594_ _1026_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2215_ _1198_ _0448_ _0458_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2146_ _1272_ _0397_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2131__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2077_ _0340_ _0341_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2000_ simon1.play1.tick_counter\[13\] _0271_ _0272_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_45_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2695_ _0124_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1646_ _0830_ _1068_ _1069_ _1070_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1715_ _1124_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1577_ _1009_ _1010_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2129_ _0368_ _0382_ _0386_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2572__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2480_ _0670_ simon1.seq\[20\]\[0\] _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1500_ _0925_ _0934_ _0937_ _0872_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1293_ simon1.score1.active_digit _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1362_ simon1.millis_counter\[4\] _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2595__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1431_ _0868_ simon1.seq\[28\]\[1\] _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2678_ _0107_ clknet_4_12_0_wb_clk_i simon1.play1.freq\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1629_ simon1.state\[6\] simon1.state\[7\] _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_41_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2747_ _0176_ clknet_4_2_0_wb_clk_i simon1.seq\[23\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2564__A1 _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2316__A1 _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1980_ _0252_ _0254_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2463_ _0634_ _0658_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2532_ _1121_ _1153_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2601_ _0039_ clknet_4_1_0_wb_clk_i simon1.seq\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1345_ _0761_ _0783_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2394_ _0597_ _0606_ _0607_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_3_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1414_ _0000_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2610__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_57_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2633__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1963_ _0228_ _0237_ _0238_ _0217_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1894_ _1262_ _1267_ simon1.play1.tick_counter\[10\] _1248_ _1268_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2446_ _0636_ _0643_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_11_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2515_ _0670_ simon1.seq\[1\]\[0\] _0694_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1328_ _0752_ _0750_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2377_ simon1.tick_counter\[6\] _0593_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_54_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2656__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2231_ _1157_ _1053_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2300_ _1025_ _1003_ _1026_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2162_ _0411_ _1018_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2093_ simon1.play1.tick_counter\[23\] _0209_ _0353_ _0355_ _0356_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_61_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1877_ simon1.play1.tick_counter\[11\] simon1.play1.tick_counter\[9\] _1250_ _1251_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1946_ _1250_ _0209_ _0223_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2679__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2429_ _0630_ _1170_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1660__A1 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2140__A2 _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1800_ simon1.score1.ones\[1\] _1184_ _1180_ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1731_ _1135_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1662_ _1084_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2214_ _0450_ _0453_ _0456_ _0995_ _0457_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_1593_ _1000_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2145_ _1272_ _0243_ _0399_ _0400_ _0390_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2076_ _1243_ _0288_ _0992_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1929_ _0200_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_33_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_42_Left_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2694_ _0123_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1576_ _0984_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1645_ _1057_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1714_ simon1.seq\[14\]\[1\] _1119_ _1122_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2717__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2059_ simon1.play1.tick_counter\[20\] _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2128_ _0385_ _0380_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2016__C _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1430_ _0852_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1292_ _0733_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1361_ simon1.millis_counter\[2\] _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2746_ _0175_ clknet_4_2_0_wb_clk_i simon1.seq\[29\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1628_ _0983_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2677_ _0106_ clknet_4_12_0_wb_clk_i simon1.play1.freq\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1559_ _0994_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2600_ _0038_ clknet_4_1_0_wb_clk_i simon1.seq\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2462_ _0404_ _0657_ _0638_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2393_ _0604_ _0601_ simon1.tick_counter\[10\] _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2531_ _1060_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1413_ _0850_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1344_ _0779_ _0750_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2729_ _0158_ clknet_4_8_0_wb_clk_i simon1.seq\[28\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2585__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1962_ _0211_ _0228_ _0229_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_34_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ simon1.play1.tick_counter\[17\] _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2376_ _0587_ _0593_ _0594_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_59_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2445_ _1009_ _0464_ _0642_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2514_ _1141_ _1148_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1327_ _0763_ _0764_ _0766_ _0768_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2230_ simon1.user_input\[0\] _0410_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1773__C _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2600__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2161_ _0410_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2092_ _0351_ _0354_ _0201_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2750__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1945_ _0991_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1876_ simon1.play1.tick_counter\[8\] _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2359_ _0583_ _0576_ _0579_ _0795_ _0573_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2428_ _1006_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2623__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1592_ _0849_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1730_ simon1.seq\[7\]\[1\] _1119_ _1133_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1661_ _1080_ simon1.seq\[12\]\[0\] _1083_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2213_ _0447_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2144_ _0394_ _0398_ _0275_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2075_ _0330_ _0334_ _0339_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1859_ simon1.play1.freq\[9\] _1232_ _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1928_ _1286_ _0206_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2646__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xurish_simon_says_80 io_oeb[35] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_45_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2669__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1713_ _1123_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2693_ _0122_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1575_ _1008_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1644_ simon1.seq_length\[2\] _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_6_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2127_ simon1.play1.tick_counter\[28\] _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2058_ _0316_ _0276_ _0324_ _0287_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_44_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1360_ _0798_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1291_ _0730_ _0731_ _0732_ simon1.score1.ena _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2676_ _0105_ clknet_4_12_0_wb_clk_i simon1.play1.freq\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2745_ _0174_ clknet_4_2_0_wb_clk_i simon1.seq\[29\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1558_ _0808_ _0811_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1627_ _0999_ _1050_ _1051_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1489_ _0856_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_61_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2707__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1348__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2530_ _0704_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1343_ _0752_ _0755_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2461_ _0795_ _0421_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2392_ _0604_ simon1.tick_counter\[10\] _0600_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1412_ _0001_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2659_ _0088_ clknet_4_3_0_wb_clk_i simon1.play1.tick_counter\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2728_ _0157_ clknet_4_0_0_wb_clk_i simon1.seq\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1745__A1 _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1961_ _0236_ _0229_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1892_ _1230_ simon1.play1.tick_counter\[5\] simon1.play1.tick_counter\[4\] simon1.play1.tick_counter\[3\]
+ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_43_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2513_ _0693_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1326_ _0754_ _0767_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2375_ simon1.tick_counter\[5\] _0591_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2444_ _0408_ _0410_ _0555_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_19_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1727__A1 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ simon1.user_input\[1\] _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2091_ _0345_ _0338_ _0194_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1957__A1 _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1944_ _0218_ _0221_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1875_ _1248_ _1229_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2427_ _0836_ _1162_ _1165_ _0384_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_24_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2358_ _0422_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1309_ _0744_ _0747_ _0750_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2289_ _0408_ _0411_ _0474_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2575__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1948__A1 _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2035__C _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1591_ _0827_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1660_ _1071_ _1082_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2212_ _0423_ _0455_ _0415_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2143_ _0394_ _0398_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2598__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2074_ _0195_ _0338_ _0201_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1858_ simon1.play1.freq\[8\] _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1927_ _0203_ _0205_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__1975__B _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1789_ simon1.score1.inc simon1.score1.ones\[0\] _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_39_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2740__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xurish_simon_says_81 io_oeb[36] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_70 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2692_ _0121_ clknet_4_7_0_wb_clk_i simon1.millis_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1643_ simon1.seq_length\[3\] _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1712_ simon1.seq\[14\]\[0\] _1116_ _1122_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1574_ simon1.state\[5\] _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2126_ _0379_ _1241_ _0383_ _0384_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2057_ _0260_ _0323_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2613__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2319__A1 _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1290_ simon1.score1.tens\[3\] _0731_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2636__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2675_ _0104_ clknet_4_12_0_wb_clk_i simon1.play1.freq\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1626_ simon1.state\[6\] simon1.state\[7\] simon1.state\[5\] _0815_ _1051_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_41_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2133__C _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2744_ _0173_ clknet_4_2_0_wb_clk_i simon1.seq\[22\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1557_ _0992_ _0993_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1488_ simon1.seq\[26\]\[0\] simon1.seq\[27\]\[0\] _0859_ _0926_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2109_ _0243_ _0366_ _0369_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_64_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2285__I _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2659__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2460_ _0650_ _0655_ _0645_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_21_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1342_ _0743_ _0781_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2391_ _0604_ _0601_ _0605_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1411_ _0848_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1609_ _0778_ _0779_ _0763_ _0780_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2589_ _0006_ clknet_4_7_0_wb_clk_i simon1.state\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2658_ _0087_ clknet_4_9_0_wb_clk_i simon1.play1.tick_counter\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2727_ _0156_ clknet_4_0_0_wb_clk_i simon1.seq\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1960_ _1232_ _1250_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1891_ _1253_ _1264_ _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2443_ _0634_ _0640_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2512_ simon1.seq\[30\]\[1\] _0668_ _0691_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1325_ _0737_ _0747_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2374_ simon1.tick_counter\[5\] _0591_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1732__I _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2090_ _0345_ _0338_ _0352_ _0289_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_61_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1874_ simon1.play1.tick_counter\[7\] _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1943_ _0219_ _0220_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2426_ _0622_ _0629_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_24_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_67_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1308_ _0734_ _0749_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2357_ _0580_ _0582_ _0998_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2288_ _0461_ _0464_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1590_ _1022_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2211_ _0821_ _0454_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2142_ _1272_ _0397_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2073_ _0337_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1788_ simon1.score1.inc simon1.score1.ones\[0\] _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1926_ _1279_ _1284_ _0204_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1857_ _1209_ simon1.play1.freq\[2\] simon1.play1.freq\[1\] _1198_ _1231_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2692__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2409_ _0987_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xurish_simon_says_82 io_oeb[37] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_71 io_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_60 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2691_ _0120_ clknet_4_7_0_wb_clk_i simon1.millis_counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1642_ _1063_ _1066_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_1711_ _1071_ _1121_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1573_ _1006_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2125_ _0789_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2056_ _0317_ _0322_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1909_ _1236_ simon1.play1.tick_counter\[5\] _1282_ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_44_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1839__A1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2264__A1 _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2588__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1915__I _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2743_ _0172_ clknet_4_2_0_wb_clk_i simon1.seq\[22\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1556_ _0807_ _0812_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1625_ _1049_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ _0103_ clknet_4_9_0_wb_clk_i simon1.play1.freq\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1487_ _0850_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2039_ _0307_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2730__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2108_ _0368_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2485__A1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1410_ _0830_ _0834_ _0842_ _0847_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_23_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1341_ _0770_ _0777_ _0781_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2390_ _0604_ _0601_ _0602_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2753__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2603__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1983__C _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2726_ _0155_ clknet_4_2_0_wb_clk_i simon1.seq\[20\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1608_ _0014_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1555__I _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2588_ _0005_ clknet_4_12_0_wb_clk_i simon1.state\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1539_ simon1.user_input\[0\] _0976_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2657_ _0086_ clknet_4_8_0_wb_clk_i simon1.play1.tick_counter\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_40_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2626__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2458__A1 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1890_ simon1.play1.tick_counter\[2\] simon1.play1.tick_counter\[1\] simon1.play1.tick_counter\[0\]
+ _1251_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2373_ _0587_ _0591_ _0592_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2442_ _0405_ _0820_ _0638_ _0639_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_59_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2511_ _0692_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1324_ _0765_ _0744_ _0747_ _0758_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_49_Left_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2649__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2709_ _0138_ clknet_4_3_0_wb_clk_i simon1.seq_length\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_58_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1942_ _0196_ _0206_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_43_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1873_ simon1.play1.tick_counter\[14\] _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2356_ _1025_ _0581_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2425_ _1088_ _0628_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_67_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1307_ _0748_ _0741_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2287_ _0448_ _0521_ _0523_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _0419_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1653__I _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2141_ simon1.play1.tick_counter\[29\] simon1.play1.tick_counter\[28\] _0380_ _0397_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2072_ _0307_ _0328_ _0332_ _0333_ _0336_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_56_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1925_ _1235_ _1229_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1787_ _1128_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1856_ _1229_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2339_ simon1.millis_counter\[4\] _0565_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2408_ _0585_ _0616_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xurish_simon_says_50 io_out[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_72 io_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_61 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2690_ _0119_ clknet_4_5_0_wb_clk_i simon1.millis_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1572_ _0788_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1641_ _1064_ _1065_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1710_ _1064_ _1099_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA_input5_I io_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2124_ _0376_ _0381_ _0382_ _0369_ _1240_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2055_ _0316_ _0318_ _0321_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1908_ _1226_ _1281_ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1839_ _1173_ _1215_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2016__A2 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2682__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2742_ _0171_ clknet_4_8_0_wb_clk_i simon1.seq\[18\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2191__B2 _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1555_ _0991_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1624_ simon1.state\[0\] simon1.state\[3\] simon1.state\[1\] _1049_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2673_ _0102_ clknet_4_9_0_wb_clk_i simon1.play1.freq\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1486_ simon1.user_input\[1\] _0923_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2107_ _0345_ _0337_ _0367_ _0289_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_37_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2038_ _0279_ _0283_ _0305_ _0306_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__2182__A1 _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1340_ _0778_ _0779_ _0780_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2656_ _0085_ clknet_4_9_0_wb_clk_i simon1.play1.tick_counter\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _0154_ clknet_4_1_0_wb_clk_i simon1.seq\[20\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1607_ _1037_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2587_ _0033_ clknet_4_15_0_wb_clk_i simon1.score1.active_digit vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2578__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1469_ _0874_ _0899_ _0906_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1538_ _0004_ _0951_ _0975_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_49_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1969__A1 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2510_ simon1.seq\[30\]\[0\] _0665_ _0691_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2720__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1323_ _0748_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2372_ simon1.tick_counter\[3\] _0588_ simon1.tick_counter\[4\] _0592_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2441_ _0803_ _0442_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2708_ _0137_ clknet_4_5_0_wb_clk_i simon1.tick_counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2639_ _0068_ clknet_4_14_0_wb_clk_i simon1.play1.tick_counter\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_53_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2743__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1872_ simon1.play1.tick_counter\[15\] _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1941_ _1277_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_16_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1306_ net3 _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2286_ _1234_ _0515_ _0522_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2355_ _0986_ _1028_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2424_ _1110_ _0623_ _1130_ _0618_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_19_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2616__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2076__B _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2639__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _0391_ _0326_ _0394_ _0396_ _0390_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2071_ _0325_ _0335_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1924_ simon1.play1.freq\[7\] simon1.play1.tick_counter\[7\] _0203_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1855_ simon1.play1.tick_counter\[6\] _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1786_ _1173_ _1020_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2338_ _0801_ _0565_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2407_ simon1.tick_counter\[15\] _0615_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2269_ _0801_ _0492_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xurish_simon_says_51 io_out[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_73 io_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xurish_simon_says_40 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xurish_simon_says_62 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_38_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1571_ _0998_ _1005_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1640_ _1057_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1664__I _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2123_ _0373_ _0374_ _0381_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_49_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2054_ _0320_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1907_ _1236_ simon1.play1.tick_counter\[5\] _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1838_ _1211_ _1214_ _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1769_ _1026_ _1008_ _0849_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2672_ _0101_ clknet_4_14_0_wb_clk_i simon1.tone_sequence_counter\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2741_ _0170_ clknet_4_3_0_wb_clk_i simon1.seq\[18\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1554_ _0990_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1623_ simon1.next_random\[0\] _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1485_ _0004_ _0888_ _0922_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
.ends

