magic
tech gf180mcuD
magscale 1 10
timestamp 1702277092
<< metal1 >>
rect 1344 56474 158592 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 81278 56474
rect 81330 56422 81382 56474
rect 81434 56422 81486 56474
rect 81538 56422 111998 56474
rect 112050 56422 112102 56474
rect 112154 56422 112206 56474
rect 112258 56422 142718 56474
rect 142770 56422 142822 56474
rect 142874 56422 142926 56474
rect 142978 56422 158592 56474
rect 1344 56388 158592 56422
rect 5070 56306 5122 56318
rect 5070 56242 5122 56254
rect 5854 56306 5906 56318
rect 5854 56242 5906 56254
rect 13470 56306 13522 56318
rect 13470 56242 13522 56254
rect 24894 56306 24946 56318
rect 24894 56242 24946 56254
rect 29710 56306 29762 56318
rect 29710 56242 29762 56254
rect 36318 56306 36370 56318
rect 36318 56242 36370 56254
rect 47742 56306 47794 56318
rect 47742 56242 47794 56254
rect 52558 56306 52610 56318
rect 52558 56242 52610 56254
rect 55358 56306 55410 56318
rect 55358 56242 55410 56254
rect 63982 56306 64034 56318
rect 63982 56242 64034 56254
rect 66782 56306 66834 56318
rect 66782 56242 66834 56254
rect 71598 56306 71650 56318
rect 71598 56242 71650 56254
rect 83022 56306 83074 56318
rect 83022 56242 83074 56254
rect 89630 56306 89682 56318
rect 89630 56242 89682 56254
rect 94446 56306 94498 56318
rect 94446 56242 94498 56254
rect 98254 56306 98306 56318
rect 98254 56242 98306 56254
rect 101054 56306 101106 56318
rect 101054 56242 101106 56254
rect 105870 56306 105922 56318
rect 105870 56242 105922 56254
rect 109678 56306 109730 56318
rect 109678 56242 109730 56254
rect 117294 56306 117346 56318
rect 117294 56242 117346 56254
rect 121102 56306 121154 56318
rect 121102 56242 121154 56254
rect 128718 56306 128770 56318
rect 128718 56242 128770 56254
rect 132526 56306 132578 56318
rect 132526 56242 132578 56254
rect 135326 56306 135378 56318
rect 135326 56242 135378 56254
rect 140142 56306 140194 56318
rect 140142 56242 140194 56254
rect 146750 56306 146802 56318
rect 146750 56242 146802 56254
rect 151566 56306 151618 56318
rect 151566 56242 151618 56254
rect 155374 56306 155426 56318
rect 155374 56242 155426 56254
rect 78206 56194 78258 56206
rect 6178 56142 6190 56194
rect 6242 56142 6254 56194
rect 67106 56142 67118 56194
rect 67170 56142 67182 56194
rect 78206 56130 78258 56142
rect 78542 56194 78594 56206
rect 89954 56142 89966 56194
rect 90018 56142 90030 56194
rect 101378 56142 101390 56194
rect 101442 56142 101454 56194
rect 112466 56142 112478 56194
rect 112530 56142 112542 56194
rect 123890 56142 123902 56194
rect 123954 56142 123966 56194
rect 144498 56142 144510 56194
rect 144562 56142 144574 56194
rect 78542 56130 78594 56142
rect 19842 56030 19854 56082
rect 19906 56030 19918 56082
rect 28690 56030 28702 56082
rect 28754 56030 28766 56082
rect 42690 56030 42702 56082
rect 42754 56030 42766 56082
rect 51538 56030 51550 56082
rect 51602 56030 51614 56082
rect 61730 56030 61742 56082
rect 61794 56030 61806 56082
rect 62962 56030 62974 56082
rect 63026 56030 63038 56082
rect 70578 56030 70590 56082
rect 70642 56030 70654 56082
rect 76962 56030 76974 56082
rect 77026 56030 77038 56082
rect 82002 56030 82014 56082
rect 82066 56030 82078 56082
rect 88386 56030 88398 56082
rect 88450 56030 88462 56082
rect 93426 56030 93438 56082
rect 93490 56030 93502 56082
rect 97570 56030 97582 56082
rect 97634 56030 97646 56082
rect 104850 56030 104862 56082
rect 104914 56030 104926 56082
rect 108658 56030 108670 56082
rect 108722 56030 108734 56082
rect 112690 56030 112702 56082
rect 112754 56030 112766 56082
rect 116274 56030 116286 56082
rect 116338 56030 116350 56082
rect 120082 56030 120094 56082
rect 120146 56030 120158 56082
rect 124114 56030 124126 56082
rect 124178 56030 124190 56082
rect 127698 56030 127710 56082
rect 127762 56030 127774 56082
rect 131506 56030 131518 56082
rect 131570 56030 131582 56082
rect 139234 56030 139246 56082
rect 139298 56030 139310 56082
rect 142930 56030 142942 56082
rect 142994 56030 143006 56082
rect 150770 56030 150782 56082
rect 150834 56030 150846 56082
rect 154578 56030 154590 56082
rect 154642 56030 154654 56082
rect 17502 55970 17554 55982
rect 17502 55906 17554 55918
rect 20974 55970 21026 55982
rect 20974 55906 21026 55918
rect 40350 55970 40402 55982
rect 40350 55906 40402 55918
rect 43822 55970 43874 55982
rect 43822 55906 43874 55918
rect 55918 55970 55970 55982
rect 55918 55906 55970 55918
rect 59390 55970 59442 55982
rect 59390 55906 59442 55918
rect 74622 55970 74674 55982
rect 74622 55906 74674 55918
rect 86046 55970 86098 55982
rect 149774 55970 149826 55982
rect 135762 55918 135774 55970
rect 135826 55918 135838 55970
rect 147186 55918 147198 55970
rect 147250 55918 147262 55970
rect 86046 55906 86098 55918
rect 149774 55906 149826 55918
rect 1344 55690 158592 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 96638 55690
rect 96690 55638 96742 55690
rect 96794 55638 96846 55690
rect 96898 55638 127358 55690
rect 127410 55638 127462 55690
rect 127514 55638 127566 55690
rect 127618 55638 158078 55690
rect 158130 55638 158182 55690
rect 158234 55638 158286 55690
rect 158338 55638 158592 55690
rect 1344 55604 158592 55638
rect 28366 55522 28418 55534
rect 28366 55458 28418 55470
rect 50094 55410 50146 55422
rect 50094 55346 50146 55358
rect 55134 55410 55186 55422
rect 55134 55346 55186 55358
rect 61294 55410 61346 55422
rect 61294 55346 61346 55358
rect 66558 55410 66610 55422
rect 66558 55346 66610 55358
rect 77982 55410 78034 55422
rect 77982 55346 78034 55358
rect 89406 55410 89458 55422
rect 89406 55346 89458 55358
rect 100830 55410 100882 55422
rect 100830 55346 100882 55358
rect 112254 55410 112306 55422
rect 112254 55346 112306 55358
rect 123678 55410 123730 55422
rect 123678 55346 123730 55358
rect 135102 55410 135154 55422
rect 135102 55346 135154 55358
rect 146862 55410 146914 55422
rect 146862 55346 146914 55358
rect 60510 55298 60562 55310
rect 60510 55234 60562 55246
rect 60958 55298 61010 55310
rect 60958 55234 61010 55246
rect 62190 55298 62242 55310
rect 62190 55234 62242 55246
rect 69806 55298 69858 55310
rect 71038 55298 71090 55310
rect 115726 55298 115778 55310
rect 70130 55246 70142 55298
rect 70194 55246 70206 55298
rect 81554 55246 81566 55298
rect 81618 55246 81630 55298
rect 92978 55246 92990 55298
rect 93042 55246 93054 55298
rect 69806 55234 69858 55246
rect 71038 55234 71090 55246
rect 115726 55234 115778 55246
rect 115950 55298 116002 55310
rect 127250 55246 127262 55298
rect 127314 55246 127326 55298
rect 139010 55246 139022 55298
rect 139074 55246 139086 55298
rect 115950 55234 116002 55246
rect 28478 55186 28530 55198
rect 28478 55122 28530 55134
rect 49982 55186 50034 55198
rect 49982 55122 50034 55134
rect 70366 55186 70418 55198
rect 71486 55186 71538 55198
rect 70690 55134 70702 55186
rect 70754 55134 70766 55186
rect 70366 55122 70418 55134
rect 71486 55122 71538 55134
rect 81118 55186 81170 55198
rect 81118 55122 81170 55134
rect 81790 55186 81842 55198
rect 81790 55122 81842 55134
rect 92542 55186 92594 55198
rect 92542 55122 92594 55134
rect 93214 55186 93266 55198
rect 93214 55122 93266 55134
rect 103966 55186 104018 55198
rect 103966 55122 104018 55134
rect 104302 55186 104354 55198
rect 104302 55122 104354 55134
rect 104638 55186 104690 55198
rect 104638 55122 104690 55134
rect 116510 55186 116562 55198
rect 116510 55122 116562 55134
rect 126814 55186 126866 55198
rect 126814 55122 126866 55134
rect 127486 55186 127538 55198
rect 127486 55122 127538 55134
rect 138350 55186 138402 55198
rect 138350 55122 138402 55134
rect 139246 55186 139298 55198
rect 139246 55122 139298 55134
rect 27918 55074 27970 55086
rect 27918 55010 27970 55022
rect 28366 55074 28418 55086
rect 28366 55010 28418 55022
rect 29374 55074 29426 55086
rect 29374 55010 29426 55022
rect 49646 55074 49698 55086
rect 49646 55010 49698 55022
rect 59950 55074 60002 55086
rect 59950 55010 60002 55022
rect 61742 55074 61794 55086
rect 61742 55010 61794 55022
rect 77198 55074 77250 55086
rect 77198 55010 77250 55022
rect 88622 55074 88674 55086
rect 88622 55010 88674 55022
rect 96910 55074 96962 55086
rect 96910 55010 96962 55022
rect 108334 55074 108386 55086
rect 108334 55010 108386 55022
rect 119758 55074 119810 55086
rect 119758 55010 119810 55022
rect 131182 55074 131234 55086
rect 131182 55010 131234 55022
rect 142606 55074 142658 55086
rect 142606 55010 142658 55022
rect 154030 55074 154082 55086
rect 154030 55010 154082 55022
rect 1344 54906 158592 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 81278 54906
rect 81330 54854 81382 54906
rect 81434 54854 81486 54906
rect 81538 54854 111998 54906
rect 112050 54854 112102 54906
rect 112154 54854 112206 54906
rect 112258 54854 142718 54906
rect 142770 54854 142822 54906
rect 142874 54854 142926 54906
rect 142978 54854 158592 54906
rect 1344 54820 158592 54854
rect 116062 54738 116114 54750
rect 116062 54674 116114 54686
rect 115826 54462 115838 54514
rect 115890 54462 115902 54514
rect 116622 54402 116674 54414
rect 116622 54338 116674 54350
rect 1344 54122 158592 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 96638 54122
rect 96690 54070 96742 54122
rect 96794 54070 96846 54122
rect 96898 54070 127358 54122
rect 127410 54070 127462 54122
rect 127514 54070 127566 54122
rect 127618 54070 158078 54122
rect 158130 54070 158182 54122
rect 158234 54070 158286 54122
rect 158338 54070 158592 54122
rect 1344 54036 158592 54070
rect 1344 53338 158592 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 81278 53338
rect 81330 53286 81382 53338
rect 81434 53286 81486 53338
rect 81538 53286 111998 53338
rect 112050 53286 112102 53338
rect 112154 53286 112206 53338
rect 112258 53286 142718 53338
rect 142770 53286 142822 53338
rect 142874 53286 142926 53338
rect 142978 53286 158592 53338
rect 1344 53252 158592 53286
rect 1344 52554 158592 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 96638 52554
rect 96690 52502 96742 52554
rect 96794 52502 96846 52554
rect 96898 52502 127358 52554
rect 127410 52502 127462 52554
rect 127514 52502 127566 52554
rect 127618 52502 158078 52554
rect 158130 52502 158182 52554
rect 158234 52502 158286 52554
rect 158338 52502 158592 52554
rect 1344 52468 158592 52502
rect 1344 51770 158592 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 81278 51770
rect 81330 51718 81382 51770
rect 81434 51718 81486 51770
rect 81538 51718 111998 51770
rect 112050 51718 112102 51770
rect 112154 51718 112206 51770
rect 112258 51718 142718 51770
rect 142770 51718 142822 51770
rect 142874 51718 142926 51770
rect 142978 51718 158592 51770
rect 1344 51684 158592 51718
rect 1344 50986 158592 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 96638 50986
rect 96690 50934 96742 50986
rect 96794 50934 96846 50986
rect 96898 50934 127358 50986
rect 127410 50934 127462 50986
rect 127514 50934 127566 50986
rect 127618 50934 158078 50986
rect 158130 50934 158182 50986
rect 158234 50934 158286 50986
rect 158338 50934 158592 50986
rect 1344 50900 158592 50934
rect 1344 50202 158592 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 81278 50202
rect 81330 50150 81382 50202
rect 81434 50150 81486 50202
rect 81538 50150 111998 50202
rect 112050 50150 112102 50202
rect 112154 50150 112206 50202
rect 112258 50150 142718 50202
rect 142770 50150 142822 50202
rect 142874 50150 142926 50202
rect 142978 50150 158592 50202
rect 1344 50116 158592 50150
rect 1344 49418 158592 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 96638 49418
rect 96690 49366 96742 49418
rect 96794 49366 96846 49418
rect 96898 49366 127358 49418
rect 127410 49366 127462 49418
rect 127514 49366 127566 49418
rect 127618 49366 158078 49418
rect 158130 49366 158182 49418
rect 158234 49366 158286 49418
rect 158338 49366 158592 49418
rect 1344 49332 158592 49366
rect 1344 48634 158592 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 81278 48634
rect 81330 48582 81382 48634
rect 81434 48582 81486 48634
rect 81538 48582 111998 48634
rect 112050 48582 112102 48634
rect 112154 48582 112206 48634
rect 112258 48582 142718 48634
rect 142770 48582 142822 48634
rect 142874 48582 142926 48634
rect 142978 48582 158592 48634
rect 1344 48548 158592 48582
rect 1344 47850 158592 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 96638 47850
rect 96690 47798 96742 47850
rect 96794 47798 96846 47850
rect 96898 47798 127358 47850
rect 127410 47798 127462 47850
rect 127514 47798 127566 47850
rect 127618 47798 158078 47850
rect 158130 47798 158182 47850
rect 158234 47798 158286 47850
rect 158338 47798 158592 47850
rect 1344 47764 158592 47798
rect 1344 47066 158592 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 81278 47066
rect 81330 47014 81382 47066
rect 81434 47014 81486 47066
rect 81538 47014 111998 47066
rect 112050 47014 112102 47066
rect 112154 47014 112206 47066
rect 112258 47014 142718 47066
rect 142770 47014 142822 47066
rect 142874 47014 142926 47066
rect 142978 47014 158592 47066
rect 1344 46980 158592 47014
rect 1344 46282 158592 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 96638 46282
rect 96690 46230 96742 46282
rect 96794 46230 96846 46282
rect 96898 46230 127358 46282
rect 127410 46230 127462 46282
rect 127514 46230 127566 46282
rect 127618 46230 158078 46282
rect 158130 46230 158182 46282
rect 158234 46230 158286 46282
rect 158338 46230 158592 46282
rect 1344 46196 158592 46230
rect 1344 45498 158592 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 81278 45498
rect 81330 45446 81382 45498
rect 81434 45446 81486 45498
rect 81538 45446 111998 45498
rect 112050 45446 112102 45498
rect 112154 45446 112206 45498
rect 112258 45446 142718 45498
rect 142770 45446 142822 45498
rect 142874 45446 142926 45498
rect 142978 45446 158592 45498
rect 1344 45412 158592 45446
rect 1344 44714 158592 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 96638 44714
rect 96690 44662 96742 44714
rect 96794 44662 96846 44714
rect 96898 44662 127358 44714
rect 127410 44662 127462 44714
rect 127514 44662 127566 44714
rect 127618 44662 158078 44714
rect 158130 44662 158182 44714
rect 158234 44662 158286 44714
rect 158338 44662 158592 44714
rect 1344 44628 158592 44662
rect 1344 43930 158592 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 81278 43930
rect 81330 43878 81382 43930
rect 81434 43878 81486 43930
rect 81538 43878 111998 43930
rect 112050 43878 112102 43930
rect 112154 43878 112206 43930
rect 112258 43878 142718 43930
rect 142770 43878 142822 43930
rect 142874 43878 142926 43930
rect 142978 43878 158592 43930
rect 1344 43844 158592 43878
rect 1344 43146 158592 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 96638 43146
rect 96690 43094 96742 43146
rect 96794 43094 96846 43146
rect 96898 43094 127358 43146
rect 127410 43094 127462 43146
rect 127514 43094 127566 43146
rect 127618 43094 158078 43146
rect 158130 43094 158182 43146
rect 158234 43094 158286 43146
rect 158338 43094 158592 43146
rect 1344 43060 158592 43094
rect 1344 42362 158592 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 81278 42362
rect 81330 42310 81382 42362
rect 81434 42310 81486 42362
rect 81538 42310 111998 42362
rect 112050 42310 112102 42362
rect 112154 42310 112206 42362
rect 112258 42310 142718 42362
rect 142770 42310 142822 42362
rect 142874 42310 142926 42362
rect 142978 42310 158592 42362
rect 1344 42276 158592 42310
rect 1344 41578 158592 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 96638 41578
rect 96690 41526 96742 41578
rect 96794 41526 96846 41578
rect 96898 41526 127358 41578
rect 127410 41526 127462 41578
rect 127514 41526 127566 41578
rect 127618 41526 158078 41578
rect 158130 41526 158182 41578
rect 158234 41526 158286 41578
rect 158338 41526 158592 41578
rect 1344 41492 158592 41526
rect 1344 40794 158592 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 81278 40794
rect 81330 40742 81382 40794
rect 81434 40742 81486 40794
rect 81538 40742 111998 40794
rect 112050 40742 112102 40794
rect 112154 40742 112206 40794
rect 112258 40742 142718 40794
rect 142770 40742 142822 40794
rect 142874 40742 142926 40794
rect 142978 40742 158592 40794
rect 1344 40708 158592 40742
rect 1344 40010 158592 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 96638 40010
rect 96690 39958 96742 40010
rect 96794 39958 96846 40010
rect 96898 39958 127358 40010
rect 127410 39958 127462 40010
rect 127514 39958 127566 40010
rect 127618 39958 158078 40010
rect 158130 39958 158182 40010
rect 158234 39958 158286 40010
rect 158338 39958 158592 40010
rect 1344 39924 158592 39958
rect 1344 39226 158592 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 81278 39226
rect 81330 39174 81382 39226
rect 81434 39174 81486 39226
rect 81538 39174 111998 39226
rect 112050 39174 112102 39226
rect 112154 39174 112206 39226
rect 112258 39174 142718 39226
rect 142770 39174 142822 39226
rect 142874 39174 142926 39226
rect 142978 39174 158592 39226
rect 1344 39140 158592 39174
rect 1344 38442 158592 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 96638 38442
rect 96690 38390 96742 38442
rect 96794 38390 96846 38442
rect 96898 38390 127358 38442
rect 127410 38390 127462 38442
rect 127514 38390 127566 38442
rect 127618 38390 158078 38442
rect 158130 38390 158182 38442
rect 158234 38390 158286 38442
rect 158338 38390 158592 38442
rect 1344 38356 158592 38390
rect 1344 37658 158592 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 81278 37658
rect 81330 37606 81382 37658
rect 81434 37606 81486 37658
rect 81538 37606 111998 37658
rect 112050 37606 112102 37658
rect 112154 37606 112206 37658
rect 112258 37606 142718 37658
rect 142770 37606 142822 37658
rect 142874 37606 142926 37658
rect 142978 37606 158592 37658
rect 1344 37572 158592 37606
rect 1344 36874 158592 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 96638 36874
rect 96690 36822 96742 36874
rect 96794 36822 96846 36874
rect 96898 36822 127358 36874
rect 127410 36822 127462 36874
rect 127514 36822 127566 36874
rect 127618 36822 158078 36874
rect 158130 36822 158182 36874
rect 158234 36822 158286 36874
rect 158338 36822 158592 36874
rect 1344 36788 158592 36822
rect 1344 36090 158592 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 81278 36090
rect 81330 36038 81382 36090
rect 81434 36038 81486 36090
rect 81538 36038 111998 36090
rect 112050 36038 112102 36090
rect 112154 36038 112206 36090
rect 112258 36038 142718 36090
rect 142770 36038 142822 36090
rect 142874 36038 142926 36090
rect 142978 36038 158592 36090
rect 1344 36004 158592 36038
rect 1344 35306 158592 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 96638 35306
rect 96690 35254 96742 35306
rect 96794 35254 96846 35306
rect 96898 35254 127358 35306
rect 127410 35254 127462 35306
rect 127514 35254 127566 35306
rect 127618 35254 158078 35306
rect 158130 35254 158182 35306
rect 158234 35254 158286 35306
rect 158338 35254 158592 35306
rect 1344 35220 158592 35254
rect 1344 34522 158592 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 81278 34522
rect 81330 34470 81382 34522
rect 81434 34470 81486 34522
rect 81538 34470 111998 34522
rect 112050 34470 112102 34522
rect 112154 34470 112206 34522
rect 112258 34470 142718 34522
rect 142770 34470 142822 34522
rect 142874 34470 142926 34522
rect 142978 34470 158592 34522
rect 1344 34436 158592 34470
rect 1344 33738 158592 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 96638 33738
rect 96690 33686 96742 33738
rect 96794 33686 96846 33738
rect 96898 33686 127358 33738
rect 127410 33686 127462 33738
rect 127514 33686 127566 33738
rect 127618 33686 158078 33738
rect 158130 33686 158182 33738
rect 158234 33686 158286 33738
rect 158338 33686 158592 33738
rect 1344 33652 158592 33686
rect 1344 32954 158592 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 81278 32954
rect 81330 32902 81382 32954
rect 81434 32902 81486 32954
rect 81538 32902 111998 32954
rect 112050 32902 112102 32954
rect 112154 32902 112206 32954
rect 112258 32902 142718 32954
rect 142770 32902 142822 32954
rect 142874 32902 142926 32954
rect 142978 32902 158592 32954
rect 1344 32868 158592 32902
rect 1344 32170 158592 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 96638 32170
rect 96690 32118 96742 32170
rect 96794 32118 96846 32170
rect 96898 32118 127358 32170
rect 127410 32118 127462 32170
rect 127514 32118 127566 32170
rect 127618 32118 158078 32170
rect 158130 32118 158182 32170
rect 158234 32118 158286 32170
rect 158338 32118 158592 32170
rect 1344 32084 158592 32118
rect 1344 31386 158592 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 81278 31386
rect 81330 31334 81382 31386
rect 81434 31334 81486 31386
rect 81538 31334 111998 31386
rect 112050 31334 112102 31386
rect 112154 31334 112206 31386
rect 112258 31334 142718 31386
rect 142770 31334 142822 31386
rect 142874 31334 142926 31386
rect 142978 31334 158592 31386
rect 1344 31300 158592 31334
rect 1344 30602 158592 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 96638 30602
rect 96690 30550 96742 30602
rect 96794 30550 96846 30602
rect 96898 30550 127358 30602
rect 127410 30550 127462 30602
rect 127514 30550 127566 30602
rect 127618 30550 158078 30602
rect 158130 30550 158182 30602
rect 158234 30550 158286 30602
rect 158338 30550 158592 30602
rect 1344 30516 158592 30550
rect 48850 30270 48862 30322
rect 48914 30270 48926 30322
rect 52098 30270 52110 30322
rect 52162 30270 52174 30322
rect 54798 30210 54850 30222
rect 61070 30210 61122 30222
rect 46050 30158 46062 30210
rect 46114 30158 46126 30210
rect 49298 30158 49310 30210
rect 49362 30158 49374 30210
rect 55234 30158 55246 30210
rect 55298 30158 55310 30210
rect 55794 30158 55806 30210
rect 55858 30158 55870 30210
rect 54798 30146 54850 30158
rect 61070 30146 61122 30158
rect 56254 30098 56306 30110
rect 46722 30046 46734 30098
rect 46786 30046 46798 30098
rect 49970 30046 49982 30098
rect 50034 30046 50046 30098
rect 56254 30034 56306 30046
rect 52782 29986 52834 29998
rect 52782 29922 52834 29934
rect 54126 29986 54178 29998
rect 54126 29922 54178 29934
rect 60510 29986 60562 29998
rect 60510 29922 60562 29934
rect 1344 29818 158592 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 81278 29818
rect 81330 29766 81382 29818
rect 81434 29766 81486 29818
rect 81538 29766 111998 29818
rect 112050 29766 112102 29818
rect 112154 29766 112206 29818
rect 112258 29766 142718 29818
rect 142770 29766 142822 29818
rect 142874 29766 142926 29818
rect 142978 29766 158592 29818
rect 1344 29732 158592 29766
rect 59502 29650 59554 29662
rect 59502 29586 59554 29598
rect 54574 29538 54626 29550
rect 43698 29486 43710 29538
rect 43762 29486 43774 29538
rect 54574 29474 54626 29486
rect 55022 29538 55074 29550
rect 55022 29474 55074 29486
rect 56590 29426 56642 29438
rect 46162 29374 46174 29426
rect 46226 29374 46238 29426
rect 46946 29374 46958 29426
rect 47010 29374 47022 29426
rect 51090 29374 51102 29426
rect 51154 29374 51166 29426
rect 56590 29362 56642 29374
rect 59390 29426 59442 29438
rect 59390 29362 59442 29374
rect 47294 29314 47346 29326
rect 47294 29250 47346 29262
rect 49086 29314 49138 29326
rect 55582 29314 55634 29326
rect 65326 29314 65378 29326
rect 51762 29262 51774 29314
rect 51826 29262 51838 29314
rect 53890 29262 53902 29314
rect 53954 29262 53966 29314
rect 57026 29262 57038 29314
rect 57090 29262 57102 29314
rect 49086 29250 49138 29262
rect 55582 29250 55634 29262
rect 65326 29250 65378 29262
rect 54462 29202 54514 29214
rect 54462 29138 54514 29150
rect 59502 29202 59554 29214
rect 59502 29138 59554 29150
rect 1344 29034 158592 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 96638 29034
rect 96690 28982 96742 29034
rect 96794 28982 96846 29034
rect 96898 28982 127358 29034
rect 127410 28982 127462 29034
rect 127514 28982 127566 29034
rect 127618 28982 158078 29034
rect 158130 28982 158182 29034
rect 158234 28982 158286 29034
rect 158338 28982 158592 29034
rect 1344 28948 158592 28982
rect 56478 28754 56530 28766
rect 32610 28702 32622 28754
rect 32674 28702 32686 28754
rect 48850 28702 48862 28754
rect 48914 28702 48926 28754
rect 56018 28702 56030 28754
rect 56082 28702 56094 28754
rect 56478 28690 56530 28702
rect 56814 28754 56866 28766
rect 56814 28690 56866 28702
rect 73390 28754 73442 28766
rect 73390 28690 73442 28702
rect 49310 28642 49362 28654
rect 50094 28642 50146 28654
rect 29810 28590 29822 28642
rect 29874 28590 29886 28642
rect 49858 28590 49870 28642
rect 49922 28590 49934 28642
rect 49310 28578 49362 28590
rect 50094 28578 50146 28590
rect 50318 28642 50370 28654
rect 50318 28578 50370 28590
rect 50542 28642 50594 28654
rect 50542 28578 50594 28590
rect 53006 28642 53058 28654
rect 57710 28642 57762 28654
rect 53442 28590 53454 28642
rect 53506 28590 53518 28642
rect 53890 28590 53902 28642
rect 53954 28590 53966 28642
rect 55906 28590 55918 28642
rect 55970 28590 55982 28642
rect 57250 28590 57262 28642
rect 57314 28590 57326 28642
rect 53006 28578 53058 28590
rect 57710 28578 57762 28590
rect 58494 28642 58546 28654
rect 58494 28578 58546 28590
rect 59054 28642 59106 28654
rect 59054 28578 59106 28590
rect 59390 28642 59442 28654
rect 59390 28578 59442 28590
rect 60734 28642 60786 28654
rect 60734 28578 60786 28590
rect 62638 28642 62690 28654
rect 62850 28590 62862 28642
rect 62914 28590 62926 28642
rect 63634 28590 63646 28642
rect 63698 28590 63710 28642
rect 69122 28590 69134 28642
rect 69186 28590 69198 28642
rect 72706 28590 72718 28642
rect 72770 28590 72782 28642
rect 62638 28578 62690 28590
rect 44830 28530 44882 28542
rect 30482 28478 30494 28530
rect 30546 28478 30558 28530
rect 44830 28466 44882 28478
rect 45166 28530 45218 28542
rect 45166 28466 45218 28478
rect 49646 28530 49698 28542
rect 55122 28478 55134 28530
rect 55186 28478 55198 28530
rect 49646 28466 49698 28478
rect 33070 28418 33122 28430
rect 51102 28418 51154 28430
rect 57822 28418 57874 28430
rect 49970 28366 49982 28418
rect 50034 28366 50046 28418
rect 54226 28366 54238 28418
rect 54290 28366 54302 28418
rect 33070 28354 33122 28366
rect 51102 28354 51154 28366
rect 57822 28354 57874 28366
rect 58046 28418 58098 28430
rect 66446 28418 66498 28430
rect 70590 28418 70642 28430
rect 59714 28366 59726 28418
rect 59778 28366 59790 28418
rect 65986 28366 65998 28418
rect 66050 28366 66062 28418
rect 69346 28366 69358 28418
rect 69410 28366 69422 28418
rect 58046 28354 58098 28366
rect 66446 28354 66498 28366
rect 70590 28354 70642 28366
rect 71038 28418 71090 28430
rect 72930 28366 72942 28418
rect 72994 28366 73006 28418
rect 71038 28354 71090 28366
rect 1344 28250 158592 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 81278 28250
rect 81330 28198 81382 28250
rect 81434 28198 81486 28250
rect 81538 28198 111998 28250
rect 112050 28198 112102 28250
rect 112154 28198 112206 28250
rect 112258 28198 142718 28250
rect 142770 28198 142822 28250
rect 142874 28198 142926 28250
rect 142978 28198 158592 28250
rect 1344 28164 158592 28198
rect 44158 28082 44210 28094
rect 44158 28018 44210 28030
rect 44718 28082 44770 28094
rect 63982 28082 64034 28094
rect 50866 28030 50878 28082
rect 50930 28030 50942 28082
rect 44718 28018 44770 28030
rect 63982 28018 64034 28030
rect 64766 28082 64818 28094
rect 64766 28018 64818 28030
rect 66110 28082 66162 28094
rect 66110 28018 66162 28030
rect 78654 28082 78706 28094
rect 78654 28018 78706 28030
rect 30942 27970 30994 27982
rect 33854 27970 33906 27982
rect 55246 27970 55298 27982
rect 63758 27970 63810 27982
rect 33170 27918 33182 27970
rect 33234 27918 33246 27970
rect 50978 27918 50990 27970
rect 51042 27918 51054 27970
rect 54002 27918 54014 27970
rect 54066 27918 54078 27970
rect 55570 27918 55582 27970
rect 55634 27918 55646 27970
rect 58034 27918 58046 27970
rect 58098 27918 58110 27970
rect 30942 27906 30994 27918
rect 33854 27906 33906 27918
rect 55246 27906 55298 27918
rect 63758 27906 63810 27918
rect 64654 27970 64706 27982
rect 64654 27906 64706 27918
rect 65326 27970 65378 27982
rect 65326 27906 65378 27918
rect 70926 27970 70978 27982
rect 73714 27918 73726 27970
rect 73778 27918 73790 27970
rect 78194 27918 78206 27970
rect 78258 27918 78270 27970
rect 70926 27906 70978 27918
rect 44606 27858 44658 27870
rect 50318 27858 50370 27870
rect 26898 27806 26910 27858
rect 26962 27806 26974 27858
rect 30706 27806 30718 27858
rect 30770 27806 30782 27858
rect 33394 27806 33406 27858
rect 33458 27806 33470 27858
rect 34178 27806 34190 27858
rect 34242 27806 34254 27858
rect 45266 27806 45278 27858
rect 45330 27806 45342 27858
rect 49410 27806 49422 27858
rect 49474 27806 49486 27858
rect 49634 27806 49646 27858
rect 49698 27806 49710 27858
rect 44606 27794 44658 27806
rect 50318 27794 50370 27806
rect 50542 27858 50594 27870
rect 53230 27858 53282 27870
rect 51202 27806 51214 27858
rect 51266 27806 51278 27858
rect 50542 27794 50594 27806
rect 53230 27794 53282 27806
rect 53342 27858 53394 27870
rect 53342 27794 53394 27806
rect 54350 27858 54402 27870
rect 57374 27858 57426 27870
rect 59278 27858 59330 27870
rect 56914 27806 56926 27858
rect 56978 27806 56990 27858
rect 57698 27806 57710 27858
rect 57762 27806 57774 27858
rect 54350 27794 54402 27806
rect 57374 27794 57426 27806
rect 59278 27794 59330 27806
rect 59502 27858 59554 27870
rect 60622 27858 60674 27870
rect 59826 27806 59838 27858
rect 59890 27806 59902 27858
rect 59502 27794 59554 27806
rect 60622 27794 60674 27806
rect 60846 27858 60898 27870
rect 63646 27858 63698 27870
rect 61058 27806 61070 27858
rect 61122 27806 61134 27858
rect 60846 27794 60898 27806
rect 63646 27794 63698 27806
rect 64542 27858 64594 27870
rect 64542 27794 64594 27806
rect 65102 27858 65154 27870
rect 65886 27858 65938 27870
rect 65650 27806 65662 27858
rect 65714 27806 65726 27858
rect 65102 27794 65154 27806
rect 65886 27794 65938 27806
rect 66222 27858 66274 27870
rect 70702 27858 70754 27870
rect 67106 27806 67118 27858
rect 67170 27806 67182 27858
rect 69682 27806 69694 27858
rect 69746 27806 69758 27858
rect 70354 27806 70366 27858
rect 70418 27806 70430 27858
rect 71138 27806 71150 27858
rect 71202 27806 71214 27858
rect 71474 27806 71486 27858
rect 71538 27806 71550 27858
rect 72706 27806 72718 27858
rect 72770 27806 72782 27858
rect 73938 27806 73950 27858
rect 74002 27806 74014 27858
rect 77634 27806 77646 27858
rect 77698 27806 77710 27858
rect 66222 27794 66274 27806
rect 70702 27794 70754 27806
rect 30158 27746 30210 27758
rect 27570 27694 27582 27746
rect 27634 27694 27646 27746
rect 29698 27694 29710 27746
rect 29762 27694 29774 27746
rect 30158 27682 30210 27694
rect 40350 27746 40402 27758
rect 40350 27682 40402 27694
rect 45054 27746 45106 27758
rect 45054 27682 45106 27694
rect 45726 27746 45778 27758
rect 51774 27746 51826 27758
rect 48962 27694 48974 27746
rect 49026 27694 49038 27746
rect 45726 27682 45778 27694
rect 51774 27682 51826 27694
rect 57150 27746 57202 27758
rect 63310 27746 63362 27758
rect 62066 27694 62078 27746
rect 62130 27694 62142 27746
rect 57150 27682 57202 27694
rect 63310 27682 63362 27694
rect 70814 27746 70866 27758
rect 70814 27682 70866 27694
rect 72270 27746 72322 27758
rect 74734 27746 74786 27758
rect 73154 27694 73166 27746
rect 73218 27694 73230 27746
rect 74274 27694 74286 27746
rect 74338 27694 74350 27746
rect 77746 27694 77758 27746
rect 77810 27694 77822 27746
rect 72270 27682 72322 27694
rect 74734 27682 74786 27694
rect 34190 27634 34242 27646
rect 34190 27570 34242 27582
rect 44830 27634 44882 27646
rect 50766 27634 50818 27646
rect 48850 27582 48862 27634
rect 48914 27582 48926 27634
rect 44830 27570 44882 27582
rect 50766 27570 50818 27582
rect 57822 27634 57874 27646
rect 57822 27570 57874 27582
rect 65662 27634 65714 27646
rect 65662 27570 65714 27582
rect 1344 27466 158592 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 96638 27466
rect 96690 27414 96742 27466
rect 96794 27414 96846 27466
rect 96898 27414 127358 27466
rect 127410 27414 127462 27466
rect 127514 27414 127566 27466
rect 127618 27414 158078 27466
rect 158130 27414 158182 27466
rect 158234 27414 158286 27466
rect 158338 27414 158592 27466
rect 1344 27380 158592 27414
rect 51774 27298 51826 27310
rect 51774 27234 51826 27246
rect 59950 27298 60002 27310
rect 59950 27234 60002 27246
rect 71598 27298 71650 27310
rect 71598 27234 71650 27246
rect 45054 27186 45106 27198
rect 59390 27186 59442 27198
rect 61630 27186 61682 27198
rect 62750 27186 62802 27198
rect 34402 27134 34414 27186
rect 34466 27134 34478 27186
rect 49858 27134 49870 27186
rect 49922 27134 49934 27186
rect 60834 27134 60846 27186
rect 60898 27134 60910 27186
rect 61954 27134 61966 27186
rect 62018 27134 62030 27186
rect 45054 27122 45106 27134
rect 59390 27122 59442 27134
rect 61630 27122 61682 27134
rect 62750 27122 62802 27134
rect 63198 27186 63250 27198
rect 63198 27122 63250 27134
rect 63646 27186 63698 27198
rect 66446 27186 66498 27198
rect 69582 27186 69634 27198
rect 64306 27134 64318 27186
rect 64370 27134 64382 27186
rect 69122 27134 69134 27186
rect 69186 27134 69198 27186
rect 63646 27122 63698 27134
rect 66446 27122 66498 27134
rect 69582 27122 69634 27134
rect 70030 27186 70082 27198
rect 75182 27186 75234 27198
rect 72818 27134 72830 27186
rect 72882 27134 72894 27186
rect 70030 27122 70082 27134
rect 75182 27122 75234 27134
rect 105758 27186 105810 27198
rect 105758 27122 105810 27134
rect 31726 27074 31778 27086
rect 36318 27074 36370 27086
rect 50094 27074 50146 27086
rect 50654 27074 50706 27086
rect 31154 27022 31166 27074
rect 31218 27022 31230 27074
rect 34738 27022 34750 27074
rect 34802 27022 34814 27074
rect 35858 27022 35870 27074
rect 35922 27022 35934 27074
rect 45938 27022 45950 27074
rect 46002 27022 46014 27074
rect 47730 27022 47742 27074
rect 47794 27022 47806 27074
rect 48626 27022 48638 27074
rect 48690 27022 48702 27074
rect 49746 27022 49758 27074
rect 49810 27022 49822 27074
rect 50418 27022 50430 27074
rect 50482 27022 50494 27074
rect 31726 27010 31778 27022
rect 36318 27010 36370 27022
rect 50094 27010 50146 27022
rect 50654 27010 50706 27022
rect 50878 27074 50930 27086
rect 50878 27010 50930 27022
rect 51438 27074 51490 27086
rect 51438 27010 51490 27022
rect 54686 27074 54738 27086
rect 57150 27074 57202 27086
rect 55010 27022 55022 27074
rect 55074 27022 55086 27074
rect 54686 27010 54738 27022
rect 57150 27010 57202 27022
rect 59614 27074 59666 27086
rect 59614 27010 59666 27022
rect 61294 27074 61346 27086
rect 61294 27010 61346 27022
rect 63982 27074 64034 27086
rect 69246 27074 69298 27086
rect 64642 27022 64654 27074
rect 64706 27022 64718 27074
rect 63982 27010 64034 27022
rect 69246 27010 69298 27022
rect 69806 27074 69858 27086
rect 69806 27010 69858 27022
rect 70254 27074 70306 27086
rect 70254 27010 70306 27022
rect 70366 27074 70418 27086
rect 70366 27010 70418 27022
rect 71710 27074 71762 27086
rect 71710 27010 71762 27022
rect 71934 27074 71986 27086
rect 71934 27010 71986 27022
rect 72270 27074 72322 27086
rect 72270 27010 72322 27022
rect 73278 27074 73330 27086
rect 73278 27010 73330 27022
rect 73614 27074 73666 27086
rect 73614 27010 73666 27022
rect 74174 27074 74226 27086
rect 74174 27010 74226 27022
rect 74958 27074 75010 27086
rect 74958 27010 75010 27022
rect 75294 27074 75346 27086
rect 75294 27010 75346 27022
rect 75518 27074 75570 27086
rect 79662 27074 79714 27086
rect 76178 27022 76190 27074
rect 76242 27022 76254 27074
rect 78530 27022 78542 27074
rect 78594 27022 78606 27074
rect 79090 27022 79102 27074
rect 79154 27022 79166 27074
rect 75518 27010 75570 27022
rect 79662 27010 79714 27022
rect 31838 26962 31890 26974
rect 31838 26898 31890 26910
rect 35310 26962 35362 26974
rect 36430 26962 36482 26974
rect 35634 26910 35646 26962
rect 35698 26910 35710 26962
rect 35310 26898 35362 26910
rect 36430 26898 36482 26910
rect 39678 26962 39730 26974
rect 39678 26898 39730 26910
rect 39902 26962 39954 26974
rect 39902 26898 39954 26910
rect 40238 26962 40290 26974
rect 40238 26898 40290 26910
rect 40574 26962 40626 26974
rect 40574 26898 40626 26910
rect 40798 26962 40850 26974
rect 40798 26898 40850 26910
rect 41022 26962 41074 26974
rect 51102 26962 51154 26974
rect 46162 26910 46174 26962
rect 46226 26910 46238 26962
rect 48738 26910 48750 26962
rect 48802 26910 48814 26962
rect 49634 26910 49646 26962
rect 49698 26910 49710 26962
rect 41022 26898 41074 26910
rect 51102 26898 51154 26910
rect 51662 26962 51714 26974
rect 61854 26962 61906 26974
rect 55122 26910 55134 26962
rect 55186 26910 55198 26962
rect 58706 26910 58718 26962
rect 58770 26910 58782 26962
rect 51662 26898 51714 26910
rect 61854 26898 61906 26910
rect 65662 26962 65714 26974
rect 65662 26898 65714 26910
rect 67566 26962 67618 26974
rect 67566 26898 67618 26910
rect 67678 26962 67730 26974
rect 67678 26898 67730 26910
rect 67902 26962 67954 26974
rect 67902 26898 67954 26910
rect 68462 26962 68514 26974
rect 68462 26898 68514 26910
rect 71262 26962 71314 26974
rect 71262 26898 71314 26910
rect 73726 26962 73778 26974
rect 73726 26898 73778 26910
rect 73950 26962 74002 26974
rect 73950 26898 74002 26910
rect 26350 26850 26402 26862
rect 26350 26786 26402 26798
rect 40014 26850 40066 26862
rect 40014 26786 40066 26798
rect 40686 26850 40738 26862
rect 55582 26850 55634 26862
rect 50530 26798 50542 26850
rect 50594 26798 50606 26850
rect 54338 26798 54350 26850
rect 54402 26798 54414 26850
rect 40686 26786 40738 26798
rect 55582 26786 55634 26798
rect 64206 26850 64258 26862
rect 64206 26786 64258 26798
rect 67006 26850 67058 26862
rect 67006 26786 67058 26798
rect 72158 26850 72210 26862
rect 72158 26786 72210 26798
rect 74286 26850 74338 26862
rect 74286 26786 74338 26798
rect 74510 26850 74562 26862
rect 74510 26786 74562 26798
rect 1344 26682 158592 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 81278 26682
rect 81330 26630 81382 26682
rect 81434 26630 81486 26682
rect 81538 26630 111998 26682
rect 112050 26630 112102 26682
rect 112154 26630 112206 26682
rect 112258 26630 142718 26682
rect 142770 26630 142822 26682
rect 142874 26630 142926 26682
rect 142978 26630 158592 26682
rect 1344 26596 158592 26630
rect 24222 26514 24274 26526
rect 24222 26450 24274 26462
rect 25790 26514 25842 26526
rect 25790 26450 25842 26462
rect 26014 26514 26066 26526
rect 26014 26450 26066 26462
rect 26686 26514 26738 26526
rect 26686 26450 26738 26462
rect 27134 26514 27186 26526
rect 27134 26450 27186 26462
rect 31726 26514 31778 26526
rect 31726 26450 31778 26462
rect 41246 26514 41298 26526
rect 41246 26450 41298 26462
rect 41694 26514 41746 26526
rect 41694 26450 41746 26462
rect 41918 26514 41970 26526
rect 41918 26450 41970 26462
rect 46062 26514 46114 26526
rect 46062 26450 46114 26462
rect 47854 26514 47906 26526
rect 47854 26450 47906 26462
rect 48862 26514 48914 26526
rect 51998 26514 52050 26526
rect 50194 26462 50206 26514
rect 50258 26462 50270 26514
rect 48862 26450 48914 26462
rect 51998 26450 52050 26462
rect 64430 26514 64482 26526
rect 64430 26450 64482 26462
rect 65438 26514 65490 26526
rect 65438 26450 65490 26462
rect 71710 26514 71762 26526
rect 71710 26450 71762 26462
rect 72494 26514 72546 26526
rect 72494 26450 72546 26462
rect 73278 26514 73330 26526
rect 73278 26450 73330 26462
rect 75294 26514 75346 26526
rect 75294 26450 75346 26462
rect 75406 26514 75458 26526
rect 75406 26450 75458 26462
rect 107102 26514 107154 26526
rect 107102 26450 107154 26462
rect 24446 26402 24498 26414
rect 24446 26338 24498 26350
rect 24558 26402 24610 26414
rect 36542 26402 36594 26414
rect 30482 26350 30494 26402
rect 30546 26350 30558 26402
rect 32050 26350 32062 26402
rect 32114 26350 32126 26402
rect 24558 26338 24610 26350
rect 36542 26338 36594 26350
rect 38334 26402 38386 26414
rect 38334 26338 38386 26350
rect 38446 26402 38498 26414
rect 38446 26338 38498 26350
rect 39454 26402 39506 26414
rect 39454 26338 39506 26350
rect 42030 26402 42082 26414
rect 42030 26338 42082 26350
rect 42590 26402 42642 26414
rect 42590 26338 42642 26350
rect 43262 26402 43314 26414
rect 48078 26402 48130 26414
rect 50766 26402 50818 26414
rect 43586 26350 43598 26402
rect 43650 26350 43662 26402
rect 49634 26350 49646 26402
rect 49698 26350 49710 26402
rect 49858 26350 49870 26402
rect 49922 26350 49934 26402
rect 43262 26338 43314 26350
rect 48078 26338 48130 26350
rect 50766 26338 50818 26350
rect 50990 26402 51042 26414
rect 50990 26338 51042 26350
rect 51886 26402 51938 26414
rect 53118 26402 53170 26414
rect 52770 26350 52782 26402
rect 52834 26350 52846 26402
rect 51886 26338 51938 26350
rect 53118 26338 53170 26350
rect 55918 26402 55970 26414
rect 58158 26402 58210 26414
rect 68350 26402 68402 26414
rect 56914 26350 56926 26402
rect 56978 26350 56990 26402
rect 63634 26350 63646 26402
rect 63698 26350 63710 26402
rect 55918 26338 55970 26350
rect 58158 26338 58210 26350
rect 68350 26338 68402 26350
rect 70142 26402 70194 26414
rect 70142 26338 70194 26350
rect 72270 26402 72322 26414
rect 72270 26338 72322 26350
rect 72718 26402 72770 26414
rect 72718 26338 72770 26350
rect 73054 26402 73106 26414
rect 75742 26402 75794 26414
rect 73938 26350 73950 26402
rect 74002 26350 74014 26402
rect 105522 26350 105534 26402
rect 105586 26350 105598 26402
rect 106530 26350 106542 26402
rect 106594 26350 106606 26402
rect 73054 26338 73106 26350
rect 75742 26338 75794 26350
rect 24782 26290 24834 26302
rect 30942 26290 30994 26302
rect 35534 26290 35586 26302
rect 25330 26238 25342 26290
rect 25394 26238 25406 26290
rect 25554 26238 25566 26290
rect 25618 26238 25630 26290
rect 30258 26238 30270 26290
rect 30322 26238 30334 26290
rect 31378 26238 31390 26290
rect 31442 26238 31454 26290
rect 24782 26226 24834 26238
rect 30942 26226 30994 26238
rect 35534 26226 35586 26238
rect 35758 26290 35810 26302
rect 35758 26226 35810 26238
rect 36206 26290 36258 26302
rect 36206 26226 36258 26238
rect 39006 26290 39058 26302
rect 39006 26226 39058 26238
rect 39118 26290 39170 26302
rect 39118 26226 39170 26238
rect 39790 26290 39842 26302
rect 39790 26226 39842 26238
rect 40014 26290 40066 26302
rect 40014 26226 40066 26238
rect 40798 26290 40850 26302
rect 40798 26226 40850 26238
rect 41470 26290 41522 26302
rect 41470 26226 41522 26238
rect 42926 26290 42978 26302
rect 42926 26226 42978 26238
rect 44270 26290 44322 26302
rect 44270 26226 44322 26238
rect 44494 26290 44546 26302
rect 48190 26290 48242 26302
rect 45490 26238 45502 26290
rect 45554 26238 45566 26290
rect 44494 26226 44546 26238
rect 48190 26226 48242 26238
rect 48974 26290 49026 26302
rect 48974 26226 49026 26238
rect 50318 26290 50370 26302
rect 50318 26226 50370 26238
rect 50878 26290 50930 26302
rect 54462 26290 54514 26302
rect 54002 26238 54014 26290
rect 54066 26238 54078 26290
rect 50878 26226 50930 26238
rect 54462 26226 54514 26238
rect 55694 26290 55746 26302
rect 55694 26226 55746 26238
rect 56030 26290 56082 26302
rect 57710 26290 57762 26302
rect 57138 26238 57150 26290
rect 57202 26238 57214 26290
rect 56030 26226 56082 26238
rect 57710 26226 57762 26238
rect 59390 26290 59442 26302
rect 59390 26226 59442 26238
rect 60510 26290 60562 26302
rect 67454 26290 67506 26302
rect 70590 26290 70642 26302
rect 62402 26238 62414 26290
rect 62466 26238 62478 26290
rect 63186 26238 63198 26290
rect 63250 26238 63262 26290
rect 63746 26238 63758 26290
rect 63810 26238 63822 26290
rect 67666 26238 67678 26290
rect 67730 26238 67742 26290
rect 60510 26226 60562 26238
rect 67454 26226 67506 26238
rect 70590 26226 70642 26238
rect 72830 26290 72882 26302
rect 72830 26226 72882 26238
rect 73614 26290 73666 26302
rect 75518 26290 75570 26302
rect 73826 26238 73838 26290
rect 73890 26238 73902 26290
rect 74722 26238 74734 26290
rect 74786 26238 74798 26290
rect 73614 26226 73666 26238
rect 75518 26226 75570 26238
rect 77198 26290 77250 26302
rect 77198 26226 77250 26238
rect 77758 26290 77810 26302
rect 86930 26238 86942 26290
rect 86994 26238 87006 26290
rect 104962 26238 104974 26290
rect 105026 26238 105038 26290
rect 105970 26238 105982 26290
rect 106034 26238 106046 26290
rect 77758 26226 77810 26238
rect 35646 26178 35698 26190
rect 25778 26126 25790 26178
rect 25842 26126 25854 26178
rect 35646 26114 35698 26126
rect 36654 26178 36706 26190
rect 36654 26114 36706 26126
rect 37998 26178 38050 26190
rect 37998 26114 38050 26126
rect 39342 26178 39394 26190
rect 39342 26114 39394 26126
rect 41358 26178 41410 26190
rect 46510 26178 46562 26190
rect 59950 26178 60002 26190
rect 61518 26178 61570 26190
rect 45378 26126 45390 26178
rect 45442 26126 45454 26178
rect 53778 26126 53790 26178
rect 53842 26126 53854 26178
rect 60946 26126 60958 26178
rect 61010 26126 61022 26178
rect 41358 26114 41410 26126
rect 46510 26114 46562 26126
rect 59950 26114 60002 26126
rect 61518 26114 61570 26126
rect 64990 26178 65042 26190
rect 64990 26114 65042 26126
rect 67790 26178 67842 26190
rect 67790 26114 67842 26126
rect 68910 26178 68962 26190
rect 76862 26178 76914 26190
rect 74162 26126 74174 26178
rect 74226 26126 74238 26178
rect 68910 26114 68962 26126
rect 76862 26114 76914 26126
rect 86158 26178 86210 26190
rect 104526 26178 104578 26190
rect 107550 26178 107602 26190
rect 86594 26126 86606 26178
rect 86658 26126 86670 26178
rect 104850 26126 104862 26178
rect 104914 26126 104926 26178
rect 86158 26114 86210 26126
rect 104526 26114 104578 26126
rect 107550 26114 107602 26126
rect 30830 26066 30882 26078
rect 30830 26002 30882 26014
rect 31166 26066 31218 26078
rect 31166 26002 31218 26014
rect 36766 26066 36818 26078
rect 36766 26002 36818 26014
rect 38446 26066 38498 26078
rect 45166 26066 45218 26078
rect 48862 26066 48914 26078
rect 40338 26014 40350 26066
rect 40402 26014 40414 26066
rect 44818 26014 44830 26066
rect 44882 26014 44894 26066
rect 45714 26014 45726 26066
rect 45778 26063 45790 26066
rect 46050 26063 46062 26066
rect 45778 26017 46062 26063
rect 45778 26014 45790 26017
rect 46050 26014 46062 26017
rect 46114 26014 46126 26066
rect 38446 26002 38498 26014
rect 45166 26002 45218 26014
rect 48862 26002 48914 26014
rect 52110 26066 52162 26078
rect 73390 26066 73442 26078
rect 54114 26014 54126 26066
rect 54178 26014 54190 26066
rect 52110 26002 52162 26014
rect 73390 26002 73442 26014
rect 106430 26066 106482 26078
rect 106430 26002 106482 26014
rect 1344 25898 158592 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 96638 25898
rect 96690 25846 96742 25898
rect 96794 25846 96846 25898
rect 96898 25846 127358 25898
rect 127410 25846 127462 25898
rect 127514 25846 127566 25898
rect 127618 25846 158078 25898
rect 158130 25846 158182 25898
rect 158234 25846 158286 25898
rect 158338 25846 158592 25898
rect 1344 25812 158592 25846
rect 35198 25730 35250 25742
rect 35198 25666 35250 25678
rect 35534 25730 35586 25742
rect 35534 25666 35586 25678
rect 36318 25730 36370 25742
rect 36318 25666 36370 25678
rect 37438 25730 37490 25742
rect 37438 25666 37490 25678
rect 37550 25730 37602 25742
rect 37550 25666 37602 25678
rect 37774 25730 37826 25742
rect 37774 25666 37826 25678
rect 62190 25730 62242 25742
rect 62190 25666 62242 25678
rect 34638 25618 34690 25630
rect 43486 25618 43538 25630
rect 31042 25566 31054 25618
rect 31106 25566 31118 25618
rect 38994 25566 39006 25618
rect 39058 25566 39070 25618
rect 34638 25554 34690 25566
rect 43486 25554 43538 25566
rect 45838 25618 45890 25630
rect 45838 25554 45890 25566
rect 48078 25618 48130 25630
rect 48078 25554 48130 25566
rect 48638 25618 48690 25630
rect 48638 25554 48690 25566
rect 48974 25618 49026 25630
rect 55918 25618 55970 25630
rect 71598 25618 71650 25630
rect 50866 25566 50878 25618
rect 50930 25566 50942 25618
rect 53106 25566 53118 25618
rect 53170 25566 53182 25618
rect 61170 25566 61182 25618
rect 61234 25566 61246 25618
rect 62626 25566 62638 25618
rect 62690 25566 62702 25618
rect 69906 25566 69918 25618
rect 69970 25566 69982 25618
rect 48974 25554 49026 25566
rect 55918 25554 55970 25566
rect 71598 25554 71650 25566
rect 87278 25618 87330 25630
rect 87278 25554 87330 25566
rect 90302 25618 90354 25630
rect 90302 25554 90354 25566
rect 101838 25618 101890 25630
rect 101838 25554 101890 25566
rect 105534 25618 105586 25630
rect 108670 25618 108722 25630
rect 106754 25566 106766 25618
rect 106818 25566 106830 25618
rect 105534 25554 105586 25566
rect 108670 25554 108722 25566
rect 31950 25506 32002 25518
rect 23426 25454 23438 25506
rect 23490 25454 23502 25506
rect 25778 25454 25790 25506
rect 25842 25454 25854 25506
rect 26562 25454 26574 25506
rect 26626 25454 26638 25506
rect 31490 25454 31502 25506
rect 31554 25454 31566 25506
rect 31950 25442 32002 25454
rect 34862 25506 34914 25518
rect 34862 25442 34914 25454
rect 35758 25506 35810 25518
rect 35758 25442 35810 25454
rect 36094 25506 36146 25518
rect 40014 25506 40066 25518
rect 38882 25454 38894 25506
rect 38946 25454 38958 25506
rect 39554 25454 39566 25506
rect 39618 25454 39630 25506
rect 36094 25442 36146 25454
rect 40014 25442 40066 25454
rect 41246 25506 41298 25518
rect 41246 25442 41298 25454
rect 41694 25506 41746 25518
rect 41694 25442 41746 25454
rect 43934 25506 43986 25518
rect 43934 25442 43986 25454
rect 44718 25506 44770 25518
rect 44718 25442 44770 25454
rect 45390 25506 45442 25518
rect 45390 25442 45442 25454
rect 47294 25506 47346 25518
rect 47294 25442 47346 25454
rect 47742 25506 47794 25518
rect 47742 25442 47794 25454
rect 48862 25506 48914 25518
rect 48862 25442 48914 25454
rect 49086 25506 49138 25518
rect 49086 25442 49138 25454
rect 49422 25506 49474 25518
rect 49422 25442 49474 25454
rect 50094 25506 50146 25518
rect 51774 25506 51826 25518
rect 53342 25506 53394 25518
rect 57598 25506 57650 25518
rect 50530 25454 50542 25506
rect 50594 25454 50606 25506
rect 50754 25454 50766 25506
rect 50818 25454 50830 25506
rect 52994 25454 53006 25506
rect 53058 25454 53070 25506
rect 53778 25454 53790 25506
rect 53842 25454 53854 25506
rect 50094 25442 50146 25454
rect 51774 25442 51826 25454
rect 53342 25442 53394 25454
rect 57598 25442 57650 25454
rect 58046 25506 58098 25518
rect 59054 25506 59106 25518
rect 61854 25506 61906 25518
rect 70478 25506 70530 25518
rect 58482 25454 58494 25506
rect 58546 25454 58558 25506
rect 59490 25454 59502 25506
rect 59554 25454 59566 25506
rect 65538 25454 65550 25506
rect 65602 25454 65614 25506
rect 68898 25454 68910 25506
rect 68962 25454 68974 25506
rect 69458 25454 69470 25506
rect 69522 25454 69534 25506
rect 58046 25442 58098 25454
rect 59054 25442 59106 25454
rect 61854 25442 61906 25454
rect 70478 25442 70530 25454
rect 70702 25506 70754 25518
rect 71150 25506 71202 25518
rect 70802 25454 70814 25506
rect 70866 25454 70878 25506
rect 70702 25442 70754 25454
rect 71150 25442 71202 25454
rect 72046 25506 72098 25518
rect 87614 25506 87666 25518
rect 72706 25454 72718 25506
rect 72770 25454 72782 25506
rect 74722 25454 74734 25506
rect 74786 25454 74798 25506
rect 77298 25454 77310 25506
rect 77362 25454 77374 25506
rect 78082 25454 78094 25506
rect 78146 25454 78158 25506
rect 72046 25442 72098 25454
rect 87614 25442 87666 25454
rect 88174 25506 88226 25518
rect 88174 25442 88226 25454
rect 88958 25506 89010 25518
rect 100494 25506 100546 25518
rect 106094 25506 106146 25518
rect 89730 25454 89742 25506
rect 89794 25454 89806 25506
rect 100930 25454 100942 25506
rect 100994 25454 101006 25506
rect 106530 25454 106542 25506
rect 106594 25454 106606 25506
rect 107650 25454 107662 25506
rect 107714 25454 107726 25506
rect 88958 25442 89010 25454
rect 100494 25442 100546 25454
rect 106094 25442 106146 25454
rect 33966 25394 34018 25406
rect 33966 25330 34018 25342
rect 34302 25394 34354 25406
rect 34302 25330 34354 25342
rect 38558 25394 38610 25406
rect 38558 25330 38610 25342
rect 39342 25394 39394 25406
rect 39342 25330 39394 25342
rect 40462 25394 40514 25406
rect 40462 25330 40514 25342
rect 43598 25394 43650 25406
rect 43598 25330 43650 25342
rect 43822 25394 43874 25406
rect 43822 25330 43874 25342
rect 45166 25394 45218 25406
rect 45166 25330 45218 25342
rect 50318 25394 50370 25406
rect 57150 25394 57202 25406
rect 61630 25394 61682 25406
rect 53890 25342 53902 25394
rect 53954 25342 53966 25394
rect 54450 25342 54462 25394
rect 54514 25342 54526 25394
rect 58818 25342 58830 25394
rect 58882 25342 58894 25394
rect 64754 25342 64766 25394
rect 64818 25342 64830 25394
rect 69906 25342 69918 25394
rect 69970 25342 69982 25394
rect 72594 25342 72606 25394
rect 72658 25342 72670 25394
rect 74834 25342 74846 25394
rect 74898 25342 74910 25394
rect 89842 25342 89854 25394
rect 89906 25342 89918 25394
rect 101378 25342 101390 25394
rect 101442 25342 101454 25394
rect 106978 25342 106990 25394
rect 107042 25342 107054 25394
rect 108210 25342 108222 25394
rect 108274 25342 108286 25394
rect 50318 25330 50370 25342
rect 57150 25330 57202 25342
rect 61630 25330 61682 25342
rect 26910 25282 26962 25294
rect 26910 25218 26962 25230
rect 33630 25282 33682 25294
rect 33630 25218 33682 25230
rect 36430 25282 36482 25294
rect 36430 25218 36482 25230
rect 37438 25282 37490 25294
rect 37438 25218 37490 25230
rect 38222 25282 38274 25294
rect 38222 25218 38274 25230
rect 38446 25282 38498 25294
rect 38446 25218 38498 25230
rect 40126 25282 40178 25294
rect 40126 25218 40178 25230
rect 40238 25282 40290 25294
rect 40238 25218 40290 25230
rect 41022 25282 41074 25294
rect 41022 25218 41074 25230
rect 41134 25282 41186 25294
rect 41134 25218 41186 25230
rect 45054 25282 45106 25294
rect 45054 25218 45106 25230
rect 46398 25282 46450 25294
rect 46398 25218 46450 25230
rect 51326 25282 51378 25294
rect 56254 25282 56306 25294
rect 54226 25230 54238 25282
rect 54290 25230 54302 25282
rect 51326 25218 51378 25230
rect 56254 25218 56306 25230
rect 60734 25282 60786 25294
rect 60734 25218 60786 25230
rect 70590 25282 70642 25294
rect 80894 25282 80946 25294
rect 80434 25230 80446 25282
rect 80498 25230 80510 25282
rect 89506 25230 89518 25282
rect 89570 25230 89582 25282
rect 100818 25230 100830 25282
rect 100882 25230 100894 25282
rect 107874 25230 107886 25282
rect 107938 25230 107950 25282
rect 70590 25218 70642 25230
rect 80894 25218 80946 25230
rect 1344 25114 158592 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 81278 25114
rect 81330 25062 81382 25114
rect 81434 25062 81486 25114
rect 81538 25062 111998 25114
rect 112050 25062 112102 25114
rect 112154 25062 112206 25114
rect 112258 25062 142718 25114
rect 142770 25062 142822 25114
rect 142874 25062 142926 25114
rect 142978 25062 158592 25114
rect 1344 25028 158592 25062
rect 23438 24946 23490 24958
rect 23438 24882 23490 24894
rect 31390 24946 31442 24958
rect 31390 24882 31442 24894
rect 36766 24946 36818 24958
rect 36766 24882 36818 24894
rect 37438 24946 37490 24958
rect 37438 24882 37490 24894
rect 39006 24946 39058 24958
rect 39006 24882 39058 24894
rect 43262 24946 43314 24958
rect 43262 24882 43314 24894
rect 46398 24946 46450 24958
rect 46398 24882 46450 24894
rect 46622 24946 46674 24958
rect 46622 24882 46674 24894
rect 49198 24946 49250 24958
rect 55806 24946 55858 24958
rect 52210 24894 52222 24946
rect 52274 24894 52286 24946
rect 49198 24882 49250 24894
rect 55806 24882 55858 24894
rect 56814 24946 56866 24958
rect 56814 24882 56866 24894
rect 62862 24946 62914 24958
rect 69470 24946 69522 24958
rect 68898 24894 68910 24946
rect 68962 24894 68974 24946
rect 62862 24882 62914 24894
rect 69470 24882 69522 24894
rect 69582 24946 69634 24958
rect 69582 24882 69634 24894
rect 69806 24946 69858 24958
rect 69806 24882 69858 24894
rect 70590 24946 70642 24958
rect 70590 24882 70642 24894
rect 70926 24946 70978 24958
rect 70926 24882 70978 24894
rect 76526 24946 76578 24958
rect 76526 24882 76578 24894
rect 78430 24946 78482 24958
rect 78430 24882 78482 24894
rect 80782 24946 80834 24958
rect 80782 24882 80834 24894
rect 107326 24946 107378 24958
rect 107326 24882 107378 24894
rect 31278 24834 31330 24846
rect 43374 24834 43426 24846
rect 55246 24834 55298 24846
rect 24546 24782 24558 24834
rect 24610 24782 24622 24834
rect 35298 24782 35310 24834
rect 35362 24782 35374 24834
rect 50642 24782 50654 24834
rect 50706 24782 50718 24834
rect 31278 24770 31330 24782
rect 43374 24770 43426 24782
rect 55246 24770 55298 24782
rect 55918 24834 55970 24846
rect 55918 24770 55970 24782
rect 56030 24834 56082 24846
rect 56030 24770 56082 24782
rect 57038 24834 57090 24846
rect 57038 24770 57090 24782
rect 57934 24834 57986 24846
rect 70030 24834 70082 24846
rect 58258 24782 58270 24834
rect 58322 24782 58334 24834
rect 64754 24782 64766 24834
rect 64818 24782 64830 24834
rect 68674 24782 68686 24834
rect 68738 24782 68750 24834
rect 57934 24770 57986 24782
rect 70030 24770 70082 24782
rect 71150 24834 71202 24846
rect 71150 24770 71202 24782
rect 71262 24834 71314 24846
rect 71262 24770 71314 24782
rect 71710 24834 71762 24846
rect 74834 24782 74846 24834
rect 74898 24782 74910 24834
rect 76850 24782 76862 24834
rect 76914 24782 76926 24834
rect 81106 24782 81118 24834
rect 81170 24782 81182 24834
rect 71710 24770 71762 24782
rect 31950 24722 32002 24734
rect 24434 24670 24446 24722
rect 24498 24670 24510 24722
rect 27234 24670 27246 24722
rect 27298 24670 27310 24722
rect 31950 24658 32002 24670
rect 32622 24722 32674 24734
rect 35534 24722 35586 24734
rect 34738 24670 34750 24722
rect 34802 24670 34814 24722
rect 32622 24658 32674 24670
rect 35534 24658 35586 24670
rect 35870 24722 35922 24734
rect 35870 24658 35922 24670
rect 36094 24722 36146 24734
rect 36094 24658 36146 24670
rect 43038 24722 43090 24734
rect 43038 24658 43090 24670
rect 44046 24722 44098 24734
rect 44046 24658 44098 24670
rect 44494 24722 44546 24734
rect 44494 24658 44546 24670
rect 45054 24722 45106 24734
rect 50430 24722 50482 24734
rect 55022 24722 55074 24734
rect 46946 24670 46958 24722
rect 47010 24670 47022 24722
rect 49410 24670 49422 24722
rect 49474 24670 49486 24722
rect 51090 24670 51102 24722
rect 51154 24670 51166 24722
rect 45054 24658 45106 24670
rect 50430 24658 50482 24670
rect 55022 24658 55074 24670
rect 55358 24722 55410 24734
rect 55358 24658 55410 24670
rect 56478 24722 56530 24734
rect 56478 24658 56530 24670
rect 57710 24722 57762 24734
rect 64430 24722 64482 24734
rect 68014 24722 68066 24734
rect 70366 24722 70418 24734
rect 58482 24670 58494 24722
rect 58546 24670 58558 24722
rect 59490 24670 59502 24722
rect 59554 24670 59566 24722
rect 67554 24670 67566 24722
rect 67618 24670 67630 24722
rect 68338 24670 68350 24722
rect 68402 24670 68414 24722
rect 57710 24658 57762 24670
rect 64430 24658 64482 24670
rect 68014 24658 68066 24670
rect 70366 24658 70418 24670
rect 72718 24722 72770 24734
rect 78206 24722 78258 24734
rect 73826 24670 73838 24722
rect 73890 24670 73902 24722
rect 74722 24670 74734 24722
rect 74786 24670 74798 24722
rect 75618 24670 75630 24722
rect 75682 24670 75694 24722
rect 78754 24670 78766 24722
rect 78818 24670 78830 24722
rect 83794 24670 83806 24722
rect 83858 24670 83870 24722
rect 84354 24670 84366 24722
rect 84418 24670 84430 24722
rect 72718 24658 72770 24670
rect 78206 24658 78258 24670
rect 30494 24610 30546 24622
rect 27906 24558 27918 24610
rect 27970 24558 27982 24610
rect 30034 24558 30046 24610
rect 30098 24558 30110 24610
rect 30494 24546 30546 24558
rect 31726 24610 31778 24622
rect 31726 24546 31778 24558
rect 35422 24610 35474 24622
rect 35422 24546 35474 24558
rect 46510 24610 46562 24622
rect 46510 24546 46562 24558
rect 49870 24610 49922 24622
rect 49870 24546 49922 24558
rect 50542 24610 50594 24622
rect 50542 24546 50594 24558
rect 51662 24610 51714 24622
rect 52782 24610 52834 24622
rect 62414 24610 62466 24622
rect 72382 24610 72434 24622
rect 78318 24610 78370 24622
rect 84926 24610 84978 24622
rect 51986 24558 51998 24610
rect 52050 24558 52062 24610
rect 57026 24558 57038 24610
rect 57090 24558 57102 24610
rect 59154 24558 59166 24610
rect 59218 24558 59230 24610
rect 69458 24558 69470 24610
rect 69522 24558 69534 24610
rect 70690 24558 70702 24610
rect 70754 24558 70766 24610
rect 74274 24558 74286 24610
rect 74338 24558 74350 24610
rect 75282 24558 75294 24610
rect 75346 24558 75358 24610
rect 81442 24558 81454 24610
rect 81506 24558 81518 24610
rect 51662 24546 51714 24558
rect 23774 24498 23826 24510
rect 23774 24434 23826 24446
rect 32174 24498 32226 24510
rect 36318 24498 36370 24510
rect 34962 24446 34974 24498
rect 35026 24446 35038 24498
rect 32174 24434 32226 24446
rect 36318 24434 36370 24446
rect 37102 24498 37154 24510
rect 37102 24434 37154 24446
rect 37326 24498 37378 24510
rect 37326 24434 37378 24446
rect 37438 24498 37490 24510
rect 37438 24434 37490 24446
rect 43822 24498 43874 24510
rect 43822 24434 43874 24446
rect 44494 24498 44546 24510
rect 44494 24434 44546 24446
rect 44606 24498 44658 24510
rect 44606 24434 44658 24446
rect 49086 24498 49138 24510
rect 49086 24434 49138 24446
rect 50878 24498 50930 24510
rect 51538 24446 51550 24498
rect 51602 24495 51614 24498
rect 52001 24495 52047 24558
rect 52782 24546 52834 24558
rect 62414 24546 62466 24558
rect 72382 24546 72434 24558
rect 78318 24546 78370 24558
rect 84926 24546 84978 24558
rect 51602 24449 52047 24495
rect 52558 24498 52610 24510
rect 51602 24446 51614 24449
rect 50878 24434 50930 24446
rect 52558 24434 52610 24446
rect 57374 24498 57426 24510
rect 62402 24446 62414 24498
rect 62466 24495 62478 24498
rect 62962 24495 62974 24498
rect 62466 24449 62974 24495
rect 62466 24446 62478 24449
rect 62962 24446 62974 24449
rect 63026 24446 63038 24498
rect 57374 24434 57426 24446
rect 1344 24330 158592 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 96638 24330
rect 96690 24278 96742 24330
rect 96794 24278 96846 24330
rect 96898 24278 127358 24330
rect 127410 24278 127462 24330
rect 127514 24278 127566 24330
rect 127618 24278 158078 24330
rect 158130 24278 158182 24330
rect 158234 24278 158286 24330
rect 158338 24278 158592 24330
rect 1344 24244 158592 24278
rect 27358 24162 27410 24174
rect 27358 24098 27410 24110
rect 46958 24162 47010 24174
rect 46958 24098 47010 24110
rect 50430 24162 50482 24174
rect 50430 24098 50482 24110
rect 53566 24162 53618 24174
rect 53566 24098 53618 24110
rect 43598 24050 43650 24062
rect 27794 23998 27806 24050
rect 27858 23998 27870 24050
rect 33954 23998 33966 24050
rect 34018 23998 34030 24050
rect 43598 23986 43650 23998
rect 48638 24050 48690 24062
rect 52782 24050 52834 24062
rect 50866 23998 50878 24050
rect 50930 23998 50942 24050
rect 48638 23986 48690 23998
rect 52782 23986 52834 23998
rect 58606 24050 58658 24062
rect 58606 23986 58658 23998
rect 64430 24050 64482 24062
rect 69246 24050 69298 24062
rect 67778 23998 67790 24050
rect 67842 23998 67854 24050
rect 64430 23986 64482 23998
rect 69246 23986 69298 23998
rect 73054 24050 73106 24062
rect 73054 23986 73106 23998
rect 34862 23938 34914 23950
rect 31154 23886 31166 23938
rect 31218 23886 31230 23938
rect 34862 23874 34914 23886
rect 35310 23938 35362 23950
rect 35310 23874 35362 23886
rect 35534 23938 35586 23950
rect 35534 23874 35586 23886
rect 39342 23938 39394 23950
rect 39342 23874 39394 23886
rect 39566 23938 39618 23950
rect 39566 23874 39618 23886
rect 40014 23938 40066 23950
rect 40014 23874 40066 23886
rect 43150 23938 43202 23950
rect 43150 23874 43202 23886
rect 45950 23938 46002 23950
rect 45950 23874 46002 23886
rect 46734 23938 46786 23950
rect 46734 23874 46786 23886
rect 47182 23938 47234 23950
rect 47182 23874 47234 23886
rect 47294 23938 47346 23950
rect 47294 23874 47346 23886
rect 47854 23938 47906 23950
rect 47854 23874 47906 23886
rect 50206 23938 50258 23950
rect 51102 23938 51154 23950
rect 50754 23886 50766 23938
rect 50818 23886 50830 23938
rect 50206 23874 50258 23886
rect 51102 23874 51154 23886
rect 51550 23938 51602 23950
rect 51550 23874 51602 23886
rect 51774 23938 51826 23950
rect 51774 23874 51826 23886
rect 52222 23938 52274 23950
rect 52222 23874 52274 23886
rect 54238 23938 54290 23950
rect 68910 23938 68962 23950
rect 54674 23886 54686 23938
rect 54738 23886 54750 23938
rect 57586 23886 57598 23938
rect 57650 23886 57662 23938
rect 58146 23886 58158 23938
rect 58210 23886 58222 23938
rect 64642 23886 64654 23938
rect 64706 23886 64718 23938
rect 65426 23886 65438 23938
rect 65490 23886 65502 23938
rect 54238 23874 54290 23886
rect 68910 23874 68962 23886
rect 73614 23938 73666 23950
rect 75630 23938 75682 23950
rect 74498 23886 74510 23938
rect 74562 23886 74574 23938
rect 74946 23886 74958 23938
rect 75010 23886 75022 23938
rect 76738 23886 76750 23938
rect 76802 23886 76814 23938
rect 78530 23886 78542 23938
rect 78594 23886 78606 23938
rect 86818 23886 86830 23938
rect 86882 23886 86894 23938
rect 73614 23874 73666 23886
rect 75630 23874 75682 23886
rect 27470 23826 27522 23838
rect 28254 23826 28306 23838
rect 28130 23774 28142 23826
rect 28194 23774 28206 23826
rect 27470 23762 27522 23774
rect 28254 23762 28306 23774
rect 28366 23826 28418 23838
rect 40462 23826 40514 23838
rect 31826 23774 31838 23826
rect 31890 23774 31902 23826
rect 28366 23762 28418 23774
rect 40462 23762 40514 23774
rect 45390 23826 45442 23838
rect 45390 23762 45442 23774
rect 45502 23826 45554 23838
rect 46286 23826 46338 23838
rect 60958 23826 61010 23838
rect 46050 23774 46062 23826
rect 46114 23774 46126 23826
rect 54786 23774 54798 23826
rect 54850 23774 54862 23826
rect 45502 23762 45554 23774
rect 46286 23762 46338 23774
rect 60958 23762 61010 23774
rect 68798 23826 68850 23838
rect 68798 23762 68850 23774
rect 69358 23826 69410 23838
rect 74162 23774 74174 23826
rect 74226 23774 74238 23826
rect 80322 23774 80334 23826
rect 80386 23774 80398 23826
rect 69358 23762 69410 23774
rect 27022 23714 27074 23726
rect 27022 23650 27074 23662
rect 27246 23714 27298 23726
rect 27246 23650 27298 23662
rect 28590 23714 28642 23726
rect 28590 23650 28642 23662
rect 34414 23714 34466 23726
rect 34414 23650 34466 23662
rect 35086 23714 35138 23726
rect 35086 23650 35138 23662
rect 39454 23714 39506 23726
rect 39454 23650 39506 23662
rect 42814 23714 42866 23726
rect 42814 23650 42866 23662
rect 45726 23714 45778 23726
rect 45726 23650 45778 23662
rect 47406 23714 47458 23726
rect 47406 23650 47458 23662
rect 48190 23714 48242 23726
rect 48190 23650 48242 23662
rect 50878 23714 50930 23726
rect 50878 23650 50930 23662
rect 51662 23714 51714 23726
rect 51662 23650 51714 23662
rect 53678 23714 53730 23726
rect 53678 23650 53730 23662
rect 53902 23714 53954 23726
rect 59390 23714 59442 23726
rect 54898 23662 54910 23714
rect 54962 23662 54974 23714
rect 53902 23650 53954 23662
rect 59390 23650 59442 23662
rect 61070 23714 61122 23726
rect 61070 23650 61122 23662
rect 61294 23714 61346 23726
rect 61294 23650 61346 23662
rect 68574 23714 68626 23726
rect 92654 23714 92706 23726
rect 75058 23662 75070 23714
rect 75122 23662 75134 23714
rect 76514 23662 76526 23714
rect 76578 23662 76590 23714
rect 86594 23662 86606 23714
rect 86658 23662 86670 23714
rect 68574 23650 68626 23662
rect 92654 23650 92706 23662
rect 93214 23714 93266 23726
rect 93214 23650 93266 23662
rect 1344 23546 158592 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 81278 23546
rect 81330 23494 81382 23546
rect 81434 23494 81486 23546
rect 81538 23494 111998 23546
rect 112050 23494 112102 23546
rect 112154 23494 112206 23546
rect 112258 23494 142718 23546
rect 142770 23494 142822 23546
rect 142874 23494 142926 23546
rect 142978 23494 158592 23546
rect 1344 23460 158592 23494
rect 25342 23378 25394 23390
rect 25342 23314 25394 23326
rect 27806 23378 27858 23390
rect 42030 23378 42082 23390
rect 38322 23326 38334 23378
rect 38386 23326 38398 23378
rect 27806 23314 27858 23326
rect 42030 23314 42082 23326
rect 43374 23378 43426 23390
rect 43374 23314 43426 23326
rect 43710 23378 43762 23390
rect 43710 23314 43762 23326
rect 44606 23378 44658 23390
rect 44606 23314 44658 23326
rect 45054 23378 45106 23390
rect 45054 23314 45106 23326
rect 45166 23378 45218 23390
rect 45166 23314 45218 23326
rect 50878 23378 50930 23390
rect 50878 23314 50930 23326
rect 51326 23378 51378 23390
rect 51326 23314 51378 23326
rect 51550 23378 51602 23390
rect 51550 23314 51602 23326
rect 78654 23378 78706 23390
rect 78654 23314 78706 23326
rect 81566 23378 81618 23390
rect 81566 23314 81618 23326
rect 82574 23378 82626 23390
rect 82574 23314 82626 23326
rect 33518 23266 33570 23278
rect 33518 23202 33570 23214
rect 34078 23266 34130 23278
rect 34078 23202 34130 23214
rect 41022 23266 41074 23278
rect 41022 23202 41074 23214
rect 42142 23266 42194 23278
rect 44158 23266 44210 23278
rect 53678 23266 53730 23278
rect 42354 23214 42366 23266
rect 42418 23214 42430 23266
rect 46386 23214 46398 23266
rect 46450 23214 46462 23266
rect 46946 23214 46958 23266
rect 47010 23214 47022 23266
rect 42142 23202 42194 23214
rect 44158 23202 44210 23214
rect 53678 23202 53730 23214
rect 53790 23266 53842 23278
rect 57822 23266 57874 23278
rect 54674 23214 54686 23266
rect 54738 23214 54750 23266
rect 53790 23202 53842 23214
rect 57822 23202 57874 23214
rect 58382 23266 58434 23278
rect 58382 23202 58434 23214
rect 59054 23266 59106 23278
rect 59054 23202 59106 23214
rect 64654 23266 64706 23278
rect 64654 23202 64706 23214
rect 65550 23266 65602 23278
rect 65550 23202 65602 23214
rect 65774 23266 65826 23278
rect 65774 23202 65826 23214
rect 80222 23266 80274 23278
rect 81790 23266 81842 23278
rect 80882 23214 80894 23266
rect 80946 23214 80958 23266
rect 80222 23202 80274 23214
rect 81790 23202 81842 23214
rect 86382 23266 86434 23278
rect 86382 23202 86434 23214
rect 93326 23266 93378 23278
rect 93326 23202 93378 23214
rect 25454 23154 25506 23166
rect 21858 23102 21870 23154
rect 21922 23102 21934 23154
rect 25454 23090 25506 23102
rect 27694 23154 27746 23166
rect 27694 23090 27746 23102
rect 33294 23154 33346 23166
rect 33294 23090 33346 23102
rect 33630 23154 33682 23166
rect 33630 23090 33682 23102
rect 33966 23154 34018 23166
rect 40798 23154 40850 23166
rect 38546 23102 38558 23154
rect 38610 23102 38622 23154
rect 33966 23090 34018 23102
rect 40798 23090 40850 23102
rect 41134 23154 41186 23166
rect 41134 23090 41186 23102
rect 41470 23154 41522 23166
rect 41470 23090 41522 23102
rect 41806 23154 41858 23166
rect 41806 23090 41858 23102
rect 43486 23154 43538 23166
rect 43486 23090 43538 23102
rect 43934 23154 43986 23166
rect 43934 23090 43986 23102
rect 45278 23154 45330 23166
rect 46622 23154 46674 23166
rect 50318 23154 50370 23166
rect 45602 23102 45614 23154
rect 45666 23102 45678 23154
rect 46274 23102 46286 23154
rect 46338 23102 46350 23154
rect 47170 23102 47182 23154
rect 47234 23102 47246 23154
rect 47730 23102 47742 23154
rect 47794 23102 47806 23154
rect 49858 23102 49870 23154
rect 49922 23102 49934 23154
rect 50082 23102 50094 23154
rect 50146 23102 50158 23154
rect 45278 23090 45330 23102
rect 46622 23090 46674 23102
rect 50318 23090 50370 23102
rect 50766 23154 50818 23166
rect 50766 23090 50818 23102
rect 50990 23154 51042 23166
rect 50990 23090 51042 23102
rect 52782 23154 52834 23166
rect 52782 23090 52834 23102
rect 52894 23154 52946 23166
rect 52894 23090 52946 23102
rect 53118 23154 53170 23166
rect 54014 23154 54066 23166
rect 56814 23154 56866 23166
rect 53330 23102 53342 23154
rect 53394 23102 53406 23154
rect 55010 23102 55022 23154
rect 55074 23102 55086 23154
rect 55682 23102 55694 23154
rect 55746 23102 55758 23154
rect 53118 23090 53170 23102
rect 54014 23090 54066 23102
rect 56814 23090 56866 23102
rect 56926 23154 56978 23166
rect 56926 23090 56978 23102
rect 58606 23154 58658 23166
rect 58606 23090 58658 23102
rect 58830 23154 58882 23166
rect 58830 23090 58882 23102
rect 59838 23154 59890 23166
rect 75742 23154 75794 23166
rect 60274 23102 60286 23154
rect 60338 23102 60350 23154
rect 72482 23102 72494 23154
rect 72546 23102 72558 23154
rect 73042 23102 73054 23154
rect 73106 23102 73118 23154
rect 59838 23090 59890 23102
rect 75742 23090 75794 23102
rect 76078 23154 76130 23166
rect 76078 23090 76130 23102
rect 76302 23154 76354 23166
rect 76302 23090 76354 23102
rect 78430 23154 78482 23166
rect 78430 23090 78482 23102
rect 78878 23154 78930 23166
rect 78878 23090 78930 23102
rect 78990 23154 79042 23166
rect 81118 23154 81170 23166
rect 80658 23102 80670 23154
rect 80722 23102 80734 23154
rect 78990 23090 79042 23102
rect 81118 23090 81170 23102
rect 82126 23154 82178 23166
rect 82126 23090 82178 23102
rect 82462 23154 82514 23166
rect 82462 23090 82514 23102
rect 82686 23154 82738 23166
rect 82686 23090 82738 23102
rect 82910 23154 82962 23166
rect 82910 23090 82962 23102
rect 83358 23154 83410 23166
rect 83358 23090 83410 23102
rect 83582 23154 83634 23166
rect 83582 23090 83634 23102
rect 86718 23154 86770 23166
rect 86718 23090 86770 23102
rect 86942 23154 86994 23166
rect 92878 23154 92930 23166
rect 89730 23102 89742 23154
rect 89794 23102 89806 23154
rect 90290 23102 90302 23154
rect 90354 23102 90366 23154
rect 86942 23090 86994 23102
rect 92878 23090 92930 23102
rect 93550 23154 93602 23166
rect 93550 23090 93602 23102
rect 25902 23042 25954 23054
rect 49086 23042 49138 23054
rect 22530 22990 22542 23042
rect 22594 22990 22606 23042
rect 24658 22990 24670 23042
rect 24722 22990 24734 23042
rect 42578 22990 42590 23042
rect 42642 22990 42654 23042
rect 25902 22978 25954 22990
rect 49086 22978 49138 22990
rect 49534 23042 49586 23054
rect 49534 22978 49586 22990
rect 50542 23042 50594 23054
rect 50542 22978 50594 22990
rect 52334 23042 52386 23054
rect 52334 22978 52386 22990
rect 53006 23042 53058 23054
rect 53006 22978 53058 22990
rect 54350 23042 54402 23054
rect 56590 23042 56642 23054
rect 55346 22990 55358 23042
rect 55410 22990 55422 23042
rect 54350 22978 54402 22990
rect 56590 22978 56642 22990
rect 59166 23042 59218 23054
rect 63086 23042 63138 23054
rect 60946 22990 60958 23042
rect 61010 22990 61022 23042
rect 59166 22978 59218 22990
rect 63086 22978 63138 22990
rect 63870 23042 63922 23054
rect 76190 23042 76242 23054
rect 64754 22990 64766 23042
rect 64818 22990 64830 23042
rect 65426 22990 65438 23042
rect 65490 22990 65502 23042
rect 75394 22990 75406 23042
rect 75458 22990 75470 23042
rect 63870 22978 63922 22990
rect 76190 22978 76242 22990
rect 79550 23042 79602 23054
rect 79550 22978 79602 22990
rect 81678 23042 81730 23054
rect 81678 22978 81730 22990
rect 83134 23042 83186 23054
rect 83134 22978 83186 22990
rect 84030 23042 84082 23054
rect 84030 22978 84082 22990
rect 84478 23042 84530 23054
rect 84478 22978 84530 22990
rect 86494 23042 86546 23054
rect 86494 22978 86546 22990
rect 87390 23042 87442 23054
rect 93102 23042 93154 23054
rect 92642 22990 92654 23042
rect 92706 22990 92718 23042
rect 87390 22978 87442 22990
rect 93102 22978 93154 22990
rect 25342 22930 25394 22942
rect 25342 22866 25394 22878
rect 27806 22930 27858 22942
rect 27806 22866 27858 22878
rect 34078 22930 34130 22942
rect 34078 22866 34130 22878
rect 51662 22930 51714 22942
rect 51662 22866 51714 22878
rect 64430 22930 64482 22942
rect 64430 22866 64482 22878
rect 80110 22930 80162 22942
rect 80110 22866 80162 22878
rect 1344 22762 158592 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 96638 22762
rect 96690 22710 96742 22762
rect 96794 22710 96846 22762
rect 96898 22710 127358 22762
rect 127410 22710 127462 22762
rect 127514 22710 127566 22762
rect 127618 22710 158078 22762
rect 158130 22710 158182 22762
rect 158234 22710 158286 22762
rect 158338 22710 158592 22762
rect 1344 22676 158592 22710
rect 51326 22594 51378 22606
rect 51326 22530 51378 22542
rect 32734 22482 32786 22494
rect 40350 22482 40402 22494
rect 23314 22430 23326 22482
rect 23378 22430 23390 22482
rect 36418 22430 36430 22482
rect 36482 22430 36494 22482
rect 36978 22430 36990 22482
rect 37042 22430 37054 22482
rect 32734 22418 32786 22430
rect 40350 22418 40402 22430
rect 42702 22482 42754 22494
rect 51438 22482 51490 22494
rect 47058 22430 47070 22482
rect 47122 22430 47134 22482
rect 42702 22418 42754 22430
rect 51438 22418 51490 22430
rect 52222 22482 52274 22494
rect 60622 22482 60674 22494
rect 74622 22482 74674 22494
rect 57026 22430 57038 22482
rect 57090 22430 57102 22482
rect 68338 22430 68350 22482
rect 68402 22430 68414 22482
rect 52222 22418 52274 22430
rect 60622 22418 60674 22430
rect 74622 22418 74674 22430
rect 75630 22482 75682 22494
rect 75630 22418 75682 22430
rect 79102 22482 79154 22494
rect 79102 22418 79154 22430
rect 84142 22482 84194 22494
rect 84142 22418 84194 22430
rect 85262 22482 85314 22494
rect 85262 22418 85314 22430
rect 90750 22482 90802 22494
rect 90750 22418 90802 22430
rect 91982 22482 92034 22494
rect 91982 22418 92034 22430
rect 29374 22370 29426 22382
rect 29374 22306 29426 22318
rect 32510 22370 32562 22382
rect 32510 22306 32562 22318
rect 32958 22370 33010 22382
rect 42590 22370 42642 22382
rect 33618 22318 33630 22370
rect 33682 22318 33694 22370
rect 39778 22318 39790 22370
rect 39842 22318 39854 22370
rect 32958 22306 33010 22318
rect 42590 22306 42642 22318
rect 43710 22370 43762 22382
rect 43710 22306 43762 22318
rect 45054 22370 45106 22382
rect 60062 22370 60114 22382
rect 50978 22318 50990 22370
rect 51042 22318 51054 22370
rect 52658 22318 52670 22370
rect 52722 22318 52734 22370
rect 45054 22306 45106 22318
rect 60062 22306 60114 22318
rect 60398 22370 60450 22382
rect 60398 22306 60450 22318
rect 60846 22370 60898 22382
rect 60846 22306 60898 22318
rect 60958 22370 61010 22382
rect 74734 22370 74786 22382
rect 71250 22318 71262 22370
rect 71314 22318 71326 22370
rect 60958 22306 61010 22318
rect 74734 22306 74786 22318
rect 75182 22370 75234 22382
rect 90526 22370 90578 22382
rect 82898 22318 82910 22370
rect 82962 22318 82974 22370
rect 83458 22318 83470 22370
rect 83522 22318 83534 22370
rect 85474 22318 85486 22370
rect 85538 22318 85550 22370
rect 86258 22318 86270 22370
rect 86322 22318 86334 22370
rect 75182 22306 75234 22318
rect 90526 22306 90578 22318
rect 91198 22370 91250 22382
rect 91198 22306 91250 22318
rect 92542 22370 92594 22382
rect 95330 22318 95342 22370
rect 95394 22318 95406 22370
rect 96114 22318 96126 22370
rect 96178 22318 96190 22370
rect 99810 22318 99822 22370
rect 99874 22318 99886 22370
rect 92542 22306 92594 22318
rect 23774 22258 23826 22270
rect 23650 22206 23662 22258
rect 23714 22206 23726 22258
rect 23774 22194 23826 22206
rect 23886 22258 23938 22270
rect 23886 22194 23938 22206
rect 28030 22258 28082 22270
rect 29038 22258 29090 22270
rect 28130 22206 28142 22258
rect 28194 22206 28206 22258
rect 28030 22194 28082 22206
rect 29038 22194 29090 22206
rect 33182 22258 33234 22270
rect 43150 22258 43202 22270
rect 34290 22206 34302 22258
rect 34354 22206 34366 22258
rect 39106 22206 39118 22258
rect 39170 22206 39182 22258
rect 33182 22194 33234 22206
rect 43150 22194 43202 22206
rect 43486 22258 43538 22270
rect 43486 22194 43538 22206
rect 51550 22258 51602 22270
rect 59726 22258 59778 22270
rect 58258 22206 58270 22258
rect 58322 22206 58334 22258
rect 51550 22194 51602 22206
rect 59726 22194 59778 22206
rect 59838 22258 59890 22270
rect 90302 22258 90354 22270
rect 70466 22206 70478 22258
rect 70530 22206 70542 22258
rect 59838 22194 59890 22206
rect 90302 22194 90354 22206
rect 90974 22258 91026 22270
rect 103506 22206 103518 22258
rect 103570 22206 103582 22258
rect 90974 22194 91026 22206
rect 24110 22146 24162 22158
rect 24110 22082 24162 22094
rect 27694 22146 27746 22158
rect 27694 22082 27746 22094
rect 27806 22146 27858 22158
rect 27806 22082 27858 22094
rect 27918 22146 27970 22158
rect 27918 22082 27970 22094
rect 29262 22146 29314 22158
rect 29262 22082 29314 22094
rect 29822 22146 29874 22158
rect 29822 22082 29874 22094
rect 42366 22146 42418 22158
rect 42366 22082 42418 22094
rect 42814 22146 42866 22158
rect 42814 22082 42866 22094
rect 43374 22146 43426 22158
rect 58606 22146 58658 22158
rect 45378 22094 45390 22146
rect 45442 22094 45454 22146
rect 43374 22082 43426 22094
rect 58606 22082 58658 22094
rect 59390 22146 59442 22158
rect 59390 22082 59442 22094
rect 65102 22146 65154 22158
rect 65102 22082 65154 22094
rect 71710 22146 71762 22158
rect 71710 22082 71762 22094
rect 74510 22146 74562 22158
rect 74510 22082 74562 22094
rect 78990 22146 79042 22158
rect 91870 22146 91922 22158
rect 80434 22094 80446 22146
rect 80498 22094 80510 22146
rect 88610 22094 88622 22146
rect 88674 22094 88686 22146
rect 78990 22082 79042 22094
rect 91870 22082 91922 22094
rect 92094 22146 92146 22158
rect 96462 22146 96514 22158
rect 92978 22094 92990 22146
rect 93042 22094 93054 22146
rect 92094 22082 92146 22094
rect 96462 22082 96514 22094
rect 1344 21978 158592 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 81278 21978
rect 81330 21926 81382 21978
rect 81434 21926 81486 21978
rect 81538 21926 111998 21978
rect 112050 21926 112102 21978
rect 112154 21926 112206 21978
rect 112258 21926 142718 21978
rect 142770 21926 142822 21978
rect 142874 21926 142926 21978
rect 142978 21926 158592 21978
rect 1344 21892 158592 21926
rect 43486 21810 43538 21822
rect 26002 21758 26014 21810
rect 26066 21758 26078 21810
rect 43486 21746 43538 21758
rect 47406 21810 47458 21822
rect 47406 21746 47458 21758
rect 47742 21810 47794 21822
rect 47742 21746 47794 21758
rect 47966 21810 48018 21822
rect 47966 21746 48018 21758
rect 49310 21810 49362 21822
rect 49310 21746 49362 21758
rect 50318 21810 50370 21822
rect 50318 21746 50370 21758
rect 52894 21810 52946 21822
rect 52894 21746 52946 21758
rect 53118 21810 53170 21822
rect 57150 21810 57202 21822
rect 55122 21758 55134 21810
rect 55186 21758 55198 21810
rect 53118 21746 53170 21758
rect 57150 21746 57202 21758
rect 59614 21810 59666 21822
rect 59614 21746 59666 21758
rect 60846 21810 60898 21822
rect 60846 21746 60898 21758
rect 80222 21810 80274 21822
rect 80222 21746 80274 21758
rect 82014 21810 82066 21822
rect 82014 21746 82066 21758
rect 82126 21810 82178 21822
rect 82126 21746 82178 21758
rect 86494 21810 86546 21822
rect 86494 21746 86546 21758
rect 86830 21810 86882 21822
rect 86830 21746 86882 21758
rect 88398 21810 88450 21822
rect 88398 21746 88450 21758
rect 93886 21810 93938 21822
rect 93886 21746 93938 21758
rect 98030 21810 98082 21822
rect 98030 21746 98082 21758
rect 24446 21698 24498 21710
rect 31614 21698 31666 21710
rect 27458 21646 27470 21698
rect 27522 21646 27534 21698
rect 24446 21634 24498 21646
rect 31614 21634 31666 21646
rect 33406 21698 33458 21710
rect 33406 21634 33458 21646
rect 34414 21698 34466 21710
rect 47294 21698 47346 21710
rect 42690 21646 42702 21698
rect 42754 21695 42766 21698
rect 42914 21695 42926 21698
rect 42754 21649 42926 21695
rect 42754 21646 42766 21649
rect 42914 21646 42926 21649
rect 42978 21646 42990 21698
rect 46610 21646 46622 21698
rect 46674 21646 46686 21698
rect 34414 21634 34466 21646
rect 47294 21634 47346 21646
rect 47630 21698 47682 21710
rect 47630 21634 47682 21646
rect 51102 21698 51154 21710
rect 60062 21698 60114 21710
rect 51102 21634 51154 21646
rect 52782 21642 52834 21654
rect 55794 21646 55806 21698
rect 55858 21646 55870 21698
rect 24222 21586 24274 21598
rect 21074 21534 21086 21586
rect 21138 21534 21150 21586
rect 24222 21522 24274 21534
rect 24558 21586 24610 21598
rect 24558 21522 24610 21534
rect 26350 21586 26402 21598
rect 31390 21586 31442 21598
rect 26674 21534 26686 21586
rect 26738 21534 26750 21586
rect 26350 21522 26402 21534
rect 31390 21522 31442 21534
rect 31726 21586 31778 21598
rect 31726 21522 31778 21534
rect 33742 21586 33794 21598
rect 33742 21522 33794 21534
rect 34078 21586 34130 21598
rect 34078 21522 34130 21534
rect 41694 21586 41746 21598
rect 46286 21586 46338 21598
rect 42018 21534 42030 21586
rect 42082 21534 42094 21586
rect 41694 21522 41746 21534
rect 46286 21522 46338 21534
rect 50542 21586 50594 21598
rect 50542 21522 50594 21534
rect 50990 21586 51042 21598
rect 50990 21522 51042 21534
rect 51214 21586 51266 21598
rect 60062 21634 60114 21646
rect 73838 21698 73890 21710
rect 88510 21698 88562 21710
rect 86146 21646 86158 21698
rect 86210 21646 86222 21698
rect 87154 21646 87166 21698
rect 87218 21646 87230 21698
rect 73838 21634 73890 21646
rect 88510 21634 88562 21646
rect 93774 21698 93826 21710
rect 93774 21634 93826 21646
rect 97470 21698 97522 21710
rect 97470 21634 97522 21646
rect 98142 21698 98194 21710
rect 108994 21646 109006 21698
rect 109058 21646 109070 21698
rect 98142 21634 98194 21646
rect 51650 21534 51662 21586
rect 51714 21534 51726 21586
rect 52322 21534 52334 21586
rect 52386 21534 52398 21586
rect 52782 21578 52834 21590
rect 54014 21586 54066 21598
rect 51214 21522 51266 21534
rect 54014 21522 54066 21534
rect 54238 21586 54290 21598
rect 56590 21586 56642 21598
rect 54898 21534 54910 21586
rect 54962 21534 54974 21586
rect 55458 21534 55470 21586
rect 55522 21534 55534 21586
rect 54238 21522 54290 21534
rect 56590 21522 56642 21534
rect 59054 21586 59106 21598
rect 59054 21522 59106 21534
rect 59502 21586 59554 21598
rect 59502 21522 59554 21534
rect 59726 21586 59778 21598
rect 60510 21586 60562 21598
rect 69470 21586 69522 21598
rect 60274 21534 60286 21586
rect 60338 21534 60350 21586
rect 60722 21534 60734 21586
rect 60786 21534 60798 21586
rect 67330 21534 67342 21586
rect 67394 21534 67406 21586
rect 59726 21522 59778 21534
rect 60510 21522 60562 21534
rect 69470 21522 69522 21534
rect 74174 21586 74226 21598
rect 74174 21522 74226 21534
rect 74398 21586 74450 21598
rect 74398 21522 74450 21534
rect 74958 21586 75010 21598
rect 81566 21586 81618 21598
rect 76402 21534 76414 21586
rect 76466 21534 76478 21586
rect 77186 21534 77198 21586
rect 77250 21534 77262 21586
rect 74958 21522 75010 21534
rect 81566 21522 81618 21534
rect 82238 21586 82290 21598
rect 82238 21522 82290 21534
rect 87838 21586 87890 21598
rect 87838 21522 87890 21534
rect 88286 21586 88338 21598
rect 93998 21586 94050 21598
rect 90514 21534 90526 21586
rect 90578 21534 90590 21586
rect 91074 21534 91086 21586
rect 91138 21534 91150 21586
rect 88286 21522 88338 21534
rect 93998 21522 94050 21534
rect 94446 21586 94498 21598
rect 94446 21522 94498 21534
rect 97694 21586 97746 21598
rect 97694 21522 97746 21534
rect 98254 21586 98306 21598
rect 108670 21586 108722 21598
rect 104402 21534 104414 21586
rect 104466 21534 104478 21586
rect 98254 21522 98306 21534
rect 108670 21522 108722 21534
rect 30046 21474 30098 21486
rect 21858 21422 21870 21474
rect 21922 21422 21934 21474
rect 23986 21422 23998 21474
rect 24050 21422 24062 21474
rect 29586 21422 29598 21474
rect 29650 21422 29662 21474
rect 30046 21410 30098 21422
rect 32286 21474 32338 21486
rect 32286 21410 32338 21422
rect 33966 21474 34018 21486
rect 33966 21410 34018 21422
rect 34862 21474 34914 21486
rect 34862 21410 34914 21422
rect 36654 21474 36706 21486
rect 36654 21410 36706 21422
rect 41470 21474 41522 21486
rect 41470 21410 41522 21422
rect 43038 21474 43090 21486
rect 43038 21410 43090 21422
rect 44046 21474 44098 21486
rect 44046 21410 44098 21422
rect 47070 21474 47122 21486
rect 47070 21410 47122 21422
rect 48862 21474 48914 21486
rect 48862 21410 48914 21422
rect 49982 21474 50034 21486
rect 67790 21474 67842 21486
rect 51762 21422 51774 21474
rect 51826 21422 51838 21474
rect 52770 21422 52782 21474
rect 52834 21422 52846 21474
rect 64418 21422 64430 21474
rect 64482 21422 64494 21474
rect 66546 21422 66558 21474
rect 66610 21422 66622 21474
rect 49982 21410 50034 21422
rect 67790 21410 67842 21422
rect 68910 21474 68962 21486
rect 68910 21410 68962 21422
rect 73950 21474 74002 21486
rect 73950 21410 74002 21422
rect 75406 21474 75458 21486
rect 103070 21474 103122 21486
rect 79538 21422 79550 21474
rect 79602 21422 79614 21474
rect 93426 21422 93438 21474
rect 93490 21422 93502 21474
rect 75406 21410 75458 21422
rect 103070 21410 103122 21422
rect 103966 21474 104018 21486
rect 103966 21410 104018 21422
rect 108334 21474 108386 21486
rect 108334 21410 108386 21422
rect 46846 21362 46898 21374
rect 51998 21362 52050 21374
rect 74846 21362 74898 21374
rect 42690 21310 42702 21362
rect 42754 21359 42766 21362
rect 43138 21359 43150 21362
rect 42754 21313 43150 21359
rect 42754 21310 42766 21313
rect 43138 21310 43150 21313
rect 43202 21310 43214 21362
rect 48962 21310 48974 21362
rect 49026 21359 49038 21362
rect 49634 21359 49646 21362
rect 49026 21313 49646 21359
rect 49026 21310 49038 21313
rect 49634 21310 49646 21313
rect 49698 21359 49710 21362
rect 49858 21359 49870 21362
rect 49698 21313 49870 21359
rect 49698 21310 49710 21313
rect 49858 21310 49870 21313
rect 49922 21310 49934 21362
rect 53666 21310 53678 21362
rect 53730 21310 53742 21362
rect 46846 21298 46898 21310
rect 51998 21298 52050 21310
rect 74846 21298 74898 21310
rect 1344 21194 158592 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 96638 21194
rect 96690 21142 96742 21194
rect 96794 21142 96846 21194
rect 96898 21142 127358 21194
rect 127410 21142 127462 21194
rect 127514 21142 127566 21194
rect 127618 21142 158078 21194
rect 158130 21142 158182 21194
rect 158234 21142 158286 21194
rect 158338 21142 158592 21194
rect 1344 21108 158592 21142
rect 27582 21026 27634 21038
rect 27582 20962 27634 20974
rect 46398 21026 46450 21038
rect 46398 20962 46450 20974
rect 50206 21026 50258 21038
rect 50206 20962 50258 20974
rect 50654 21026 50706 21038
rect 50654 20962 50706 20974
rect 24558 20914 24610 20926
rect 23314 20862 23326 20914
rect 23378 20862 23390 20914
rect 24558 20850 24610 20862
rect 25006 20914 25058 20926
rect 25006 20850 25058 20862
rect 38558 20914 38610 20926
rect 53678 20914 53730 20926
rect 42018 20862 42030 20914
rect 42082 20862 42094 20914
rect 52098 20862 52110 20914
rect 52162 20862 52174 20914
rect 38558 20850 38610 20862
rect 53678 20850 53730 20862
rect 57374 20914 57426 20926
rect 57374 20850 57426 20862
rect 58270 20914 58322 20926
rect 58270 20850 58322 20862
rect 59838 20914 59890 20926
rect 59838 20850 59890 20862
rect 59950 20914 60002 20926
rect 59950 20850 60002 20862
rect 60510 20914 60562 20926
rect 60510 20850 60562 20862
rect 77534 20914 77586 20926
rect 77534 20850 77586 20862
rect 78430 20914 78482 20926
rect 78430 20850 78482 20862
rect 79326 20914 79378 20926
rect 79326 20850 79378 20862
rect 81454 20914 81506 20926
rect 81454 20850 81506 20862
rect 88734 20914 88786 20926
rect 88734 20850 88786 20862
rect 91310 20914 91362 20926
rect 91310 20850 91362 20862
rect 91982 20914 92034 20926
rect 91982 20850 92034 20862
rect 24110 20802 24162 20814
rect 30046 20802 30098 20814
rect 36878 20802 36930 20814
rect 26674 20750 26686 20802
rect 26738 20750 26750 20802
rect 28578 20750 28590 20802
rect 28642 20750 28654 20802
rect 29362 20750 29374 20802
rect 29426 20750 29438 20802
rect 31826 20750 31838 20802
rect 31890 20750 31902 20802
rect 24110 20738 24162 20750
rect 30046 20738 30098 20750
rect 36878 20738 36930 20750
rect 37326 20802 37378 20814
rect 37326 20738 37378 20750
rect 37774 20802 37826 20814
rect 42702 20802 42754 20814
rect 41794 20750 41806 20802
rect 41858 20750 41870 20802
rect 37774 20738 37826 20750
rect 42702 20738 42754 20750
rect 45054 20802 45106 20814
rect 45054 20738 45106 20750
rect 45390 20802 45442 20814
rect 45390 20738 45442 20750
rect 45614 20802 45666 20814
rect 47406 20802 47458 20814
rect 49534 20802 49586 20814
rect 51326 20802 51378 20814
rect 45938 20750 45950 20802
rect 46002 20750 46014 20802
rect 47730 20750 47742 20802
rect 47794 20750 47806 20802
rect 48962 20750 48974 20802
rect 49026 20750 49038 20802
rect 49298 20750 49310 20802
rect 49362 20750 49374 20802
rect 49858 20750 49870 20802
rect 49922 20750 49934 20802
rect 45614 20738 45666 20750
rect 47406 20738 47458 20750
rect 49534 20738 49586 20750
rect 51326 20738 51378 20750
rect 52558 20802 52610 20814
rect 54798 20802 54850 20814
rect 54338 20750 54350 20802
rect 54402 20750 54414 20802
rect 52558 20738 52610 20750
rect 54798 20738 54850 20750
rect 55918 20802 55970 20814
rect 59054 20802 59106 20814
rect 56354 20750 56366 20802
rect 56418 20750 56430 20802
rect 55918 20738 55970 20750
rect 59054 20738 59106 20750
rect 59390 20802 59442 20814
rect 60622 20802 60674 20814
rect 63310 20802 63362 20814
rect 63870 20802 63922 20814
rect 59602 20750 59614 20802
rect 59666 20750 59678 20802
rect 60946 20750 60958 20802
rect 61010 20750 61022 20802
rect 63634 20750 63646 20802
rect 63698 20750 63710 20802
rect 59390 20738 59442 20750
rect 60622 20738 60674 20750
rect 63310 20738 63362 20750
rect 63870 20738 63922 20750
rect 64094 20802 64146 20814
rect 65214 20802 65266 20814
rect 77086 20802 77138 20814
rect 64754 20750 64766 20802
rect 64818 20750 64830 20802
rect 65538 20750 65550 20802
rect 65602 20750 65614 20802
rect 66994 20750 67006 20802
rect 67058 20750 67070 20802
rect 72034 20750 72046 20802
rect 72098 20750 72110 20802
rect 72818 20750 72830 20802
rect 72882 20750 72894 20802
rect 64094 20738 64146 20750
rect 65214 20738 65266 20750
rect 77086 20738 77138 20750
rect 77758 20802 77810 20814
rect 77758 20738 77810 20750
rect 77982 20802 78034 20814
rect 77982 20738 78034 20750
rect 78542 20802 78594 20814
rect 91870 20802 91922 20814
rect 87602 20750 87614 20802
rect 87666 20750 87678 20802
rect 88386 20750 88398 20802
rect 88450 20750 88462 20802
rect 78542 20738 78594 20750
rect 91870 20738 91922 20750
rect 92094 20802 92146 20814
rect 92094 20738 92146 20750
rect 92430 20802 92482 20814
rect 92430 20738 92482 20750
rect 92878 20802 92930 20814
rect 92878 20738 92930 20750
rect 93438 20802 93490 20814
rect 95554 20750 95566 20802
rect 95618 20750 95630 20802
rect 96338 20750 96350 20802
rect 96402 20750 96414 20802
rect 103506 20750 103518 20802
rect 103570 20750 103582 20802
rect 104290 20750 104302 20802
rect 104354 20750 104366 20802
rect 108210 20750 108222 20802
rect 108274 20750 108286 20802
rect 108994 20750 109006 20802
rect 109058 20750 109070 20802
rect 111682 20750 111694 20802
rect 111746 20750 111758 20802
rect 112354 20750 112366 20802
rect 112418 20750 112430 20802
rect 93438 20738 93490 20750
rect 23774 20690 23826 20702
rect 37550 20690 37602 20702
rect 23650 20638 23662 20690
rect 23714 20638 23726 20690
rect 29138 20638 29150 20690
rect 29202 20638 29214 20690
rect 34738 20638 34750 20690
rect 34802 20638 34814 20690
rect 23774 20626 23826 20638
rect 37550 20626 37602 20638
rect 37998 20690 38050 20702
rect 37998 20626 38050 20638
rect 38110 20690 38162 20702
rect 46846 20690 46898 20702
rect 50094 20690 50146 20702
rect 45826 20638 45838 20690
rect 45890 20638 45902 20690
rect 48178 20638 48190 20690
rect 48242 20638 48254 20690
rect 48514 20638 48526 20690
rect 48578 20638 48590 20690
rect 38110 20626 38162 20638
rect 46846 20626 46898 20638
rect 50094 20626 50146 20638
rect 51662 20690 51714 20702
rect 53006 20690 53058 20702
rect 51762 20638 51774 20690
rect 51826 20638 51838 20690
rect 51662 20626 51714 20638
rect 53006 20626 53058 20638
rect 53230 20690 53282 20702
rect 64318 20690 64370 20702
rect 66558 20690 66610 20702
rect 55122 20638 55134 20690
rect 55186 20638 55198 20690
rect 65762 20638 65774 20690
rect 65826 20638 65838 20690
rect 66210 20638 66222 20690
rect 66274 20638 66286 20690
rect 53230 20626 53282 20638
rect 64318 20626 64370 20638
rect 66558 20626 66610 20638
rect 77422 20690 77474 20702
rect 77422 20626 77474 20638
rect 78766 20690 78818 20702
rect 78766 20626 78818 20638
rect 23886 20578 23938 20590
rect 30606 20578 30658 20590
rect 26450 20526 26462 20578
rect 26514 20526 26526 20578
rect 23886 20514 23938 20526
rect 30606 20514 30658 20526
rect 37214 20578 37266 20590
rect 37214 20514 37266 20526
rect 47070 20578 47122 20590
rect 47070 20514 47122 20526
rect 47294 20578 47346 20590
rect 47294 20514 47346 20526
rect 50766 20578 50818 20590
rect 50766 20514 50818 20526
rect 50878 20578 50930 20590
rect 50878 20514 50930 20526
rect 51550 20578 51602 20590
rect 51550 20514 51602 20526
rect 52894 20578 52946 20590
rect 56814 20578 56866 20590
rect 54114 20526 54126 20578
rect 54178 20526 54190 20578
rect 52894 20514 52946 20526
rect 56814 20514 56866 20526
rect 58830 20578 58882 20590
rect 58830 20514 58882 20526
rect 59166 20578 59218 20590
rect 59166 20514 59218 20526
rect 64430 20578 64482 20590
rect 75630 20578 75682 20590
rect 75170 20526 75182 20578
rect 75234 20526 75246 20578
rect 64430 20514 64482 20526
rect 75630 20514 75682 20526
rect 76526 20578 76578 20590
rect 76526 20514 76578 20526
rect 78318 20578 78370 20590
rect 78318 20514 78370 20526
rect 81566 20578 81618 20590
rect 92766 20578 92818 20590
rect 85250 20526 85262 20578
rect 85314 20526 85326 20578
rect 81566 20514 81618 20526
rect 92766 20514 92818 20526
rect 92990 20578 93042 20590
rect 92990 20514 93042 20526
rect 93774 20578 93826 20590
rect 99150 20578 99202 20590
rect 98690 20526 98702 20578
rect 98754 20526 98766 20578
rect 93774 20514 93826 20526
rect 99150 20514 99202 20526
rect 103294 20578 103346 20590
rect 107998 20578 108050 20590
rect 106642 20526 106654 20578
rect 106706 20526 106718 20578
rect 111346 20526 111358 20578
rect 111410 20526 111422 20578
rect 114818 20526 114830 20578
rect 114882 20526 114894 20578
rect 103294 20514 103346 20526
rect 107998 20514 108050 20526
rect 1344 20410 158592 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 81278 20410
rect 81330 20358 81382 20410
rect 81434 20358 81486 20410
rect 81538 20358 111998 20410
rect 112050 20358 112102 20410
rect 112154 20358 112206 20410
rect 112258 20358 142718 20410
rect 142770 20358 142822 20410
rect 142874 20358 142926 20410
rect 142978 20358 158592 20410
rect 1344 20324 158592 20358
rect 52558 20242 52610 20254
rect 52558 20178 52610 20190
rect 52782 20242 52834 20254
rect 52782 20178 52834 20190
rect 56478 20242 56530 20254
rect 56478 20178 56530 20190
rect 59390 20242 59442 20254
rect 59390 20178 59442 20190
rect 64430 20242 64482 20254
rect 64430 20178 64482 20190
rect 69694 20242 69746 20254
rect 69694 20178 69746 20190
rect 74734 20242 74786 20254
rect 74734 20178 74786 20190
rect 86270 20242 86322 20254
rect 86270 20178 86322 20190
rect 86942 20242 86994 20254
rect 86942 20178 86994 20190
rect 93662 20242 93714 20254
rect 93662 20178 93714 20190
rect 96574 20242 96626 20254
rect 96574 20178 96626 20190
rect 97582 20242 97634 20254
rect 97582 20178 97634 20190
rect 104750 20242 104802 20254
rect 104750 20178 104802 20190
rect 109006 20242 109058 20254
rect 109006 20178 109058 20190
rect 111582 20242 111634 20254
rect 111582 20178 111634 20190
rect 23326 20130 23378 20142
rect 26798 20130 26850 20142
rect 26450 20078 26462 20130
rect 26514 20078 26526 20130
rect 23326 20066 23378 20078
rect 26798 20066 26850 20078
rect 26910 20130 26962 20142
rect 26910 20066 26962 20078
rect 31390 20130 31442 20142
rect 34078 20130 34130 20142
rect 32274 20078 32286 20130
rect 32338 20078 32350 20130
rect 31390 20066 31442 20078
rect 34078 20066 34130 20078
rect 34190 20130 34242 20142
rect 34190 20066 34242 20078
rect 38334 20130 38386 20142
rect 38334 20066 38386 20078
rect 38446 20130 38498 20142
rect 38446 20066 38498 20078
rect 44270 20130 44322 20142
rect 44270 20066 44322 20078
rect 52894 20130 52946 20142
rect 56702 20130 56754 20142
rect 60958 20130 61010 20142
rect 52994 20078 53006 20130
rect 53058 20078 53070 20130
rect 60162 20078 60174 20130
rect 60226 20078 60238 20130
rect 52894 20066 52946 20078
rect 56702 20066 56754 20078
rect 60958 20066 61010 20078
rect 70366 20130 70418 20142
rect 70366 20066 70418 20078
rect 74062 20130 74114 20142
rect 74062 20066 74114 20078
rect 74622 20130 74674 20142
rect 74622 20066 74674 20078
rect 78094 20130 78146 20142
rect 78094 20066 78146 20078
rect 81790 20130 81842 20142
rect 81790 20066 81842 20078
rect 82238 20130 82290 20142
rect 82238 20066 82290 20078
rect 82574 20130 82626 20142
rect 82574 20066 82626 20078
rect 86046 20130 86098 20142
rect 95230 20130 95282 20142
rect 96798 20130 96850 20142
rect 87266 20078 87278 20130
rect 87330 20078 87342 20130
rect 96114 20078 96126 20130
rect 96178 20078 96190 20130
rect 86046 20066 86098 20078
rect 95230 20066 95282 20078
rect 96798 20066 96850 20078
rect 97806 20130 97858 20142
rect 97806 20066 97858 20078
rect 101838 20130 101890 20142
rect 101838 20066 101890 20078
rect 105870 20130 105922 20142
rect 105870 20066 105922 20078
rect 106094 20130 106146 20142
rect 107774 20130 107826 20142
rect 109454 20130 109506 20142
rect 106754 20078 106766 20130
rect 106818 20078 106830 20130
rect 108546 20078 108558 20130
rect 108610 20078 108622 20130
rect 106094 20066 106146 20078
rect 107774 20066 107826 20078
rect 109454 20066 109506 20078
rect 109902 20130 109954 20142
rect 109902 20066 109954 20078
rect 110238 20130 110290 20142
rect 110238 20066 110290 20078
rect 113374 20130 113426 20142
rect 113374 20066 113426 20078
rect 23102 20018 23154 20030
rect 19170 19966 19182 20018
rect 19234 19966 19246 20018
rect 23102 19954 23154 19966
rect 23438 20018 23490 20030
rect 30942 20018 30994 20030
rect 26226 19966 26238 20018
rect 26290 19966 26302 20018
rect 27794 19966 27806 20018
rect 27858 19966 27870 20018
rect 23438 19954 23490 19966
rect 30942 19954 30994 19966
rect 31614 20018 31666 20030
rect 31614 19954 31666 19966
rect 31950 20018 32002 20030
rect 31950 19954 32002 19966
rect 32958 20018 33010 20030
rect 32958 19954 33010 19966
rect 33406 20018 33458 20030
rect 33406 19954 33458 19966
rect 33630 20018 33682 20030
rect 33630 19954 33682 19966
rect 33854 20018 33906 20030
rect 33854 19954 33906 19966
rect 34750 20018 34802 20030
rect 41022 20018 41074 20030
rect 56814 20018 56866 20030
rect 69134 20018 69186 20030
rect 74510 20018 74562 20030
rect 35186 19966 35198 20018
rect 35250 19966 35262 20018
rect 43698 19966 43710 20018
rect 43762 19966 43774 20018
rect 51986 19966 51998 20018
rect 52050 19966 52062 20018
rect 59714 19966 59726 20018
rect 59778 19966 59790 20018
rect 61170 19966 61182 20018
rect 61234 19966 61246 20018
rect 67890 19966 67902 20018
rect 67954 19966 67966 20018
rect 70130 19966 70142 20018
rect 70194 19966 70206 20018
rect 34750 19954 34802 19966
rect 41022 19954 41074 19966
rect 56814 19954 56866 19966
rect 69134 19954 69186 19966
rect 74510 19954 74562 19966
rect 75182 20018 75234 20030
rect 75182 19954 75234 19966
rect 75406 20018 75458 20030
rect 75406 19954 75458 19966
rect 75966 20018 76018 20030
rect 75966 19954 76018 19966
rect 76302 20018 76354 20030
rect 80894 20018 80946 20030
rect 77298 19966 77310 20018
rect 77362 19966 77374 20018
rect 76302 19954 76354 19966
rect 80894 19954 80946 19966
rect 81230 20018 81282 20030
rect 81230 19954 81282 19966
rect 81566 20018 81618 20030
rect 81566 19954 81618 19966
rect 82126 20018 82178 20030
rect 82126 19954 82178 19966
rect 82350 20018 82402 20030
rect 82350 19954 82402 19966
rect 86382 20018 86434 20030
rect 86382 19954 86434 19966
rect 86606 20018 86658 20030
rect 95790 20018 95842 20030
rect 90290 19966 90302 20018
rect 90354 19966 90366 20018
rect 90850 19966 90862 20018
rect 90914 19966 90926 20018
rect 86606 19954 86658 19966
rect 95790 19954 95842 19966
rect 96462 20018 96514 20030
rect 96462 19954 96514 19966
rect 97022 20018 97074 20030
rect 97022 19954 97074 19966
rect 97358 20018 97410 20030
rect 97358 19954 97410 19966
rect 97470 20018 97522 20030
rect 104638 20018 104690 20030
rect 100818 19966 100830 20018
rect 100882 19966 100894 20018
rect 101266 19966 101278 20018
rect 101330 19966 101342 20018
rect 97470 19954 97522 19966
rect 104638 19954 104690 19966
rect 104974 20018 105026 20030
rect 104974 19954 105026 19966
rect 105198 20018 105250 20030
rect 105198 19954 105250 19966
rect 105422 20018 105474 20030
rect 105422 19954 105474 19966
rect 105982 20018 106034 20030
rect 105982 19954 106034 19966
rect 106430 20018 106482 20030
rect 106430 19954 106482 19966
rect 107214 20018 107266 20030
rect 107214 19954 107266 19966
rect 108222 20018 108274 20030
rect 108222 19954 108274 19966
rect 108782 20018 108834 20030
rect 108782 19954 108834 19966
rect 109118 20018 109170 20030
rect 109118 19954 109170 19966
rect 109790 20018 109842 20030
rect 109790 19954 109842 19966
rect 110014 20018 110066 20030
rect 110014 19954 110066 19966
rect 111918 20018 111970 20030
rect 111918 19954 111970 19966
rect 112366 20018 112418 20030
rect 112366 19954 112418 19966
rect 112590 20018 112642 20030
rect 112590 19954 112642 19966
rect 112926 20018 112978 20030
rect 112926 19954 112978 19966
rect 113262 20018 113314 20030
rect 113262 19954 113314 19966
rect 113486 20018 113538 20030
rect 113486 19954 113538 19966
rect 113934 20018 113986 20030
rect 113934 19954 113986 19966
rect 22430 19906 22482 19918
rect 31166 19906 31218 19918
rect 19842 19854 19854 19906
rect 19906 19854 19918 19906
rect 21970 19854 21982 19906
rect 22034 19854 22046 19906
rect 28578 19854 28590 19906
rect 28642 19854 28654 19906
rect 30706 19854 30718 19906
rect 30770 19854 30782 19906
rect 22430 19842 22482 19854
rect 31166 19842 31218 19854
rect 33182 19906 33234 19918
rect 39006 19906 39058 19918
rect 35858 19854 35870 19906
rect 35922 19854 35934 19906
rect 37986 19854 37998 19906
rect 38050 19854 38062 19906
rect 33182 19842 33234 19854
rect 39006 19842 39058 19854
rect 41582 19906 41634 19918
rect 53902 19906 53954 19918
rect 64542 19906 64594 19918
rect 68350 19906 68402 19918
rect 43362 19854 43374 19906
rect 43426 19854 43438 19906
rect 50978 19854 50990 19906
rect 51042 19854 51054 19906
rect 53330 19854 53342 19906
rect 53394 19854 53406 19906
rect 59826 19854 59838 19906
rect 59890 19854 59902 19906
rect 64978 19854 64990 19906
rect 65042 19854 65054 19906
rect 67106 19854 67118 19906
rect 67170 19854 67182 19906
rect 41582 19842 41634 19854
rect 53902 19842 53954 19854
rect 64542 19842 64594 19854
rect 68350 19842 68402 19854
rect 73166 19906 73218 19918
rect 73166 19842 73218 19854
rect 73614 19906 73666 19918
rect 81342 19906 81394 19918
rect 76738 19854 76750 19906
rect 76802 19854 76814 19906
rect 77634 19854 77646 19906
rect 77698 19854 77710 19906
rect 73614 19842 73666 19854
rect 81342 19842 81394 19854
rect 85374 19906 85426 19918
rect 85374 19842 85426 19854
rect 85710 19906 85762 19918
rect 94894 19906 94946 19918
rect 110910 19906 110962 19918
rect 93202 19854 93214 19906
rect 93266 19854 93278 19906
rect 98354 19854 98366 19906
rect 98418 19854 98430 19906
rect 85710 19842 85762 19854
rect 94894 19842 94946 19854
rect 110910 19842 110962 19854
rect 112478 19906 112530 19918
rect 112478 19842 112530 19854
rect 26910 19794 26962 19806
rect 26910 19730 26962 19742
rect 38446 19794 38498 19806
rect 38446 19730 38498 19742
rect 74174 19794 74226 19806
rect 74174 19730 74226 19742
rect 78206 19794 78258 19806
rect 78206 19730 78258 19742
rect 107886 19794 107938 19806
rect 107886 19730 107938 19742
rect 1344 19626 158592 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 96638 19626
rect 96690 19574 96742 19626
rect 96794 19574 96846 19626
rect 96898 19574 127358 19626
rect 127410 19574 127462 19626
rect 127514 19574 127566 19626
rect 127618 19574 158078 19626
rect 158130 19574 158182 19626
rect 158234 19574 158286 19626
rect 158338 19574 158592 19626
rect 1344 19540 158592 19574
rect 22766 19458 22818 19470
rect 22766 19394 22818 19406
rect 43262 19458 43314 19470
rect 43262 19394 43314 19406
rect 52110 19458 52162 19470
rect 52110 19394 52162 19406
rect 53118 19458 53170 19470
rect 85698 19406 85710 19458
rect 85762 19455 85774 19458
rect 86370 19455 86382 19458
rect 85762 19409 86382 19455
rect 85762 19406 85774 19409
rect 86370 19406 86382 19409
rect 86434 19406 86446 19458
rect 94322 19406 94334 19458
rect 94386 19455 94398 19458
rect 94882 19455 94894 19458
rect 94386 19409 94894 19455
rect 94386 19406 94398 19409
rect 94882 19406 94894 19409
rect 94946 19406 94958 19458
rect 53118 19394 53170 19406
rect 37102 19346 37154 19358
rect 49870 19346 49922 19358
rect 28466 19294 28478 19346
rect 28530 19294 28542 19346
rect 40786 19294 40798 19346
rect 40850 19294 40862 19346
rect 37102 19282 37154 19294
rect 49870 19282 49922 19294
rect 52894 19346 52946 19358
rect 52894 19282 52946 19294
rect 55246 19346 55298 19358
rect 66782 19346 66834 19358
rect 71934 19346 71986 19358
rect 74286 19346 74338 19358
rect 58594 19294 58606 19346
rect 58658 19294 58670 19346
rect 68450 19294 68462 19346
rect 68514 19294 68526 19346
rect 70578 19294 70590 19346
rect 70642 19294 70654 19346
rect 73714 19294 73726 19346
rect 73778 19294 73790 19346
rect 55246 19282 55298 19294
rect 66782 19282 66834 19294
rect 71934 19282 71986 19294
rect 74286 19282 74338 19294
rect 82014 19346 82066 19358
rect 82014 19282 82066 19294
rect 86270 19346 86322 19358
rect 86270 19282 86322 19294
rect 86718 19346 86770 19358
rect 86718 19282 86770 19294
rect 90862 19346 90914 19358
rect 90862 19282 90914 19294
rect 94334 19346 94386 19358
rect 94334 19282 94386 19294
rect 95230 19346 95282 19358
rect 95230 19282 95282 19294
rect 95790 19346 95842 19358
rect 95790 19282 95842 19294
rect 98142 19346 98194 19358
rect 98142 19282 98194 19294
rect 105422 19346 105474 19358
rect 105422 19282 105474 19294
rect 108670 19346 108722 19358
rect 108670 19282 108722 19294
rect 112366 19346 112418 19358
rect 112366 19282 112418 19294
rect 114046 19346 114098 19358
rect 114046 19282 114098 19294
rect 23886 19234 23938 19246
rect 37326 19234 37378 19246
rect 23090 19182 23102 19234
rect 23154 19182 23166 19234
rect 25442 19182 25454 19234
rect 25506 19182 25518 19234
rect 33842 19182 33854 19234
rect 33906 19182 33918 19234
rect 23886 19170 23938 19182
rect 37326 19170 37378 19182
rect 37550 19234 37602 19246
rect 37550 19170 37602 19182
rect 37998 19234 38050 19246
rect 51326 19234 51378 19246
rect 51998 19234 52050 19246
rect 56030 19234 56082 19246
rect 63870 19234 63922 19246
rect 66334 19234 66386 19246
rect 67566 19234 67618 19246
rect 86830 19234 86882 19246
rect 39106 19182 39118 19234
rect 39170 19182 39182 19234
rect 41346 19182 41358 19234
rect 41410 19182 41422 19234
rect 43586 19182 43598 19234
rect 43650 19182 43662 19234
rect 47618 19182 47630 19234
rect 47682 19182 47694 19234
rect 48402 19182 48414 19234
rect 48466 19182 48478 19234
rect 48962 19182 48974 19234
rect 49026 19182 49038 19234
rect 51090 19182 51102 19234
rect 51154 19182 51166 19234
rect 51426 19182 51438 19234
rect 51490 19182 51502 19234
rect 53330 19182 53342 19234
rect 53394 19182 53406 19234
rect 55122 19182 55134 19234
rect 55186 19182 55198 19234
rect 58706 19182 58718 19234
rect 58770 19182 58782 19234
rect 60722 19182 60734 19234
rect 60786 19182 60798 19234
rect 61170 19182 61182 19234
rect 61234 19182 61246 19234
rect 64194 19182 64206 19234
rect 64258 19182 64270 19234
rect 66994 19182 67006 19234
rect 67058 19182 67070 19234
rect 71362 19182 71374 19234
rect 71426 19182 71438 19234
rect 77186 19182 77198 19234
rect 77250 19182 77262 19234
rect 37998 19170 38050 19182
rect 51326 19170 51378 19182
rect 51998 19170 52050 19182
rect 56030 19170 56082 19182
rect 63870 19170 63922 19182
rect 66334 19170 66386 19182
rect 67566 19170 67618 19182
rect 86830 19170 86882 19182
rect 87278 19234 87330 19246
rect 87278 19170 87330 19182
rect 90638 19234 90690 19246
rect 90638 19170 90690 19182
rect 96014 19234 96066 19246
rect 109454 19234 109506 19246
rect 97234 19182 97246 19234
rect 97298 19182 97310 19234
rect 106082 19182 106094 19234
rect 106146 19182 106158 19234
rect 96014 19170 96066 19182
rect 109454 19170 109506 19182
rect 112702 19234 112754 19246
rect 112702 19170 112754 19182
rect 23326 19122 23378 19134
rect 23326 19058 23378 19070
rect 23774 19122 23826 19134
rect 36990 19122 37042 19134
rect 26226 19070 26238 19122
rect 26290 19070 26302 19122
rect 30258 19070 30270 19122
rect 30322 19070 30334 19122
rect 23774 19058 23826 19070
rect 36990 19058 37042 19070
rect 39790 19122 39842 19134
rect 46734 19122 46786 19134
rect 42802 19070 42814 19122
rect 42866 19070 42878 19122
rect 39790 19058 39842 19070
rect 46734 19058 46786 19070
rect 46846 19122 46898 19134
rect 50206 19122 50258 19134
rect 47506 19070 47518 19122
rect 47570 19070 47582 19122
rect 48290 19070 48302 19122
rect 48354 19070 48366 19122
rect 46846 19058 46898 19070
rect 50206 19058 50258 19070
rect 52670 19122 52722 19134
rect 52670 19058 52722 19070
rect 53566 19122 53618 19134
rect 53566 19058 53618 19070
rect 54014 19122 54066 19134
rect 54014 19058 54066 19070
rect 55358 19122 55410 19134
rect 55358 19058 55410 19070
rect 55694 19122 55746 19134
rect 55694 19058 55746 19070
rect 58270 19122 58322 19134
rect 64766 19122 64818 19134
rect 75294 19122 75346 19134
rect 62290 19070 62302 19122
rect 62354 19070 62366 19122
rect 66546 19070 66558 19122
rect 66610 19070 66622 19122
rect 72930 19070 72942 19122
rect 72994 19070 73006 19122
rect 58270 19058 58322 19070
rect 64766 19058 64818 19070
rect 75294 19058 75346 19070
rect 75518 19122 75570 19134
rect 87614 19122 87666 19134
rect 78978 19070 78990 19122
rect 79042 19070 79054 19122
rect 75518 19058 75570 19070
rect 87614 19058 87666 19070
rect 91086 19122 91138 19134
rect 91086 19058 91138 19070
rect 91310 19122 91362 19134
rect 91310 19058 91362 19070
rect 97806 19122 97858 19134
rect 97806 19058 97858 19070
rect 99934 19122 99986 19134
rect 99934 19058 99986 19070
rect 104974 19122 105026 19134
rect 107886 19122 107938 19134
rect 105858 19070 105870 19122
rect 105922 19070 105934 19122
rect 104974 19058 105026 19070
rect 107886 19058 107938 19070
rect 113150 19122 113202 19134
rect 113150 19058 113202 19070
rect 22878 19010 22930 19022
rect 22878 18946 22930 18958
rect 23550 19010 23602 19022
rect 23550 18946 23602 18958
rect 24446 19010 24498 19022
rect 24446 18946 24498 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 43374 19010 43426 19022
rect 43374 18946 43426 18958
rect 46510 19010 46562 19022
rect 46510 18946 46562 18958
rect 49534 19010 49586 19022
rect 49534 18946 49586 18958
rect 49758 19010 49810 19022
rect 49758 18946 49810 18958
rect 49982 19010 50034 19022
rect 49982 18946 50034 18958
rect 50878 19010 50930 19022
rect 50878 18946 50930 18958
rect 51662 19010 51714 19022
rect 51662 18946 51714 18958
rect 52558 19010 52610 19022
rect 52558 18946 52610 18958
rect 54686 19010 54738 19022
rect 54686 18946 54738 18958
rect 54910 19010 54962 19022
rect 54910 18946 54962 18958
rect 55918 19010 55970 19022
rect 55918 18946 55970 18958
rect 61294 19010 61346 19022
rect 67118 19010 67170 19022
rect 62402 18958 62414 19010
rect 62466 18958 62478 19010
rect 61294 18946 61346 18958
rect 67118 18946 67170 18958
rect 73278 19010 73330 19022
rect 73278 18946 73330 18958
rect 74846 19010 74898 19022
rect 74846 18946 74898 18958
rect 75070 19010 75122 19022
rect 75070 18946 75122 18958
rect 75182 19010 75234 19022
rect 75182 18946 75234 18958
rect 85038 19010 85090 19022
rect 85038 18946 85090 18958
rect 85486 19010 85538 19022
rect 85486 18946 85538 18958
rect 85822 19010 85874 19022
rect 85822 18946 85874 18958
rect 86606 19010 86658 19022
rect 86606 18946 86658 18958
rect 87838 19010 87890 19022
rect 87838 18946 87890 18958
rect 87950 19010 88002 19022
rect 87950 18946 88002 18958
rect 88062 19010 88114 19022
rect 88062 18946 88114 18958
rect 88622 19010 88674 19022
rect 88622 18946 88674 18958
rect 91982 19010 92034 19022
rect 91982 18946 92034 18958
rect 92430 19010 92482 19022
rect 92430 18946 92482 18958
rect 93550 19010 93602 19022
rect 93550 18946 93602 18958
rect 94782 19010 94834 19022
rect 96686 19010 96738 19022
rect 96338 18958 96350 19010
rect 96402 18958 96414 19010
rect 94782 18946 94834 18958
rect 96686 18946 96738 18958
rect 96798 19010 96850 19022
rect 96798 18946 96850 18958
rect 96910 19010 96962 19022
rect 96910 18946 96962 18958
rect 98030 19010 98082 19022
rect 98030 18946 98082 18958
rect 98254 19010 98306 19022
rect 98254 18946 98306 18958
rect 98814 19010 98866 19022
rect 98814 18946 98866 18958
rect 99262 19010 99314 19022
rect 99262 18946 99314 18958
rect 100270 19010 100322 19022
rect 100270 18946 100322 18958
rect 112814 19010 112866 19022
rect 112814 18946 112866 18958
rect 112926 19010 112978 19022
rect 112926 18946 112978 18958
rect 114158 19010 114210 19022
rect 114158 18946 114210 18958
rect 1344 18842 158592 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 81278 18842
rect 81330 18790 81382 18842
rect 81434 18790 81486 18842
rect 81538 18790 111998 18842
rect 112050 18790 112102 18842
rect 112154 18790 112206 18842
rect 112258 18790 142718 18842
rect 142770 18790 142822 18842
rect 142874 18790 142926 18842
rect 142978 18790 158592 18842
rect 1344 18756 158592 18790
rect 26350 18674 26402 18686
rect 26350 18610 26402 18622
rect 26686 18674 26738 18686
rect 26686 18610 26738 18622
rect 32174 18674 32226 18686
rect 32174 18610 32226 18622
rect 34302 18674 34354 18686
rect 34302 18610 34354 18622
rect 34862 18674 34914 18686
rect 53454 18674 53506 18686
rect 49522 18622 49534 18674
rect 49586 18622 49598 18674
rect 34862 18610 34914 18622
rect 53454 18610 53506 18622
rect 56702 18674 56754 18686
rect 86158 18674 86210 18686
rect 60050 18622 60062 18674
rect 60114 18622 60126 18674
rect 66770 18622 66782 18674
rect 66834 18622 66846 18674
rect 70130 18622 70142 18674
rect 70194 18622 70206 18674
rect 56702 18610 56754 18622
rect 86158 18610 86210 18622
rect 91534 18674 91586 18686
rect 91534 18610 91586 18622
rect 91646 18674 91698 18686
rect 91646 18610 91698 18622
rect 91758 18674 91810 18686
rect 91758 18610 91810 18622
rect 25342 18562 25394 18574
rect 25342 18498 25394 18510
rect 26462 18562 26514 18574
rect 26462 18498 26514 18510
rect 52446 18562 52498 18574
rect 52446 18498 52498 18510
rect 58606 18562 58658 18574
rect 58606 18498 58658 18510
rect 58718 18562 58770 18574
rect 62526 18562 62578 18574
rect 61954 18510 61966 18562
rect 62018 18510 62030 18562
rect 58718 18498 58770 18510
rect 62526 18498 62578 18510
rect 62638 18562 62690 18574
rect 62638 18498 62690 18510
rect 65102 18562 65154 18574
rect 65102 18498 65154 18510
rect 67678 18562 67730 18574
rect 67678 18498 67730 18510
rect 74622 18562 74674 18574
rect 74622 18498 74674 18510
rect 93550 18562 93602 18574
rect 93550 18498 93602 18510
rect 95790 18562 95842 18574
rect 95790 18498 95842 18510
rect 96350 18562 96402 18574
rect 114942 18562 114994 18574
rect 100370 18510 100382 18562
rect 100434 18510 100446 18562
rect 106418 18510 106430 18562
rect 106482 18510 106494 18562
rect 96350 18498 96402 18510
rect 114942 18498 114994 18510
rect 28814 18450 28866 18462
rect 21522 18398 21534 18450
rect 21586 18398 21598 18450
rect 26898 18398 26910 18450
rect 26962 18398 26974 18450
rect 28814 18386 28866 18398
rect 29822 18450 29874 18462
rect 29822 18386 29874 18398
rect 30046 18450 30098 18462
rect 30046 18386 30098 18398
rect 30270 18450 30322 18462
rect 30270 18386 30322 18398
rect 30494 18450 30546 18462
rect 30494 18386 30546 18398
rect 31838 18450 31890 18462
rect 31838 18386 31890 18398
rect 32510 18450 32562 18462
rect 32510 18386 32562 18398
rect 34638 18450 34690 18462
rect 34638 18386 34690 18398
rect 34750 18450 34802 18462
rect 34750 18386 34802 18398
rect 35310 18450 35362 18462
rect 42590 18450 42642 18462
rect 46286 18450 46338 18462
rect 37314 18398 37326 18450
rect 37378 18398 37390 18450
rect 42130 18398 42142 18450
rect 42194 18398 42206 18450
rect 43586 18398 43598 18450
rect 43650 18398 43662 18450
rect 45378 18398 45390 18450
rect 45442 18398 45454 18450
rect 35310 18386 35362 18398
rect 42590 18386 42642 18398
rect 46286 18386 46338 18398
rect 47518 18450 47570 18462
rect 47518 18386 47570 18398
rect 47630 18450 47682 18462
rect 47630 18386 47682 18398
rect 47742 18450 47794 18462
rect 48862 18450 48914 18462
rect 49982 18450 50034 18462
rect 52110 18450 52162 18462
rect 53118 18450 53170 18462
rect 48178 18398 48190 18450
rect 48242 18398 48254 18450
rect 49298 18398 49310 18450
rect 49362 18398 49374 18450
rect 50306 18398 50318 18450
rect 50370 18398 50382 18450
rect 51202 18398 51214 18450
rect 51266 18398 51278 18450
rect 51874 18398 51886 18450
rect 51938 18398 51950 18450
rect 52658 18398 52670 18450
rect 52722 18398 52734 18450
rect 47742 18386 47794 18398
rect 48862 18386 48914 18398
rect 49982 18386 50034 18398
rect 52110 18386 52162 18398
rect 53118 18386 53170 18398
rect 53342 18450 53394 18462
rect 58382 18450 58434 18462
rect 56914 18398 56926 18450
rect 56978 18398 56990 18450
rect 53342 18386 53394 18398
rect 58382 18386 58434 18398
rect 59502 18450 59554 18462
rect 62862 18450 62914 18462
rect 60722 18398 60734 18450
rect 60786 18398 60798 18450
rect 61618 18398 61630 18450
rect 61682 18398 61694 18450
rect 59502 18386 59554 18398
rect 62862 18386 62914 18398
rect 63422 18450 63474 18462
rect 66558 18450 66610 18462
rect 64418 18398 64430 18450
rect 64482 18398 64494 18450
rect 63422 18386 63474 18398
rect 66558 18386 66610 18398
rect 69022 18450 69074 18462
rect 69022 18386 69074 18398
rect 69470 18450 69522 18462
rect 69470 18386 69522 18398
rect 69582 18450 69634 18462
rect 69582 18386 69634 18398
rect 69694 18450 69746 18462
rect 69694 18386 69746 18398
rect 70702 18450 70754 18462
rect 74062 18450 74114 18462
rect 73266 18398 73278 18450
rect 73330 18398 73342 18450
rect 70702 18386 70754 18398
rect 74062 18386 74114 18398
rect 74174 18450 74226 18462
rect 74174 18386 74226 18398
rect 74286 18450 74338 18462
rect 85822 18450 85874 18462
rect 76066 18398 76078 18450
rect 76130 18398 76142 18450
rect 77746 18398 77758 18450
rect 77810 18398 77822 18450
rect 79538 18398 79550 18450
rect 79602 18398 79614 18450
rect 80434 18398 80446 18450
rect 80498 18398 80510 18450
rect 81106 18398 81118 18450
rect 81170 18398 81182 18450
rect 83458 18398 83470 18450
rect 83522 18398 83534 18450
rect 74286 18386 74338 18398
rect 85822 18386 85874 18398
rect 86382 18450 86434 18462
rect 86382 18386 86434 18398
rect 86830 18450 86882 18462
rect 92206 18450 92258 18462
rect 90290 18398 90302 18450
rect 90354 18398 90366 18450
rect 91074 18398 91086 18450
rect 91138 18398 91150 18450
rect 86830 18386 86882 18398
rect 92206 18386 92258 18398
rect 92542 18450 92594 18462
rect 92542 18386 92594 18398
rect 93102 18450 93154 18462
rect 93102 18386 93154 18398
rect 95342 18450 95394 18462
rect 95342 18386 95394 18398
rect 96126 18450 96178 18462
rect 99710 18450 99762 18462
rect 96674 18398 96686 18450
rect 96738 18398 96750 18450
rect 96126 18386 96178 18398
rect 99710 18386 99762 18398
rect 100046 18450 100098 18462
rect 100046 18386 100098 18398
rect 101390 18450 101442 18462
rect 101390 18386 101442 18398
rect 101726 18450 101778 18462
rect 101726 18386 101778 18398
rect 101950 18450 102002 18462
rect 101950 18386 102002 18398
rect 102510 18450 102562 18462
rect 102510 18386 102562 18398
rect 106094 18450 106146 18462
rect 106094 18386 106146 18398
rect 106990 18450 107042 18462
rect 106990 18386 107042 18398
rect 108670 18450 108722 18462
rect 108670 18386 108722 18398
rect 108894 18450 108946 18462
rect 108894 18386 108946 18398
rect 109342 18450 109394 18462
rect 109342 18386 109394 18398
rect 109566 18450 109618 18462
rect 109566 18386 109618 18398
rect 111694 18450 111746 18462
rect 111694 18386 111746 18398
rect 112142 18450 112194 18462
rect 112142 18386 112194 18398
rect 112366 18450 112418 18462
rect 112366 18386 112418 18398
rect 27358 18338 27410 18350
rect 22194 18286 22206 18338
rect 22258 18286 22270 18338
rect 24322 18286 24334 18338
rect 24386 18286 24398 18338
rect 27358 18274 27410 18286
rect 33742 18338 33794 18350
rect 33742 18274 33794 18286
rect 35646 18338 35698 18350
rect 35646 18274 35698 18286
rect 36206 18338 36258 18350
rect 36206 18274 36258 18286
rect 36990 18338 37042 18350
rect 42702 18338 42754 18350
rect 38098 18286 38110 18338
rect 38162 18286 38174 18338
rect 40226 18286 40238 18338
rect 40290 18286 40302 18338
rect 36990 18274 37042 18286
rect 42702 18274 42754 18286
rect 43150 18338 43202 18350
rect 57374 18338 57426 18350
rect 45714 18286 45726 18338
rect 45778 18286 45790 18338
rect 51762 18286 51774 18338
rect 51826 18286 51838 18338
rect 43150 18274 43202 18286
rect 57374 18274 57426 18286
rect 57822 18338 57874 18350
rect 63086 18338 63138 18350
rect 71598 18338 71650 18350
rect 61058 18286 61070 18338
rect 61122 18286 61134 18338
rect 63746 18286 63758 18338
rect 63810 18286 63822 18338
rect 57822 18274 57874 18286
rect 63086 18274 63138 18286
rect 71598 18274 71650 18286
rect 75630 18338 75682 18350
rect 75630 18274 75682 18286
rect 76638 18338 76690 18350
rect 76638 18274 76690 18286
rect 84030 18338 84082 18350
rect 84030 18274 84082 18286
rect 84478 18338 84530 18350
rect 84478 18274 84530 18286
rect 85038 18338 85090 18350
rect 85038 18274 85090 18286
rect 85486 18338 85538 18350
rect 85486 18274 85538 18286
rect 86270 18338 86322 18350
rect 86270 18274 86322 18286
rect 87166 18338 87218 18350
rect 94446 18338 94498 18350
rect 87938 18286 87950 18338
rect 88002 18286 88014 18338
rect 87166 18274 87218 18286
rect 94446 18274 94498 18286
rect 94782 18338 94834 18350
rect 94782 18274 94834 18286
rect 95902 18338 95954 18350
rect 100830 18338 100882 18350
rect 98914 18286 98926 18338
rect 98978 18286 98990 18338
rect 95902 18274 95954 18286
rect 100830 18274 100882 18286
rect 101838 18338 101890 18350
rect 101838 18274 101890 18286
rect 105758 18338 105810 18350
rect 105758 18274 105810 18286
rect 109118 18338 109170 18350
rect 109118 18274 109170 18286
rect 111022 18338 111074 18350
rect 111022 18274 111074 18286
rect 111918 18338 111970 18350
rect 111918 18274 111970 18286
rect 33182 18226 33234 18238
rect 33182 18162 33234 18174
rect 33518 18226 33570 18238
rect 52894 18226 52946 18238
rect 35410 18174 35422 18226
rect 35474 18223 35486 18226
rect 35634 18223 35646 18226
rect 35474 18177 35646 18223
rect 35474 18174 35486 18177
rect 35634 18174 35646 18177
rect 35698 18174 35710 18226
rect 33518 18162 33570 18174
rect 52894 18162 52946 18174
rect 56590 18226 56642 18238
rect 56590 18162 56642 18174
rect 57262 18226 57314 18238
rect 57262 18162 57314 18174
rect 59726 18226 59778 18238
rect 59726 18162 59778 18174
rect 62078 18226 62130 18238
rect 62078 18162 62130 18174
rect 72942 18226 72994 18238
rect 72942 18162 72994 18174
rect 115054 18226 115106 18238
rect 115054 18162 115106 18174
rect 1344 18058 158592 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 96638 18058
rect 96690 18006 96742 18058
rect 96794 18006 96846 18058
rect 96898 18006 127358 18058
rect 127410 18006 127462 18058
rect 127514 18006 127566 18058
rect 127618 18006 158078 18058
rect 158130 18006 158182 18058
rect 158234 18006 158286 18058
rect 158338 18006 158592 18058
rect 1344 17972 158592 18006
rect 22654 17890 22706 17902
rect 22654 17826 22706 17838
rect 23214 17890 23266 17902
rect 23214 17826 23266 17838
rect 41918 17890 41970 17902
rect 41918 17826 41970 17838
rect 42142 17890 42194 17902
rect 42142 17826 42194 17838
rect 42254 17890 42306 17902
rect 42254 17826 42306 17838
rect 50990 17890 51042 17902
rect 50990 17826 51042 17838
rect 64430 17890 64482 17902
rect 64430 17826 64482 17838
rect 24558 17778 24610 17790
rect 35422 17778 35474 17790
rect 64318 17778 64370 17790
rect 84254 17778 84306 17790
rect 88174 17778 88226 17790
rect 32050 17726 32062 17778
rect 32114 17726 32126 17778
rect 34178 17726 34190 17778
rect 34242 17726 34254 17778
rect 45378 17726 45390 17778
rect 45442 17726 45454 17778
rect 56130 17726 56142 17778
rect 56194 17726 56206 17778
rect 58370 17726 58382 17778
rect 58434 17726 58446 17778
rect 60610 17726 60622 17778
rect 60674 17726 60686 17778
rect 71362 17726 71374 17778
rect 71426 17726 71438 17778
rect 72258 17726 72270 17778
rect 72322 17726 72334 17778
rect 73042 17726 73054 17778
rect 73106 17726 73118 17778
rect 77186 17726 77198 17778
rect 77250 17726 77262 17778
rect 86930 17726 86942 17778
rect 86994 17726 87006 17778
rect 24558 17714 24610 17726
rect 35422 17714 35474 17726
rect 64318 17714 64370 17726
rect 84254 17714 84306 17726
rect 88174 17714 88226 17726
rect 89630 17778 89682 17790
rect 89630 17714 89682 17726
rect 93214 17778 93266 17790
rect 97694 17778 97746 17790
rect 97234 17726 97246 17778
rect 97298 17726 97310 17778
rect 93214 17714 93266 17726
rect 97694 17714 97746 17726
rect 98142 17778 98194 17790
rect 98142 17714 98194 17726
rect 22766 17666 22818 17678
rect 22766 17602 22818 17614
rect 22990 17666 23042 17678
rect 23774 17666 23826 17678
rect 23314 17614 23326 17666
rect 23378 17614 23390 17666
rect 22990 17602 23042 17614
rect 23774 17602 23826 17614
rect 24110 17666 24162 17678
rect 24110 17602 24162 17614
rect 31054 17666 31106 17678
rect 34526 17666 34578 17678
rect 45838 17666 45890 17678
rect 47294 17666 47346 17678
rect 31378 17614 31390 17666
rect 31442 17614 31454 17666
rect 41682 17614 41694 17666
rect 41746 17614 41758 17666
rect 46498 17614 46510 17666
rect 46562 17614 46574 17666
rect 31054 17602 31106 17614
rect 34526 17602 34578 17614
rect 45838 17602 45890 17614
rect 47294 17602 47346 17614
rect 47966 17666 48018 17678
rect 47966 17602 48018 17614
rect 48862 17666 48914 17678
rect 48862 17602 48914 17614
rect 49534 17666 49586 17678
rect 70030 17666 70082 17678
rect 70926 17666 70978 17678
rect 55458 17614 55470 17666
rect 55522 17614 55534 17666
rect 62178 17614 62190 17666
rect 62242 17614 62254 17666
rect 63410 17614 63422 17666
rect 63474 17614 63486 17666
rect 63858 17614 63870 17666
rect 63922 17614 63934 17666
rect 65650 17614 65662 17666
rect 65714 17614 65726 17666
rect 68898 17614 68910 17666
rect 68962 17614 68974 17666
rect 69570 17614 69582 17666
rect 69634 17614 69646 17666
rect 70466 17614 70478 17666
rect 70530 17614 70542 17666
rect 49534 17602 49586 17614
rect 70030 17602 70082 17614
rect 70926 17602 70978 17614
rect 71822 17666 71874 17678
rect 85374 17666 85426 17678
rect 76850 17614 76862 17666
rect 76914 17614 76926 17666
rect 79986 17614 79998 17666
rect 80050 17614 80062 17666
rect 80770 17614 80782 17666
rect 80834 17614 80846 17666
rect 71822 17602 71874 17614
rect 85374 17602 85426 17614
rect 85598 17666 85650 17678
rect 85598 17602 85650 17614
rect 86046 17666 86098 17678
rect 87838 17666 87890 17678
rect 87266 17614 87278 17666
rect 87330 17614 87342 17666
rect 86046 17602 86098 17614
rect 87838 17602 87890 17614
rect 87950 17666 88002 17678
rect 87950 17602 88002 17614
rect 88286 17666 88338 17678
rect 106206 17666 106258 17678
rect 94322 17614 94334 17666
rect 94386 17614 94398 17666
rect 94882 17614 94894 17666
rect 94946 17614 94958 17666
rect 99810 17614 99822 17666
rect 99874 17614 99886 17666
rect 88286 17602 88338 17614
rect 106206 17602 106258 17614
rect 106542 17666 106594 17678
rect 106542 17602 106594 17614
rect 107550 17666 107602 17678
rect 109106 17614 109118 17666
rect 109170 17614 109182 17666
rect 109778 17614 109790 17666
rect 109842 17614 109854 17666
rect 107550 17602 107602 17614
rect 23550 17554 23602 17566
rect 23550 17490 23602 17502
rect 23998 17554 24050 17566
rect 30718 17554 30770 17566
rect 29586 17502 29598 17554
rect 29650 17502 29662 17554
rect 23998 17490 24050 17502
rect 30718 17490 30770 17502
rect 39454 17554 39506 17566
rect 39454 17490 39506 17502
rect 39566 17554 39618 17566
rect 39566 17490 39618 17502
rect 41022 17554 41074 17566
rect 41022 17490 41074 17502
rect 41134 17554 41186 17566
rect 41134 17490 41186 17502
rect 46286 17554 46338 17566
rect 46286 17490 46338 17502
rect 48078 17554 48130 17566
rect 50990 17554 51042 17566
rect 49186 17502 49198 17554
rect 49250 17502 49262 17554
rect 49858 17502 49870 17554
rect 49922 17502 49934 17554
rect 50530 17502 50542 17554
rect 50594 17502 50606 17554
rect 48078 17490 48130 17502
rect 50990 17490 51042 17502
rect 51102 17554 51154 17566
rect 51102 17490 51154 17502
rect 58830 17554 58882 17566
rect 58830 17490 58882 17502
rect 58942 17554 58994 17566
rect 58942 17490 58994 17502
rect 59502 17554 59554 17566
rect 67006 17554 67058 17566
rect 69358 17554 69410 17566
rect 61954 17502 61966 17554
rect 62018 17502 62030 17554
rect 65426 17502 65438 17554
rect 65490 17502 65502 17554
rect 68674 17502 68686 17554
rect 68738 17502 68750 17554
rect 59502 17490 59554 17502
rect 67006 17490 67058 17502
rect 69358 17490 69410 17502
rect 72718 17554 72770 17566
rect 72718 17490 72770 17502
rect 88734 17554 88786 17566
rect 88734 17490 88786 17502
rect 92206 17554 92258 17566
rect 106766 17554 106818 17566
rect 101714 17502 101726 17554
rect 101778 17502 101790 17554
rect 92206 17490 92258 17502
rect 106766 17490 106818 17502
rect 107662 17554 107714 17566
rect 107662 17490 107714 17502
rect 107998 17554 108050 17566
rect 107998 17490 108050 17502
rect 22318 17442 22370 17454
rect 22318 17378 22370 17390
rect 22654 17442 22706 17454
rect 22654 17378 22706 17390
rect 29934 17442 29986 17454
rect 29934 17378 29986 17390
rect 30830 17442 30882 17454
rect 39230 17442 39282 17454
rect 34850 17390 34862 17442
rect 34914 17390 34926 17442
rect 30830 17378 30882 17390
rect 39230 17378 39282 17390
rect 41358 17442 41410 17454
rect 48302 17442 48354 17454
rect 46946 17390 46958 17442
rect 47010 17390 47022 17442
rect 41358 17378 41410 17390
rect 48302 17378 48354 17390
rect 50206 17442 50258 17454
rect 50206 17378 50258 17390
rect 52782 17442 52834 17454
rect 52782 17378 52834 17390
rect 59166 17442 59218 17454
rect 59166 17378 59218 17390
rect 59950 17442 60002 17454
rect 59950 17378 60002 17390
rect 61070 17442 61122 17454
rect 61070 17378 61122 17390
rect 67790 17442 67842 17454
rect 67790 17378 67842 17390
rect 73726 17442 73778 17454
rect 73726 17378 73778 17390
rect 74174 17442 74226 17454
rect 74174 17378 74226 17390
rect 79326 17442 79378 17454
rect 79326 17378 79378 17390
rect 79774 17442 79826 17454
rect 84366 17442 84418 17454
rect 83122 17390 83134 17442
rect 83186 17390 83198 17442
rect 79774 17378 79826 17390
rect 84366 17378 84418 17390
rect 85150 17442 85202 17454
rect 85150 17378 85202 17390
rect 85822 17442 85874 17454
rect 85822 17378 85874 17390
rect 86382 17442 86434 17454
rect 86382 17378 86434 17390
rect 89294 17442 89346 17454
rect 89294 17378 89346 17390
rect 90078 17442 90130 17454
rect 90078 17378 90130 17390
rect 90862 17442 90914 17454
rect 90862 17378 90914 17390
rect 91198 17442 91250 17454
rect 91198 17378 91250 17390
rect 92766 17442 92818 17454
rect 92766 17378 92818 17390
rect 93662 17442 93714 17454
rect 93662 17378 93714 17390
rect 97806 17442 97858 17454
rect 97806 17378 97858 17390
rect 98254 17442 98306 17454
rect 98254 17378 98306 17390
rect 98702 17442 98754 17454
rect 98702 17378 98754 17390
rect 99262 17442 99314 17454
rect 99262 17378 99314 17390
rect 106318 17442 106370 17454
rect 106318 17378 106370 17390
rect 107774 17442 107826 17454
rect 107774 17378 107826 17390
rect 108894 17442 108946 17454
rect 112242 17390 112254 17442
rect 112306 17390 112318 17442
rect 108894 17378 108946 17390
rect 1344 17274 158592 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 81278 17274
rect 81330 17222 81382 17274
rect 81434 17222 81486 17274
rect 81538 17222 111998 17274
rect 112050 17222 112102 17274
rect 112154 17222 112206 17274
rect 112258 17222 142718 17274
rect 142770 17222 142822 17274
rect 142874 17222 142926 17274
rect 142978 17222 158592 17274
rect 1344 17188 158592 17222
rect 19630 17106 19682 17118
rect 19630 17042 19682 17054
rect 23550 17106 23602 17118
rect 23550 17042 23602 17054
rect 25342 17106 25394 17118
rect 25342 17042 25394 17054
rect 28254 17106 28306 17118
rect 28254 17042 28306 17054
rect 30046 17106 30098 17118
rect 30046 17042 30098 17054
rect 36094 17106 36146 17118
rect 36094 17042 36146 17054
rect 38110 17106 38162 17118
rect 38110 17042 38162 17054
rect 44270 17106 44322 17118
rect 44270 17042 44322 17054
rect 49870 17106 49922 17118
rect 49870 17042 49922 17054
rect 51102 17106 51154 17118
rect 51102 17042 51154 17054
rect 51214 17106 51266 17118
rect 51214 17042 51266 17054
rect 51326 17106 51378 17118
rect 51326 17042 51378 17054
rect 51886 17106 51938 17118
rect 51886 17042 51938 17054
rect 52334 17106 52386 17118
rect 52334 17042 52386 17054
rect 56702 17106 56754 17118
rect 56702 17042 56754 17054
rect 58718 17106 58770 17118
rect 58718 17042 58770 17054
rect 60398 17106 60450 17118
rect 64542 17106 64594 17118
rect 63074 17054 63086 17106
rect 63138 17054 63150 17106
rect 60398 17042 60450 17054
rect 64542 17042 64594 17054
rect 75742 17106 75794 17118
rect 75742 17042 75794 17054
rect 79214 17106 79266 17118
rect 79214 17042 79266 17054
rect 80110 17106 80162 17118
rect 80110 17042 80162 17054
rect 80894 17106 80946 17118
rect 80894 17042 80946 17054
rect 81230 17106 81282 17118
rect 81230 17042 81282 17054
rect 82126 17106 82178 17118
rect 82126 17042 82178 17054
rect 83246 17106 83298 17118
rect 87390 17106 87442 17118
rect 83906 17054 83918 17106
rect 83970 17054 83982 17106
rect 83246 17042 83298 17054
rect 87390 17042 87442 17054
rect 89070 17106 89122 17118
rect 89070 17042 89122 17054
rect 89630 17106 89682 17118
rect 89630 17042 89682 17054
rect 90862 17106 90914 17118
rect 90862 17042 90914 17054
rect 92318 17106 92370 17118
rect 92318 17042 92370 17054
rect 92542 17106 92594 17118
rect 92542 17042 92594 17054
rect 93662 17106 93714 17118
rect 93662 17042 93714 17054
rect 93886 17106 93938 17118
rect 93886 17042 93938 17054
rect 95006 17106 95058 17118
rect 95006 17042 95058 17054
rect 96238 17106 96290 17118
rect 96238 17042 96290 17054
rect 97358 17106 97410 17118
rect 97358 17042 97410 17054
rect 99598 17106 99650 17118
rect 99598 17042 99650 17054
rect 99822 17106 99874 17118
rect 99822 17042 99874 17054
rect 100942 17106 100994 17118
rect 100942 17042 100994 17054
rect 102510 17106 102562 17118
rect 102510 17042 102562 17054
rect 105422 17106 105474 17118
rect 105422 17042 105474 17054
rect 109790 17106 109842 17118
rect 109790 17042 109842 17054
rect 109902 17106 109954 17118
rect 115266 17054 115278 17106
rect 115330 17054 115342 17106
rect 109902 17042 109954 17054
rect 28030 16994 28082 17006
rect 21634 16942 21646 16994
rect 21698 16942 21710 16994
rect 28030 16930 28082 16942
rect 30270 16994 30322 17006
rect 30270 16930 30322 16942
rect 31054 16994 31106 17006
rect 31054 16930 31106 16942
rect 31502 16994 31554 17006
rect 38222 16994 38274 17006
rect 32162 16942 32174 16994
rect 32226 16942 32238 16994
rect 33842 16942 33854 16994
rect 33906 16942 33918 16994
rect 31502 16930 31554 16942
rect 38222 16930 38274 16942
rect 38894 16994 38946 17006
rect 38894 16930 38946 16942
rect 39006 16994 39058 17006
rect 39006 16930 39058 16942
rect 45950 16994 46002 17006
rect 45950 16930 46002 16942
rect 47406 16994 47458 17006
rect 47406 16930 47458 16942
rect 47630 16994 47682 17006
rect 57598 16994 57650 17006
rect 48738 16942 48750 16994
rect 48802 16942 48814 16994
rect 53554 16942 53566 16994
rect 53618 16942 53630 16994
rect 47630 16930 47682 16942
rect 57598 16930 57650 16942
rect 63758 16994 63810 17006
rect 81118 16994 81170 17006
rect 68898 16942 68910 16994
rect 68962 16942 68974 16994
rect 79538 16942 79550 16994
rect 79602 16942 79614 16994
rect 80434 16942 80446 16994
rect 80498 16942 80510 16994
rect 63758 16930 63810 16942
rect 81118 16930 81170 16942
rect 81678 16994 81730 17006
rect 81678 16930 81730 16942
rect 81902 16994 81954 17006
rect 81902 16930 81954 16942
rect 82238 16994 82290 17006
rect 82238 16930 82290 16942
rect 82686 16994 82738 17006
rect 82686 16930 82738 16942
rect 94446 16994 94498 17006
rect 94446 16930 94498 16942
rect 98254 16994 98306 17006
rect 101726 16994 101778 17006
rect 100146 16942 100158 16994
rect 100210 16942 100222 16994
rect 98254 16930 98306 16942
rect 101726 16930 101778 16942
rect 104974 16994 105026 17006
rect 104974 16930 105026 16942
rect 105310 16994 105362 17006
rect 105310 16930 105362 16942
rect 115614 16994 115666 17006
rect 115614 16930 115666 16942
rect 19294 16882 19346 16894
rect 26462 16882 26514 16894
rect 20178 16830 20190 16882
rect 20242 16830 20254 16882
rect 19294 16818 19346 16830
rect 26462 16818 26514 16830
rect 26686 16882 26738 16894
rect 26686 16818 26738 16830
rect 27134 16882 27186 16894
rect 27134 16818 27186 16830
rect 27918 16882 27970 16894
rect 27918 16818 27970 16830
rect 30382 16882 30434 16894
rect 30382 16818 30434 16830
rect 30718 16882 30770 16894
rect 30718 16818 30770 16830
rect 31838 16882 31890 16894
rect 37774 16882 37826 16894
rect 32386 16830 32398 16882
rect 32450 16830 32462 16882
rect 35634 16830 35646 16882
rect 35698 16830 35710 16882
rect 31838 16818 31890 16830
rect 37774 16818 37826 16830
rect 38334 16882 38386 16894
rect 38334 16818 38386 16830
rect 38670 16882 38722 16894
rect 47854 16882 47906 16894
rect 40898 16830 40910 16882
rect 40962 16830 40974 16882
rect 38670 16818 38722 16830
rect 47854 16818 47906 16830
rect 48078 16882 48130 16894
rect 48078 16818 48130 16830
rect 49086 16882 49138 16894
rect 49086 16818 49138 16830
rect 50878 16882 50930 16894
rect 57038 16882 57090 16894
rect 52882 16830 52894 16882
rect 52946 16830 52958 16882
rect 50878 16818 50930 16830
rect 57038 16818 57090 16830
rect 60734 16882 60786 16894
rect 66222 16882 66274 16894
rect 76190 16882 76242 16894
rect 60946 16830 60958 16882
rect 61010 16830 61022 16882
rect 62178 16830 62190 16882
rect 62242 16830 62254 16882
rect 62402 16830 62414 16882
rect 62466 16830 62478 16882
rect 63410 16830 63422 16882
rect 63474 16830 63486 16882
rect 66434 16830 66446 16882
rect 66498 16830 66510 16882
rect 72482 16830 72494 16882
rect 72546 16830 72558 16882
rect 60734 16818 60786 16830
rect 66222 16818 66274 16830
rect 76190 16818 76242 16830
rect 76414 16882 76466 16894
rect 76414 16818 76466 16830
rect 76862 16882 76914 16894
rect 76862 16818 76914 16830
rect 81342 16882 81394 16894
rect 81342 16818 81394 16830
rect 83582 16882 83634 16894
rect 89294 16882 89346 16894
rect 86258 16830 86270 16882
rect 86322 16830 86334 16882
rect 87042 16830 87054 16882
rect 87106 16830 87118 16882
rect 83582 16818 83634 16830
rect 89294 16818 89346 16830
rect 89742 16882 89794 16894
rect 89742 16818 89794 16830
rect 89966 16882 90018 16894
rect 89966 16818 90018 16830
rect 93102 16882 93154 16894
rect 93102 16818 93154 16830
rect 96350 16882 96402 16894
rect 96350 16818 96402 16830
rect 96686 16882 96738 16894
rect 96686 16818 96738 16830
rect 97022 16882 97074 16894
rect 97022 16818 97074 16830
rect 97582 16882 97634 16894
rect 100382 16882 100434 16894
rect 97906 16830 97918 16882
rect 97970 16830 97982 16882
rect 97582 16818 97634 16830
rect 100382 16818 100434 16830
rect 100830 16882 100882 16894
rect 100830 16818 100882 16830
rect 101054 16882 101106 16894
rect 101054 16818 101106 16830
rect 101390 16882 101442 16894
rect 101390 16818 101442 16830
rect 101950 16882 102002 16894
rect 109230 16882 109282 16894
rect 105634 16830 105646 16882
rect 105698 16830 105710 16882
rect 106306 16830 106318 16882
rect 106370 16830 106382 16882
rect 108770 16830 108782 16882
rect 108834 16830 108846 16882
rect 101950 16818 102002 16830
rect 109230 16818 109282 16830
rect 109678 16882 109730 16894
rect 109678 16818 109730 16830
rect 111918 16882 111970 16894
rect 112130 16830 112142 16882
rect 112194 16830 112206 16882
rect 112802 16830 112814 16882
rect 112866 16830 112878 16882
rect 111918 16818 111970 16830
rect 26574 16770 26626 16782
rect 61518 16770 61570 16782
rect 76302 16770 76354 16782
rect 20290 16718 20302 16770
rect 20354 16718 20366 16770
rect 41682 16718 41694 16770
rect 41746 16718 41758 16770
rect 43810 16718 43822 16770
rect 43874 16718 43886 16770
rect 55682 16718 55694 16770
rect 55746 16718 55758 16770
rect 62066 16718 62078 16770
rect 62130 16718 62142 16770
rect 73154 16718 73166 16770
rect 73218 16718 73230 16770
rect 75282 16718 75294 16770
rect 75346 16718 75358 16770
rect 26574 16706 26626 16718
rect 61518 16706 61570 16718
rect 76302 16706 76354 16718
rect 77198 16770 77250 16782
rect 77198 16706 77250 16718
rect 77646 16770 77698 16782
rect 77646 16706 77698 16718
rect 78206 16770 78258 16782
rect 78206 16706 78258 16718
rect 78990 16770 79042 16782
rect 78990 16706 79042 16718
rect 88398 16770 88450 16782
rect 88398 16706 88450 16718
rect 90414 16770 90466 16782
rect 90414 16706 90466 16718
rect 91646 16770 91698 16782
rect 91646 16706 91698 16718
rect 96574 16770 96626 16782
rect 96574 16706 96626 16718
rect 97470 16770 97522 16782
rect 97470 16706 97522 16718
rect 98814 16770 98866 16782
rect 98814 16706 98866 16718
rect 101502 16770 101554 16782
rect 101502 16706 101554 16718
rect 102958 16770 103010 16782
rect 102958 16706 103010 16718
rect 103854 16770 103906 16782
rect 103854 16706 103906 16718
rect 104190 16770 104242 16782
rect 104190 16706 104242 16718
rect 50654 16658 50706 16670
rect 50654 16594 50706 16606
rect 82574 16658 82626 16670
rect 82574 16594 82626 16606
rect 98366 16658 98418 16670
rect 98366 16594 98418 16606
rect 115726 16658 115778 16670
rect 115726 16594 115778 16606
rect 1344 16490 158592 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 96638 16490
rect 96690 16438 96742 16490
rect 96794 16438 96846 16490
rect 96898 16438 127358 16490
rect 127410 16438 127462 16490
rect 127514 16438 127566 16490
rect 127618 16438 158078 16490
rect 158130 16438 158182 16490
rect 158234 16438 158286 16490
rect 158338 16438 158592 16490
rect 1344 16404 158592 16438
rect 31166 16322 31218 16334
rect 31166 16258 31218 16270
rect 31950 16322 32002 16334
rect 31950 16258 32002 16270
rect 32622 16322 32674 16334
rect 32622 16258 32674 16270
rect 33406 16322 33458 16334
rect 33406 16258 33458 16270
rect 33742 16322 33794 16334
rect 62078 16322 62130 16334
rect 48402 16270 48414 16322
rect 48466 16270 48478 16322
rect 78530 16270 78542 16322
rect 78594 16319 78606 16322
rect 79314 16319 79326 16322
rect 78594 16273 79326 16319
rect 78594 16270 78606 16273
rect 79314 16270 79326 16273
rect 79378 16270 79390 16322
rect 84130 16270 84142 16322
rect 84194 16319 84206 16322
rect 84914 16319 84926 16322
rect 84194 16273 84926 16319
rect 84194 16270 84206 16273
rect 84914 16270 84926 16273
rect 84978 16270 84990 16322
rect 87378 16270 87390 16322
rect 87442 16270 87454 16322
rect 95330 16319 95342 16322
rect 94785 16273 95342 16319
rect 33742 16258 33794 16270
rect 62078 16258 62130 16270
rect 34974 16210 35026 16222
rect 20738 16158 20750 16210
rect 20802 16158 20814 16210
rect 24546 16158 24558 16210
rect 24610 16158 24622 16210
rect 28466 16158 28478 16210
rect 28530 16158 28542 16210
rect 34974 16146 35026 16158
rect 36430 16210 36482 16222
rect 40910 16210 40962 16222
rect 39890 16158 39902 16210
rect 39954 16158 39966 16210
rect 36430 16146 36482 16158
rect 40910 16146 40962 16158
rect 47518 16210 47570 16222
rect 47518 16146 47570 16158
rect 53006 16210 53058 16222
rect 53006 16146 53058 16158
rect 53566 16210 53618 16222
rect 53566 16146 53618 16158
rect 55918 16210 55970 16222
rect 55918 16146 55970 16158
rect 61070 16210 61122 16222
rect 61070 16146 61122 16158
rect 64318 16210 64370 16222
rect 72046 16210 72098 16222
rect 71250 16158 71262 16210
rect 71314 16158 71326 16210
rect 64318 16146 64370 16158
rect 72046 16146 72098 16158
rect 72494 16210 72546 16222
rect 72494 16146 72546 16158
rect 73166 16210 73218 16222
rect 73166 16146 73218 16158
rect 74286 16210 74338 16222
rect 74286 16146 74338 16158
rect 77982 16210 78034 16222
rect 77982 16146 78034 16158
rect 78430 16210 78482 16222
rect 78430 16146 78482 16158
rect 79998 16210 80050 16222
rect 79998 16146 80050 16158
rect 82126 16210 82178 16222
rect 82126 16146 82178 16158
rect 84142 16210 84194 16222
rect 90750 16210 90802 16222
rect 87154 16158 87166 16210
rect 87218 16158 87230 16210
rect 88946 16158 88958 16210
rect 89010 16158 89022 16210
rect 84142 16146 84194 16158
rect 90750 16146 90802 16158
rect 91982 16210 92034 16222
rect 91982 16146 92034 16158
rect 92878 16210 92930 16222
rect 92878 16146 92930 16158
rect 93998 16210 94050 16222
rect 93998 16146 94050 16158
rect 24894 16098 24946 16110
rect 30494 16098 30546 16110
rect 31838 16098 31890 16110
rect 17938 16046 17950 16098
rect 18002 16046 18014 16098
rect 21634 16046 21646 16098
rect 21698 16046 21710 16098
rect 25554 16046 25566 16098
rect 25618 16046 25630 16098
rect 29810 16046 29822 16098
rect 29874 16046 29886 16098
rect 30034 16046 30046 16098
rect 30098 16046 30110 16098
rect 30818 16046 30830 16098
rect 30882 16046 30894 16098
rect 24894 16034 24946 16046
rect 30494 16034 30546 16046
rect 31838 16034 31890 16046
rect 32510 16098 32562 16110
rect 32510 16034 32562 16046
rect 34078 16098 34130 16110
rect 40238 16098 40290 16110
rect 36978 16046 36990 16098
rect 37042 16046 37054 16098
rect 34078 16034 34130 16046
rect 40238 16034 40290 16046
rect 40574 16098 40626 16110
rect 40574 16034 40626 16046
rect 41134 16098 41186 16110
rect 41134 16034 41186 16046
rect 41358 16098 41410 16110
rect 41358 16034 41410 16046
rect 42030 16098 42082 16110
rect 42030 16034 42082 16046
rect 42142 16098 42194 16110
rect 49534 16098 49586 16110
rect 46834 16046 46846 16098
rect 46898 16046 46910 16098
rect 48066 16046 48078 16098
rect 48130 16046 48142 16098
rect 48626 16046 48638 16098
rect 48690 16046 48702 16098
rect 49186 16046 49198 16098
rect 49250 16046 49262 16098
rect 42142 16034 42194 16046
rect 49534 16034 49586 16046
rect 49870 16098 49922 16110
rect 57486 16098 57538 16110
rect 61966 16098 62018 16110
rect 73278 16098 73330 16110
rect 52882 16046 52894 16098
rect 52946 16046 52958 16098
rect 61394 16046 61406 16098
rect 61458 16046 61470 16098
rect 64530 16046 64542 16098
rect 64594 16046 64606 16098
rect 68450 16046 68462 16098
rect 68514 16046 68526 16098
rect 49870 16034 49922 16046
rect 57486 16034 57538 16046
rect 61966 16034 62018 16046
rect 73278 16034 73330 16046
rect 73614 16098 73666 16110
rect 73614 16034 73666 16046
rect 74846 16098 74898 16110
rect 74846 16034 74898 16046
rect 75070 16098 75122 16110
rect 75070 16034 75122 16046
rect 75294 16098 75346 16110
rect 75294 16034 75346 16046
rect 77086 16098 77138 16110
rect 77086 16034 77138 16046
rect 77646 16098 77698 16110
rect 77646 16034 77698 16046
rect 80558 16098 80610 16110
rect 80558 16034 80610 16046
rect 80782 16098 80834 16110
rect 80782 16034 80834 16046
rect 81342 16098 81394 16110
rect 90638 16098 90690 16110
rect 86930 16046 86942 16098
rect 86994 16046 87006 16098
rect 88834 16046 88846 16098
rect 88898 16046 88910 16098
rect 81342 16034 81394 16046
rect 90638 16034 90690 16046
rect 93550 16098 93602 16110
rect 93550 16034 93602 16046
rect 25230 15986 25282 15998
rect 33630 15986 33682 15998
rect 18610 15934 18622 15986
rect 18674 15934 18686 15986
rect 22418 15934 22430 15986
rect 22482 15934 22494 15986
rect 26338 15934 26350 15986
rect 26402 15934 26414 15986
rect 25230 15922 25282 15934
rect 33630 15922 33682 15934
rect 35758 15986 35810 15998
rect 40798 15986 40850 15998
rect 37762 15934 37774 15986
rect 37826 15934 37838 15986
rect 35758 15922 35810 15934
rect 40798 15922 40850 15934
rect 41694 15986 41746 15998
rect 41694 15922 41746 15934
rect 42814 15986 42866 15998
rect 42814 15922 42866 15934
rect 43150 15986 43202 15998
rect 43150 15922 43202 15934
rect 43598 15986 43650 15998
rect 43598 15922 43650 15934
rect 47294 15986 47346 15998
rect 47294 15922 47346 15934
rect 49758 15986 49810 15998
rect 49758 15922 49810 15934
rect 53118 15986 53170 15998
rect 56926 15986 56978 15998
rect 56578 15934 56590 15986
rect 56642 15934 56654 15986
rect 53118 15922 53170 15934
rect 56926 15922 56978 15934
rect 62078 15986 62130 15998
rect 62078 15922 62130 15934
rect 65102 15986 65154 15998
rect 73054 15986 73106 15998
rect 69122 15934 69134 15986
rect 69186 15934 69198 15986
rect 65102 15922 65154 15934
rect 73054 15922 73106 15934
rect 75630 15986 75682 15998
rect 75630 15922 75682 15934
rect 80334 15986 80386 15998
rect 80334 15922 80386 15934
rect 91086 15986 91138 15998
rect 94785 15986 94831 16273
rect 95330 16270 95342 16273
rect 95394 16270 95406 16322
rect 104626 16270 104638 16322
rect 104690 16319 104702 16322
rect 105298 16319 105310 16322
rect 104690 16273 105310 16319
rect 104690 16270 104702 16273
rect 105298 16270 105310 16273
rect 105362 16270 105374 16322
rect 95342 16210 95394 16222
rect 100270 16210 100322 16222
rect 104862 16210 104914 16222
rect 98802 16158 98814 16210
rect 98866 16158 98878 16210
rect 104402 16158 104414 16210
rect 104466 16158 104478 16210
rect 95342 16146 95394 16158
rect 100270 16146 100322 16158
rect 104862 16146 104914 16158
rect 105310 16210 105362 16222
rect 105310 16146 105362 16158
rect 107886 16098 107938 16110
rect 95778 16046 95790 16098
rect 95842 16046 95854 16098
rect 96450 16046 96462 16098
rect 96514 16046 96526 16098
rect 101490 16046 101502 16098
rect 101554 16046 101566 16098
rect 101938 16046 101950 16098
rect 102002 16046 102014 16098
rect 107886 16034 107938 16046
rect 108558 16098 108610 16110
rect 108558 16034 108610 16046
rect 110238 16098 110290 16110
rect 110238 16034 110290 16046
rect 112366 16098 112418 16110
rect 112366 16034 112418 16046
rect 94770 15934 94782 15986
rect 94834 15934 94846 15986
rect 91086 15922 91138 15934
rect 25118 15874 25170 15886
rect 25118 15810 25170 15822
rect 29598 15874 29650 15886
rect 29598 15810 29650 15822
rect 30270 15874 30322 15886
rect 30270 15810 30322 15822
rect 30382 15874 30434 15886
rect 30382 15810 30434 15822
rect 31054 15874 31106 15886
rect 31054 15810 31106 15822
rect 31950 15874 32002 15886
rect 31950 15810 32002 15822
rect 32622 15874 32674 15886
rect 32622 15810 32674 15822
rect 34414 15874 34466 15886
rect 34414 15810 34466 15822
rect 35534 15874 35586 15886
rect 35534 15810 35586 15822
rect 35870 15874 35922 15886
rect 35870 15810 35922 15822
rect 36094 15874 36146 15886
rect 36094 15810 36146 15822
rect 40350 15874 40402 15886
rect 40350 15810 40402 15822
rect 41806 15874 41858 15886
rect 41806 15810 41858 15822
rect 47406 15874 47458 15886
rect 47406 15810 47458 15822
rect 47630 15874 47682 15886
rect 47630 15810 47682 15822
rect 51774 15874 51826 15886
rect 51774 15810 51826 15822
rect 52222 15874 52274 15886
rect 52222 15810 52274 15822
rect 52670 15874 52722 15886
rect 52670 15810 52722 15822
rect 54126 15874 54178 15886
rect 54126 15810 54178 15822
rect 56254 15874 56306 15886
rect 56254 15810 56306 15822
rect 61518 15874 61570 15886
rect 61518 15810 61570 15822
rect 62638 15874 62690 15886
rect 75182 15874 75234 15886
rect 64082 15822 64094 15874
rect 64146 15822 64158 15874
rect 62638 15810 62690 15822
rect 75182 15810 75234 15822
rect 76302 15874 76354 15886
rect 76302 15810 76354 15822
rect 76974 15874 77026 15886
rect 76974 15810 77026 15822
rect 77198 15874 77250 15886
rect 77198 15810 77250 15822
rect 78990 15874 79042 15886
rect 78990 15810 79042 15822
rect 79438 15874 79490 15886
rect 79438 15810 79490 15822
rect 80558 15874 80610 15886
rect 82686 15874 82738 15886
rect 81666 15822 81678 15874
rect 81730 15822 81742 15874
rect 80558 15810 80610 15822
rect 82686 15810 82738 15822
rect 83134 15874 83186 15886
rect 83134 15810 83186 15822
rect 83582 15874 83634 15886
rect 83582 15810 83634 15822
rect 84590 15874 84642 15886
rect 84590 15810 84642 15822
rect 85150 15874 85202 15886
rect 85150 15810 85202 15822
rect 85598 15874 85650 15886
rect 85598 15810 85650 15822
rect 85934 15874 85986 15886
rect 85934 15810 85986 15822
rect 86494 15874 86546 15886
rect 86494 15810 86546 15822
rect 90862 15874 90914 15886
rect 90862 15810 90914 15822
rect 92430 15874 92482 15886
rect 92430 15810 92482 15822
rect 94558 15874 94610 15886
rect 94558 15810 94610 15822
rect 94894 15874 94946 15886
rect 94894 15810 94946 15822
rect 99822 15874 99874 15886
rect 99822 15810 99874 15822
rect 100830 15874 100882 15886
rect 100830 15810 100882 15822
rect 105758 15874 105810 15886
rect 105758 15810 105810 15822
rect 106318 15874 106370 15886
rect 106318 15810 106370 15822
rect 106990 15874 107042 15886
rect 106990 15810 107042 15822
rect 107998 15874 108050 15886
rect 107998 15810 108050 15822
rect 108110 15874 108162 15886
rect 108110 15810 108162 15822
rect 108894 15874 108946 15886
rect 108894 15810 108946 15822
rect 110350 15874 110402 15886
rect 110350 15810 110402 15822
rect 112478 15874 112530 15886
rect 112478 15810 112530 15822
rect 1344 15706 158592 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 81278 15706
rect 81330 15654 81382 15706
rect 81434 15654 81486 15706
rect 81538 15654 111998 15706
rect 112050 15654 112102 15706
rect 112154 15654 112206 15706
rect 112258 15654 142718 15706
rect 142770 15654 142822 15706
rect 142874 15654 142926 15706
rect 142978 15654 158592 15706
rect 1344 15620 158592 15654
rect 20414 15538 20466 15550
rect 20414 15474 20466 15486
rect 20750 15538 20802 15550
rect 20750 15474 20802 15486
rect 22318 15538 22370 15550
rect 22318 15474 22370 15486
rect 22766 15538 22818 15550
rect 22766 15474 22818 15486
rect 26014 15538 26066 15550
rect 26014 15474 26066 15486
rect 27582 15538 27634 15550
rect 27582 15474 27634 15486
rect 27918 15538 27970 15550
rect 27918 15474 27970 15486
rect 28814 15538 28866 15550
rect 28814 15474 28866 15486
rect 34078 15538 34130 15550
rect 34078 15474 34130 15486
rect 35982 15538 36034 15550
rect 35982 15474 36034 15486
rect 36542 15538 36594 15550
rect 36542 15474 36594 15486
rect 37326 15538 37378 15550
rect 37326 15474 37378 15486
rect 38334 15538 38386 15550
rect 38334 15474 38386 15486
rect 44270 15538 44322 15550
rect 44270 15474 44322 15486
rect 48862 15538 48914 15550
rect 48862 15474 48914 15486
rect 49422 15538 49474 15550
rect 49422 15474 49474 15486
rect 54126 15538 54178 15550
rect 54126 15474 54178 15486
rect 54350 15538 54402 15550
rect 54350 15474 54402 15486
rect 55134 15538 55186 15550
rect 55134 15474 55186 15486
rect 57150 15538 57202 15550
rect 57150 15474 57202 15486
rect 57374 15538 57426 15550
rect 57374 15474 57426 15486
rect 60510 15538 60562 15550
rect 60510 15474 60562 15486
rect 68350 15538 68402 15550
rect 68350 15474 68402 15486
rect 69694 15538 69746 15550
rect 69694 15474 69746 15486
rect 70142 15538 70194 15550
rect 70142 15474 70194 15486
rect 71486 15538 71538 15550
rect 71486 15474 71538 15486
rect 73838 15538 73890 15550
rect 73838 15474 73890 15486
rect 78430 15538 78482 15550
rect 78430 15474 78482 15486
rect 79550 15538 79602 15550
rect 79550 15474 79602 15486
rect 87278 15538 87330 15550
rect 92094 15538 92146 15550
rect 87938 15486 87950 15538
rect 88002 15486 88014 15538
rect 87278 15474 87330 15486
rect 92094 15474 92146 15486
rect 94334 15538 94386 15550
rect 94334 15474 94386 15486
rect 100270 15538 100322 15550
rect 100270 15474 100322 15486
rect 101726 15538 101778 15550
rect 101726 15474 101778 15486
rect 102062 15538 102114 15550
rect 102062 15474 102114 15486
rect 102174 15538 102226 15550
rect 102174 15474 102226 15486
rect 102510 15538 102562 15550
rect 102510 15474 102562 15486
rect 107550 15538 107602 15550
rect 107550 15474 107602 15486
rect 108222 15538 108274 15550
rect 108222 15474 108274 15486
rect 108782 15538 108834 15550
rect 108782 15474 108834 15486
rect 109230 15538 109282 15550
rect 109230 15474 109282 15486
rect 20862 15426 20914 15438
rect 20862 15362 20914 15374
rect 21982 15426 22034 15438
rect 21982 15362 22034 15374
rect 22206 15426 22258 15438
rect 22206 15362 22258 15374
rect 22878 15426 22930 15438
rect 22878 15362 22930 15374
rect 23326 15426 23378 15438
rect 23326 15362 23378 15374
rect 25230 15426 25282 15438
rect 25230 15362 25282 15374
rect 26126 15426 26178 15438
rect 26126 15362 26178 15374
rect 35758 15426 35810 15438
rect 35758 15362 35810 15374
rect 36318 15426 36370 15438
rect 36318 15362 36370 15374
rect 37662 15426 37714 15438
rect 37662 15362 37714 15374
rect 38110 15426 38162 15438
rect 48974 15426 49026 15438
rect 70926 15426 70978 15438
rect 41682 15374 41694 15426
rect 41746 15374 41758 15426
rect 46050 15374 46062 15426
rect 46114 15374 46126 15426
rect 57698 15374 57710 15426
rect 57762 15374 57774 15426
rect 38110 15362 38162 15374
rect 48974 15362 49026 15374
rect 70926 15362 70978 15374
rect 72494 15426 72546 15438
rect 72494 15362 72546 15374
rect 74286 15426 74338 15438
rect 83470 15426 83522 15438
rect 100382 15426 100434 15438
rect 75842 15374 75854 15426
rect 75906 15374 75918 15426
rect 80882 15374 80894 15426
rect 80946 15374 80958 15426
rect 89394 15374 89406 15426
rect 89458 15374 89470 15426
rect 74286 15362 74338 15374
rect 83470 15362 83522 15374
rect 100382 15362 100434 15374
rect 101614 15426 101666 15438
rect 101614 15362 101666 15374
rect 108446 15426 108498 15438
rect 108446 15362 108498 15374
rect 108894 15426 108946 15438
rect 108894 15362 108946 15374
rect 20638 15314 20690 15326
rect 22430 15314 22482 15326
rect 21186 15262 21198 15314
rect 21250 15262 21262 15314
rect 20638 15250 20690 15262
rect 22430 15250 22482 15262
rect 25342 15314 25394 15326
rect 27470 15314 27522 15326
rect 25778 15262 25790 15314
rect 25842 15262 25854 15314
rect 25342 15250 25394 15262
rect 27470 15250 27522 15262
rect 27694 15314 27746 15326
rect 27694 15250 27746 15262
rect 35646 15314 35698 15326
rect 35646 15250 35698 15262
rect 36206 15314 36258 15326
rect 36206 15250 36258 15262
rect 36990 15314 37042 15326
rect 36990 15250 37042 15262
rect 37326 15314 37378 15326
rect 37326 15250 37378 15262
rect 37998 15314 38050 15326
rect 54798 15314 54850 15326
rect 63198 15314 63250 15326
rect 41010 15262 41022 15314
rect 41074 15262 41086 15314
rect 45266 15262 45278 15314
rect 45330 15262 45342 15314
rect 53778 15262 53790 15314
rect 53842 15262 53854 15314
rect 61394 15262 61406 15314
rect 61458 15262 61470 15314
rect 37998 15250 38050 15262
rect 54798 15250 54850 15262
rect 63198 15250 63250 15262
rect 63758 15314 63810 15326
rect 68014 15314 68066 15326
rect 64418 15262 64430 15314
rect 64482 15262 64494 15314
rect 63758 15250 63810 15262
rect 68014 15250 68066 15262
rect 68462 15314 68514 15326
rect 68462 15250 68514 15262
rect 68686 15314 68738 15326
rect 68686 15250 68738 15262
rect 70702 15314 70754 15326
rect 70702 15250 70754 15262
rect 71038 15314 71090 15326
rect 100046 15314 100098 15326
rect 75170 15262 75182 15314
rect 75234 15262 75246 15314
rect 80098 15262 80110 15314
rect 80162 15262 80174 15314
rect 86818 15262 86830 15314
rect 86882 15262 86894 15314
rect 88162 15262 88174 15314
rect 88226 15262 88238 15314
rect 88722 15262 88734 15314
rect 88786 15262 88798 15314
rect 93314 15262 93326 15314
rect 93378 15262 93390 15314
rect 96002 15262 96014 15314
rect 96066 15262 96078 15314
rect 97570 15262 97582 15314
rect 97634 15262 97646 15314
rect 97906 15262 97918 15314
rect 97970 15262 97982 15314
rect 71038 15250 71090 15262
rect 100046 15250 100098 15262
rect 100606 15314 100658 15326
rect 100606 15250 100658 15262
rect 101054 15314 101106 15326
rect 101054 15250 101106 15262
rect 101502 15314 101554 15326
rect 101502 15250 101554 15262
rect 102286 15314 102338 15326
rect 107998 15314 108050 15326
rect 103506 15262 103518 15314
rect 103570 15262 103582 15314
rect 104178 15262 104190 15314
rect 104242 15262 104254 15314
rect 106642 15262 106654 15314
rect 106706 15262 106718 15314
rect 102286 15250 102338 15262
rect 107998 15250 108050 15262
rect 108110 15314 108162 15326
rect 108110 15250 108162 15262
rect 109006 15314 109058 15326
rect 109006 15250 109058 15262
rect 24670 15202 24722 15214
rect 24670 15138 24722 15150
rect 39006 15202 39058 15214
rect 39006 15138 39058 15150
rect 39454 15202 39506 15214
rect 54238 15202 54290 15214
rect 43810 15150 43822 15202
rect 43874 15150 43886 15202
rect 48178 15150 48190 15202
rect 48242 15150 48254 15202
rect 50866 15150 50878 15202
rect 50930 15150 50942 15202
rect 52994 15150 53006 15202
rect 53058 15150 53070 15202
rect 39454 15138 39506 15150
rect 54238 15138 54290 15150
rect 58270 15202 58322 15214
rect 58270 15138 58322 15150
rect 58718 15202 58770 15214
rect 58718 15138 58770 15150
rect 59502 15202 59554 15214
rect 59502 15138 59554 15150
rect 60286 15202 60338 15214
rect 60286 15138 60338 15150
rect 61070 15202 61122 15214
rect 69134 15202 69186 15214
rect 62178 15150 62190 15202
rect 62242 15150 62254 15202
rect 65202 15150 65214 15202
rect 65266 15150 65278 15202
rect 67330 15150 67342 15202
rect 67394 15150 67406 15202
rect 61070 15138 61122 15150
rect 69134 15138 69186 15150
rect 70590 15202 70642 15214
rect 70590 15138 70642 15150
rect 73166 15202 73218 15214
rect 73166 15138 73218 15150
rect 74734 15202 74786 15214
rect 79102 15202 79154 15214
rect 103070 15202 103122 15214
rect 77970 15150 77982 15202
rect 78034 15150 78046 15202
rect 83010 15150 83022 15202
rect 83074 15150 83086 15202
rect 83906 15150 83918 15202
rect 83970 15150 83982 15202
rect 86034 15150 86046 15202
rect 86098 15150 86110 15202
rect 91522 15150 91534 15202
rect 91586 15150 91598 15202
rect 93986 15150 93998 15202
rect 94050 15150 94062 15202
rect 95106 15150 95118 15202
rect 95170 15150 95182 15202
rect 95890 15150 95902 15202
rect 95954 15150 95966 15202
rect 74734 15138 74786 15150
rect 79102 15138 79154 15150
rect 103070 15138 103122 15150
rect 107102 15202 107154 15214
rect 107102 15138 107154 15150
rect 109790 15202 109842 15214
rect 109790 15138 109842 15150
rect 48862 15090 48914 15102
rect 48862 15026 48914 15038
rect 92878 15090 92930 15102
rect 98802 15038 98814 15090
rect 98866 15038 98878 15090
rect 92878 15026 92930 15038
rect 1344 14922 158592 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 96638 14922
rect 96690 14870 96742 14922
rect 96794 14870 96846 14922
rect 96898 14870 127358 14922
rect 127410 14870 127462 14922
rect 127514 14870 127566 14922
rect 127618 14870 158078 14922
rect 158130 14870 158182 14922
rect 158234 14870 158286 14922
rect 158338 14870 158592 14922
rect 1344 14836 158592 14870
rect 44942 14754 44994 14766
rect 81454 14754 81506 14766
rect 37538 14702 37550 14754
rect 37602 14751 37614 14754
rect 37874 14751 37886 14754
rect 37602 14705 37886 14751
rect 37602 14702 37614 14705
rect 37874 14702 37886 14705
rect 37938 14751 37950 14754
rect 38322 14751 38334 14754
rect 37938 14705 38334 14751
rect 37938 14702 37950 14705
rect 38322 14702 38334 14705
rect 38386 14702 38398 14754
rect 38994 14702 39006 14754
rect 39058 14751 39070 14754
rect 39330 14751 39342 14754
rect 39058 14705 39342 14751
rect 39058 14702 39070 14705
rect 39330 14702 39342 14705
rect 39394 14751 39406 14754
rect 39778 14751 39790 14754
rect 39394 14705 39790 14751
rect 39394 14702 39406 14705
rect 39778 14702 39790 14705
rect 39842 14702 39854 14754
rect 57698 14702 57710 14754
rect 57762 14751 57774 14754
rect 57762 14705 58207 14751
rect 57762 14702 57774 14705
rect 44942 14690 44994 14702
rect 37550 14642 37602 14654
rect 19954 14590 19966 14642
rect 20018 14590 20030 14642
rect 33954 14590 33966 14642
rect 34018 14590 34030 14642
rect 37550 14578 37602 14590
rect 39006 14642 39058 14654
rect 39006 14578 39058 14590
rect 42142 14642 42194 14654
rect 42142 14578 42194 14590
rect 48638 14642 48690 14654
rect 48638 14578 48690 14590
rect 57822 14642 57874 14654
rect 58161 14639 58207 14705
rect 62514 14702 62526 14754
rect 62578 14751 62590 14754
rect 63410 14751 63422 14754
rect 62578 14705 63422 14751
rect 62578 14702 62590 14705
rect 63410 14702 63422 14705
rect 63474 14702 63486 14754
rect 73490 14751 73502 14754
rect 72497 14705 73502 14751
rect 62526 14642 62578 14654
rect 58370 14639 58382 14642
rect 58161 14593 58382 14639
rect 58370 14590 58382 14593
rect 58434 14590 58446 14642
rect 59378 14590 59390 14642
rect 59442 14590 59454 14642
rect 57822 14578 57874 14590
rect 62526 14578 62578 14590
rect 62862 14642 62914 14654
rect 62862 14578 62914 14590
rect 63310 14642 63362 14654
rect 72382 14642 72434 14654
rect 71810 14590 71822 14642
rect 71874 14590 71886 14642
rect 63310 14578 63362 14590
rect 72382 14578 72434 14590
rect 37102 14530 37154 14542
rect 17154 14478 17166 14530
rect 17218 14478 17230 14530
rect 31042 14478 31054 14530
rect 31106 14478 31118 14530
rect 37102 14466 37154 14478
rect 47966 14530 48018 14542
rect 47966 14466 48018 14478
rect 52670 14530 52722 14542
rect 52670 14466 52722 14478
rect 52894 14530 52946 14542
rect 52894 14466 52946 14478
rect 53230 14530 53282 14542
rect 61406 14530 61458 14542
rect 58370 14478 58382 14530
rect 58434 14478 58446 14530
rect 53230 14466 53282 14478
rect 61406 14466 61458 14478
rect 61630 14530 61682 14542
rect 61630 14466 61682 14478
rect 62078 14530 62130 14542
rect 72497 14530 72543 14705
rect 73490 14702 73502 14705
rect 73554 14751 73566 14754
rect 74386 14751 74398 14754
rect 73554 14705 74398 14751
rect 73554 14702 73566 14705
rect 74386 14702 74398 14705
rect 74450 14702 74462 14754
rect 89058 14702 89070 14754
rect 89122 14702 89134 14754
rect 94434 14702 94446 14754
rect 94498 14702 94510 14754
rect 81454 14690 81506 14702
rect 72942 14642 72994 14654
rect 72942 14578 72994 14590
rect 76750 14642 76802 14654
rect 76750 14578 76802 14590
rect 83134 14642 83186 14654
rect 83134 14578 83186 14590
rect 85262 14642 85314 14654
rect 85262 14578 85314 14590
rect 92094 14642 92146 14654
rect 98254 14642 98306 14654
rect 95218 14590 95230 14642
rect 95282 14590 95294 14642
rect 92094 14578 92146 14590
rect 98254 14578 98306 14590
rect 98702 14642 98754 14654
rect 98702 14578 98754 14590
rect 99038 14642 99090 14654
rect 106082 14590 106094 14642
rect 106146 14590 106158 14642
rect 110562 14590 110574 14642
rect 110626 14590 110638 14642
rect 99038 14578 99090 14590
rect 82686 14530 82738 14542
rect 88174 14530 88226 14542
rect 92878 14530 92930 14542
rect 106430 14530 106482 14542
rect 69010 14478 69022 14530
rect 69074 14478 69086 14530
rect 72482 14478 72494 14530
rect 72546 14478 72558 14530
rect 77074 14478 77086 14530
rect 77138 14478 77150 14530
rect 79202 14478 79214 14530
rect 79266 14478 79278 14530
rect 80770 14478 80782 14530
rect 80834 14478 80846 14530
rect 84690 14478 84702 14530
rect 84754 14478 84766 14530
rect 86818 14478 86830 14530
rect 86882 14478 86894 14530
rect 88834 14478 88846 14530
rect 88898 14478 88910 14530
rect 90066 14478 90078 14530
rect 90130 14478 90142 14530
rect 93090 14478 93102 14530
rect 93154 14478 93166 14530
rect 94882 14478 94894 14530
rect 94946 14478 94958 14530
rect 99586 14478 99598 14530
rect 99650 14478 99662 14530
rect 100258 14478 100270 14530
rect 100322 14478 100334 14530
rect 103170 14478 103182 14530
rect 103234 14478 103246 14530
rect 103730 14478 103742 14530
rect 103794 14478 103806 14530
rect 62078 14466 62130 14478
rect 82686 14466 82738 14478
rect 88174 14466 88226 14478
rect 92878 14466 92930 14478
rect 106430 14466 106482 14478
rect 106654 14530 106706 14542
rect 106654 14466 106706 14478
rect 106990 14530 107042 14542
rect 107650 14478 107662 14530
rect 107714 14478 107726 14530
rect 108098 14478 108110 14530
rect 108162 14478 108174 14530
rect 106990 14466 107042 14478
rect 29150 14418 29202 14430
rect 17826 14366 17838 14418
rect 17890 14366 17902 14418
rect 29150 14354 29202 14366
rect 29262 14418 29314 14430
rect 38446 14418 38498 14430
rect 31826 14366 31838 14418
rect 31890 14366 31902 14418
rect 29262 14354 29314 14366
rect 38446 14354 38498 14366
rect 44830 14418 44882 14430
rect 44830 14354 44882 14366
rect 64990 14418 65042 14430
rect 64990 14354 65042 14366
rect 65326 14418 65378 14430
rect 65326 14354 65378 14366
rect 65550 14418 65602 14430
rect 65550 14354 65602 14366
rect 65886 14418 65938 14430
rect 65886 14354 65938 14366
rect 66446 14418 66498 14430
rect 66446 14354 66498 14366
rect 66670 14418 66722 14430
rect 66670 14354 66722 14366
rect 66782 14418 66834 14430
rect 75182 14418 75234 14430
rect 81566 14418 81618 14430
rect 69682 14366 69694 14418
rect 69746 14366 69758 14418
rect 77858 14366 77870 14418
rect 77922 14366 77934 14418
rect 81106 14366 81118 14418
rect 81170 14366 81182 14418
rect 66782 14354 66834 14366
rect 75182 14354 75234 14366
rect 81566 14354 81618 14366
rect 20414 14306 20466 14318
rect 20414 14242 20466 14254
rect 25230 14306 25282 14318
rect 25230 14242 25282 14254
rect 29710 14306 29762 14318
rect 29710 14242 29762 14254
rect 34414 14306 34466 14318
rect 34414 14242 34466 14254
rect 34862 14306 34914 14318
rect 34862 14242 34914 14254
rect 35310 14306 35362 14318
rect 35310 14242 35362 14254
rect 35758 14306 35810 14318
rect 35758 14242 35810 14254
rect 38110 14306 38162 14318
rect 38110 14242 38162 14254
rect 39454 14306 39506 14318
rect 39454 14242 39506 14254
rect 39902 14306 39954 14318
rect 39902 14242 39954 14254
rect 41806 14306 41858 14318
rect 41806 14242 41858 14254
rect 42702 14306 42754 14318
rect 42702 14242 42754 14254
rect 46062 14306 46114 14318
rect 46062 14242 46114 14254
rect 47742 14306 47794 14318
rect 47742 14242 47794 14254
rect 48078 14306 48130 14318
rect 48078 14242 48130 14254
rect 49422 14306 49474 14318
rect 49422 14242 49474 14254
rect 49758 14306 49810 14318
rect 49758 14242 49810 14254
rect 53006 14306 53058 14318
rect 53006 14242 53058 14254
rect 54014 14306 54066 14318
rect 54014 14242 54066 14254
rect 54574 14306 54626 14318
rect 54574 14242 54626 14254
rect 57038 14306 57090 14318
rect 57038 14242 57090 14254
rect 57486 14306 57538 14318
rect 57486 14242 57538 14254
rect 60734 14306 60786 14318
rect 60734 14242 60786 14254
rect 61070 14306 61122 14318
rect 61070 14242 61122 14254
rect 61518 14306 61570 14318
rect 61518 14242 61570 14254
rect 64094 14306 64146 14318
rect 64094 14242 64146 14254
rect 64542 14306 64594 14318
rect 64542 14242 64594 14254
rect 65214 14306 65266 14318
rect 65214 14242 65266 14254
rect 66222 14306 66274 14318
rect 66222 14242 66274 14254
rect 68574 14306 68626 14318
rect 68574 14242 68626 14254
rect 73390 14306 73442 14318
rect 73390 14242 73442 14254
rect 73950 14306 74002 14318
rect 73950 14242 74002 14254
rect 74286 14306 74338 14318
rect 74286 14242 74338 14254
rect 74846 14306 74898 14318
rect 74846 14242 74898 14254
rect 75294 14306 75346 14318
rect 75294 14242 75346 14254
rect 81230 14306 81282 14318
rect 81230 14242 81282 14254
rect 81902 14306 81954 14318
rect 81902 14242 81954 14254
rect 84030 14306 84082 14318
rect 84030 14242 84082 14254
rect 85822 14306 85874 14318
rect 85822 14242 85874 14254
rect 86270 14306 86322 14318
rect 86270 14242 86322 14254
rect 90750 14306 90802 14318
rect 90750 14242 90802 14254
rect 91086 14306 91138 14318
rect 91086 14242 91138 14254
rect 92430 14306 92482 14318
rect 92430 14242 92482 14254
rect 96910 14306 96962 14318
rect 96910 14242 96962 14254
rect 97470 14306 97522 14318
rect 97470 14242 97522 14254
rect 97806 14306 97858 14318
rect 97806 14242 97858 14254
rect 99150 14306 99202 14318
rect 106654 14306 106706 14318
rect 102722 14254 102734 14306
rect 102786 14254 102798 14306
rect 99150 14242 99202 14254
rect 106654 14242 106706 14254
rect 1344 14138 158592 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 81278 14138
rect 81330 14086 81382 14138
rect 81434 14086 81486 14138
rect 81538 14086 111998 14138
rect 112050 14086 112102 14138
rect 112154 14086 112206 14138
rect 112258 14086 142718 14138
rect 142770 14086 142822 14138
rect 142874 14086 142926 14138
rect 142978 14086 158592 14138
rect 1344 14052 158592 14086
rect 24558 13970 24610 13982
rect 24558 13906 24610 13918
rect 25678 13970 25730 13982
rect 25678 13906 25730 13918
rect 30158 13970 30210 13982
rect 30158 13906 30210 13918
rect 32510 13970 32562 13982
rect 37102 13970 37154 13982
rect 34178 13918 34190 13970
rect 34242 13918 34254 13970
rect 32510 13906 32562 13918
rect 37102 13906 37154 13918
rect 41694 13970 41746 13982
rect 41694 13906 41746 13918
rect 42142 13970 42194 13982
rect 42142 13906 42194 13918
rect 42590 13970 42642 13982
rect 42590 13906 42642 13918
rect 44494 13970 44546 13982
rect 44494 13906 44546 13918
rect 44942 13970 44994 13982
rect 44942 13906 44994 13918
rect 46398 13970 46450 13982
rect 46398 13906 46450 13918
rect 49198 13970 49250 13982
rect 49198 13906 49250 13918
rect 50206 13970 50258 13982
rect 50206 13906 50258 13918
rect 50766 13970 50818 13982
rect 63758 13970 63810 13982
rect 62850 13918 62862 13970
rect 62914 13918 62926 13970
rect 50766 13906 50818 13918
rect 63758 13906 63810 13918
rect 64542 13970 64594 13982
rect 64542 13906 64594 13918
rect 66670 13970 66722 13982
rect 66670 13906 66722 13918
rect 68910 13970 68962 13982
rect 68910 13906 68962 13918
rect 69470 13970 69522 13982
rect 69470 13906 69522 13918
rect 70814 13970 70866 13982
rect 70814 13906 70866 13918
rect 71262 13970 71314 13982
rect 71262 13906 71314 13918
rect 72382 13970 72434 13982
rect 72382 13906 72434 13918
rect 73502 13970 73554 13982
rect 79214 13970 79266 13982
rect 78642 13918 78654 13970
rect 78706 13918 78718 13970
rect 73502 13906 73554 13918
rect 79214 13906 79266 13918
rect 80334 13970 80386 13982
rect 86942 13970 86994 13982
rect 85922 13918 85934 13970
rect 85986 13918 85998 13970
rect 80334 13906 80386 13918
rect 86942 13906 86994 13918
rect 87390 13970 87442 13982
rect 87390 13906 87442 13918
rect 93102 13970 93154 13982
rect 93102 13906 93154 13918
rect 93886 13970 93938 13982
rect 93886 13906 93938 13918
rect 103742 13970 103794 13982
rect 103742 13906 103794 13918
rect 107214 13970 107266 13982
rect 110562 13918 110574 13970
rect 110626 13918 110638 13970
rect 107214 13906 107266 13918
rect 31166 13858 31218 13870
rect 31166 13794 31218 13806
rect 62526 13858 62578 13870
rect 62526 13794 62578 13806
rect 65662 13858 65714 13870
rect 65662 13794 65714 13806
rect 65774 13858 65826 13870
rect 93550 13858 93602 13870
rect 75506 13806 75518 13858
rect 75570 13806 75582 13858
rect 84578 13806 84590 13858
rect 84642 13806 84654 13858
rect 65774 13794 65826 13806
rect 93550 13794 93602 13806
rect 103630 13858 103682 13870
rect 103630 13794 103682 13806
rect 103966 13858 104018 13870
rect 103966 13794 104018 13806
rect 104190 13858 104242 13870
rect 104190 13794 104242 13806
rect 104638 13858 104690 13870
rect 104638 13794 104690 13806
rect 105198 13858 105250 13870
rect 105198 13794 105250 13806
rect 105534 13858 105586 13870
rect 105534 13794 105586 13806
rect 106094 13858 106146 13870
rect 106094 13794 106146 13806
rect 106654 13858 106706 13870
rect 106654 13794 106706 13806
rect 111470 13858 111522 13870
rect 111470 13794 111522 13806
rect 29710 13746 29762 13758
rect 20066 13694 20078 13746
rect 20130 13694 20142 13746
rect 26674 13694 26686 13746
rect 26738 13694 26750 13746
rect 29710 13682 29762 13694
rect 30382 13746 30434 13758
rect 34302 13746 34354 13758
rect 33842 13694 33854 13746
rect 33906 13694 33918 13746
rect 30382 13682 30434 13694
rect 34302 13682 34354 13694
rect 34638 13746 34690 13758
rect 41022 13746 41074 13758
rect 55134 13746 55186 13758
rect 35298 13694 35310 13746
rect 35362 13694 35374 13746
rect 37426 13694 37438 13746
rect 37490 13694 37502 13746
rect 45826 13694 45838 13746
rect 45890 13694 45902 13746
rect 52658 13694 52670 13746
rect 52722 13694 52734 13746
rect 34638 13682 34690 13694
rect 41022 13682 41074 13694
rect 55134 13682 55186 13694
rect 56590 13746 56642 13758
rect 56590 13682 56642 13694
rect 56814 13746 56866 13758
rect 64430 13746 64482 13758
rect 57138 13694 57150 13746
rect 57202 13694 57214 13746
rect 59378 13694 59390 13746
rect 59442 13694 59454 13746
rect 56814 13682 56866 13694
rect 64430 13682 64482 13694
rect 64654 13746 64706 13758
rect 65438 13746 65490 13758
rect 64978 13694 64990 13746
rect 65042 13694 65054 13746
rect 64654 13682 64706 13694
rect 65438 13682 65490 13694
rect 66222 13746 66274 13758
rect 66222 13682 66274 13694
rect 69134 13746 69186 13758
rect 69134 13682 69186 13694
rect 69582 13746 69634 13758
rect 69582 13682 69634 13694
rect 69806 13746 69858 13758
rect 69806 13682 69858 13694
rect 71038 13746 71090 13758
rect 71038 13682 71090 13694
rect 71374 13746 71426 13758
rect 71374 13682 71426 13694
rect 72494 13746 72546 13758
rect 77422 13746 77474 13758
rect 102734 13746 102786 13758
rect 74946 13694 74958 13746
rect 75010 13694 75022 13746
rect 76402 13694 76414 13746
rect 76466 13694 76478 13746
rect 78194 13694 78206 13746
rect 78258 13694 78270 13746
rect 81106 13694 81118 13746
rect 81170 13694 81182 13746
rect 82562 13694 82574 13746
rect 82626 13694 82638 13746
rect 82898 13694 82910 13746
rect 82962 13694 82974 13746
rect 83906 13694 83918 13746
rect 83970 13694 83982 13746
rect 85698 13694 85710 13746
rect 85762 13694 85774 13746
rect 89058 13694 89070 13746
rect 89122 13694 89134 13746
rect 90738 13694 90750 13746
rect 90802 13694 90814 13746
rect 96002 13694 96014 13746
rect 96066 13694 96078 13746
rect 97794 13694 97806 13746
rect 97858 13694 97870 13746
rect 100258 13694 100270 13746
rect 100322 13694 100334 13746
rect 72494 13682 72546 13694
rect 77422 13682 77474 13694
rect 102734 13682 102786 13694
rect 104526 13746 104578 13758
rect 104526 13682 104578 13694
rect 104862 13746 104914 13758
rect 104862 13682 104914 13694
rect 106206 13746 106258 13758
rect 107650 13694 107662 13746
rect 107714 13694 107726 13746
rect 108210 13694 108222 13746
rect 108274 13694 108286 13746
rect 106206 13682 106258 13694
rect 19742 13634 19794 13646
rect 20974 13634 21026 13646
rect 20178 13582 20190 13634
rect 20242 13582 20254 13634
rect 19742 13570 19794 13582
rect 20974 13570 21026 13582
rect 21422 13634 21474 13646
rect 21422 13570 21474 13582
rect 24670 13634 24722 13646
rect 30270 13634 30322 13646
rect 27346 13582 27358 13634
rect 27410 13582 27422 13634
rect 29474 13582 29486 13634
rect 29538 13582 29550 13634
rect 24670 13570 24722 13582
rect 30270 13570 30322 13582
rect 31614 13634 31666 13646
rect 31614 13570 31666 13582
rect 32174 13634 32226 13646
rect 32174 13570 32226 13582
rect 33518 13634 33570 13646
rect 33518 13570 33570 13582
rect 35086 13634 35138 13646
rect 35086 13570 35138 13582
rect 35758 13634 35810 13646
rect 35758 13570 35810 13582
rect 36206 13634 36258 13646
rect 36206 13570 36258 13582
rect 36766 13634 36818 13646
rect 43150 13634 43202 13646
rect 38210 13582 38222 13634
rect 38274 13582 38286 13634
rect 40338 13582 40350 13634
rect 40402 13582 40414 13634
rect 36766 13570 36818 13582
rect 43150 13570 43202 13582
rect 43710 13634 43762 13646
rect 43710 13570 43762 13582
rect 44158 13634 44210 13646
rect 44158 13570 44210 13582
rect 45614 13634 45666 13646
rect 45614 13570 45666 13582
rect 46846 13634 46898 13646
rect 46846 13570 46898 13582
rect 47406 13634 47458 13646
rect 47406 13570 47458 13582
rect 47742 13634 47794 13646
rect 47742 13570 47794 13582
rect 48190 13634 48242 13646
rect 48190 13570 48242 13582
rect 49646 13634 49698 13646
rect 49646 13570 49698 13582
rect 50878 13634 50930 13646
rect 50878 13570 50930 13582
rect 51886 13634 51938 13646
rect 55918 13634 55970 13646
rect 54450 13582 54462 13634
rect 54514 13582 54526 13634
rect 51886 13570 51938 13582
rect 55918 13570 55970 13582
rect 56702 13634 56754 13646
rect 56702 13570 56754 13582
rect 57598 13634 57650 13646
rect 57598 13570 57650 13582
rect 58046 13634 58098 13646
rect 58046 13570 58098 13582
rect 58606 13634 58658 13646
rect 58606 13570 58658 13582
rect 58942 13634 58994 13646
rect 63310 13634 63362 13646
rect 67230 13634 67282 13646
rect 60050 13582 60062 13634
rect 60114 13582 60126 13634
rect 62178 13582 62190 13634
rect 62242 13582 62254 13634
rect 64978 13582 64990 13634
rect 65042 13631 65054 13634
rect 65042 13585 65263 13631
rect 65042 13582 65054 13585
rect 58942 13570 58994 13582
rect 63310 13570 63362 13582
rect 20414 13522 20466 13534
rect 34190 13522 34242 13534
rect 31266 13470 31278 13522
rect 31330 13519 31342 13522
rect 31602 13519 31614 13522
rect 31330 13473 31614 13519
rect 31330 13470 31342 13473
rect 31602 13470 31614 13473
rect 31666 13470 31678 13522
rect 20414 13458 20466 13470
rect 34190 13458 34242 13470
rect 34974 13522 35026 13534
rect 45502 13522 45554 13534
rect 48078 13522 48130 13534
rect 65217 13522 65263 13585
rect 67230 13570 67282 13582
rect 67678 13634 67730 13646
rect 67678 13570 67730 13582
rect 68126 13634 68178 13646
rect 68126 13570 68178 13582
rect 70366 13634 70418 13646
rect 70366 13570 70418 13582
rect 72942 13634 72994 13646
rect 72942 13570 72994 13582
rect 73950 13634 74002 13646
rect 73950 13570 74002 13582
rect 74398 13634 74450 13646
rect 74398 13570 74450 13582
rect 79326 13634 79378 13646
rect 79326 13570 79378 13582
rect 80782 13634 80834 13646
rect 80782 13570 80834 13582
rect 86494 13634 86546 13646
rect 86494 13570 86546 13582
rect 88062 13634 88114 13646
rect 92654 13634 92706 13646
rect 88834 13582 88846 13634
rect 88898 13582 88910 13634
rect 90514 13582 90526 13634
rect 90578 13582 90590 13634
rect 88062 13570 88114 13582
rect 92654 13570 92706 13582
rect 95230 13634 95282 13646
rect 105086 13634 105138 13646
rect 95890 13582 95902 13634
rect 95954 13582 95966 13634
rect 98018 13582 98030 13634
rect 98082 13582 98094 13634
rect 102050 13582 102062 13634
rect 102114 13582 102126 13634
rect 95230 13570 95282 13582
rect 105086 13570 105138 13582
rect 112030 13634 112082 13646
rect 112030 13570 112082 13582
rect 72382 13522 72434 13534
rect 94670 13522 94722 13534
rect 105646 13522 105698 13534
rect 35522 13470 35534 13522
rect 35586 13519 35598 13522
rect 36306 13519 36318 13522
rect 35586 13473 36318 13519
rect 35586 13470 35598 13473
rect 36306 13470 36318 13473
rect 36370 13470 36382 13522
rect 41794 13470 41806 13522
rect 41858 13519 41870 13522
rect 43138 13519 43150 13522
rect 41858 13473 43150 13519
rect 41858 13470 41870 13473
rect 43138 13470 43150 13473
rect 43202 13470 43214 13522
rect 43922 13470 43934 13522
rect 43986 13519 43998 13522
rect 44818 13519 44830 13522
rect 43986 13473 44830 13519
rect 43986 13470 43998 13473
rect 44818 13470 44830 13473
rect 44882 13470 44894 13522
rect 46050 13470 46062 13522
rect 46114 13519 46126 13522
rect 47058 13519 47070 13522
rect 46114 13473 47070 13519
rect 46114 13470 46126 13473
rect 47058 13470 47070 13473
rect 47122 13519 47134 13522
rect 47730 13519 47742 13522
rect 47122 13473 47742 13519
rect 47122 13470 47134 13473
rect 47730 13470 47742 13473
rect 47794 13470 47806 13522
rect 49298 13470 49310 13522
rect 49362 13519 49374 13522
rect 49746 13519 49758 13522
rect 49362 13473 49758 13519
rect 49362 13470 49374 13473
rect 49746 13470 49758 13473
rect 49810 13470 49822 13522
rect 63074 13470 63086 13522
rect 63138 13519 63150 13522
rect 63298 13519 63310 13522
rect 63138 13473 63310 13519
rect 63138 13470 63150 13473
rect 63298 13470 63310 13473
rect 63362 13470 63374 13522
rect 65202 13470 65214 13522
rect 65266 13470 65278 13522
rect 73378 13470 73390 13522
rect 73442 13519 73454 13522
rect 73826 13519 73838 13522
rect 73442 13473 73838 13519
rect 73442 13470 73454 13473
rect 73826 13470 73838 13473
rect 73890 13470 73902 13522
rect 89170 13470 89182 13522
rect 89234 13470 89246 13522
rect 92642 13470 92654 13522
rect 92706 13519 92718 13522
rect 93426 13519 93438 13522
rect 92706 13473 93438 13519
rect 92706 13470 92718 13473
rect 93426 13470 93438 13473
rect 93490 13470 93502 13522
rect 98802 13470 98814 13522
rect 98866 13470 98878 13522
rect 102610 13470 102622 13522
rect 102674 13519 102686 13522
rect 103170 13519 103182 13522
rect 102674 13473 103182 13519
rect 102674 13470 102686 13473
rect 103170 13470 103182 13473
rect 103234 13470 103246 13522
rect 34974 13458 35026 13470
rect 45502 13458 45554 13470
rect 48078 13458 48130 13470
rect 72382 13458 72434 13470
rect 94670 13458 94722 13470
rect 105646 13458 105698 13470
rect 106094 13522 106146 13534
rect 106094 13458 106146 13470
rect 111582 13522 111634 13534
rect 111582 13458 111634 13470
rect 1344 13354 158592 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 96638 13354
rect 96690 13302 96742 13354
rect 96794 13302 96846 13354
rect 96898 13302 127358 13354
rect 127410 13302 127462 13354
rect 127514 13302 127566 13354
rect 127618 13302 158078 13354
rect 158130 13302 158182 13354
rect 158234 13302 158286 13354
rect 158338 13302 158592 13354
rect 1344 13268 158592 13302
rect 20190 13186 20242 13198
rect 32510 13186 32562 13198
rect 61742 13186 61794 13198
rect 100158 13186 100210 13198
rect 27010 13134 27022 13186
rect 27074 13134 27086 13186
rect 31938 13134 31950 13186
rect 32002 13134 32014 13186
rect 39106 13134 39118 13186
rect 39170 13183 39182 13186
rect 39666 13183 39678 13186
rect 39170 13137 39678 13183
rect 39170 13134 39182 13137
rect 39666 13134 39678 13137
rect 39730 13134 39742 13186
rect 97346 13134 97358 13186
rect 97410 13134 97422 13186
rect 20190 13122 20242 13134
rect 32510 13122 32562 13134
rect 61742 13122 61794 13134
rect 100158 13122 100210 13134
rect 19854 13074 19906 13086
rect 19854 13010 19906 13022
rect 21870 13074 21922 13086
rect 26126 13074 26178 13086
rect 25442 13022 25454 13074
rect 25506 13022 25518 13074
rect 21870 13010 21922 13022
rect 26126 13010 26178 13022
rect 26574 13074 26626 13086
rect 38222 13074 38274 13086
rect 34290 13022 34302 13074
rect 34354 13022 34366 13074
rect 36418 13022 36430 13074
rect 36482 13022 36494 13074
rect 26574 13010 26626 13022
rect 38222 13010 38274 13022
rect 38782 13074 38834 13086
rect 38782 13010 38834 13022
rect 39678 13074 39730 13086
rect 39678 13010 39730 13022
rect 40686 13074 40738 13086
rect 50430 13074 50482 13086
rect 43922 13022 43934 13074
rect 43986 13022 43998 13074
rect 44818 13022 44830 13074
rect 44882 13022 44894 13074
rect 48850 13022 48862 13074
rect 48914 13022 48926 13074
rect 40686 13010 40738 13022
rect 50430 13010 50482 13022
rect 58718 13074 58770 13086
rect 58718 13010 58770 13022
rect 59502 13074 59554 13086
rect 59502 13010 59554 13022
rect 60622 13074 60674 13086
rect 60622 13010 60674 13022
rect 62302 13074 62354 13086
rect 62302 13010 62354 13022
rect 62750 13074 62802 13086
rect 62750 13010 62802 13022
rect 63422 13074 63474 13086
rect 68798 13074 68850 13086
rect 74174 13074 74226 13086
rect 66658 13022 66670 13074
rect 66722 13022 66734 13074
rect 72706 13022 72718 13074
rect 72770 13022 72782 13074
rect 63422 13010 63474 13022
rect 68798 13010 68850 13022
rect 74174 13010 74226 13022
rect 92318 13074 92370 13086
rect 92318 13010 92370 13022
rect 100718 13074 100770 13086
rect 108222 13074 108274 13086
rect 103506 13022 103518 13074
rect 103570 13022 103582 13074
rect 100718 13010 100770 13022
rect 108222 13010 108274 13022
rect 108670 13074 108722 13086
rect 108670 13010 108722 13022
rect 109118 13074 109170 13086
rect 109118 13010 109170 13022
rect 19742 12962 19794 12974
rect 19742 12898 19794 12910
rect 20078 12962 20130 12974
rect 29822 12962 29874 12974
rect 30830 12962 30882 12974
rect 20290 12910 20302 12962
rect 20354 12910 20366 12962
rect 22642 12910 22654 12962
rect 22706 12910 22718 12962
rect 26674 12910 26686 12962
rect 26738 12910 26750 12962
rect 27122 12910 27134 12962
rect 27186 12910 27198 12962
rect 29362 12910 29374 12962
rect 29426 12910 29438 12962
rect 30370 12910 30382 12962
rect 30434 12910 30446 12962
rect 20078 12898 20130 12910
rect 29822 12898 29874 12910
rect 30830 12898 30882 12910
rect 31390 12962 31442 12974
rect 38110 12962 38162 12974
rect 31602 12910 31614 12962
rect 31666 12910 31678 12962
rect 31938 12910 31950 12962
rect 32002 12910 32014 12962
rect 32498 12910 32510 12962
rect 32562 12910 32574 12962
rect 33618 12910 33630 12962
rect 33682 12910 33694 12962
rect 37202 12910 37214 12962
rect 37266 12910 37278 12962
rect 37762 12910 37774 12962
rect 37826 12910 37838 12962
rect 31390 12898 31442 12910
rect 38110 12898 38162 12910
rect 38334 12962 38386 12974
rect 48750 12962 48802 12974
rect 41010 12910 41022 12962
rect 41074 12910 41086 12962
rect 47730 12910 47742 12962
rect 47794 12910 47806 12962
rect 48290 12910 48302 12962
rect 48354 12910 48366 12962
rect 38334 12898 38386 12910
rect 48750 12898 48802 12910
rect 49758 12962 49810 12974
rect 53006 12962 53058 12974
rect 49970 12910 49982 12962
rect 50034 12910 50046 12962
rect 49758 12898 49810 12910
rect 53006 12898 53058 12910
rect 53790 12962 53842 12974
rect 58382 12962 58434 12974
rect 54338 12910 54350 12962
rect 54402 12910 54414 12962
rect 53790 12898 53842 12910
rect 58382 12898 58434 12910
rect 60510 12962 60562 12974
rect 60510 12898 60562 12910
rect 60846 12962 60898 12974
rect 60846 12898 60898 12910
rect 61070 12962 61122 12974
rect 88734 12962 88786 12974
rect 63858 12910 63870 12962
rect 63922 12910 63934 12962
rect 69906 12910 69918 12962
rect 69970 12910 69982 12962
rect 77186 12910 77198 12962
rect 77250 12910 77262 12962
rect 78530 12910 78542 12962
rect 78594 12910 78606 12962
rect 79874 12910 79886 12962
rect 79938 12910 79950 12962
rect 80210 12910 80222 12962
rect 80274 12910 80286 12962
rect 81554 12910 81566 12962
rect 81618 12910 81630 12962
rect 83122 12910 83134 12962
rect 83186 12910 83198 12962
rect 84802 12910 84814 12962
rect 84866 12910 84878 12962
rect 86034 12910 86046 12962
rect 86098 12910 86110 12962
rect 88274 12910 88286 12962
rect 88338 12910 88350 12962
rect 61070 12898 61122 12910
rect 88734 12898 88786 12910
rect 88958 12962 89010 12974
rect 92542 12962 92594 12974
rect 90514 12910 90526 12962
rect 90578 12910 90590 12962
rect 88958 12898 89010 12910
rect 92542 12898 92594 12910
rect 93998 12962 94050 12974
rect 95902 12962 95954 12974
rect 94546 12910 94558 12962
rect 94610 12910 94622 12962
rect 93998 12898 94050 12910
rect 95902 12898 95954 12910
rect 96238 12962 96290 12974
rect 100606 12962 100658 12974
rect 96338 12910 96350 12962
rect 96402 12910 96414 12962
rect 96238 12898 96290 12910
rect 100606 12898 100658 12910
rect 100830 12962 100882 12974
rect 107550 12962 107602 12974
rect 102386 12910 102398 12962
rect 102450 12910 102462 12962
rect 100830 12898 100882 12910
rect 107550 12898 107602 12910
rect 109566 12962 109618 12974
rect 109566 12898 109618 12910
rect 110014 12962 110066 12974
rect 110014 12898 110066 12910
rect 110686 12962 110738 12974
rect 110686 12898 110738 12910
rect 112142 12962 112194 12974
rect 112142 12898 112194 12910
rect 26462 12850 26514 12862
rect 19394 12798 19406 12850
rect 19458 12798 19470 12850
rect 23314 12798 23326 12850
rect 23378 12798 23390 12850
rect 26462 12786 26514 12798
rect 29934 12850 29986 12862
rect 29934 12786 29986 12798
rect 30942 12850 30994 12862
rect 30942 12786 30994 12798
rect 32846 12850 32898 12862
rect 49310 12850 49362 12862
rect 57710 12850 57762 12862
rect 36978 12798 36990 12850
rect 37042 12798 37054 12850
rect 41794 12798 41806 12850
rect 41858 12798 41870 12850
rect 46946 12798 46958 12850
rect 47010 12798 47022 12850
rect 55010 12798 55022 12850
rect 55074 12798 55086 12850
rect 32846 12786 32898 12798
rect 49310 12786 49362 12798
rect 57710 12786 57762 12798
rect 57934 12850 57986 12862
rect 57934 12786 57986 12798
rect 61630 12850 61682 12862
rect 76190 12850 76242 12862
rect 93102 12850 93154 12862
rect 64530 12798 64542 12850
rect 64594 12798 64606 12850
rect 70578 12798 70590 12850
rect 70642 12798 70654 12850
rect 74946 12798 74958 12850
rect 75010 12798 75022 12850
rect 78082 12798 78094 12850
rect 78146 12798 78158 12850
rect 82786 12798 82798 12850
rect 82850 12798 82862 12850
rect 84242 12798 84254 12850
rect 84306 12798 84318 12850
rect 87714 12798 87726 12850
rect 87778 12798 87790 12850
rect 90066 12798 90078 12850
rect 90130 12798 90142 12850
rect 91074 12798 91086 12850
rect 91138 12798 91150 12850
rect 61630 12786 61682 12798
rect 76190 12786 76242 12798
rect 93102 12786 93154 12798
rect 100158 12850 100210 12862
rect 100158 12786 100210 12798
rect 100270 12850 100322 12862
rect 100270 12786 100322 12798
rect 101054 12850 101106 12862
rect 101054 12786 101106 12798
rect 111694 12850 111746 12862
rect 111694 12786 111746 12798
rect 112702 12850 112754 12862
rect 112702 12786 112754 12798
rect 19070 12738 19122 12750
rect 19070 12674 19122 12686
rect 29598 12738 29650 12750
rect 29598 12674 29650 12686
rect 29710 12738 29762 12750
rect 29710 12674 29762 12686
rect 30606 12738 30658 12750
rect 30606 12674 30658 12686
rect 30718 12738 30770 12750
rect 39342 12738 39394 12750
rect 31826 12686 31838 12738
rect 31890 12686 31902 12738
rect 30718 12674 30770 12686
rect 39342 12674 39394 12686
rect 40350 12738 40402 12750
rect 40350 12674 40402 12686
rect 48526 12738 48578 12750
rect 48526 12674 48578 12686
rect 48862 12738 48914 12750
rect 48862 12674 48914 12686
rect 49534 12738 49586 12750
rect 49534 12674 49586 12686
rect 49646 12738 49698 12750
rect 49646 12674 49698 12686
rect 51102 12738 51154 12750
rect 51102 12674 51154 12686
rect 51662 12738 51714 12750
rect 51662 12674 51714 12686
rect 52222 12738 52274 12750
rect 52222 12674 52274 12686
rect 53454 12738 53506 12750
rect 53454 12674 53506 12686
rect 53678 12738 53730 12750
rect 53678 12674 53730 12686
rect 53902 12738 53954 12750
rect 58046 12738 58098 12750
rect 57250 12686 57262 12738
rect 57314 12686 57326 12738
rect 53902 12674 53954 12686
rect 58046 12674 58098 12686
rect 60062 12738 60114 12750
rect 60062 12674 60114 12686
rect 61742 12738 61794 12750
rect 61742 12674 61794 12686
rect 67566 12738 67618 12750
rect 67566 12674 67618 12686
rect 69134 12738 69186 12750
rect 69134 12674 69186 12686
rect 73278 12738 73330 12750
rect 73278 12674 73330 12686
rect 73726 12738 73778 12750
rect 73726 12674 73778 12686
rect 74622 12738 74674 12750
rect 74622 12674 74674 12686
rect 75294 12738 75346 12750
rect 75294 12674 75346 12686
rect 76302 12738 76354 12750
rect 89742 12738 89794 12750
rect 92766 12738 92818 12750
rect 83458 12686 83470 12738
rect 83522 12686 83534 12738
rect 87938 12686 87950 12738
rect 88002 12686 88014 12738
rect 89282 12686 89294 12738
rect 89346 12686 89358 12738
rect 90514 12686 90526 12738
rect 90578 12686 90590 12738
rect 91970 12686 91982 12738
rect 92034 12686 92046 12738
rect 76302 12674 76354 12686
rect 89742 12674 89794 12686
rect 92766 12674 92818 12686
rect 92990 12738 93042 12750
rect 92990 12674 93042 12686
rect 93550 12738 93602 12750
rect 93550 12674 93602 12686
rect 98366 12738 98418 12750
rect 98366 12674 98418 12686
rect 98814 12738 98866 12750
rect 98814 12674 98866 12686
rect 107662 12738 107714 12750
rect 107662 12674 107714 12686
rect 107886 12738 107938 12750
rect 107886 12674 107938 12686
rect 110798 12738 110850 12750
rect 110798 12674 110850 12686
rect 111246 12738 111298 12750
rect 111246 12674 111298 12686
rect 113038 12738 113090 12750
rect 113038 12674 113090 12686
rect 1344 12570 158592 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 81278 12570
rect 81330 12518 81382 12570
rect 81434 12518 81486 12570
rect 81538 12518 111998 12570
rect 112050 12518 112102 12570
rect 112154 12518 112206 12570
rect 112258 12518 142718 12570
rect 142770 12518 142822 12570
rect 142874 12518 142926 12570
rect 142978 12518 158592 12570
rect 1344 12484 158592 12518
rect 18174 12402 18226 12414
rect 18174 12338 18226 12350
rect 18622 12402 18674 12414
rect 18622 12338 18674 12350
rect 18958 12402 19010 12414
rect 18958 12338 19010 12350
rect 21198 12402 21250 12414
rect 21198 12338 21250 12350
rect 21982 12402 22034 12414
rect 21982 12338 22034 12350
rect 23998 12402 24050 12414
rect 23998 12338 24050 12350
rect 24110 12402 24162 12414
rect 24110 12338 24162 12350
rect 27246 12402 27298 12414
rect 27246 12338 27298 12350
rect 27358 12402 27410 12414
rect 27358 12338 27410 12350
rect 29486 12402 29538 12414
rect 37774 12402 37826 12414
rect 36642 12350 36654 12402
rect 36706 12350 36718 12402
rect 29486 12338 29538 12350
rect 37774 12338 37826 12350
rect 39902 12402 39954 12414
rect 39902 12338 39954 12350
rect 40798 12402 40850 12414
rect 45614 12402 45666 12414
rect 43810 12350 43822 12402
rect 43874 12350 43886 12402
rect 40798 12338 40850 12350
rect 45614 12338 45666 12350
rect 46398 12402 46450 12414
rect 46398 12338 46450 12350
rect 47182 12402 47234 12414
rect 47182 12338 47234 12350
rect 47518 12402 47570 12414
rect 47518 12338 47570 12350
rect 47966 12402 48018 12414
rect 54462 12402 54514 12414
rect 49634 12350 49646 12402
rect 49698 12350 49710 12402
rect 47966 12338 48018 12350
rect 19518 12290 19570 12302
rect 21310 12290 21362 12302
rect 19730 12238 19742 12290
rect 19794 12238 19806 12290
rect 19518 12226 19570 12238
rect 21310 12226 21362 12238
rect 21534 12290 21586 12302
rect 21534 12226 21586 12238
rect 22430 12290 22482 12302
rect 22430 12226 22482 12238
rect 25790 12290 25842 12302
rect 25790 12226 25842 12238
rect 26238 12290 26290 12302
rect 26238 12226 26290 12238
rect 29150 12290 29202 12302
rect 29150 12226 29202 12238
rect 29710 12290 29762 12302
rect 37326 12290 37378 12302
rect 31714 12238 31726 12290
rect 31778 12238 31790 12290
rect 32386 12238 32398 12290
rect 32450 12238 32462 12290
rect 29710 12226 29762 12238
rect 37326 12226 37378 12238
rect 37886 12290 37938 12302
rect 45950 12290 46002 12302
rect 42354 12238 42366 12290
rect 42418 12238 42430 12290
rect 42690 12238 42702 12290
rect 42754 12238 42766 12290
rect 48738 12238 48750 12290
rect 48802 12238 48814 12290
rect 37886 12226 37938 12238
rect 45950 12226 46002 12238
rect 19630 12178 19682 12190
rect 20974 12178 21026 12190
rect 20178 12126 20190 12178
rect 20242 12126 20254 12178
rect 19630 12114 19682 12126
rect 20974 12114 21026 12126
rect 21758 12178 21810 12190
rect 21758 12114 21810 12126
rect 22206 12178 22258 12190
rect 22206 12114 22258 12126
rect 22878 12178 22930 12190
rect 22878 12114 22930 12126
rect 23886 12178 23938 12190
rect 23886 12114 23938 12126
rect 24558 12178 24610 12190
rect 24558 12114 24610 12126
rect 25230 12178 25282 12190
rect 25230 12114 25282 12126
rect 25342 12178 25394 12190
rect 25342 12114 25394 12126
rect 25566 12178 25618 12190
rect 25566 12114 25618 12126
rect 29374 12178 29426 12190
rect 36990 12178 37042 12190
rect 30258 12126 30270 12178
rect 30322 12126 30334 12178
rect 31378 12126 31390 12178
rect 31442 12126 31454 12178
rect 32162 12126 32174 12178
rect 32226 12126 32238 12178
rect 35970 12126 35982 12178
rect 36034 12126 36046 12178
rect 29374 12114 29426 12126
rect 36990 12114 37042 12126
rect 37662 12178 37714 12190
rect 44270 12178 44322 12190
rect 40898 12126 40910 12178
rect 40962 12126 40974 12178
rect 41906 12126 41918 12178
rect 41970 12126 41982 12178
rect 42802 12126 42814 12178
rect 42866 12126 42878 12178
rect 43586 12126 43598 12178
rect 43650 12126 43662 12178
rect 44034 12126 44046 12178
rect 44098 12126 44110 12178
rect 37662 12114 37714 12126
rect 44270 12114 44322 12126
rect 44830 12178 44882 12190
rect 44830 12114 44882 12126
rect 45166 12178 45218 12190
rect 46174 12178 46226 12190
rect 49086 12178 49138 12190
rect 45602 12126 45614 12178
rect 45666 12126 45678 12178
rect 46610 12126 46622 12178
rect 46674 12126 46686 12178
rect 45166 12114 45218 12126
rect 46174 12114 46226 12126
rect 49086 12114 49138 12126
rect 49310 12178 49362 12190
rect 49310 12114 49362 12126
rect 19966 12066 20018 12078
rect 18946 12014 18958 12066
rect 19010 12014 19022 12066
rect 19966 12002 20018 12014
rect 28702 12066 28754 12078
rect 38782 12066 38834 12078
rect 32498 12014 32510 12066
rect 32562 12014 32574 12066
rect 34402 12014 34414 12066
rect 34466 12014 34478 12066
rect 28702 12002 28754 12014
rect 38782 12002 38834 12014
rect 39454 12066 39506 12078
rect 39454 12002 39506 12014
rect 40238 12066 40290 12078
rect 40238 12002 40290 12014
rect 46286 12066 46338 12078
rect 46286 12002 46338 12014
rect 19182 11954 19234 11966
rect 19182 11890 19234 11902
rect 27134 11954 27186 11966
rect 27134 11890 27186 11902
rect 40350 11954 40402 11966
rect 43698 11902 43710 11954
rect 43762 11902 43774 11954
rect 45378 11902 45390 11954
rect 45442 11902 45454 11954
rect 49649 11951 49695 12350
rect 54462 12338 54514 12350
rect 54910 12402 54962 12414
rect 54910 12338 54962 12350
rect 56030 12402 56082 12414
rect 60846 12402 60898 12414
rect 59826 12350 59838 12402
rect 59890 12350 59902 12402
rect 60498 12350 60510 12402
rect 60562 12350 60574 12402
rect 56030 12338 56082 12350
rect 60846 12338 60898 12350
rect 64878 12402 64930 12414
rect 64878 12338 64930 12350
rect 70366 12402 70418 12414
rect 70366 12338 70418 12350
rect 73726 12402 73778 12414
rect 85710 12402 85762 12414
rect 78418 12350 78430 12402
rect 78482 12350 78494 12402
rect 84914 12350 84926 12402
rect 84978 12350 84990 12402
rect 73726 12338 73778 12350
rect 85710 12338 85762 12350
rect 88062 12402 88114 12414
rect 104862 12402 104914 12414
rect 90290 12350 90302 12402
rect 90354 12350 90366 12402
rect 90962 12350 90974 12402
rect 91026 12350 91038 12402
rect 88062 12338 88114 12350
rect 104862 12338 104914 12350
rect 105982 12402 106034 12414
rect 105982 12338 106034 12350
rect 109342 12402 109394 12414
rect 109342 12338 109394 12350
rect 110350 12402 110402 12414
rect 110350 12338 110402 12350
rect 110798 12402 110850 12414
rect 110798 12338 110850 12350
rect 113822 12402 113874 12414
rect 113822 12338 113874 12350
rect 49758 12290 49810 12302
rect 49758 12226 49810 12238
rect 50206 12290 50258 12302
rect 50206 12226 50258 12238
rect 50542 12290 50594 12302
rect 50542 12226 50594 12238
rect 54686 12290 54738 12302
rect 54686 12226 54738 12238
rect 55246 12290 55298 12302
rect 61294 12290 61346 12302
rect 57586 12238 57598 12290
rect 57650 12238 57662 12290
rect 55246 12226 55298 12238
rect 61294 12226 61346 12238
rect 65102 12290 65154 12302
rect 79438 12290 79490 12302
rect 85822 12290 85874 12302
rect 75394 12238 75406 12290
rect 75458 12238 75470 12290
rect 77858 12238 77870 12290
rect 77922 12238 77934 12290
rect 83234 12238 83246 12290
rect 83298 12238 83310 12290
rect 84354 12238 84366 12290
rect 84418 12238 84430 12290
rect 65102 12226 65154 12238
rect 79438 12226 79490 12238
rect 85822 12226 85874 12238
rect 88510 12290 88562 12302
rect 90414 12290 90466 12302
rect 104078 12290 104130 12302
rect 106654 12290 106706 12302
rect 89394 12238 89406 12290
rect 89458 12238 89470 12290
rect 93986 12238 93998 12290
rect 94050 12238 94062 12290
rect 105634 12238 105646 12290
rect 105698 12238 105710 12290
rect 106306 12238 106318 12290
rect 106370 12238 106382 12290
rect 88510 12226 88562 12238
rect 90414 12226 90466 12238
rect 104078 12226 104130 12238
rect 106654 12226 106706 12238
rect 106990 12290 107042 12302
rect 106990 12226 107042 12238
rect 107438 12290 107490 12302
rect 107438 12226 107490 12238
rect 107998 12290 108050 12302
rect 107998 12226 108050 12238
rect 108558 12290 108610 12302
rect 108558 12226 108610 12238
rect 54910 12178 54962 12190
rect 64654 12178 64706 12190
rect 51090 12126 51102 12178
rect 51154 12126 51166 12178
rect 56914 12126 56926 12178
rect 56978 12126 56990 12178
rect 54910 12114 54962 12126
rect 64654 12114 64706 12126
rect 65214 12178 65266 12190
rect 69918 12178 69970 12190
rect 68898 12126 68910 12178
rect 68962 12126 68974 12178
rect 65214 12114 65266 12126
rect 69918 12114 69970 12126
rect 70254 12178 70306 12190
rect 70254 12114 70306 12126
rect 70478 12178 70530 12190
rect 79214 12178 79266 12190
rect 74498 12126 74510 12178
rect 74562 12126 74574 12178
rect 76290 12126 76302 12178
rect 76354 12126 76366 12178
rect 78194 12126 78206 12178
rect 78258 12126 78270 12178
rect 70478 12114 70530 12126
rect 79214 12114 79266 12126
rect 79550 12178 79602 12190
rect 91310 12178 91362 12190
rect 80098 12126 80110 12178
rect 80162 12126 80174 12178
rect 81442 12126 81454 12178
rect 81506 12126 81518 12178
rect 83010 12126 83022 12178
rect 83074 12126 83086 12178
rect 84690 12126 84702 12178
rect 84754 12126 84766 12178
rect 86146 12126 86158 12178
rect 86210 12126 86222 12178
rect 89170 12126 89182 12178
rect 89234 12126 89246 12178
rect 90626 12126 90638 12178
rect 90690 12126 90702 12178
rect 79550 12114 79602 12126
rect 91310 12114 91362 12126
rect 91534 12178 91586 12190
rect 102958 12178 103010 12190
rect 94770 12126 94782 12178
rect 94834 12126 94846 12178
rect 96114 12126 96126 12178
rect 96178 12126 96190 12178
rect 97794 12126 97806 12178
rect 97858 12126 97870 12178
rect 102610 12126 102622 12178
rect 102674 12126 102686 12178
rect 91534 12114 91586 12126
rect 102958 12114 103010 12126
rect 103966 12178 104018 12190
rect 103966 12114 104018 12126
rect 104302 12178 104354 12190
rect 105310 12178 105362 12190
rect 104626 12126 104638 12178
rect 104690 12126 104702 12178
rect 104302 12114 104354 12126
rect 105310 12114 105362 12126
rect 107326 12178 107378 12190
rect 107326 12114 107378 12126
rect 107662 12178 107714 12190
rect 107662 12114 107714 12126
rect 108110 12178 108162 12190
rect 108110 12114 108162 12126
rect 108446 12178 108498 12190
rect 108446 12114 108498 12126
rect 109454 12178 109506 12190
rect 109454 12114 109506 12126
rect 61742 12066 61794 12078
rect 51762 12014 51774 12066
rect 51826 12014 51838 12066
rect 53890 12014 53902 12066
rect 53954 12014 53966 12066
rect 61742 12002 61794 12014
rect 62638 12066 62690 12078
rect 62638 12002 62690 12014
rect 62974 12066 63026 12078
rect 62974 12002 63026 12014
rect 63422 12066 63474 12078
rect 63422 12002 63474 12014
rect 63870 12066 63922 12078
rect 69582 12066 69634 12078
rect 65986 12014 65998 12066
rect 66050 12014 66062 12066
rect 68114 12014 68126 12066
rect 68178 12014 68190 12066
rect 63870 12002 63922 12014
rect 69582 12002 69634 12014
rect 71262 12066 71314 12078
rect 71262 12002 71314 12014
rect 71710 12066 71762 12078
rect 71710 12002 71762 12014
rect 72382 12066 72434 12078
rect 72382 12002 72434 12014
rect 72830 12066 72882 12078
rect 72830 12002 72882 12014
rect 73390 12066 73442 12078
rect 73390 12002 73442 12014
rect 74286 12066 74338 12078
rect 95230 12066 95282 12078
rect 103070 12066 103122 12078
rect 87266 12014 87278 12066
rect 87330 12014 87342 12066
rect 91858 12014 91870 12066
rect 91922 12014 91934 12066
rect 95890 12014 95902 12066
rect 95954 12014 95966 12066
rect 98130 12014 98142 12066
rect 98194 12014 98206 12066
rect 99698 12014 99710 12066
rect 99762 12014 99774 12066
rect 101826 12014 101838 12066
rect 101890 12014 101902 12066
rect 74286 12002 74338 12014
rect 95230 12002 95282 12014
rect 103070 12002 103122 12014
rect 109902 12066 109954 12078
rect 109902 12002 109954 12014
rect 111582 12066 111634 12078
rect 111582 12002 111634 12014
rect 112030 12066 112082 12078
rect 112030 12002 112082 12014
rect 112478 12066 112530 12078
rect 112478 12002 112530 12014
rect 112926 12066 112978 12078
rect 112926 12002 112978 12014
rect 113374 12066 113426 12078
rect 113374 12002 113426 12014
rect 85710 11954 85762 11966
rect 107998 11954 108050 11966
rect 49746 11951 49758 11954
rect 49649 11905 49758 11951
rect 49746 11902 49758 11905
rect 49810 11902 49822 11954
rect 61170 11902 61182 11954
rect 61234 11951 61246 11954
rect 61730 11951 61742 11954
rect 61234 11905 61742 11951
rect 61234 11902 61246 11905
rect 61730 11902 61742 11905
rect 61794 11902 61806 11954
rect 64306 11902 64318 11954
rect 64370 11951 64382 11954
rect 64530 11951 64542 11954
rect 64370 11905 64542 11951
rect 64370 11902 64382 11905
rect 64530 11902 64542 11905
rect 64594 11902 64606 11954
rect 72370 11902 72382 11954
rect 72434 11951 72446 11954
rect 72930 11951 72942 11954
rect 72434 11905 72942 11951
rect 72434 11902 72446 11905
rect 72930 11902 72942 11905
rect 72994 11902 73006 11954
rect 98802 11902 98814 11954
rect 98866 11902 98878 11954
rect 40350 11890 40402 11902
rect 85710 11890 85762 11902
rect 107998 11890 108050 11902
rect 108558 11954 108610 11966
rect 108558 11890 108610 11902
rect 109342 11954 109394 11966
rect 111570 11902 111582 11954
rect 111634 11951 111646 11954
rect 112578 11951 112590 11954
rect 111634 11905 112590 11951
rect 111634 11902 111646 11905
rect 112578 11902 112590 11905
rect 112642 11951 112654 11954
rect 113362 11951 113374 11954
rect 112642 11905 113374 11951
rect 112642 11902 112654 11905
rect 113362 11902 113374 11905
rect 113426 11902 113438 11954
rect 109342 11890 109394 11902
rect 1344 11786 158592 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 96638 11786
rect 96690 11734 96742 11786
rect 96794 11734 96846 11786
rect 96898 11734 127358 11786
rect 127410 11734 127462 11786
rect 127514 11734 127566 11786
rect 127618 11734 158078 11786
rect 158130 11734 158182 11786
rect 158234 11734 158286 11786
rect 158338 11734 158592 11786
rect 1344 11700 158592 11734
rect 27582 11618 27634 11630
rect 20290 11566 20302 11618
rect 20354 11566 20366 11618
rect 27582 11554 27634 11566
rect 42926 11618 42978 11630
rect 60622 11618 60674 11630
rect 67006 11618 67058 11630
rect 93550 11618 93602 11630
rect 45938 11566 45950 11618
rect 46002 11615 46014 11618
rect 46386 11615 46398 11618
rect 46002 11569 46398 11615
rect 46002 11566 46014 11569
rect 46386 11566 46398 11569
rect 46450 11566 46462 11618
rect 62962 11566 62974 11618
rect 63026 11615 63038 11618
rect 63298 11615 63310 11618
rect 63026 11569 63310 11615
rect 63026 11566 63038 11569
rect 63298 11566 63310 11569
rect 63362 11566 63374 11618
rect 63522 11566 63534 11618
rect 63586 11615 63598 11618
rect 63970 11615 63982 11618
rect 63586 11569 63982 11615
rect 63586 11566 63598 11569
rect 63970 11566 63982 11569
rect 64034 11615 64046 11618
rect 64642 11615 64654 11618
rect 64034 11569 64654 11615
rect 64034 11566 64046 11569
rect 64642 11566 64654 11569
rect 64706 11566 64718 11618
rect 68898 11566 68910 11618
rect 68962 11615 68974 11618
rect 69122 11615 69134 11618
rect 68962 11569 69134 11615
rect 68962 11566 68974 11569
rect 69122 11566 69134 11569
rect 69186 11566 69198 11618
rect 73266 11566 73278 11618
rect 73330 11566 73342 11618
rect 112690 11566 112702 11618
rect 112754 11615 112766 11618
rect 113474 11615 113486 11618
rect 112754 11569 113486 11615
rect 112754 11566 112766 11569
rect 113474 11566 113486 11569
rect 113538 11615 113550 11618
rect 114370 11615 114382 11618
rect 113538 11569 114382 11615
rect 113538 11566 113550 11569
rect 114370 11566 114382 11569
rect 114434 11615 114446 11618
rect 114818 11615 114830 11618
rect 114434 11569 114830 11615
rect 114434 11566 114446 11569
rect 114818 11566 114830 11569
rect 114882 11566 114894 11618
rect 42926 11554 42978 11566
rect 60622 11554 60674 11566
rect 67006 11554 67058 11566
rect 22542 11506 22594 11518
rect 15586 11454 15598 11506
rect 15650 11454 15662 11506
rect 17714 11454 17726 11506
rect 17778 11454 17790 11506
rect 21298 11454 21310 11506
rect 21362 11454 21374 11506
rect 22542 11442 22594 11454
rect 28702 11506 28754 11518
rect 47854 11506 47906 11518
rect 33506 11454 33518 11506
rect 33570 11454 33582 11506
rect 41794 11454 41806 11506
rect 41858 11454 41870 11506
rect 28702 11442 28754 11454
rect 47854 11442 47906 11454
rect 50766 11506 50818 11518
rect 50766 11442 50818 11454
rect 51662 11506 51714 11518
rect 51662 11442 51714 11454
rect 52110 11506 52162 11518
rect 52110 11442 52162 11454
rect 52782 11506 52834 11518
rect 63534 11506 63586 11518
rect 58706 11454 58718 11506
rect 58770 11454 58782 11506
rect 52782 11442 52834 11454
rect 63534 11442 63586 11454
rect 64878 11506 64930 11518
rect 64878 11442 64930 11454
rect 71038 11506 71090 11518
rect 71038 11442 71090 11454
rect 19742 11394 19794 11406
rect 18498 11342 18510 11394
rect 18562 11342 18574 11394
rect 19742 11330 19794 11342
rect 20078 11394 20130 11406
rect 24782 11394 24834 11406
rect 48526 11394 48578 11406
rect 52670 11394 52722 11406
rect 20514 11342 20526 11394
rect 20578 11342 20590 11394
rect 34402 11342 34414 11394
rect 34466 11342 34478 11394
rect 41122 11342 41134 11394
rect 41186 11342 41198 11394
rect 42242 11342 42254 11394
rect 42306 11342 42318 11394
rect 42914 11342 42926 11394
rect 42978 11342 42990 11394
rect 50082 11342 50094 11394
rect 50146 11342 50158 11394
rect 20078 11330 20130 11342
rect 24782 11330 24834 11342
rect 48526 11330 48578 11342
rect 52670 11330 52722 11342
rect 53006 11394 53058 11406
rect 53006 11330 53058 11342
rect 53230 11394 53282 11406
rect 53230 11330 53282 11342
rect 53566 11394 53618 11406
rect 53566 11330 53618 11342
rect 53790 11394 53842 11406
rect 65438 11394 65490 11406
rect 54562 11342 54574 11394
rect 54626 11342 54638 11394
rect 61394 11342 61406 11394
rect 61458 11342 61470 11394
rect 53790 11330 53842 11342
rect 65438 11330 65490 11342
rect 65886 11394 65938 11406
rect 65886 11330 65938 11342
rect 66334 11394 66386 11406
rect 66334 11330 66386 11342
rect 66446 11394 66498 11406
rect 66446 11330 66498 11342
rect 70142 11394 70194 11406
rect 70142 11330 70194 11342
rect 71598 11394 71650 11406
rect 71598 11330 71650 11342
rect 73054 11394 73106 11406
rect 73281 11394 73327 11566
rect 93550 11554 93602 11566
rect 77086 11506 77138 11518
rect 99150 11506 99202 11518
rect 89058 11454 89070 11506
rect 89122 11454 89134 11506
rect 95218 11454 95230 11506
rect 95282 11454 95294 11506
rect 77086 11442 77138 11454
rect 99150 11442 99202 11454
rect 100606 11506 100658 11518
rect 112590 11506 112642 11518
rect 102946 11454 102958 11506
rect 103010 11454 103022 11506
rect 100606 11442 100658 11454
rect 112590 11442 112642 11454
rect 113486 11506 113538 11518
rect 113486 11442 113538 11454
rect 114382 11506 114434 11518
rect 114382 11442 114434 11454
rect 114830 11506 114882 11518
rect 114830 11442 114882 11454
rect 74398 11394 74450 11406
rect 73266 11342 73278 11394
rect 73330 11342 73342 11394
rect 73054 11330 73106 11342
rect 74398 11330 74450 11342
rect 74846 11394 74898 11406
rect 74846 11330 74898 11342
rect 74958 11394 75010 11406
rect 74958 11330 75010 11342
rect 76078 11394 76130 11406
rect 76974 11394 77026 11406
rect 76738 11342 76750 11394
rect 76802 11342 76814 11394
rect 76078 11330 76130 11342
rect 76974 11330 77026 11342
rect 77198 11394 77250 11406
rect 84142 11394 84194 11406
rect 91982 11394 92034 11406
rect 77410 11342 77422 11394
rect 77474 11342 77486 11394
rect 81890 11342 81902 11394
rect 81954 11342 81966 11394
rect 84802 11342 84814 11394
rect 84866 11342 84878 11394
rect 86258 11342 86270 11394
rect 86322 11342 86334 11394
rect 88498 11342 88510 11394
rect 88562 11342 88574 11394
rect 89170 11342 89182 11394
rect 89234 11342 89246 11394
rect 89842 11342 89854 11394
rect 89906 11342 89918 11394
rect 77198 11330 77250 11342
rect 84142 11330 84194 11342
rect 91982 11330 92034 11342
rect 92318 11394 92370 11406
rect 92318 11330 92370 11342
rect 92654 11394 92706 11406
rect 92654 11330 92706 11342
rect 94110 11394 94162 11406
rect 95566 11394 95618 11406
rect 94546 11342 94558 11394
rect 94610 11342 94622 11394
rect 94110 11330 94162 11342
rect 95566 11330 95618 11342
rect 96910 11394 96962 11406
rect 96910 11330 96962 11342
rect 100270 11394 100322 11406
rect 100270 11330 100322 11342
rect 100382 11394 100434 11406
rect 100382 11330 100434 11342
rect 101278 11394 101330 11406
rect 107774 11394 107826 11406
rect 111022 11394 111074 11406
rect 101278 11330 101330 11342
rect 102622 11338 102674 11350
rect 105858 11342 105870 11394
rect 105922 11342 105934 11394
rect 106418 11342 106430 11394
rect 106482 11342 106494 11394
rect 108546 11342 108558 11394
rect 108610 11342 108622 11394
rect 109218 11342 109230 11394
rect 109282 11342 109294 11394
rect 109890 11342 109902 11394
rect 109954 11342 109966 11394
rect 19406 11282 19458 11294
rect 19058 11230 19070 11282
rect 19122 11230 19134 11282
rect 19406 11218 19458 11230
rect 21422 11282 21474 11294
rect 21422 11218 21474 11230
rect 21646 11282 21698 11294
rect 21646 11218 21698 11230
rect 36318 11282 36370 11294
rect 36318 11218 36370 11230
rect 36430 11282 36482 11294
rect 39006 11282 39058 11294
rect 37314 11230 37326 11282
rect 37378 11230 37390 11282
rect 37650 11230 37662 11282
rect 37714 11230 37726 11282
rect 36430 11218 36482 11230
rect 39006 11218 39058 11230
rect 39118 11282 39170 11294
rect 39118 11218 39170 11230
rect 39342 11282 39394 11294
rect 39342 11218 39394 11230
rect 40686 11282 40738 11294
rect 42590 11282 42642 11294
rect 41234 11230 41246 11282
rect 41298 11230 41310 11282
rect 40686 11218 40738 11230
rect 42590 11218 42642 11230
rect 48190 11282 48242 11294
rect 54126 11282 54178 11294
rect 48738 11230 48750 11282
rect 48802 11230 48814 11282
rect 49522 11230 49534 11282
rect 49586 11230 49598 11282
rect 48190 11218 48242 11230
rect 54126 11218 54178 11230
rect 60510 11282 60562 11294
rect 60510 11218 60562 11230
rect 61630 11282 61682 11294
rect 61630 11218 61682 11230
rect 66894 11282 66946 11294
rect 66894 11218 66946 11230
rect 67006 11282 67058 11294
rect 67006 11218 67058 11230
rect 71934 11282 71986 11294
rect 71934 11218 71986 11230
rect 72718 11282 72770 11294
rect 72718 11218 72770 11230
rect 76302 11282 76354 11294
rect 76302 11218 76354 11230
rect 76414 11282 76466 11294
rect 84030 11282 84082 11294
rect 90974 11282 91026 11294
rect 78978 11230 78990 11282
rect 79042 11230 79054 11282
rect 84466 11230 84478 11282
rect 84530 11230 84542 11282
rect 86930 11230 86942 11282
rect 86994 11230 87006 11282
rect 87714 11230 87726 11282
rect 87778 11230 87790 11282
rect 89394 11230 89406 11282
rect 89458 11230 89470 11282
rect 76414 11218 76466 11230
rect 84030 11218 84082 11230
rect 90974 11218 91026 11230
rect 93102 11282 93154 11294
rect 93102 11218 93154 11230
rect 93662 11282 93714 11294
rect 93662 11218 93714 11230
rect 97246 11282 97298 11294
rect 97246 11218 97298 11230
rect 100718 11282 100770 11294
rect 100718 11218 100770 11230
rect 102510 11282 102562 11294
rect 107774 11330 107826 11342
rect 111022 11330 111074 11342
rect 112142 11394 112194 11406
rect 112142 11330 112194 11342
rect 102622 11274 102674 11286
rect 107550 11282 107602 11294
rect 105074 11230 105086 11282
rect 105138 11230 105150 11282
rect 106194 11230 106206 11282
rect 106258 11230 106270 11282
rect 102510 11218 102562 11230
rect 107550 11218 107602 11230
rect 108110 11282 108162 11294
rect 110686 11282 110738 11294
rect 108770 11230 108782 11282
rect 108834 11230 108846 11282
rect 108110 11218 108162 11230
rect 110686 11218 110738 11230
rect 111470 11282 111522 11294
rect 111470 11218 111522 11230
rect 22094 11170 22146 11182
rect 20178 11118 20190 11170
rect 20242 11118 20254 11170
rect 22094 11106 22146 11118
rect 24446 11170 24498 11182
rect 24446 11106 24498 11118
rect 25342 11170 25394 11182
rect 25342 11106 25394 11118
rect 26014 11170 26066 11182
rect 26014 11106 26066 11118
rect 27694 11170 27746 11182
rect 27694 11106 27746 11118
rect 27806 11170 27858 11182
rect 27806 11106 27858 11118
rect 29262 11170 29314 11182
rect 29262 11106 29314 11118
rect 29934 11170 29986 11182
rect 29934 11106 29986 11118
rect 30270 11170 30322 11182
rect 30270 11106 30322 11118
rect 36094 11170 36146 11182
rect 36094 11106 36146 11118
rect 36990 11170 37042 11182
rect 36990 11106 37042 11118
rect 37998 11170 38050 11182
rect 37998 11106 38050 11118
rect 38334 11170 38386 11182
rect 39790 11170 39842 11182
rect 40350 11170 40402 11182
rect 38658 11118 38670 11170
rect 38722 11118 38734 11170
rect 40114 11118 40126 11170
rect 40178 11118 40190 11170
rect 38334 11106 38386 11118
rect 39790 11106 39842 11118
rect 40350 11106 40402 11118
rect 40574 11170 40626 11182
rect 40574 11106 40626 11118
rect 43822 11170 43874 11182
rect 43822 11106 43874 11118
rect 44270 11170 44322 11182
rect 44270 11106 44322 11118
rect 45054 11170 45106 11182
rect 45054 11106 45106 11118
rect 45502 11170 45554 11182
rect 45502 11106 45554 11118
rect 45838 11170 45890 11182
rect 45838 11106 45890 11118
rect 46286 11170 46338 11182
rect 46286 11106 46338 11118
rect 46958 11170 47010 11182
rect 46958 11106 47010 11118
rect 47406 11170 47458 11182
rect 51214 11170 51266 11182
rect 49074 11118 49086 11170
rect 49138 11118 49150 11170
rect 50306 11118 50318 11170
rect 50370 11118 50382 11170
rect 47406 11106 47458 11118
rect 51214 11106 51266 11118
rect 53678 11170 53730 11182
rect 53678 11106 53730 11118
rect 61966 11170 62018 11182
rect 61966 11106 62018 11118
rect 62078 11170 62130 11182
rect 62078 11106 62130 11118
rect 62190 11170 62242 11182
rect 62190 11106 62242 11118
rect 62414 11170 62466 11182
rect 62414 11106 62466 11118
rect 62974 11170 63026 11182
rect 62974 11106 63026 11118
rect 63982 11170 64034 11182
rect 63982 11106 64034 11118
rect 64318 11170 64370 11182
rect 64318 11106 64370 11118
rect 65102 11170 65154 11182
rect 65102 11106 65154 11118
rect 66222 11170 66274 11182
rect 66222 11106 66274 11118
rect 67902 11170 67954 11182
rect 67902 11106 67954 11118
rect 68574 11170 68626 11182
rect 68574 11106 68626 11118
rect 69022 11170 69074 11182
rect 69022 11106 69074 11118
rect 69358 11170 69410 11182
rect 69358 11106 69410 11118
rect 69806 11170 69858 11182
rect 69806 11106 69858 11118
rect 70478 11170 70530 11182
rect 70478 11106 70530 11118
rect 71262 11170 71314 11182
rect 71262 11106 71314 11118
rect 71486 11170 71538 11182
rect 71486 11106 71538 11118
rect 72046 11170 72098 11182
rect 72046 11106 72098 11118
rect 72270 11170 72322 11182
rect 72270 11106 72322 11118
rect 72830 11170 72882 11182
rect 72830 11106 72882 11118
rect 73614 11170 73666 11182
rect 74622 11170 74674 11182
rect 73938 11118 73950 11170
rect 74002 11118 74014 11170
rect 73614 11106 73666 11118
rect 74622 11106 74674 11118
rect 75630 11170 75682 11182
rect 75630 11106 75682 11118
rect 90190 11170 90242 11182
rect 90190 11106 90242 11118
rect 90638 11170 90690 11182
rect 90638 11106 90690 11118
rect 90862 11170 90914 11182
rect 90862 11106 90914 11118
rect 92430 11170 92482 11182
rect 92430 11106 92482 11118
rect 92766 11170 92818 11182
rect 92766 11106 92818 11118
rect 92990 11170 93042 11182
rect 92990 11106 93042 11118
rect 93550 11170 93602 11182
rect 93550 11106 93602 11118
rect 96350 11170 96402 11182
rect 96350 11106 96402 11118
rect 96574 11170 96626 11182
rect 96574 11106 96626 11118
rect 96798 11170 96850 11182
rect 96798 11106 96850 11118
rect 97358 11170 97410 11182
rect 97358 11106 97410 11118
rect 97806 11170 97858 11182
rect 97806 11106 97858 11118
rect 98254 11170 98306 11182
rect 98254 11106 98306 11118
rect 98702 11170 98754 11182
rect 98702 11106 98754 11118
rect 99822 11170 99874 11182
rect 99822 11106 99874 11118
rect 100942 11170 100994 11182
rect 100942 11106 100994 11118
rect 101166 11170 101218 11182
rect 101950 11170 102002 11182
rect 101602 11118 101614 11170
rect 101666 11118 101678 11170
rect 101166 11106 101218 11118
rect 101950 11106 102002 11118
rect 102286 11170 102338 11182
rect 102286 11106 102338 11118
rect 106990 11170 107042 11182
rect 106990 11106 107042 11118
rect 107998 11170 108050 11182
rect 107998 11106 108050 11118
rect 109454 11170 109506 11182
rect 109454 11106 109506 11118
rect 110126 11170 110178 11182
rect 110126 11106 110178 11118
rect 110798 11170 110850 11182
rect 110798 11106 110850 11118
rect 111582 11170 111634 11182
rect 111582 11106 111634 11118
rect 111806 11170 111858 11182
rect 111806 11106 111858 11118
rect 113038 11170 113090 11182
rect 113038 11106 113090 11118
rect 114046 11170 114098 11182
rect 114046 11106 114098 11118
rect 1344 11002 158592 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 81278 11002
rect 81330 10950 81382 11002
rect 81434 10950 81486 11002
rect 81538 10950 111998 11002
rect 112050 10950 112102 11002
rect 112154 10950 112206 11002
rect 112258 10950 142718 11002
rect 142770 10950 142822 11002
rect 142874 10950 142926 11002
rect 142978 10950 158592 11002
rect 1344 10916 158592 10950
rect 21646 10834 21698 10846
rect 21646 10770 21698 10782
rect 22878 10834 22930 10846
rect 22878 10770 22930 10782
rect 23886 10834 23938 10846
rect 23886 10770 23938 10782
rect 28366 10834 28418 10846
rect 35198 10834 35250 10846
rect 31490 10782 31502 10834
rect 31554 10782 31566 10834
rect 33954 10782 33966 10834
rect 34018 10782 34030 10834
rect 28366 10770 28418 10782
rect 35198 10770 35250 10782
rect 35422 10834 35474 10846
rect 35422 10770 35474 10782
rect 35534 10834 35586 10846
rect 35534 10770 35586 10782
rect 37550 10834 37602 10846
rect 37550 10770 37602 10782
rect 41358 10834 41410 10846
rect 41358 10770 41410 10782
rect 42590 10834 42642 10846
rect 42590 10770 42642 10782
rect 43038 10834 43090 10846
rect 54126 10834 54178 10846
rect 54798 10834 54850 10846
rect 46834 10782 46846 10834
rect 46898 10782 46910 10834
rect 54450 10782 54462 10834
rect 54514 10782 54526 10834
rect 43038 10770 43090 10782
rect 54126 10770 54178 10782
rect 54798 10770 54850 10782
rect 55470 10834 55522 10846
rect 55470 10770 55522 10782
rect 55582 10834 55634 10846
rect 55582 10770 55634 10782
rect 56702 10834 56754 10846
rect 56702 10770 56754 10782
rect 56814 10834 56866 10846
rect 56814 10770 56866 10782
rect 56926 10834 56978 10846
rect 56926 10770 56978 10782
rect 58046 10834 58098 10846
rect 58046 10770 58098 10782
rect 58158 10834 58210 10846
rect 58158 10770 58210 10782
rect 59278 10834 59330 10846
rect 76974 10834 77026 10846
rect 59278 10770 59330 10782
rect 63422 10778 63474 10790
rect 66322 10782 66334 10834
rect 66386 10782 66398 10834
rect 20638 10722 20690 10734
rect 18162 10670 18174 10722
rect 18226 10670 18238 10722
rect 20638 10658 20690 10670
rect 20974 10722 21026 10734
rect 20974 10658 21026 10670
rect 24670 10722 24722 10734
rect 24670 10658 24722 10670
rect 25342 10722 25394 10734
rect 25342 10658 25394 10670
rect 26910 10722 26962 10734
rect 34974 10722 35026 10734
rect 31602 10670 31614 10722
rect 31666 10670 31678 10722
rect 32386 10670 32398 10722
rect 32450 10670 32462 10722
rect 33394 10670 33406 10722
rect 33458 10670 33470 10722
rect 26910 10658 26962 10670
rect 34974 10658 35026 10670
rect 38782 10722 38834 10734
rect 38782 10658 38834 10670
rect 38894 10722 38946 10734
rect 40350 10722 40402 10734
rect 42142 10722 42194 10734
rect 53790 10722 53842 10734
rect 39666 10670 39678 10722
rect 39730 10670 39742 10722
rect 41906 10670 41918 10722
rect 41970 10670 41982 10722
rect 46162 10670 46174 10722
rect 46226 10670 46238 10722
rect 38894 10658 38946 10670
rect 40350 10658 40402 10670
rect 42142 10658 42194 10670
rect 53790 10658 53842 10670
rect 57598 10722 57650 10734
rect 57598 10658 57650 10670
rect 58718 10722 58770 10734
rect 58718 10658 58770 10670
rect 58830 10722 58882 10734
rect 76974 10770 77026 10782
rect 77198 10834 77250 10846
rect 77198 10770 77250 10782
rect 77310 10834 77362 10846
rect 77310 10770 77362 10782
rect 77870 10834 77922 10846
rect 78766 10834 78818 10846
rect 83918 10834 83970 10846
rect 78194 10782 78206 10834
rect 78258 10782 78270 10834
rect 80434 10782 80446 10834
rect 80498 10782 80510 10834
rect 77870 10770 77922 10782
rect 78766 10770 78818 10782
rect 83918 10770 83970 10782
rect 85038 10834 85090 10846
rect 85038 10770 85090 10782
rect 85822 10834 85874 10846
rect 85822 10770 85874 10782
rect 86382 10834 86434 10846
rect 93662 10834 93714 10846
rect 88274 10782 88286 10834
rect 88338 10782 88350 10834
rect 86382 10770 86434 10782
rect 93662 10770 93714 10782
rect 95678 10834 95730 10846
rect 109790 10834 109842 10846
rect 102834 10782 102846 10834
rect 102898 10782 102910 10834
rect 95678 10770 95730 10782
rect 109790 10770 109842 10782
rect 110910 10834 110962 10846
rect 110910 10770 110962 10782
rect 63422 10714 63474 10726
rect 64878 10722 64930 10734
rect 58830 10658 58882 10670
rect 64878 10658 64930 10670
rect 64990 10722 65042 10734
rect 79214 10722 79266 10734
rect 67218 10670 67230 10722
rect 67282 10670 67294 10722
rect 74386 10670 74398 10722
rect 74450 10670 74462 10722
rect 64990 10658 65042 10670
rect 79214 10658 79266 10670
rect 84478 10722 84530 10734
rect 84478 10658 84530 10670
rect 84590 10722 84642 10734
rect 92654 10722 92706 10734
rect 102174 10722 102226 10734
rect 91298 10670 91310 10722
rect 91362 10670 91374 10722
rect 95778 10670 95790 10722
rect 95842 10670 95854 10722
rect 99810 10670 99822 10722
rect 99874 10670 99886 10722
rect 101490 10670 101502 10722
rect 101554 10670 101566 10722
rect 84590 10658 84642 10670
rect 92654 10658 92706 10670
rect 102174 10658 102226 10670
rect 109454 10722 109506 10734
rect 109454 10658 109506 10670
rect 109678 10722 109730 10734
rect 109678 10658 109730 10670
rect 110014 10722 110066 10734
rect 110014 10658 110066 10670
rect 22094 10610 22146 10622
rect 17490 10558 17502 10610
rect 17554 10558 17566 10610
rect 21410 10558 21422 10610
rect 21474 10558 21486 10610
rect 22094 10546 22146 10558
rect 23550 10610 23602 10622
rect 26574 10610 26626 10622
rect 24098 10558 24110 10610
rect 24162 10558 24174 10610
rect 24434 10558 24446 10610
rect 24498 10558 24510 10610
rect 23550 10546 23602 10558
rect 26574 10546 26626 10558
rect 27246 10610 27298 10622
rect 28030 10610 28082 10622
rect 35982 10610 36034 10622
rect 27570 10558 27582 10610
rect 27634 10558 27646 10610
rect 30370 10558 30382 10610
rect 30434 10558 30446 10610
rect 31378 10558 31390 10610
rect 31442 10558 31454 10610
rect 32050 10558 32062 10610
rect 32114 10558 32126 10610
rect 33058 10558 33070 10610
rect 33122 10558 33134 10610
rect 34178 10558 34190 10610
rect 34242 10558 34254 10610
rect 27246 10546 27298 10558
rect 28030 10546 28082 10558
rect 35982 10546 36034 10558
rect 36542 10610 36594 10622
rect 36542 10546 36594 10558
rect 39118 10610 39170 10622
rect 44270 10610 44322 10622
rect 39442 10558 39454 10610
rect 39506 10558 39518 10610
rect 40002 10558 40014 10610
rect 40066 10558 40078 10610
rect 41346 10558 41358 10610
rect 41410 10558 41422 10610
rect 39118 10546 39170 10558
rect 44270 10546 44322 10558
rect 44606 10610 44658 10622
rect 47630 10610 47682 10622
rect 44818 10558 44830 10610
rect 44882 10558 44894 10610
rect 46050 10558 46062 10610
rect 46114 10558 46126 10610
rect 46722 10558 46734 10610
rect 46786 10558 46798 10610
rect 44606 10546 44658 10558
rect 47630 10546 47682 10558
rect 48190 10610 48242 10622
rect 49198 10610 49250 10622
rect 48962 10558 48974 10610
rect 49026 10558 49038 10610
rect 48190 10546 48242 10558
rect 49198 10546 49250 10558
rect 49982 10610 50034 10622
rect 55694 10610 55746 10622
rect 50194 10558 50206 10610
rect 50258 10558 50270 10610
rect 49982 10546 50034 10558
rect 55694 10546 55746 10558
rect 56142 10610 56194 10622
rect 57822 10610 57874 10622
rect 57250 10558 57262 10610
rect 57314 10558 57326 10610
rect 56142 10546 56194 10558
rect 57822 10546 57874 10558
rect 59390 10610 59442 10622
rect 63310 10610 63362 10622
rect 60050 10558 60062 10610
rect 60114 10558 60126 10610
rect 59390 10546 59442 10558
rect 63310 10546 63362 10558
rect 64654 10610 64706 10622
rect 72494 10610 72546 10622
rect 65426 10558 65438 10610
rect 65490 10558 65502 10610
rect 66546 10558 66558 10610
rect 66610 10558 66622 10610
rect 67554 10558 67566 10610
rect 67618 10558 67630 10610
rect 68898 10558 68910 10610
rect 68962 10558 68974 10610
rect 64654 10546 64706 10558
rect 72494 10546 72546 10558
rect 72718 10610 72770 10622
rect 77086 10610 77138 10622
rect 79102 10610 79154 10622
rect 73714 10558 73726 10610
rect 73778 10558 73790 10610
rect 77522 10558 77534 10610
rect 77586 10558 77598 10610
rect 72718 10546 72770 10558
rect 77086 10546 77138 10558
rect 79102 10546 79154 10558
rect 79662 10610 79714 10622
rect 79662 10546 79714 10558
rect 80110 10610 80162 10622
rect 83806 10610 83858 10622
rect 82898 10558 82910 10610
rect 82962 10558 82974 10610
rect 80110 10546 80162 10558
rect 83806 10546 83858 10558
rect 85486 10610 85538 10622
rect 85486 10546 85538 10558
rect 85710 10610 85762 10622
rect 85710 10546 85762 10558
rect 86046 10610 86098 10622
rect 89518 10610 89570 10622
rect 92430 10610 92482 10622
rect 86930 10558 86942 10610
rect 86994 10558 87006 10610
rect 88722 10558 88734 10610
rect 88786 10558 88798 10610
rect 90066 10558 90078 10610
rect 90130 10558 90142 10610
rect 92194 10558 92206 10610
rect 92258 10558 92270 10610
rect 86046 10546 86098 10558
rect 89518 10546 89570 10558
rect 92430 10546 92482 10558
rect 92766 10610 92818 10622
rect 95342 10610 95394 10622
rect 100382 10610 100434 10622
rect 94322 10558 94334 10610
rect 94386 10558 94398 10610
rect 94546 10558 94558 10610
rect 94610 10558 94622 10610
rect 96114 10558 96126 10610
rect 96178 10558 96190 10610
rect 97458 10558 97470 10610
rect 97522 10558 97534 10610
rect 99250 10558 99262 10610
rect 99314 10558 99326 10610
rect 92766 10546 92818 10558
rect 95342 10546 95394 10558
rect 100382 10546 100434 10558
rect 100606 10610 100658 10622
rect 100606 10546 100658 10558
rect 100942 10610 100994 10622
rect 100942 10546 100994 10558
rect 101166 10610 101218 10622
rect 101166 10546 101218 10558
rect 101838 10610 101890 10622
rect 111582 10610 111634 10622
rect 102610 10558 102622 10610
rect 102674 10558 102686 10610
rect 103618 10558 103630 10610
rect 103682 10558 103694 10610
rect 112690 10558 112702 10610
rect 112754 10558 112766 10610
rect 101838 10546 101890 10558
rect 111582 10546 111634 10558
rect 26126 10498 26178 10510
rect 20290 10446 20302 10498
rect 20354 10446 20366 10498
rect 26126 10434 26178 10446
rect 27022 10498 27074 10510
rect 27022 10434 27074 10446
rect 29150 10498 29202 10510
rect 29150 10434 29202 10446
rect 29598 10498 29650 10510
rect 29598 10434 29650 10446
rect 30046 10498 30098 10510
rect 30046 10434 30098 10446
rect 34638 10498 34690 10510
rect 34638 10434 34690 10446
rect 35310 10498 35362 10510
rect 35310 10434 35362 10446
rect 36990 10498 37042 10510
rect 36990 10434 37042 10446
rect 38446 10498 38498 10510
rect 38446 10434 38498 10446
rect 40238 10498 40290 10510
rect 40238 10434 40290 10446
rect 41134 10498 41186 10510
rect 41134 10434 41186 10446
rect 43486 10498 43538 10510
rect 43486 10434 43538 10446
rect 43822 10498 43874 10510
rect 43822 10434 43874 10446
rect 44382 10498 44434 10510
rect 44382 10434 44434 10446
rect 45614 10498 45666 10510
rect 45614 10434 45666 10446
rect 48862 10498 48914 10510
rect 48862 10434 48914 10446
rect 51550 10498 51602 10510
rect 51550 10434 51602 10446
rect 51886 10498 51938 10510
rect 51886 10434 51938 10446
rect 52334 10498 52386 10510
rect 52334 10434 52386 10446
rect 52894 10498 52946 10510
rect 52894 10434 52946 10446
rect 53342 10498 53394 10510
rect 53342 10434 53394 10446
rect 57934 10498 57986 10510
rect 65886 10498 65938 10510
rect 68574 10498 68626 10510
rect 73278 10498 73330 10510
rect 79438 10498 79490 10510
rect 84926 10498 84978 10510
rect 93102 10498 93154 10510
rect 100718 10498 100770 10510
rect 110350 10498 110402 10510
rect 60834 10446 60846 10498
rect 60898 10446 60910 10498
rect 62962 10446 62974 10498
rect 63026 10446 63038 10498
rect 66994 10446 67006 10498
rect 67058 10446 67070 10498
rect 69570 10446 69582 10498
rect 69634 10446 69646 10498
rect 71698 10446 71710 10498
rect 71762 10446 71774 10498
rect 76514 10446 76526 10498
rect 76578 10446 76590 10498
rect 81890 10446 81902 10498
rect 81954 10446 81966 10498
rect 87266 10446 87278 10498
rect 87330 10446 87342 10498
rect 94210 10446 94222 10498
rect 94274 10446 94286 10498
rect 105970 10446 105982 10498
rect 106034 10446 106046 10498
rect 57934 10434 57986 10446
rect 65886 10434 65938 10446
rect 68574 10434 68626 10446
rect 73278 10434 73330 10446
rect 79438 10434 79490 10446
rect 84926 10434 84978 10446
rect 93102 10434 93154 10446
rect 100718 10434 100770 10446
rect 110350 10434 110402 10446
rect 112142 10498 112194 10510
rect 115950 10498 116002 10510
rect 113362 10446 113374 10498
rect 113426 10446 113438 10498
rect 115490 10446 115502 10498
rect 115554 10446 115566 10498
rect 112142 10434 112194 10446
rect 115950 10434 116002 10446
rect 116398 10498 116450 10510
rect 116398 10434 116450 10446
rect 24222 10386 24274 10398
rect 24222 10322 24274 10334
rect 25230 10386 25282 10398
rect 25230 10322 25282 10334
rect 25566 10386 25618 10398
rect 38222 10386 38274 10398
rect 43934 10386 43986 10398
rect 58718 10386 58770 10398
rect 27458 10334 27470 10386
rect 27522 10334 27534 10386
rect 29250 10334 29262 10386
rect 29314 10383 29326 10386
rect 29810 10383 29822 10386
rect 29314 10337 29822 10383
rect 29314 10334 29326 10337
rect 29810 10334 29822 10337
rect 29874 10334 29886 10386
rect 37874 10334 37886 10386
rect 37938 10334 37950 10386
rect 41570 10334 41582 10386
rect 41634 10334 41646 10386
rect 42354 10334 42366 10386
rect 42418 10383 42430 10386
rect 43138 10383 43150 10386
rect 42418 10337 43150 10383
rect 42418 10334 42430 10337
rect 43138 10334 43150 10337
rect 43202 10334 43214 10386
rect 44818 10334 44830 10386
rect 44882 10334 44894 10386
rect 50642 10334 50654 10386
rect 50706 10334 50718 10386
rect 25566 10322 25618 10334
rect 38222 10322 38274 10334
rect 43934 10322 43986 10334
rect 58718 10322 58770 10334
rect 59278 10386 59330 10398
rect 59278 10322 59330 10334
rect 63422 10386 63474 10398
rect 63422 10322 63474 10334
rect 83918 10386 83970 10398
rect 83918 10322 83970 10334
rect 84478 10386 84530 10398
rect 84478 10322 84530 10334
rect 1344 10218 158592 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 96638 10218
rect 96690 10166 96742 10218
rect 96794 10166 96846 10218
rect 96898 10166 127358 10218
rect 127410 10166 127462 10218
rect 127514 10166 127566 10218
rect 127618 10166 158078 10218
rect 158130 10166 158182 10218
rect 158234 10166 158286 10218
rect 158338 10166 158592 10218
rect 1344 10132 158592 10166
rect 45054 10050 45106 10062
rect 19394 9998 19406 10050
rect 19458 10047 19470 10050
rect 19618 10047 19630 10050
rect 19458 10001 19630 10047
rect 19458 9998 19470 10001
rect 19618 9998 19630 10001
rect 19682 9998 19694 10050
rect 45054 9986 45106 9998
rect 45950 10050 46002 10062
rect 45950 9986 46002 9998
rect 59838 10050 59890 10062
rect 59838 9986 59890 9998
rect 64094 10050 64146 10062
rect 66098 9998 66110 10050
rect 66162 10047 66174 10050
rect 67890 10047 67902 10050
rect 66162 10001 67902 10047
rect 66162 9998 66174 10001
rect 67890 9998 67902 10001
rect 67954 9998 67966 10050
rect 116050 9998 116062 10050
rect 116114 10047 116126 10050
rect 117058 10047 117070 10050
rect 116114 10001 117070 10047
rect 116114 9998 116126 10001
rect 117058 9998 117070 10001
rect 117122 9998 117134 10050
rect 64094 9986 64146 9998
rect 18846 9938 18898 9950
rect 18846 9874 18898 9886
rect 19630 9938 19682 9950
rect 19630 9874 19682 9886
rect 20302 9938 20354 9950
rect 20302 9874 20354 9886
rect 21534 9938 21586 9950
rect 30494 9938 30546 9950
rect 40798 9938 40850 9950
rect 43150 9938 43202 9950
rect 22978 9886 22990 9938
rect 23042 9886 23054 9938
rect 25106 9886 25118 9938
rect 25170 9886 25182 9938
rect 26226 9886 26238 9938
rect 26290 9886 26302 9938
rect 31154 9886 31166 9938
rect 31218 9886 31230 9938
rect 42578 9886 42590 9938
rect 42642 9886 42654 9938
rect 21534 9874 21586 9886
rect 30494 9874 30546 9886
rect 40798 9874 40850 9886
rect 43150 9874 43202 9886
rect 45166 9938 45218 9950
rect 45166 9874 45218 9886
rect 47742 9938 47794 9950
rect 47742 9874 47794 9886
rect 50206 9938 50258 9950
rect 56702 9938 56754 9950
rect 59054 9938 59106 9950
rect 53554 9886 53566 9938
rect 53618 9886 53630 9938
rect 55682 9886 55694 9938
rect 55746 9886 55758 9938
rect 58258 9886 58270 9938
rect 58322 9886 58334 9938
rect 50206 9874 50258 9886
rect 56702 9874 56754 9886
rect 59054 9874 59106 9886
rect 60846 9938 60898 9950
rect 60846 9874 60898 9886
rect 66110 9938 66162 9950
rect 66110 9874 66162 9886
rect 67790 9938 67842 9950
rect 67790 9874 67842 9886
rect 70254 9938 70306 9950
rect 70254 9874 70306 9886
rect 75182 9938 75234 9950
rect 81902 9938 81954 9950
rect 78530 9886 78542 9938
rect 78594 9886 78606 9938
rect 80658 9886 80670 9938
rect 80722 9886 80734 9938
rect 75182 9874 75234 9886
rect 81902 9874 81954 9886
rect 85486 9938 85538 9950
rect 97582 9938 97634 9950
rect 104862 9938 104914 9950
rect 116062 9938 116114 9950
rect 94210 9886 94222 9938
rect 94274 9886 94286 9938
rect 99698 9886 99710 9938
rect 99762 9886 99774 9938
rect 101826 9886 101838 9938
rect 101890 9886 101902 9938
rect 109218 9886 109230 9938
rect 109282 9886 109294 9938
rect 85486 9874 85538 9886
rect 97582 9874 97634 9886
rect 104862 9874 104914 9886
rect 116062 9874 116114 9886
rect 30270 9826 30322 9838
rect 37326 9826 37378 9838
rect 22306 9774 22318 9826
rect 22370 9774 22382 9826
rect 25442 9774 25454 9826
rect 25506 9774 25518 9826
rect 29922 9774 29934 9826
rect 29986 9774 29998 9826
rect 30818 9774 30830 9826
rect 30882 9774 30894 9826
rect 31826 9774 31838 9826
rect 31890 9774 31902 9826
rect 32386 9774 32398 9826
rect 32450 9774 32462 9826
rect 33506 9774 33518 9826
rect 33570 9774 33582 9826
rect 34066 9774 34078 9826
rect 34130 9774 34142 9826
rect 35522 9774 35534 9826
rect 35586 9774 35598 9826
rect 36306 9774 36318 9826
rect 36370 9774 36382 9826
rect 30270 9762 30322 9774
rect 37326 9762 37378 9774
rect 37662 9826 37714 9838
rect 46734 9826 46786 9838
rect 38098 9774 38110 9826
rect 38162 9774 38174 9826
rect 43586 9774 43598 9826
rect 43650 9774 43662 9826
rect 45378 9774 45390 9826
rect 45442 9774 45454 9826
rect 37662 9762 37714 9774
rect 46734 9762 46786 9774
rect 48526 9826 48578 9838
rect 48526 9762 48578 9774
rect 48638 9826 48690 9838
rect 50542 9826 50594 9838
rect 56814 9826 56866 9838
rect 49186 9774 49198 9826
rect 49250 9774 49262 9826
rect 49746 9774 49758 9826
rect 49810 9774 49822 9826
rect 52770 9774 52782 9826
rect 52834 9774 52846 9826
rect 48638 9762 48690 9774
rect 50542 9762 50594 9774
rect 56814 9762 56866 9774
rect 57038 9826 57090 9838
rect 57038 9762 57090 9774
rect 57934 9826 57986 9838
rect 57934 9762 57986 9774
rect 58158 9826 58210 9838
rect 58158 9762 58210 9774
rect 59950 9826 60002 9838
rect 59950 9762 60002 9774
rect 61294 9826 61346 9838
rect 61294 9762 61346 9774
rect 62526 9826 62578 9838
rect 62526 9762 62578 9774
rect 63422 9826 63474 9838
rect 63422 9762 63474 9774
rect 63758 9826 63810 9838
rect 63758 9762 63810 9774
rect 67454 9826 67506 9838
rect 67454 9762 67506 9774
rect 70590 9826 70642 9838
rect 70590 9762 70642 9774
rect 72942 9826 72994 9838
rect 72942 9762 72994 9774
rect 73390 9826 73442 9838
rect 73390 9762 73442 9774
rect 73726 9826 73778 9838
rect 75294 9826 75346 9838
rect 74834 9774 74846 9826
rect 74898 9774 74910 9826
rect 73726 9762 73778 9774
rect 75294 9762 75346 9774
rect 75406 9826 75458 9838
rect 75406 9762 75458 9774
rect 76190 9826 76242 9838
rect 83246 9826 83298 9838
rect 81442 9774 81454 9826
rect 81506 9774 81518 9826
rect 82338 9774 82350 9826
rect 82402 9774 82414 9826
rect 76190 9762 76242 9774
rect 83246 9762 83298 9774
rect 83582 9826 83634 9838
rect 83582 9762 83634 9774
rect 84590 9826 84642 9838
rect 84590 9762 84642 9774
rect 86158 9826 86210 9838
rect 86158 9762 86210 9774
rect 86830 9826 86882 9838
rect 91870 9826 91922 9838
rect 87826 9774 87838 9826
rect 87890 9774 87902 9826
rect 89618 9774 89630 9826
rect 89682 9774 89694 9826
rect 91186 9774 91198 9826
rect 91250 9774 91262 9826
rect 86830 9762 86882 9774
rect 91870 9762 91922 9774
rect 92206 9826 92258 9838
rect 92206 9762 92258 9774
rect 92542 9826 92594 9838
rect 92542 9762 92594 9774
rect 92654 9826 92706 9838
rect 104526 9826 104578 9838
rect 93762 9774 93774 9826
rect 93826 9774 93838 9826
rect 93986 9774 93998 9826
rect 94050 9774 94062 9826
rect 95218 9774 95230 9826
rect 95282 9774 95294 9826
rect 96674 9774 96686 9826
rect 96738 9774 96750 9826
rect 99138 9774 99150 9826
rect 99202 9774 99214 9826
rect 102610 9774 102622 9826
rect 102674 9774 102686 9826
rect 103058 9774 103070 9826
rect 103122 9774 103134 9826
rect 103730 9774 103742 9826
rect 103794 9774 103806 9826
rect 92654 9762 92706 9774
rect 104526 9762 104578 9774
rect 104638 9826 104690 9838
rect 104638 9762 104690 9774
rect 105870 9826 105922 9838
rect 105870 9762 105922 9774
rect 106766 9826 106818 9838
rect 106766 9762 106818 9774
rect 107102 9826 107154 9838
rect 107998 9826 108050 9838
rect 113150 9826 113202 9838
rect 107650 9774 107662 9826
rect 107714 9774 107726 9826
rect 108210 9774 108222 9826
rect 108274 9774 108286 9826
rect 112130 9774 112142 9826
rect 112194 9774 112206 9826
rect 107102 9762 107154 9774
rect 107998 9762 108050 9774
rect 113150 9762 113202 9774
rect 113710 9826 113762 9838
rect 113710 9762 113762 9774
rect 114158 9826 114210 9838
rect 114158 9762 114210 9774
rect 114494 9826 114546 9838
rect 114494 9762 114546 9774
rect 115614 9826 115666 9838
rect 115614 9762 115666 9774
rect 29262 9714 29314 9726
rect 44046 9714 44098 9726
rect 31266 9662 31278 9714
rect 31330 9662 31342 9714
rect 32722 9662 32734 9714
rect 32786 9662 32798 9714
rect 33282 9662 33294 9714
rect 33346 9662 33358 9714
rect 35298 9662 35310 9714
rect 35362 9662 35374 9714
rect 38658 9662 38670 9714
rect 38722 9662 38734 9714
rect 41682 9662 41694 9714
rect 41746 9662 41758 9714
rect 29262 9650 29314 9662
rect 44046 9650 44098 9662
rect 44158 9714 44210 9726
rect 44158 9650 44210 9662
rect 45838 9714 45890 9726
rect 45838 9650 45890 9662
rect 45950 9714 46002 9726
rect 45950 9650 46002 9662
rect 46622 9714 46674 9726
rect 46622 9650 46674 9662
rect 48750 9714 48802 9726
rect 48750 9650 48802 9662
rect 51662 9714 51714 9726
rect 51662 9650 51714 9662
rect 56030 9714 56082 9726
rect 56030 9650 56082 9662
rect 56366 9714 56418 9726
rect 56366 9650 56418 9662
rect 56590 9714 56642 9726
rect 56590 9650 56642 9662
rect 57710 9714 57762 9726
rect 59838 9714 59890 9726
rect 59378 9662 59390 9714
rect 59442 9662 59454 9714
rect 57710 9650 57762 9662
rect 59838 9650 59890 9662
rect 60734 9714 60786 9726
rect 60734 9650 60786 9662
rect 61070 9714 61122 9726
rect 61070 9650 61122 9662
rect 61966 9714 62018 9726
rect 61966 9650 62018 9662
rect 62638 9714 62690 9726
rect 62638 9650 62690 9662
rect 63534 9714 63586 9726
rect 63534 9650 63586 9662
rect 64206 9714 64258 9726
rect 64206 9650 64258 9662
rect 65214 9714 65266 9726
rect 65214 9650 65266 9662
rect 69358 9714 69410 9726
rect 69358 9650 69410 9662
rect 69470 9714 69522 9726
rect 69470 9650 69522 9662
rect 70142 9714 70194 9726
rect 70142 9650 70194 9662
rect 70478 9714 70530 9726
rect 70478 9650 70530 9662
rect 70926 9714 70978 9726
rect 70926 9650 70978 9662
rect 71150 9714 71202 9726
rect 71150 9650 71202 9662
rect 71262 9714 71314 9726
rect 71262 9650 71314 9662
rect 72046 9714 72098 9726
rect 72046 9650 72098 9662
rect 72606 9714 72658 9726
rect 72606 9650 72658 9662
rect 73166 9714 73218 9726
rect 73166 9650 73218 9662
rect 73278 9714 73330 9726
rect 73278 9650 73330 9662
rect 74174 9714 74226 9726
rect 74174 9650 74226 9662
rect 82910 9714 82962 9726
rect 82910 9650 82962 9662
rect 85038 9714 85090 9726
rect 85038 9650 85090 9662
rect 85934 9714 85986 9726
rect 85934 9650 85986 9662
rect 86606 9714 86658 9726
rect 92990 9714 93042 9726
rect 103966 9714 104018 9726
rect 87938 9662 87950 9714
rect 88002 9662 88014 9714
rect 88946 9662 88958 9714
rect 89010 9662 89022 9714
rect 90402 9662 90414 9714
rect 90466 9662 90478 9714
rect 95778 9662 95790 9714
rect 95842 9662 95854 9714
rect 99026 9662 99038 9714
rect 99090 9662 99102 9714
rect 103282 9662 103294 9714
rect 103346 9662 103358 9714
rect 86606 9650 86658 9662
rect 92990 9650 93042 9662
rect 103966 9650 104018 9662
rect 104974 9714 105026 9726
rect 104974 9650 105026 9662
rect 106430 9714 106482 9726
rect 112478 9714 112530 9726
rect 111346 9662 111358 9714
rect 111410 9662 111422 9714
rect 106430 9650 106482 9662
rect 112478 9650 112530 9662
rect 112702 9714 112754 9726
rect 112702 9650 112754 9662
rect 113374 9714 113426 9726
rect 113374 9650 113426 9662
rect 113934 9714 113986 9726
rect 113934 9650 113986 9662
rect 114382 9714 114434 9726
rect 114382 9650 114434 9662
rect 20750 9602 20802 9614
rect 20750 9538 20802 9550
rect 21982 9602 22034 9614
rect 29374 9602 29426 9614
rect 44382 9602 44434 9614
rect 28466 9550 28478 9602
rect 28530 9550 28542 9602
rect 33394 9550 33406 9602
rect 33458 9550 33470 9602
rect 36194 9550 36206 9602
rect 36258 9550 36270 9602
rect 36978 9550 36990 9602
rect 37042 9550 37054 9602
rect 21982 9538 22034 9550
rect 29374 9538 29426 9550
rect 44382 9538 44434 9550
rect 46398 9602 46450 9614
rect 46398 9538 46450 9550
rect 47182 9602 47234 9614
rect 47182 9538 47234 9550
rect 48190 9602 48242 9614
rect 52222 9602 52274 9614
rect 50866 9550 50878 9602
rect 50930 9550 50942 9602
rect 48190 9538 48242 9550
rect 52222 9538 52274 9550
rect 56142 9602 56194 9614
rect 56142 9538 56194 9550
rect 58270 9602 58322 9614
rect 62862 9602 62914 9614
rect 61618 9550 61630 9602
rect 61682 9550 61694 9602
rect 58270 9538 58322 9550
rect 62862 9538 62914 9550
rect 64094 9602 64146 9614
rect 64094 9538 64146 9550
rect 64878 9602 64930 9614
rect 64878 9538 64930 9550
rect 65326 9602 65378 9614
rect 65326 9538 65378 9550
rect 65550 9602 65602 9614
rect 65550 9538 65602 9550
rect 66446 9602 66498 9614
rect 66446 9538 66498 9550
rect 67006 9602 67058 9614
rect 67006 9538 67058 9550
rect 68462 9602 68514 9614
rect 68462 9538 68514 9550
rect 69022 9602 69074 9614
rect 69022 9538 69074 9550
rect 69134 9602 69186 9614
rect 69134 9538 69186 9550
rect 71710 9602 71762 9614
rect 71710 9538 71762 9550
rect 72158 9602 72210 9614
rect 72158 9538 72210 9550
rect 72382 9602 72434 9614
rect 72382 9538 72434 9550
rect 72718 9602 72770 9614
rect 72718 9538 72770 9550
rect 74510 9602 74562 9614
rect 74510 9538 74562 9550
rect 75070 9602 75122 9614
rect 75070 9538 75122 9550
rect 76750 9602 76802 9614
rect 77422 9602 77474 9614
rect 77074 9550 77086 9602
rect 77138 9550 77150 9602
rect 76750 9538 76802 9550
rect 77422 9538 77474 9550
rect 77870 9602 77922 9614
rect 83358 9602 83410 9614
rect 78194 9550 78206 9602
rect 78258 9550 78270 9602
rect 82562 9550 82574 9602
rect 82626 9550 82638 9602
rect 77870 9538 77922 9550
rect 83358 9538 83410 9550
rect 84478 9602 84530 9614
rect 84478 9538 84530 9550
rect 84702 9602 84754 9614
rect 84702 9538 84754 9550
rect 84814 9602 84866 9614
rect 84814 9538 84866 9550
rect 86494 9602 86546 9614
rect 86494 9538 86546 9550
rect 92318 9602 92370 9614
rect 92318 9538 92370 9550
rect 92878 9602 92930 9614
rect 105310 9602 105362 9614
rect 93762 9550 93774 9602
rect 93826 9550 93838 9602
rect 92878 9538 92930 9550
rect 105310 9538 105362 9550
rect 106766 9602 106818 9614
rect 106766 9538 106818 9550
rect 108894 9602 108946 9614
rect 108894 9538 108946 9550
rect 112926 9602 112978 9614
rect 112926 9538 112978 9550
rect 113710 9602 113762 9614
rect 113710 9538 113762 9550
rect 115278 9602 115330 9614
rect 115278 9538 115330 9550
rect 115502 9602 115554 9614
rect 115502 9538 115554 9550
rect 116510 9602 116562 9614
rect 116510 9538 116562 9550
rect 116958 9602 117010 9614
rect 116958 9538 117010 9550
rect 1344 9434 158592 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 81278 9434
rect 81330 9382 81382 9434
rect 81434 9382 81486 9434
rect 81538 9382 111998 9434
rect 112050 9382 112102 9434
rect 112154 9382 112206 9434
rect 112258 9382 142718 9434
rect 142770 9382 142822 9434
rect 142874 9382 142926 9434
rect 142978 9382 158592 9434
rect 1344 9348 158592 9382
rect 20974 9266 21026 9278
rect 20974 9202 21026 9214
rect 22878 9266 22930 9278
rect 39678 9266 39730 9278
rect 26786 9214 26798 9266
rect 26850 9214 26862 9266
rect 27458 9214 27470 9266
rect 27522 9214 27534 9266
rect 22878 9202 22930 9214
rect 39678 9202 39730 9214
rect 40798 9266 40850 9278
rect 40798 9202 40850 9214
rect 48302 9266 48354 9278
rect 48302 9202 48354 9214
rect 48974 9266 49026 9278
rect 48974 9202 49026 9214
rect 49310 9266 49362 9278
rect 49310 9202 49362 9214
rect 49758 9266 49810 9278
rect 49758 9202 49810 9214
rect 50318 9266 50370 9278
rect 50318 9202 50370 9214
rect 51998 9266 52050 9278
rect 51998 9202 52050 9214
rect 52558 9266 52610 9278
rect 61182 9266 61234 9278
rect 63086 9266 63138 9278
rect 60386 9214 60398 9266
rect 60450 9214 60462 9266
rect 60834 9214 60846 9266
rect 60898 9214 60910 9266
rect 62402 9214 62414 9266
rect 62466 9214 62478 9266
rect 52558 9202 52610 9214
rect 61182 9202 61234 9214
rect 63086 9202 63138 9214
rect 65886 9266 65938 9278
rect 65886 9202 65938 9214
rect 66110 9266 66162 9278
rect 66110 9202 66162 9214
rect 66670 9266 66722 9278
rect 72494 9266 72546 9278
rect 71698 9214 71710 9266
rect 71762 9214 71774 9266
rect 66670 9202 66722 9214
rect 72494 9202 72546 9214
rect 73390 9266 73442 9278
rect 73390 9202 73442 9214
rect 75854 9266 75906 9278
rect 75854 9202 75906 9214
rect 80446 9266 80498 9278
rect 80446 9202 80498 9214
rect 81230 9266 81282 9278
rect 86158 9266 86210 9278
rect 81230 9202 81282 9214
rect 85822 9210 85874 9222
rect 21422 9154 21474 9166
rect 21422 9090 21474 9102
rect 21758 9154 21810 9166
rect 21758 9090 21810 9102
rect 22430 9154 22482 9166
rect 28366 9154 28418 9166
rect 40910 9154 40962 9166
rect 47518 9154 47570 9166
rect 23986 9102 23998 9154
rect 24050 9102 24062 9154
rect 32162 9102 32174 9154
rect 32226 9102 32238 9154
rect 35634 9102 35646 9154
rect 35698 9102 35710 9154
rect 38658 9102 38670 9154
rect 38722 9102 38734 9154
rect 41906 9102 41918 9154
rect 41970 9102 41982 9154
rect 44482 9102 44494 9154
rect 44546 9102 44558 9154
rect 22430 9090 22482 9102
rect 28366 9090 28418 9102
rect 40910 9090 40962 9102
rect 47518 9090 47570 9102
rect 47630 9154 47682 9166
rect 52894 9154 52946 9166
rect 55358 9154 55410 9166
rect 51314 9102 51326 9154
rect 51378 9102 51390 9154
rect 54338 9102 54350 9154
rect 54402 9102 54414 9154
rect 47630 9090 47682 9102
rect 21870 9042 21922 9054
rect 21870 8978 21922 8990
rect 27134 9042 27186 9054
rect 27134 8978 27186 8990
rect 27806 9042 27858 9054
rect 29486 9042 29538 9054
rect 28914 8990 28926 9042
rect 28978 8990 28990 9042
rect 27806 8978 27858 8990
rect 29486 8978 29538 8990
rect 30046 9042 30098 9054
rect 30046 8978 30098 8990
rect 30382 9042 30434 9054
rect 32510 9042 32562 9054
rect 39790 9042 39842 9054
rect 31490 8990 31502 9042
rect 31554 8990 31566 9042
rect 34402 8990 34414 9042
rect 34466 8990 34478 9042
rect 30382 8978 30434 8990
rect 32510 8978 32562 8990
rect 39790 8978 39842 8990
rect 40014 9042 40066 9054
rect 47294 9042 47346 9054
rect 41122 8990 41134 9042
rect 41186 8990 41198 9042
rect 41346 8990 41358 9042
rect 41410 8990 41422 9042
rect 43810 8990 43822 9042
rect 43874 8990 43886 9042
rect 40014 8978 40066 8990
rect 47294 8978 47346 8990
rect 51214 9042 51266 9054
rect 51214 8978 51266 8990
rect 20414 8930 20466 8942
rect 20414 8866 20466 8878
rect 21534 8930 21586 8942
rect 21534 8866 21586 8878
rect 23438 8930 23490 8942
rect 23438 8866 23490 8878
rect 23662 8930 23714 8942
rect 23662 8866 23714 8878
rect 24670 8930 24722 8942
rect 24670 8866 24722 8878
rect 25566 8930 25618 8942
rect 25566 8866 25618 8878
rect 26126 8930 26178 8942
rect 26126 8866 26178 8878
rect 26574 8930 26626 8942
rect 39230 8930 39282 8942
rect 47182 8930 47234 8942
rect 30818 8878 30830 8930
rect 30882 8878 30894 8930
rect 31826 8878 31838 8930
rect 31890 8878 31902 8930
rect 43026 8878 43038 8930
rect 43090 8878 43102 8930
rect 46610 8878 46622 8930
rect 46674 8878 46686 8930
rect 26574 8866 26626 8878
rect 39230 8866 39282 8878
rect 47182 8866 47234 8878
rect 50654 8930 50706 8942
rect 50654 8866 50706 8878
rect 28142 8818 28194 8830
rect 22306 8766 22318 8818
rect 22370 8815 22382 8818
rect 23314 8815 23326 8818
rect 22370 8769 23326 8815
rect 22370 8766 22382 8769
rect 23314 8766 23326 8769
rect 23378 8766 23390 8818
rect 25554 8766 25566 8818
rect 25618 8815 25630 8818
rect 26450 8815 26462 8818
rect 25618 8769 26462 8815
rect 25618 8766 25630 8769
rect 26450 8766 26462 8769
rect 26514 8766 26526 8818
rect 28142 8754 28194 8766
rect 28478 8818 28530 8830
rect 28478 8754 28530 8766
rect 29038 8818 29090 8830
rect 29038 8754 29090 8766
rect 39006 8818 39058 8830
rect 39006 8754 39058 8766
rect 39678 8818 39730 8830
rect 50978 8766 50990 8818
rect 51042 8815 51054 8818
rect 51329 8815 51375 9102
rect 52894 9090 52946 9102
rect 55358 9090 55410 9102
rect 55806 9154 55858 9166
rect 55806 9090 55858 9102
rect 55918 9154 55970 9166
rect 55918 9090 55970 9102
rect 56926 9154 56978 9166
rect 61742 9154 61794 9166
rect 58258 9102 58270 9154
rect 58322 9102 58334 9154
rect 59154 9102 59166 9154
rect 59218 9102 59230 9154
rect 56926 9090 56978 9102
rect 61742 9090 61794 9102
rect 62078 9154 62130 9166
rect 62078 9090 62130 9102
rect 66446 9154 66498 9166
rect 66446 9090 66498 9102
rect 67342 9154 67394 9166
rect 73726 9154 73778 9166
rect 80110 9154 80162 9166
rect 86158 9202 86210 9214
rect 94446 9266 94498 9278
rect 94446 9202 94498 9214
rect 105534 9266 105586 9278
rect 105534 9202 105586 9214
rect 114830 9266 114882 9278
rect 114830 9202 114882 9214
rect 115390 9266 115442 9278
rect 115390 9202 115442 9214
rect 115950 9266 116002 9278
rect 115950 9202 116002 9214
rect 117182 9266 117234 9278
rect 117182 9202 117234 9214
rect 67890 9102 67902 9154
rect 67954 9102 67966 9154
rect 70578 9102 70590 9154
rect 70642 9102 70654 9154
rect 75394 9102 75406 9154
rect 75458 9102 75470 9154
rect 76178 9102 76190 9154
rect 76242 9102 76254 9154
rect 83346 9102 83358 9154
rect 83410 9102 83422 9154
rect 85822 9146 85874 9158
rect 85934 9154 85986 9166
rect 67342 9090 67394 9102
rect 73726 9090 73778 9102
rect 80110 9090 80162 9102
rect 85934 9090 85986 9102
rect 86494 9154 86546 9166
rect 86494 9090 86546 9102
rect 87278 9154 87330 9166
rect 87278 9090 87330 9102
rect 87390 9154 87442 9166
rect 102286 9154 102338 9166
rect 88722 9102 88734 9154
rect 88786 9102 88798 9154
rect 93314 9102 93326 9154
rect 93378 9102 93390 9154
rect 96338 9102 96350 9154
rect 96402 9102 96414 9154
rect 98130 9102 98142 9154
rect 98194 9102 98206 9154
rect 100370 9102 100382 9154
rect 100434 9102 100446 9154
rect 87390 9090 87442 9102
rect 102286 9090 102338 9102
rect 102846 9154 102898 9166
rect 102846 9090 102898 9102
rect 105422 9154 105474 9166
rect 105422 9090 105474 9102
rect 105758 9154 105810 9166
rect 113150 9154 113202 9166
rect 108322 9102 108334 9154
rect 108386 9102 108398 9154
rect 105758 9090 105810 9102
rect 113150 9090 113202 9102
rect 114158 9154 114210 9166
rect 114158 9090 114210 9102
rect 115614 9154 115666 9166
rect 115614 9090 115666 9102
rect 115726 9154 115778 9166
rect 115726 9090 115778 9102
rect 116174 9154 116226 9166
rect 116174 9090 116226 9102
rect 52782 9042 52834 9054
rect 52782 8978 52834 8990
rect 53118 9042 53170 9054
rect 53118 8978 53170 8990
rect 55246 9042 55298 9054
rect 55246 8978 55298 8990
rect 55582 9042 55634 9054
rect 55582 8978 55634 8990
rect 56142 9042 56194 9054
rect 56142 8978 56194 8990
rect 56590 9042 56642 9054
rect 62750 9042 62802 9054
rect 59042 8990 59054 9042
rect 59106 8990 59118 9042
rect 60386 8990 60398 9042
rect 60450 8990 60462 9042
rect 56590 8978 56642 8990
rect 62750 8978 62802 8990
rect 63422 9042 63474 9054
rect 63422 8978 63474 8990
rect 64318 9042 64370 9054
rect 64318 8978 64370 8990
rect 64654 9042 64706 9054
rect 64654 8978 64706 8990
rect 64990 9042 65042 9054
rect 64990 8978 65042 8990
rect 65774 9042 65826 9054
rect 65774 8978 65826 8990
rect 66334 9042 66386 9054
rect 66334 8978 66386 8990
rect 67230 9042 67282 9054
rect 67230 8978 67282 8990
rect 71374 9042 71426 9054
rect 73054 9042 73106 9054
rect 72706 8990 72718 9042
rect 72770 8990 72782 9042
rect 71374 8978 71426 8990
rect 73054 8978 73106 8990
rect 73390 9042 73442 9054
rect 80334 9042 80386 9054
rect 77522 8990 77534 9042
rect 77586 8990 77598 9042
rect 78418 8990 78430 9042
rect 78482 8990 78494 9042
rect 78754 8990 78766 9042
rect 78818 8990 78830 9042
rect 73390 8978 73442 8990
rect 80334 8978 80386 8990
rect 80782 9042 80834 9054
rect 86270 9042 86322 9054
rect 81890 8990 81902 9042
rect 81954 8990 81966 9042
rect 82674 8990 82686 9042
rect 82738 8990 82750 9042
rect 80782 8978 80834 8990
rect 86270 8978 86322 8990
rect 86606 9042 86658 9054
rect 102510 9042 102562 9054
rect 105198 9042 105250 9054
rect 112926 9042 112978 9054
rect 87938 8990 87950 9042
rect 88002 8990 88014 9042
rect 94098 8990 94110 9042
rect 94162 8990 94174 9042
rect 96562 8990 96574 9042
rect 96626 8990 96638 9042
rect 97906 8990 97918 9042
rect 97970 8990 97982 9042
rect 99698 8990 99710 9042
rect 99762 8990 99774 9042
rect 101042 8990 101054 9042
rect 101106 8990 101118 9042
rect 101266 8990 101278 9042
rect 101330 8990 101342 9042
rect 103618 8990 103630 9042
rect 103682 8990 103694 9042
rect 108994 8990 109006 9042
rect 109058 8990 109070 9042
rect 109666 8990 109678 9042
rect 109730 8990 109742 9042
rect 111570 8990 111582 9042
rect 111634 8990 111646 9042
rect 86606 8978 86658 8990
rect 102510 8978 102562 8990
rect 105198 8978 105250 8990
rect 112926 8978 112978 8990
rect 113262 9042 113314 9054
rect 113262 8978 113314 8990
rect 113486 9042 113538 9054
rect 113486 8978 113538 8990
rect 113934 9042 113986 9054
rect 113934 8978 113986 8990
rect 114606 9042 114658 9054
rect 114606 8978 114658 8990
rect 115166 9042 115218 9054
rect 115166 8978 115218 8990
rect 116286 9042 116338 9054
rect 116286 8978 116338 8990
rect 51550 8930 51602 8942
rect 63982 8930 64034 8942
rect 53554 8878 53566 8930
rect 53618 8878 53630 8930
rect 57474 8878 57486 8930
rect 57538 8878 57550 8930
rect 59266 8878 59278 8930
rect 59330 8878 59342 8930
rect 51550 8866 51602 8878
rect 63982 8866 64034 8878
rect 64542 8930 64594 8942
rect 64542 8866 64594 8878
rect 65438 8930 65490 8942
rect 81454 8930 81506 8942
rect 95790 8930 95842 8942
rect 102398 8930 102450 8942
rect 114382 8930 114434 8942
rect 69234 8878 69246 8930
rect 69298 8878 69310 8930
rect 69570 8878 69582 8930
rect 69634 8878 69646 8930
rect 74050 8878 74062 8930
rect 74114 8878 74126 8930
rect 76626 8878 76638 8930
rect 76690 8878 76702 8930
rect 78306 8878 78318 8930
rect 78370 8878 78382 8930
rect 85474 8878 85486 8930
rect 85538 8878 85550 8930
rect 90850 8878 90862 8930
rect 90914 8878 90926 8930
rect 91186 8878 91198 8930
rect 91250 8878 91262 8930
rect 94882 8878 94894 8930
rect 94946 8878 94958 8930
rect 101602 8878 101614 8930
rect 101666 8878 101678 8930
rect 104514 8878 104526 8930
rect 104578 8878 104590 8930
rect 106194 8878 106206 8930
rect 106258 8878 106270 8930
rect 110562 8878 110574 8930
rect 110626 8878 110638 8930
rect 112130 8878 112142 8930
rect 112194 8878 112206 8930
rect 65438 8866 65490 8878
rect 81454 8866 81506 8878
rect 95790 8866 95842 8878
rect 102398 8866 102450 8878
rect 114382 8866 114434 8878
rect 116734 8930 116786 8942
rect 116734 8866 116786 8878
rect 117630 8930 117682 8942
rect 117630 8866 117682 8878
rect 118078 8930 118130 8942
rect 118078 8866 118130 8878
rect 118638 8930 118690 8942
rect 118638 8866 118690 8878
rect 67342 8818 67394 8830
rect 87278 8818 87330 8830
rect 51042 8769 51375 8815
rect 51042 8766 51054 8769
rect 52210 8766 52222 8818
rect 52274 8815 52286 8818
rect 52546 8815 52558 8818
rect 52274 8769 52558 8815
rect 52274 8766 52286 8769
rect 52546 8766 52558 8769
rect 52610 8766 52622 8818
rect 78642 8766 78654 8818
rect 78706 8766 78718 8818
rect 39678 8754 39730 8766
rect 67342 8754 67394 8766
rect 87278 8754 87330 8766
rect 95902 8818 95954 8830
rect 100818 8766 100830 8818
rect 100882 8766 100894 8818
rect 95902 8754 95954 8766
rect 1344 8650 158592 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 96638 8650
rect 96690 8598 96742 8650
rect 96794 8598 96846 8650
rect 96898 8598 127358 8650
rect 127410 8598 127462 8650
rect 127514 8598 127566 8650
rect 127618 8598 158078 8650
rect 158130 8598 158182 8650
rect 158234 8598 158286 8650
rect 158338 8598 158592 8650
rect 1344 8564 158592 8598
rect 29934 8482 29986 8494
rect 29934 8418 29986 8430
rect 94110 8482 94162 8494
rect 117618 8430 117630 8482
rect 117682 8479 117694 8482
rect 118178 8479 118190 8482
rect 117682 8433 118190 8479
rect 117682 8430 117694 8433
rect 118178 8430 118190 8433
rect 118242 8430 118254 8482
rect 94110 8418 94162 8430
rect 23438 8370 23490 8382
rect 20178 8318 20190 8370
rect 20242 8318 20254 8370
rect 23438 8306 23490 8318
rect 27134 8370 27186 8382
rect 27134 8306 27186 8318
rect 28142 8370 28194 8382
rect 28142 8306 28194 8318
rect 29486 8370 29538 8382
rect 29486 8306 29538 8318
rect 32958 8370 33010 8382
rect 37102 8370 37154 8382
rect 34850 8318 34862 8370
rect 34914 8318 34926 8370
rect 32958 8306 33010 8318
rect 37102 8306 37154 8318
rect 37662 8370 37714 8382
rect 37662 8306 37714 8318
rect 37774 8370 37826 8382
rect 48862 8370 48914 8382
rect 57710 8370 57762 8382
rect 38546 8318 38558 8370
rect 38610 8318 38622 8370
rect 40674 8318 40686 8370
rect 40738 8318 40750 8370
rect 41906 8318 41918 8370
rect 41970 8318 41982 8370
rect 47506 8318 47518 8370
rect 47570 8318 47582 8370
rect 50866 8318 50878 8370
rect 50930 8318 50942 8370
rect 55010 8318 55022 8370
rect 55074 8318 55086 8370
rect 57138 8318 57150 8370
rect 57202 8318 57214 8370
rect 37774 8306 37826 8318
rect 48862 8306 48914 8318
rect 57710 8306 57762 8318
rect 60622 8370 60674 8382
rect 71710 8370 71762 8382
rect 90750 8370 90802 8382
rect 62850 8318 62862 8370
rect 62914 8318 62926 8370
rect 63970 8318 63982 8370
rect 64034 8318 64046 8370
rect 66098 8318 66110 8370
rect 66162 8318 66174 8370
rect 66546 8367 66558 8370
rect 66337 8321 66558 8367
rect 60622 8306 60674 8318
rect 20750 8258 20802 8270
rect 17378 8206 17390 8258
rect 17442 8206 17454 8258
rect 20750 8194 20802 8206
rect 21870 8258 21922 8270
rect 21870 8194 21922 8206
rect 22094 8258 22146 8270
rect 22094 8194 22146 8206
rect 22542 8258 22594 8270
rect 22542 8194 22594 8206
rect 23886 8258 23938 8270
rect 23886 8194 23938 8206
rect 25566 8258 25618 8270
rect 25566 8194 25618 8206
rect 29262 8258 29314 8270
rect 29262 8194 29314 8206
rect 29934 8258 29986 8270
rect 33070 8258 33122 8270
rect 37214 8258 37266 8270
rect 30706 8206 30718 8258
rect 30770 8206 30782 8258
rect 32610 8206 32622 8258
rect 32674 8206 32686 8258
rect 33842 8206 33854 8258
rect 33906 8206 33918 8258
rect 29934 8194 29986 8206
rect 33070 8194 33122 8206
rect 37214 8194 37266 8206
rect 37438 8258 37490 8270
rect 45054 8258 45106 8270
rect 41346 8206 41358 8258
rect 41410 8206 41422 8258
rect 37438 8194 37490 8206
rect 45054 8194 45106 8206
rect 45502 8258 45554 8270
rect 45502 8194 45554 8206
rect 45726 8258 45778 8270
rect 45726 8194 45778 8206
rect 49422 8258 49474 8270
rect 49422 8194 49474 8206
rect 53566 8258 53618 8270
rect 60734 8258 60786 8270
rect 66337 8258 66383 8321
rect 66546 8318 66558 8321
rect 66610 8318 66622 8370
rect 72930 8318 72942 8370
rect 72994 8318 73006 8370
rect 75058 8318 75070 8370
rect 75122 8318 75134 8370
rect 76962 8318 76974 8370
rect 77026 8318 77038 8370
rect 78082 8318 78094 8370
rect 78146 8318 78158 8370
rect 80210 8318 80222 8370
rect 80274 8318 80286 8370
rect 85138 8318 85150 8370
rect 85202 8318 85214 8370
rect 86258 8318 86270 8370
rect 86322 8318 86334 8370
rect 71710 8306 71762 8318
rect 90750 8306 90802 8318
rect 90974 8370 91026 8382
rect 90974 8306 91026 8318
rect 91422 8370 91474 8382
rect 101390 8370 101442 8382
rect 93314 8318 93326 8370
rect 93378 8318 93390 8370
rect 96226 8318 96238 8370
rect 96290 8318 96302 8370
rect 100594 8318 100606 8370
rect 100658 8318 100670 8370
rect 104626 8318 104638 8370
rect 104690 8318 104702 8370
rect 106194 8318 106206 8370
rect 106258 8318 106270 8370
rect 111346 8318 111358 8370
rect 111410 8318 111422 8370
rect 113474 8318 113486 8370
rect 113538 8318 113550 8370
rect 115378 8318 115390 8370
rect 115442 8318 115454 8370
rect 91422 8306 91474 8318
rect 101390 8306 101442 8318
rect 66670 8258 66722 8270
rect 54338 8206 54350 8258
rect 54402 8206 54414 8258
rect 63186 8206 63198 8258
rect 63250 8206 63262 8258
rect 66322 8206 66334 8258
rect 66386 8206 66398 8258
rect 53566 8194 53618 8206
rect 60734 8194 60786 8206
rect 66670 8194 66722 8206
rect 67006 8258 67058 8270
rect 67006 8194 67058 8206
rect 67230 8258 67282 8270
rect 67230 8194 67282 8206
rect 67454 8258 67506 8270
rect 67454 8194 67506 8206
rect 67790 8258 67842 8270
rect 75406 8258 75458 8270
rect 72258 8206 72270 8258
rect 72322 8206 72334 8258
rect 67790 8194 67842 8206
rect 75406 8194 75458 8206
rect 75742 8258 75794 8270
rect 77534 8258 77586 8270
rect 82910 8258 82962 8270
rect 84254 8258 84306 8270
rect 85486 8258 85538 8270
rect 77074 8206 77086 8258
rect 77138 8206 77150 8258
rect 80994 8206 81006 8258
rect 81058 8206 81070 8258
rect 81442 8206 81454 8258
rect 81506 8206 81518 8258
rect 81890 8206 81902 8258
rect 81954 8206 81966 8258
rect 82226 8206 82238 8258
rect 82290 8206 82302 8258
rect 84018 8206 84030 8258
rect 84082 8206 84094 8258
rect 84690 8206 84702 8258
rect 84754 8206 84766 8258
rect 85026 8206 85038 8258
rect 85090 8206 85102 8258
rect 75742 8194 75794 8206
rect 77534 8194 77586 8206
rect 82910 8194 82962 8206
rect 84254 8194 84306 8206
rect 85486 8194 85538 8206
rect 86158 8258 86210 8270
rect 86158 8194 86210 8206
rect 88286 8258 88338 8270
rect 88286 8194 88338 8206
rect 88846 8258 88898 8270
rect 88846 8194 88898 8206
rect 88958 8258 89010 8270
rect 88958 8194 89010 8206
rect 89294 8258 89346 8270
rect 90526 8258 90578 8270
rect 89954 8206 89966 8258
rect 90018 8206 90030 8258
rect 89294 8194 89346 8206
rect 90526 8194 90578 8206
rect 93886 8258 93938 8270
rect 93886 8194 93938 8206
rect 94334 8258 94386 8270
rect 94334 8194 94386 8206
rect 95230 8258 95282 8270
rect 95230 8194 95282 8206
rect 95566 8258 95618 8270
rect 105198 8258 105250 8270
rect 106542 8258 106594 8270
rect 99138 8206 99150 8258
rect 99202 8206 99214 8258
rect 100034 8206 100046 8258
rect 100098 8206 100110 8258
rect 100258 8206 100270 8258
rect 100322 8206 100334 8258
rect 101714 8206 101726 8258
rect 101778 8206 101790 8258
rect 106082 8206 106094 8258
rect 106146 8206 106158 8258
rect 95566 8194 95618 8206
rect 105198 8194 105250 8206
rect 106542 8194 106594 8206
rect 110686 8258 110738 8270
rect 117182 8258 117234 8270
rect 114258 8206 114270 8258
rect 114322 8206 114334 8258
rect 110686 8194 110738 8206
rect 117182 8194 117234 8206
rect 117518 8258 117570 8270
rect 117518 8194 117570 8206
rect 118302 8258 118354 8270
rect 118302 8194 118354 8206
rect 118750 8258 118802 8270
rect 118750 8194 118802 8206
rect 20414 8146 20466 8158
rect 18050 8094 18062 8146
rect 18114 8094 18126 8146
rect 20414 8082 20466 8094
rect 21422 8146 21474 8158
rect 21422 8082 21474 8094
rect 21534 8146 21586 8158
rect 21534 8082 21586 8094
rect 22766 8146 22818 8158
rect 22766 8082 22818 8094
rect 22878 8146 22930 8158
rect 22878 8082 22930 8094
rect 25230 8146 25282 8158
rect 25230 8082 25282 8094
rect 25342 8146 25394 8158
rect 25342 8082 25394 8094
rect 25790 8146 25842 8158
rect 25790 8082 25842 8094
rect 25902 8146 25954 8158
rect 25902 8082 25954 8094
rect 27022 8146 27074 8158
rect 27022 8082 27074 8094
rect 27246 8146 27298 8158
rect 27246 8082 27298 8094
rect 28702 8146 28754 8158
rect 28702 8082 28754 8094
rect 30046 8146 30098 8158
rect 38110 8146 38162 8158
rect 47854 8146 47906 8158
rect 30370 8094 30382 8146
rect 30434 8094 30446 8146
rect 36194 8094 36206 8146
rect 36258 8094 36270 8146
rect 43810 8094 43822 8146
rect 43874 8094 43886 8146
rect 46274 8094 46286 8146
rect 46338 8094 46350 8146
rect 30046 8082 30098 8094
rect 38110 8082 38162 8094
rect 47854 8082 47906 8094
rect 47966 8146 48018 8158
rect 51886 8146 51938 8158
rect 49746 8094 49758 8146
rect 49810 8094 49822 8146
rect 47966 8082 48018 8094
rect 51886 8082 51938 8094
rect 52670 8146 52722 8158
rect 52670 8082 52722 8094
rect 53006 8146 53058 8158
rect 53006 8082 53058 8094
rect 53230 8146 53282 8158
rect 60510 8146 60562 8158
rect 59490 8094 59502 8146
rect 59554 8094 59566 8146
rect 53230 8082 53282 8094
rect 60510 8082 60562 8094
rect 61070 8146 61122 8158
rect 85710 8146 85762 8158
rect 61506 8094 61518 8146
rect 61570 8094 61582 8146
rect 70354 8094 70366 8146
rect 70418 8094 70430 8146
rect 83234 8094 83246 8146
rect 83298 8094 83310 8146
rect 61070 8082 61122 8094
rect 85710 8082 85762 8094
rect 86270 8146 86322 8158
rect 86270 8082 86322 8094
rect 86494 8146 86546 8158
rect 86494 8082 86546 8094
rect 86718 8146 86770 8158
rect 86718 8082 86770 8094
rect 87502 8146 87554 8158
rect 87502 8082 87554 8094
rect 88398 8146 88450 8158
rect 88398 8082 88450 8094
rect 89182 8146 89234 8158
rect 93662 8146 93714 8158
rect 91970 8094 91982 8146
rect 92034 8094 92046 8146
rect 89182 8082 89234 8094
rect 93662 8082 93714 8094
rect 95678 8146 95730 8158
rect 95678 8082 95730 8094
rect 95790 8146 95842 8158
rect 110910 8146 110962 8158
rect 98354 8094 98366 8146
rect 98418 8094 98430 8146
rect 102498 8094 102510 8146
rect 102562 8094 102574 8146
rect 110226 8094 110238 8146
rect 110290 8094 110302 8146
rect 95790 8082 95842 8094
rect 110910 8082 110962 8094
rect 111022 8146 111074 8158
rect 111022 8082 111074 8094
rect 114606 8146 114658 8158
rect 114606 8082 114658 8094
rect 114942 8146 114994 8158
rect 116610 8094 116622 8146
rect 116674 8094 116686 8146
rect 114942 8082 114994 8094
rect 20638 8034 20690 8046
rect 20638 7970 20690 7982
rect 21198 8034 21250 8046
rect 21198 7970 21250 7982
rect 22318 8034 22370 8046
rect 22318 7970 22370 7982
rect 23102 8034 23154 8046
rect 23102 7970 23154 7982
rect 24334 8034 24386 8046
rect 24334 7970 24386 7982
rect 24782 8034 24834 8046
rect 24782 7970 24834 7982
rect 25006 8034 25058 8046
rect 26574 8034 26626 8046
rect 26226 7982 26238 8034
rect 26290 7982 26302 8034
rect 25006 7970 25058 7982
rect 26574 7970 26626 7982
rect 27582 8034 27634 8046
rect 27582 7970 27634 7982
rect 38222 8034 38274 8046
rect 38222 7970 38274 7982
rect 45278 8034 45330 8046
rect 45278 7970 45330 7982
rect 48190 8034 48242 8046
rect 48190 7970 48242 7982
rect 51550 8034 51602 8046
rect 51550 7970 51602 7982
rect 51998 8034 52050 8046
rect 51998 7970 52050 7982
rect 52222 8034 52274 8046
rect 52222 7970 52274 7982
rect 52782 8034 52834 8046
rect 52782 7970 52834 7982
rect 53902 8034 53954 8046
rect 53902 7970 53954 7982
rect 67118 8034 67170 8046
rect 67118 7970 67170 7982
rect 67678 8034 67730 8046
rect 67678 7970 67730 7982
rect 68238 8034 68290 8046
rect 68238 7970 68290 7982
rect 71150 8034 71202 8046
rect 71150 7970 71202 7982
rect 75518 8034 75570 8046
rect 84366 8034 84418 8046
rect 77410 7982 77422 8034
rect 77474 7982 77486 8034
rect 82114 7982 82126 8034
rect 82178 7982 82190 8034
rect 75518 7970 75570 7982
rect 84366 7970 84418 7982
rect 84478 8034 84530 8046
rect 84478 7970 84530 7982
rect 85262 8034 85314 8046
rect 85262 7970 85314 7982
rect 87166 8034 87218 8046
rect 87166 7970 87218 7982
rect 87390 8034 87442 8046
rect 87390 7970 87442 7982
rect 88622 8034 88674 8046
rect 88622 7970 88674 7982
rect 90190 8034 90242 8046
rect 90190 7970 90242 7982
rect 94782 8034 94834 8046
rect 94782 7970 94834 7982
rect 99598 8034 99650 8046
rect 99598 7970 99650 7982
rect 104862 8034 104914 8046
rect 104862 7970 104914 7982
rect 105086 8034 105138 8046
rect 107662 8034 107714 8046
rect 106418 7982 106430 8034
rect 106482 7982 106494 8034
rect 105086 7970 105138 7982
rect 107662 7970 107714 7982
rect 107886 8034 107938 8046
rect 107886 7970 107938 7982
rect 114718 8034 114770 8046
rect 114718 7970 114770 7982
rect 117294 8034 117346 8046
rect 117294 7970 117346 7982
rect 117854 8034 117906 8046
rect 117854 7970 117906 7982
rect 119198 8034 119250 8046
rect 119198 7970 119250 7982
rect 1344 7866 158592 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 81278 7866
rect 81330 7814 81382 7866
rect 81434 7814 81486 7866
rect 81538 7814 111998 7866
rect 112050 7814 112102 7866
rect 112154 7814 112206 7866
rect 112258 7814 142718 7866
rect 142770 7814 142822 7866
rect 142874 7814 142926 7866
rect 142978 7814 158592 7866
rect 1344 7780 158592 7814
rect 23102 7698 23154 7710
rect 23102 7634 23154 7646
rect 24558 7698 24610 7710
rect 24558 7634 24610 7646
rect 26014 7698 26066 7710
rect 29486 7698 29538 7710
rect 28018 7646 28030 7698
rect 28082 7646 28094 7698
rect 26014 7634 26066 7646
rect 29486 7634 29538 7646
rect 32174 7698 32226 7710
rect 40238 7698 40290 7710
rect 35634 7646 35646 7698
rect 35698 7646 35710 7698
rect 32174 7634 32226 7646
rect 40238 7634 40290 7646
rect 41022 7698 41074 7710
rect 41022 7634 41074 7646
rect 49534 7698 49586 7710
rect 49534 7634 49586 7646
rect 50654 7698 50706 7710
rect 50654 7634 50706 7646
rect 51438 7698 51490 7710
rect 51438 7634 51490 7646
rect 56702 7698 56754 7710
rect 56702 7634 56754 7646
rect 57262 7698 57314 7710
rect 57262 7634 57314 7646
rect 64430 7698 64482 7710
rect 64430 7634 64482 7646
rect 65326 7698 65378 7710
rect 66558 7698 66610 7710
rect 65650 7646 65662 7698
rect 65714 7646 65726 7698
rect 65326 7634 65378 7646
rect 66558 7634 66610 7646
rect 85934 7698 85986 7710
rect 94670 7698 94722 7710
rect 87378 7646 87390 7698
rect 87442 7646 87454 7698
rect 85934 7634 85986 7646
rect 94670 7634 94722 7646
rect 95902 7698 95954 7710
rect 95902 7634 95954 7646
rect 110574 7698 110626 7710
rect 111470 7698 111522 7710
rect 110898 7646 110910 7698
rect 110962 7646 110974 7698
rect 110574 7634 110626 7646
rect 111470 7634 111522 7646
rect 118750 7698 118802 7710
rect 118750 7634 118802 7646
rect 119870 7698 119922 7710
rect 119870 7634 119922 7646
rect 23998 7586 24050 7598
rect 23998 7522 24050 7534
rect 24334 7586 24386 7598
rect 24334 7522 24386 7534
rect 24670 7586 24722 7598
rect 28702 7586 28754 7598
rect 37214 7586 37266 7598
rect 49198 7586 49250 7598
rect 27234 7534 27246 7586
rect 27298 7534 27310 7586
rect 31042 7534 31054 7586
rect 31106 7534 31118 7586
rect 34290 7534 34302 7586
rect 34354 7534 34366 7586
rect 34738 7534 34750 7586
rect 34802 7534 34814 7586
rect 39218 7534 39230 7586
rect 39282 7534 39294 7586
rect 39554 7534 39566 7586
rect 39618 7534 39630 7586
rect 42802 7534 42814 7586
rect 42866 7534 42878 7586
rect 24670 7522 24722 7534
rect 28702 7522 28754 7534
rect 37214 7522 37266 7534
rect 49198 7522 49250 7534
rect 49310 7586 49362 7598
rect 49310 7522 49362 7534
rect 54462 7586 54514 7598
rect 54462 7522 54514 7534
rect 56590 7586 56642 7598
rect 56590 7522 56642 7534
rect 57374 7586 57426 7598
rect 72270 7586 72322 7598
rect 58706 7534 58718 7586
rect 58770 7534 58782 7586
rect 63522 7534 63534 7586
rect 63586 7534 63598 7586
rect 67778 7534 67790 7586
rect 67842 7534 67854 7586
rect 71474 7534 71486 7586
rect 71538 7534 71550 7586
rect 57374 7522 57426 7534
rect 72270 7522 72322 7534
rect 72606 7586 72658 7598
rect 72606 7522 72658 7534
rect 73166 7586 73218 7598
rect 92094 7586 92146 7598
rect 94894 7586 94946 7598
rect 74610 7534 74622 7586
rect 74674 7534 74686 7586
rect 78418 7534 78430 7586
rect 78482 7534 78494 7586
rect 82674 7534 82686 7586
rect 82738 7534 82750 7586
rect 88722 7534 88734 7586
rect 88786 7534 88798 7586
rect 92754 7534 92766 7586
rect 92818 7534 92830 7586
rect 73166 7522 73218 7534
rect 92094 7522 92146 7534
rect 94894 7522 94946 7534
rect 95790 7586 95842 7598
rect 120318 7586 120370 7598
rect 96338 7534 96350 7586
rect 96402 7534 96414 7586
rect 98018 7534 98030 7586
rect 98082 7534 98094 7586
rect 100370 7534 100382 7586
rect 100434 7534 100446 7586
rect 102050 7534 102062 7586
rect 102114 7534 102126 7586
rect 106306 7534 106318 7586
rect 106370 7534 106382 7586
rect 108882 7534 108894 7586
rect 108946 7534 108958 7586
rect 114594 7534 114606 7586
rect 114658 7534 114670 7586
rect 116386 7534 116398 7586
rect 116450 7534 116462 7586
rect 95790 7522 95842 7534
rect 120318 7522 120370 7534
rect 22878 7474 22930 7486
rect 19842 7422 19854 7474
rect 19906 7422 19918 7474
rect 22878 7410 22930 7422
rect 23214 7474 23266 7486
rect 23214 7410 23266 7422
rect 23886 7474 23938 7486
rect 23886 7410 23938 7422
rect 28366 7474 28418 7486
rect 29150 7474 29202 7486
rect 32622 7474 32674 7486
rect 39902 7474 39954 7486
rect 28914 7422 28926 7474
rect 28978 7422 28990 7474
rect 29250 7422 29262 7474
rect 29314 7422 29326 7474
rect 33170 7422 33182 7474
rect 33234 7422 33246 7474
rect 33730 7422 33742 7474
rect 33794 7422 33806 7474
rect 34626 7422 34638 7474
rect 34690 7422 34702 7474
rect 38434 7422 38446 7474
rect 38498 7422 38510 7474
rect 28366 7410 28418 7422
rect 29150 7410 29202 7422
rect 32622 7410 32674 7422
rect 39902 7410 39954 7422
rect 41358 7474 41410 7486
rect 54014 7474 54066 7486
rect 42018 7422 42030 7474
rect 42082 7422 42094 7474
rect 45378 7422 45390 7474
rect 45442 7422 45454 7474
rect 50194 7422 50206 7474
rect 50258 7422 50270 7474
rect 52098 7422 52110 7474
rect 52162 7422 52174 7474
rect 52546 7422 52558 7474
rect 52610 7422 52622 7474
rect 53554 7422 53566 7474
rect 53618 7422 53630 7474
rect 41358 7410 41410 7422
rect 54014 7410 54066 7422
rect 54686 7474 54738 7486
rect 54686 7410 54738 7422
rect 55134 7474 55186 7486
rect 55134 7410 55186 7422
rect 55694 7474 55746 7486
rect 55694 7410 55746 7422
rect 56926 7474 56978 7486
rect 56926 7410 56978 7422
rect 57598 7474 57650 7486
rect 66446 7474 66498 7486
rect 72942 7474 72994 7486
rect 58034 7422 58046 7474
rect 58098 7422 58110 7474
rect 67106 7422 67118 7474
rect 67170 7422 67182 7474
rect 57598 7410 57650 7422
rect 66446 7410 66498 7422
rect 72942 7410 72994 7422
rect 73614 7474 73666 7486
rect 86718 7474 86770 7486
rect 73938 7422 73950 7474
rect 74002 7422 74014 7474
rect 78978 7422 78990 7474
rect 79042 7422 79054 7474
rect 81554 7422 81566 7474
rect 81618 7422 81630 7474
rect 73614 7410 73666 7422
rect 86718 7410 86770 7422
rect 87054 7474 87106 7486
rect 91422 7474 91474 7486
rect 87938 7422 87950 7474
rect 88002 7422 88014 7474
rect 87054 7410 87106 7422
rect 91422 7410 91474 7422
rect 91646 7474 91698 7486
rect 91646 7410 91698 7422
rect 93998 7474 94050 7486
rect 93998 7410 94050 7422
rect 94558 7474 94610 7486
rect 94558 7410 94610 7422
rect 95006 7474 95058 7486
rect 102510 7474 102562 7486
rect 96226 7422 96238 7474
rect 96290 7422 96302 7474
rect 97906 7422 97918 7474
rect 97970 7422 97982 7474
rect 99698 7422 99710 7474
rect 99762 7422 99774 7474
rect 95006 7410 95058 7422
rect 102510 7410 102562 7422
rect 103070 7474 103122 7486
rect 117742 7474 117794 7486
rect 103954 7422 103966 7474
rect 104018 7422 104030 7474
rect 104290 7422 104302 7474
rect 104354 7422 104366 7474
rect 105522 7422 105534 7474
rect 105586 7422 105598 7474
rect 115266 7422 115278 7474
rect 115330 7422 115342 7474
rect 103070 7410 103122 7422
rect 117742 7410 117794 7422
rect 25454 7362 25506 7374
rect 48750 7362 48802 7374
rect 20514 7310 20526 7362
rect 20578 7310 20590 7362
rect 22642 7310 22654 7362
rect 22706 7310 22718 7362
rect 26226 7310 26238 7362
rect 26290 7310 26302 7362
rect 29810 7310 29822 7362
rect 29874 7310 29886 7362
rect 33618 7310 33630 7362
rect 33682 7310 33694 7362
rect 44930 7310 44942 7362
rect 44994 7310 45006 7362
rect 46050 7310 46062 7362
rect 46114 7310 46126 7362
rect 48178 7310 48190 7362
rect 48242 7310 48254 7362
rect 25454 7298 25506 7310
rect 48750 7298 48802 7310
rect 49870 7362 49922 7374
rect 49870 7298 49922 7310
rect 54238 7362 54290 7374
rect 64990 7362 65042 7374
rect 60834 7310 60846 7362
rect 60898 7310 60910 7362
rect 61506 7310 61518 7362
rect 61570 7310 61582 7362
rect 54238 7298 54290 7310
rect 64990 7298 65042 7310
rect 66222 7362 66274 7374
rect 73390 7362 73442 7374
rect 79438 7362 79490 7374
rect 69906 7310 69918 7362
rect 69970 7310 69982 7362
rect 70466 7310 70478 7362
rect 70530 7310 70542 7362
rect 76738 7310 76750 7362
rect 76802 7310 76814 7362
rect 77074 7310 77086 7362
rect 77138 7310 77150 7362
rect 66222 7298 66274 7310
rect 73390 7298 73442 7310
rect 79438 7298 79490 7310
rect 86158 7362 86210 7374
rect 91198 7362 91250 7374
rect 112030 7362 112082 7374
rect 119422 7362 119474 7374
rect 90850 7310 90862 7362
rect 90914 7310 90926 7362
rect 92978 7310 92990 7362
rect 93042 7310 93054 7362
rect 100706 7310 100718 7362
rect 100770 7310 100782 7362
rect 104738 7310 104750 7362
rect 104802 7310 104814 7362
rect 108434 7310 108446 7362
rect 108498 7310 108510 7362
rect 110226 7310 110238 7362
rect 110290 7310 110302 7362
rect 112466 7310 112478 7362
rect 112530 7310 112542 7362
rect 117394 7310 117406 7362
rect 117458 7310 117470 7362
rect 118178 7310 118190 7362
rect 118242 7310 118254 7362
rect 86158 7298 86210 7310
rect 91198 7298 91250 7310
rect 112030 7298 112082 7310
rect 119422 7298 119474 7310
rect 23998 7250 24050 7262
rect 23998 7186 24050 7198
rect 41022 7250 41074 7262
rect 41022 7186 41074 7198
rect 41134 7250 41186 7262
rect 41134 7186 41186 7198
rect 48862 7250 48914 7262
rect 48862 7186 48914 7198
rect 66558 7250 66610 7262
rect 66558 7186 66610 7198
rect 94334 7250 94386 7262
rect 103954 7198 103966 7250
rect 104018 7198 104030 7250
rect 94334 7186 94386 7198
rect 1344 7082 158592 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 96638 7082
rect 96690 7030 96742 7082
rect 96794 7030 96846 7082
rect 96898 7030 127358 7082
rect 127410 7030 127462 7082
rect 127514 7030 127566 7082
rect 127618 7030 158078 7082
rect 158130 7030 158182 7082
rect 158234 7030 158286 7082
rect 158338 7030 158592 7082
rect 1344 6996 158592 7030
rect 21982 6914 22034 6926
rect 21982 6850 22034 6862
rect 29486 6914 29538 6926
rect 29486 6850 29538 6862
rect 29598 6914 29650 6926
rect 29598 6850 29650 6862
rect 30382 6914 30434 6926
rect 30382 6850 30434 6862
rect 30606 6914 30658 6926
rect 30606 6850 30658 6862
rect 61070 6914 61122 6926
rect 61070 6850 61122 6862
rect 61294 6914 61346 6926
rect 61294 6850 61346 6862
rect 75742 6914 75794 6926
rect 75742 6850 75794 6862
rect 117294 6914 117346 6926
rect 117294 6850 117346 6862
rect 28590 6802 28642 6814
rect 18610 6750 18622 6802
rect 18674 6750 18686 6802
rect 21634 6750 21646 6802
rect 21698 6750 21710 6802
rect 22306 6750 22318 6802
rect 22370 6750 22382 6802
rect 25106 6750 25118 6802
rect 25170 6750 25182 6802
rect 27234 6750 27246 6802
rect 27298 6750 27310 6802
rect 28590 6738 28642 6750
rect 29262 6802 29314 6814
rect 29262 6738 29314 6750
rect 30830 6802 30882 6814
rect 39006 6802 39058 6814
rect 34962 6750 34974 6802
rect 35026 6750 35038 6802
rect 38434 6750 38446 6802
rect 38498 6750 38510 6802
rect 30830 6738 30882 6750
rect 39006 6738 39058 6750
rect 45614 6802 45666 6814
rect 45614 6738 45666 6750
rect 48638 6802 48690 6814
rect 61854 6802 61906 6814
rect 69918 6802 69970 6814
rect 52098 6750 52110 6802
rect 52162 6750 52174 6802
rect 57698 6750 57710 6802
rect 57762 6750 57774 6802
rect 59938 6750 59950 6802
rect 60002 6750 60014 6802
rect 61618 6750 61630 6802
rect 61682 6750 61694 6802
rect 68898 6750 68910 6802
rect 68962 6750 68974 6802
rect 48638 6738 48690 6750
rect 61854 6738 61906 6750
rect 69918 6738 69970 6750
rect 78206 6802 78258 6814
rect 104862 6802 104914 6814
rect 118190 6802 118242 6814
rect 80098 6750 80110 6802
rect 80162 6750 80174 6802
rect 82338 6750 82350 6802
rect 82402 6750 82414 6802
rect 84690 6750 84702 6802
rect 84754 6750 84766 6802
rect 89394 6750 89406 6802
rect 89458 6750 89470 6802
rect 91970 6750 91982 6802
rect 92034 6750 92046 6802
rect 96002 6750 96014 6802
rect 96066 6750 96078 6802
rect 100258 6750 100270 6802
rect 100322 6750 100334 6802
rect 107538 6750 107550 6802
rect 107602 6750 107614 6802
rect 116834 6750 116846 6802
rect 116898 6750 116910 6802
rect 78206 6738 78258 6750
rect 104862 6738 104914 6750
rect 118190 6738 118242 6750
rect 19854 6690 19906 6702
rect 31390 6690 31442 6702
rect 20290 6638 20302 6690
rect 20354 6638 20366 6690
rect 24322 6638 24334 6690
rect 24386 6638 24398 6690
rect 28130 6638 28142 6690
rect 28194 6638 28206 6690
rect 19854 6626 19906 6638
rect 31390 6626 31442 6638
rect 31726 6690 31778 6702
rect 33518 6690 33570 6702
rect 33170 6638 33182 6690
rect 33234 6638 33246 6690
rect 31726 6626 31778 6638
rect 33518 6626 33570 6638
rect 33854 6690 33906 6702
rect 45390 6690 45442 6702
rect 34066 6638 34078 6690
rect 34130 6638 34142 6690
rect 39554 6638 39566 6690
rect 39618 6638 39630 6690
rect 41570 6638 41582 6690
rect 41634 6638 41646 6690
rect 45042 6638 45054 6690
rect 45106 6638 45118 6690
rect 33854 6626 33906 6638
rect 45390 6626 45442 6638
rect 45838 6690 45890 6702
rect 45838 6626 45890 6638
rect 45950 6690 46002 6702
rect 60734 6690 60786 6702
rect 49186 6638 49198 6690
rect 49250 6638 49262 6690
rect 53666 6638 53678 6690
rect 53730 6638 53742 6690
rect 45950 6626 46002 6638
rect 60734 6626 60786 6638
rect 61742 6690 61794 6702
rect 61742 6626 61794 6638
rect 62302 6690 62354 6702
rect 62302 6626 62354 6638
rect 64318 6690 64370 6702
rect 64318 6626 64370 6638
rect 66558 6690 66610 6702
rect 66558 6626 66610 6638
rect 67230 6690 67282 6702
rect 67230 6626 67282 6638
rect 67790 6690 67842 6702
rect 67790 6626 67842 6638
rect 69358 6690 69410 6702
rect 91310 6690 91362 6702
rect 99710 6690 99762 6702
rect 103742 6690 103794 6702
rect 117182 6690 117234 6702
rect 76402 6638 76414 6690
rect 76466 6638 76478 6690
rect 79538 6638 79550 6690
rect 79602 6638 79614 6690
rect 82226 6638 82238 6690
rect 82290 6638 82302 6690
rect 82450 6638 82462 6690
rect 82514 6638 82526 6690
rect 84130 6638 84142 6690
rect 84194 6638 84206 6690
rect 95442 6638 95454 6690
rect 95506 6638 95518 6690
rect 98130 6638 98142 6690
rect 98194 6638 98206 6690
rect 98914 6638 98926 6690
rect 98978 6638 98990 6690
rect 102386 6638 102398 6690
rect 102450 6638 102462 6690
rect 103058 6638 103070 6690
rect 103122 6638 103134 6690
rect 106642 6638 106654 6690
rect 106706 6638 106718 6690
rect 109666 6638 109678 6690
rect 109730 6638 109742 6690
rect 110338 6638 110350 6690
rect 110402 6638 110414 6690
rect 110898 6638 110910 6690
rect 110962 6638 110974 6690
rect 69358 6626 69410 6638
rect 91310 6626 91362 6638
rect 99710 6626 99762 6638
rect 103742 6626 103794 6638
rect 117182 6626 117234 6638
rect 21758 6578 21810 6590
rect 27694 6578 27746 6590
rect 23538 6526 23550 6578
rect 23602 6526 23614 6578
rect 21758 6514 21810 6526
rect 27694 6514 27746 6526
rect 29150 6578 29202 6590
rect 29150 6514 29202 6526
rect 29934 6578 29986 6590
rect 29934 6514 29986 6526
rect 34638 6578 34690 6590
rect 38894 6578 38946 6590
rect 36082 6526 36094 6578
rect 36146 6526 36158 6578
rect 37426 6526 37438 6578
rect 37490 6526 37502 6578
rect 34638 6514 34690 6526
rect 38894 6514 38946 6526
rect 39118 6578 39170 6590
rect 39118 6514 39170 6526
rect 40686 6578 40738 6590
rect 44046 6578 44098 6590
rect 43362 6526 43374 6578
rect 43426 6526 43438 6578
rect 40686 6514 40738 6526
rect 44046 6514 44098 6526
rect 44158 6578 44210 6590
rect 44158 6514 44210 6526
rect 44382 6578 44434 6590
rect 63422 6578 63474 6590
rect 46498 6526 46510 6578
rect 46562 6526 46574 6578
rect 49970 6526 49982 6578
rect 50034 6526 50046 6578
rect 58594 6526 58606 6578
rect 58658 6526 58670 6578
rect 44382 6514 44434 6526
rect 63422 6514 63474 6526
rect 64878 6578 64930 6590
rect 64878 6514 64930 6526
rect 66334 6578 66386 6590
rect 66334 6514 66386 6526
rect 66894 6578 66946 6590
rect 72830 6578 72882 6590
rect 76974 6578 77026 6590
rect 91198 6578 91250 6590
rect 99822 6578 99874 6590
rect 71698 6526 71710 6578
rect 71762 6526 71774 6578
rect 72482 6526 72494 6578
rect 72546 6526 72558 6578
rect 73378 6526 73390 6578
rect 73442 6526 73454 6578
rect 81106 6526 81118 6578
rect 81170 6526 81182 6578
rect 84354 6526 84366 6578
rect 84418 6526 84430 6578
rect 85922 6526 85934 6578
rect 85986 6526 85998 6578
rect 86594 6526 86606 6578
rect 86658 6526 86670 6578
rect 90626 6526 90638 6578
rect 90690 6526 90702 6578
rect 94210 6526 94222 6578
rect 94274 6526 94286 6578
rect 95218 6526 95230 6578
rect 95282 6526 95294 6578
rect 66894 6514 66946 6526
rect 72830 6514 72882 6526
rect 76974 6514 77026 6526
rect 91198 6514 91250 6526
rect 99822 6514 99874 6526
rect 103406 6578 103458 6590
rect 103406 6514 103458 6526
rect 106094 6578 106146 6590
rect 106094 6514 106146 6526
rect 111358 6578 111410 6590
rect 114718 6578 114770 6590
rect 112354 6526 112366 6578
rect 112418 6526 112430 6578
rect 115490 6526 115502 6578
rect 115554 6526 115566 6578
rect 120306 6526 120318 6578
rect 120370 6526 120382 6578
rect 111358 6514 111410 6526
rect 114718 6514 114770 6526
rect 17838 6466 17890 6478
rect 17838 6402 17890 6414
rect 19070 6466 19122 6478
rect 19070 6402 19122 6414
rect 19630 6466 19682 6478
rect 19630 6402 19682 6414
rect 27582 6466 27634 6478
rect 66782 6466 66834 6478
rect 39778 6414 39790 6466
rect 39842 6414 39854 6466
rect 44818 6414 44830 6466
rect 44882 6414 44894 6466
rect 64978 6414 64990 6466
rect 65042 6414 65054 6466
rect 27582 6402 27634 6414
rect 66782 6402 66834 6414
rect 68462 6466 68514 6478
rect 68462 6402 68514 6414
rect 77982 6466 78034 6478
rect 77982 6402 78034 6414
rect 79774 6466 79826 6478
rect 79774 6402 79826 6414
rect 81790 6466 81842 6478
rect 81790 6402 81842 6414
rect 89070 6466 89122 6478
rect 100046 6466 100098 6478
rect 94882 6414 94894 6466
rect 94946 6414 94958 6466
rect 89070 6402 89122 6414
rect 100046 6402 100098 6414
rect 103630 6466 103682 6478
rect 103630 6402 103682 6414
rect 106542 6466 106594 6478
rect 106542 6402 106594 6414
rect 111806 6466 111858 6478
rect 111806 6402 111858 6414
rect 117294 6466 117346 6478
rect 117294 6402 117346 6414
rect 120878 6466 120930 6478
rect 120878 6402 120930 6414
rect 121662 6466 121714 6478
rect 121662 6402 121714 6414
rect 122558 6466 122610 6478
rect 122558 6402 122610 6414
rect 123790 6466 123842 6478
rect 123790 6402 123842 6414
rect 125806 6466 125858 6478
rect 125806 6402 125858 6414
rect 1344 6298 158592 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 81278 6298
rect 81330 6246 81382 6298
rect 81434 6246 81486 6298
rect 81538 6246 111998 6298
rect 112050 6246 112102 6298
rect 112154 6246 112206 6298
rect 112258 6246 142718 6298
rect 142770 6246 142822 6298
rect 142874 6246 142926 6298
rect 142978 6246 158592 6298
rect 1344 6212 158592 6246
rect 20078 6130 20130 6142
rect 20078 6066 20130 6078
rect 21086 6130 21138 6142
rect 21086 6066 21138 6078
rect 22878 6130 22930 6142
rect 22878 6066 22930 6078
rect 30270 6130 30322 6142
rect 30270 6066 30322 6078
rect 35198 6130 35250 6142
rect 42366 6130 42418 6142
rect 39890 6078 39902 6130
rect 39954 6078 39966 6130
rect 35198 6066 35250 6078
rect 42366 6066 42418 6078
rect 43262 6130 43314 6142
rect 43262 6066 43314 6078
rect 71822 6130 71874 6142
rect 71822 6066 71874 6078
rect 79438 6130 79490 6142
rect 79438 6066 79490 6078
rect 88062 6130 88114 6142
rect 88062 6066 88114 6078
rect 94222 6130 94274 6142
rect 94222 6066 94274 6078
rect 95230 6130 95282 6142
rect 95230 6066 95282 6078
rect 102622 6130 102674 6142
rect 102622 6066 102674 6078
rect 108782 6130 108834 6142
rect 108782 6066 108834 6078
rect 109006 6130 109058 6142
rect 109006 6066 109058 6078
rect 114382 6130 114434 6142
rect 114382 6066 114434 6078
rect 21310 6018 21362 6030
rect 25118 6018 25170 6030
rect 39342 6018 39394 6030
rect 53006 6018 53058 6030
rect 18162 5966 18174 6018
rect 18226 5966 18238 6018
rect 24546 5966 24558 6018
rect 24610 5966 24622 6018
rect 27234 5966 27246 6018
rect 27298 5966 27310 6018
rect 29362 5966 29374 6018
rect 29426 5966 29438 6018
rect 32050 5966 32062 6018
rect 32114 5966 32126 6018
rect 34066 5966 34078 6018
rect 34130 5966 34142 6018
rect 37538 5966 37550 6018
rect 37602 5966 37614 6018
rect 47842 5966 47854 6018
rect 47906 5966 47918 6018
rect 51874 5966 51886 6018
rect 51938 5966 51950 6018
rect 21310 5954 21362 5966
rect 25118 5954 25170 5966
rect 39342 5954 39394 5966
rect 53006 5954 53058 5966
rect 53118 6018 53170 6030
rect 53118 5954 53170 5966
rect 53342 6018 53394 6030
rect 56814 6018 56866 6030
rect 68014 6018 68066 6030
rect 87166 6018 87218 6030
rect 55570 5966 55582 6018
rect 55634 5966 55646 6018
rect 60610 5966 60622 6018
rect 60674 5966 60686 6018
rect 61506 5966 61518 6018
rect 61570 5966 61582 6018
rect 64978 5966 64990 6018
rect 65042 5966 65054 6018
rect 73378 5966 73390 6018
rect 73442 5966 73454 6018
rect 76962 5966 76974 6018
rect 77026 5966 77038 6018
rect 80322 5966 80334 6018
rect 80386 5966 80398 6018
rect 53342 5954 53394 5966
rect 56814 5954 56866 5966
rect 68014 5954 68066 5966
rect 87166 5954 87218 5966
rect 87278 6018 87330 6030
rect 87278 5954 87330 5966
rect 88174 6018 88226 6030
rect 95118 6018 95170 6030
rect 98702 6018 98754 6030
rect 102510 6018 102562 6030
rect 91858 5966 91870 6018
rect 91922 5966 91934 6018
rect 96226 5966 96238 6018
rect 96290 5966 96302 6018
rect 99026 5966 99038 6018
rect 99090 5966 99102 6018
rect 101714 5966 101726 6018
rect 101778 5966 101790 6018
rect 88174 5954 88226 5966
rect 95118 5954 95170 5966
rect 98702 5954 98754 5966
rect 102510 5954 102562 5966
rect 102846 6018 102898 6030
rect 105758 6018 105810 6030
rect 109118 6018 109170 6030
rect 111358 6018 111410 6030
rect 121214 6018 121266 6030
rect 124350 6018 124402 6030
rect 105410 5966 105422 6018
rect 105474 5966 105486 6018
rect 107874 5966 107886 6018
rect 107938 5966 107950 6018
rect 110674 5966 110686 6018
rect 110738 5966 110750 6018
rect 113474 5966 113486 6018
rect 113538 5966 113550 6018
rect 115154 5966 115166 6018
rect 115218 5966 115230 6018
rect 123218 5966 123230 6018
rect 123282 5966 123294 6018
rect 125570 5966 125582 6018
rect 125634 5966 125646 6018
rect 102846 5954 102898 5966
rect 105758 5954 105810 5966
rect 109118 5954 109170 5966
rect 111358 5954 111410 5966
rect 121214 5954 121266 5966
rect 124350 5954 124402 5966
rect 21870 5906 21922 5918
rect 30270 5906 30322 5918
rect 22642 5854 22654 5906
rect 22706 5854 22718 5906
rect 21870 5842 21922 5854
rect 30270 5842 30322 5854
rect 30606 5906 30658 5918
rect 38446 5906 38498 5918
rect 34962 5854 34974 5906
rect 35026 5854 35038 5906
rect 36418 5854 36430 5906
rect 36482 5854 36494 5906
rect 37874 5854 37886 5906
rect 37938 5854 37950 5906
rect 30606 5842 30658 5854
rect 38446 5842 38498 5854
rect 39006 5906 39058 5918
rect 39006 5842 39058 5854
rect 39566 5906 39618 5918
rect 39566 5842 39618 5854
rect 39790 5906 39842 5918
rect 39790 5842 39842 5854
rect 39902 5906 39954 5918
rect 40910 5906 40962 5918
rect 40226 5854 40238 5906
rect 40290 5854 40302 5906
rect 39902 5842 39954 5854
rect 40910 5842 40962 5854
rect 41022 5906 41074 5918
rect 41806 5906 41858 5918
rect 57038 5906 57090 5918
rect 41458 5854 41470 5906
rect 41522 5854 41534 5906
rect 43698 5854 43710 5906
rect 43762 5854 43774 5906
rect 48850 5854 48862 5906
rect 48914 5854 48926 5906
rect 52658 5854 52670 5906
rect 52722 5854 52734 5906
rect 41022 5842 41074 5854
rect 41806 5842 41858 5854
rect 57038 5842 57090 5854
rect 57262 5906 57314 5918
rect 57262 5842 57314 5854
rect 58270 5906 58322 5918
rect 66782 5906 66834 5918
rect 64418 5854 64430 5906
rect 64482 5854 64494 5906
rect 58270 5842 58322 5854
rect 66782 5842 66834 5854
rect 67342 5906 67394 5918
rect 67342 5842 67394 5854
rect 67566 5906 67618 5918
rect 67566 5842 67618 5854
rect 67678 5906 67730 5918
rect 85262 5906 85314 5918
rect 68450 5854 68462 5906
rect 68514 5854 68526 5906
rect 69122 5854 69134 5906
rect 69186 5854 69198 5906
rect 72258 5854 72270 5906
rect 72322 5854 72334 5906
rect 76402 5854 76414 5906
rect 76466 5854 76478 5906
rect 82114 5854 82126 5906
rect 82178 5854 82190 5906
rect 67678 5842 67730 5854
rect 85262 5842 85314 5854
rect 85822 5906 85874 5918
rect 85822 5842 85874 5854
rect 86046 5906 86098 5918
rect 86046 5842 86098 5854
rect 86494 5906 86546 5918
rect 86494 5842 86546 5854
rect 86718 5906 86770 5918
rect 86718 5842 86770 5854
rect 86942 5906 86994 5918
rect 86942 5842 86994 5854
rect 87838 5906 87890 5918
rect 102958 5906 103010 5918
rect 120654 5906 120706 5918
rect 124014 5906 124066 5918
rect 89058 5854 89070 5906
rect 89122 5854 89134 5906
rect 89842 5854 89854 5906
rect 89906 5854 89918 5906
rect 90514 5854 90526 5906
rect 90578 5854 90590 5906
rect 117842 5854 117854 5906
rect 117906 5854 117918 5906
rect 118066 5854 118078 5906
rect 118130 5854 118142 5906
rect 119634 5854 119646 5906
rect 119698 5854 119710 5906
rect 119970 5854 119982 5906
rect 120034 5854 120046 5906
rect 120978 5854 120990 5906
rect 121042 5854 121054 5906
rect 87838 5842 87890 5854
rect 102958 5842 103010 5854
rect 120654 5842 120706 5854
rect 124014 5842 124066 5854
rect 17838 5794 17890 5806
rect 20638 5794 20690 5806
rect 56926 5794 56978 5806
rect 19282 5742 19294 5794
rect 19346 5742 19358 5794
rect 23202 5742 23214 5794
rect 23266 5742 23278 5794
rect 28466 5742 28478 5794
rect 28530 5742 28542 5794
rect 31266 5742 31278 5794
rect 31330 5742 31342 5794
rect 33282 5742 33294 5794
rect 33346 5742 33358 5794
rect 37986 5742 37998 5794
rect 38050 5742 38062 5794
rect 42802 5742 42814 5794
rect 42866 5742 42878 5794
rect 46498 5742 46510 5794
rect 46562 5742 46574 5794
rect 49186 5742 49198 5794
rect 49250 5742 49262 5794
rect 49746 5742 49758 5794
rect 49810 5742 49822 5794
rect 53554 5742 53566 5794
rect 53618 5742 53630 5794
rect 17838 5730 17890 5742
rect 20638 5730 20690 5742
rect 56926 5730 56978 5742
rect 57710 5794 57762 5806
rect 86270 5794 86322 5806
rect 103742 5794 103794 5806
rect 116958 5794 117010 5806
rect 121662 5794 121714 5806
rect 127710 5794 127762 5806
rect 58594 5742 58606 5794
rect 58658 5742 58670 5794
rect 63746 5742 63758 5794
rect 63810 5742 63822 5794
rect 65538 5742 65550 5794
rect 65602 5742 65614 5794
rect 71250 5742 71262 5794
rect 71314 5742 71326 5794
rect 81666 5742 81678 5794
rect 81730 5742 81742 5794
rect 82786 5742 82798 5794
rect 82850 5742 82862 5794
rect 84914 5742 84926 5794
rect 84978 5742 84990 5794
rect 89730 5742 89742 5794
rect 89794 5742 89806 5794
rect 93874 5742 93886 5794
rect 93938 5742 93950 5794
rect 94658 5742 94670 5794
rect 94722 5742 94734 5794
rect 100370 5742 100382 5794
rect 100434 5742 100446 5794
rect 100706 5742 100718 5794
rect 100770 5742 100782 5794
rect 104290 5742 104302 5794
rect 104354 5742 104366 5794
rect 109442 5742 109454 5794
rect 109506 5742 109518 5794
rect 117618 5742 117630 5794
rect 117682 5742 117694 5794
rect 119410 5742 119422 5794
rect 119474 5742 119486 5794
rect 122210 5742 122222 5794
rect 122274 5742 122286 5794
rect 126578 5742 126590 5794
rect 126642 5742 126654 5794
rect 57710 5730 57762 5742
rect 86270 5730 86322 5742
rect 103742 5730 103794 5742
rect 116958 5730 117010 5742
rect 121662 5730 121714 5742
rect 127710 5730 127762 5742
rect 138910 5794 138962 5806
rect 138910 5730 138962 5742
rect 143838 5794 143890 5806
rect 143838 5730 143890 5742
rect 144174 5794 144226 5806
rect 144174 5730 144226 5742
rect 30382 5682 30434 5694
rect 30382 5618 30434 5630
rect 41246 5682 41298 5694
rect 41246 5618 41298 5630
rect 44606 5682 44658 5694
rect 44606 5618 44658 5630
rect 74174 5682 74226 5694
rect 139022 5682 139074 5694
rect 118626 5630 118638 5682
rect 118690 5630 118702 5682
rect 74174 5618 74226 5630
rect 139022 5618 139074 5630
rect 1344 5514 158592 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 96638 5514
rect 96690 5462 96742 5514
rect 96794 5462 96846 5514
rect 96898 5462 127358 5514
rect 127410 5462 127462 5514
rect 127514 5462 127566 5514
rect 127618 5462 158078 5514
rect 158130 5462 158182 5514
rect 158234 5462 158286 5514
rect 158338 5462 158592 5514
rect 1344 5428 158592 5462
rect 21646 5346 21698 5358
rect 15922 5294 15934 5346
rect 15986 5294 15998 5346
rect 21646 5282 21698 5294
rect 32286 5346 32338 5358
rect 32286 5282 32338 5294
rect 36878 5346 36930 5358
rect 45278 5346 45330 5358
rect 40450 5294 40462 5346
rect 40514 5294 40526 5346
rect 36878 5282 36930 5294
rect 45278 5282 45330 5294
rect 45390 5346 45442 5358
rect 45390 5282 45442 5294
rect 45614 5346 45666 5358
rect 45614 5282 45666 5294
rect 52782 5346 52834 5358
rect 52782 5282 52834 5294
rect 60622 5346 60674 5358
rect 98702 5346 98754 5358
rect 68450 5294 68462 5346
rect 68514 5294 68526 5346
rect 60622 5282 60674 5294
rect 98702 5282 98754 5294
rect 99038 5346 99090 5358
rect 99038 5282 99090 5294
rect 102510 5346 102562 5358
rect 102510 5282 102562 5294
rect 125918 5346 125970 5358
rect 125918 5282 125970 5294
rect 16382 5234 16434 5246
rect 19070 5234 19122 5246
rect 32958 5234 33010 5246
rect 46286 5234 46338 5246
rect 76974 5234 77026 5246
rect 17490 5182 17502 5234
rect 17554 5182 17566 5234
rect 19282 5182 19294 5234
rect 19346 5182 19358 5234
rect 23650 5182 23662 5234
rect 23714 5182 23726 5234
rect 25778 5182 25790 5234
rect 25842 5182 25854 5234
rect 26338 5182 26350 5234
rect 26402 5182 26414 5234
rect 27122 5182 27134 5234
rect 27186 5182 27198 5234
rect 34738 5182 34750 5234
rect 34802 5182 34814 5234
rect 39890 5182 39902 5234
rect 39954 5182 39966 5234
rect 43250 5182 43262 5234
rect 43314 5182 43326 5234
rect 48738 5182 48750 5234
rect 48802 5182 48814 5234
rect 57026 5182 57038 5234
rect 57090 5182 57102 5234
rect 61618 5182 61630 5234
rect 61682 5182 61694 5234
rect 64418 5182 64430 5234
rect 64482 5182 64494 5234
rect 69458 5182 69470 5234
rect 69522 5182 69534 5234
rect 74162 5182 74174 5234
rect 74226 5182 74238 5234
rect 16382 5170 16434 5182
rect 19070 5170 19122 5182
rect 32958 5170 33010 5182
rect 46286 5170 46338 5182
rect 76974 5170 77026 5182
rect 79214 5234 79266 5246
rect 79214 5170 79266 5182
rect 80334 5234 80386 5246
rect 110126 5234 110178 5246
rect 85362 5182 85374 5234
rect 85426 5182 85438 5234
rect 89506 5182 89518 5234
rect 89570 5182 89582 5234
rect 89954 5182 89966 5234
rect 90018 5182 90030 5234
rect 92418 5182 92430 5234
rect 92482 5182 92494 5234
rect 102834 5182 102846 5234
rect 102898 5182 102910 5234
rect 108770 5182 108782 5234
rect 108834 5182 108846 5234
rect 80334 5170 80386 5182
rect 110126 5170 110178 5182
rect 113038 5234 113090 5246
rect 113038 5170 113090 5182
rect 116174 5234 116226 5246
rect 116174 5170 116226 5182
rect 120542 5234 120594 5246
rect 121090 5182 121102 5234
rect 121154 5182 121166 5234
rect 123218 5182 123230 5234
rect 123282 5182 123294 5234
rect 134978 5182 134990 5234
rect 135042 5182 135054 5234
rect 140130 5182 140142 5234
rect 140194 5182 140206 5234
rect 142930 5182 142942 5234
rect 142994 5182 143006 5234
rect 150658 5182 150670 5234
rect 150722 5182 150734 5234
rect 120542 5170 120594 5182
rect 15374 5122 15426 5134
rect 15374 5058 15426 5070
rect 15598 5122 15650 5134
rect 26798 5122 26850 5134
rect 16818 5070 16830 5122
rect 16882 5070 16894 5122
rect 21298 5070 21310 5122
rect 21362 5070 21374 5122
rect 21858 5070 21870 5122
rect 21922 5070 21934 5122
rect 22866 5070 22878 5122
rect 22930 5070 22942 5122
rect 15598 5058 15650 5070
rect 26798 5058 26850 5070
rect 29486 5122 29538 5134
rect 45726 5122 45778 5134
rect 52670 5122 52722 5134
rect 33170 5070 33182 5122
rect 33234 5070 33246 5122
rect 35746 5070 35758 5122
rect 35810 5070 35822 5122
rect 40338 5070 40350 5122
rect 40402 5070 40414 5122
rect 42242 5070 42254 5122
rect 42306 5070 42318 5122
rect 43698 5070 43710 5122
rect 43762 5070 43774 5122
rect 50418 5070 50430 5122
rect 50482 5070 50494 5122
rect 51762 5070 51774 5122
rect 51826 5070 51838 5122
rect 29486 5058 29538 5070
rect 45726 5058 45778 5070
rect 52670 5058 52722 5070
rect 53342 5122 53394 5134
rect 53342 5058 53394 5070
rect 53454 5122 53506 5134
rect 53454 5058 53506 5070
rect 53678 5122 53730 5134
rect 53678 5058 53730 5070
rect 53790 5122 53842 5134
rect 60734 5122 60786 5134
rect 71598 5122 71650 5134
rect 54226 5070 54238 5122
rect 54290 5070 54302 5122
rect 54898 5070 54910 5122
rect 54962 5070 54974 5122
rect 63634 5070 63646 5122
rect 63698 5070 63710 5122
rect 65762 5070 65774 5122
rect 65826 5070 65838 5122
rect 67778 5070 67790 5122
rect 67842 5070 67854 5122
rect 68674 5070 68686 5122
rect 68738 5070 68750 5122
rect 69010 5070 69022 5122
rect 69074 5070 69086 5122
rect 53790 5058 53842 5070
rect 60734 5058 60786 5070
rect 71598 5058 71650 5070
rect 72046 5122 72098 5134
rect 82910 5122 82962 5134
rect 77186 5070 77198 5122
rect 77250 5070 77262 5122
rect 79650 5070 79662 5122
rect 79714 5070 79726 5122
rect 72046 5058 72098 5070
rect 82910 5058 82962 5070
rect 83246 5122 83298 5134
rect 83246 5058 83298 5070
rect 83582 5122 83634 5134
rect 98926 5122 98978 5134
rect 103518 5122 103570 5134
rect 84130 5070 84142 5122
rect 84194 5070 84206 5122
rect 85250 5070 85262 5122
rect 85314 5070 85326 5122
rect 85586 5070 85598 5122
rect 85650 5070 85662 5122
rect 86706 5070 86718 5122
rect 86770 5070 86782 5122
rect 94210 5070 94222 5122
rect 94274 5070 94286 5122
rect 95554 5070 95566 5122
rect 95618 5070 95630 5122
rect 103170 5070 103182 5122
rect 103234 5070 103246 5122
rect 83582 5058 83634 5070
rect 98926 5058 98978 5070
rect 103518 5058 103570 5070
rect 103854 5122 103906 5134
rect 129166 5122 129218 5134
rect 111906 5070 111918 5122
rect 111970 5070 111982 5122
rect 113250 5070 113262 5122
rect 113314 5070 113326 5122
rect 116386 5070 116398 5122
rect 116450 5070 116462 5122
rect 103854 5058 103906 5070
rect 129166 5058 129218 5070
rect 132302 5122 132354 5134
rect 132302 5058 132354 5070
rect 137454 5122 137506 5134
rect 137454 5058 137506 5070
rect 138238 5122 138290 5134
rect 138238 5058 138290 5070
rect 142718 5122 142770 5134
rect 142718 5058 142770 5070
rect 147646 5122 147698 5134
rect 149214 5122 149266 5134
rect 148082 5070 148094 5122
rect 148146 5070 148158 5122
rect 147646 5058 147698 5070
rect 149214 5058 149266 5070
rect 22094 5010 22146 5022
rect 52782 5010 52834 5022
rect 60622 5010 60674 5022
rect 17042 4958 17054 5010
rect 17106 4958 17118 5010
rect 20290 4958 20302 5010
rect 20354 4958 20366 5010
rect 28130 4958 28142 5010
rect 28194 4958 28206 5010
rect 29810 4958 29822 5010
rect 29874 4958 29886 5010
rect 34738 4958 34750 5010
rect 34802 4958 34814 5010
rect 35522 4958 35534 5010
rect 35586 4958 35598 5010
rect 38994 4958 39006 5010
rect 39058 4958 39070 5010
rect 48066 4958 48078 5010
rect 48130 4958 48142 5010
rect 50306 4958 50318 5010
rect 50370 4958 50382 5010
rect 51538 4958 51550 5010
rect 51602 4958 51614 5010
rect 59714 4958 59726 5010
rect 59778 4958 59790 5010
rect 22094 4946 22146 4958
rect 52782 4946 52834 4958
rect 60622 4946 60674 4958
rect 64654 5010 64706 5022
rect 71150 5010 71202 5022
rect 67666 4958 67678 5010
rect 67730 4958 67742 5010
rect 64654 4946 64706 4958
rect 71150 4946 71202 4958
rect 72606 5010 72658 5022
rect 77758 5010 77810 5022
rect 84366 5010 84418 5022
rect 91982 5010 92034 5022
rect 75506 4958 75518 5010
rect 75570 4958 75582 5010
rect 82450 4958 82462 5010
rect 82514 4958 82526 5010
rect 87378 4958 87390 5010
rect 87442 4958 87454 5010
rect 90850 4958 90862 5010
rect 90914 4958 90926 5010
rect 72606 4946 72658 4958
rect 77758 4946 77810 4958
rect 84366 4946 84418 4958
rect 91982 4946 92034 4958
rect 92094 5010 92146 5022
rect 99038 5010 99090 5022
rect 103742 5010 103794 5022
rect 106766 5010 106818 5022
rect 111358 5010 111410 5022
rect 93986 4958 93998 5010
rect 94050 4958 94062 5010
rect 95218 4958 95230 5010
rect 95282 4958 95294 5010
rect 96226 4958 96238 5010
rect 96290 4958 96302 5010
rect 100034 4958 100046 5010
rect 100098 4958 100110 5010
rect 104626 4958 104638 5010
rect 104690 4958 104702 5010
rect 107650 4958 107662 5010
rect 107714 4958 107726 5010
rect 92094 4946 92146 4958
rect 99038 4946 99090 4958
rect 103742 4946 103794 4958
rect 106766 4946 106818 4958
rect 111358 4946 111410 4958
rect 113822 5010 113874 5022
rect 113822 4946 113874 4958
rect 116958 5010 117010 5022
rect 128830 5010 128882 5022
rect 144734 5010 144786 5022
rect 118738 4958 118750 5010
rect 118802 4958 118814 5010
rect 122098 4958 122110 5010
rect 122162 4958 122174 5010
rect 125234 4958 125246 5010
rect 125298 4958 125310 5010
rect 128034 4958 128046 5010
rect 128098 4958 128110 5010
rect 133858 4958 133870 5010
rect 133922 4958 133934 5010
rect 141362 4958 141374 5010
rect 141426 4958 141438 5010
rect 143938 4958 143950 5010
rect 144002 4958 144014 5010
rect 116958 4946 117010 4958
rect 128830 4946 128882 4958
rect 144734 4946 144786 4958
rect 145070 5010 145122 5022
rect 149538 4958 149550 5010
rect 149602 4958 149614 5010
rect 145070 4946 145122 4958
rect 17950 4898 18002 4910
rect 17950 4834 18002 4846
rect 18622 4898 18674 4910
rect 22542 4898 22594 4910
rect 21746 4846 21758 4898
rect 21810 4846 21822 4898
rect 18622 4834 18674 4846
rect 22542 4834 22594 4846
rect 57374 4898 57426 4910
rect 57374 4834 57426 4846
rect 70702 4898 70754 4910
rect 70702 4834 70754 4846
rect 76414 4898 76466 4910
rect 76414 4834 76466 4846
rect 83358 4898 83410 4910
rect 91758 4898 91810 4910
rect 85586 4846 85598 4898
rect 85650 4846 85662 4898
rect 83358 4834 83410 4846
rect 91758 4834 91810 4846
rect 111806 4898 111858 4910
rect 111806 4834 111858 4846
rect 113374 4898 113426 4910
rect 113374 4834 113426 4846
rect 117854 4898 117906 4910
rect 117854 4834 117906 4846
rect 133534 4898 133586 4910
rect 133534 4834 133586 4846
rect 135998 4898 136050 4910
rect 135998 4834 136050 4846
rect 138350 4898 138402 4910
rect 138350 4834 138402 4846
rect 147870 4898 147922 4910
rect 147870 4834 147922 4846
rect 1344 4730 158592 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 81278 4730
rect 81330 4678 81382 4730
rect 81434 4678 81486 4730
rect 81538 4678 111998 4730
rect 112050 4678 112102 4730
rect 112154 4678 112206 4730
rect 112258 4678 142718 4730
rect 142770 4678 142822 4730
rect 142874 4678 142926 4730
rect 142978 4678 158592 4730
rect 1344 4644 158592 4678
rect 19070 4562 19122 4574
rect 19070 4498 19122 4510
rect 23886 4562 23938 4574
rect 23886 4498 23938 4510
rect 25342 4562 25394 4574
rect 25342 4498 25394 4510
rect 26686 4562 26738 4574
rect 26686 4498 26738 4510
rect 30718 4562 30770 4574
rect 39118 4562 39170 4574
rect 38658 4510 38670 4562
rect 38722 4510 38734 4562
rect 30718 4498 30770 4510
rect 39118 4498 39170 4510
rect 39342 4562 39394 4574
rect 39342 4498 39394 4510
rect 42590 4562 42642 4574
rect 42590 4498 42642 4510
rect 48078 4562 48130 4574
rect 48078 4498 48130 4510
rect 48302 4562 48354 4574
rect 48302 4498 48354 4510
rect 50430 4562 50482 4574
rect 50430 4498 50482 4510
rect 56030 4562 56082 4574
rect 68574 4562 68626 4574
rect 64530 4510 64542 4562
rect 64594 4510 64606 4562
rect 56030 4498 56082 4510
rect 68574 4498 68626 4510
rect 72494 4562 72546 4574
rect 72494 4498 72546 4510
rect 72718 4562 72770 4574
rect 72718 4498 72770 4510
rect 76302 4562 76354 4574
rect 76302 4498 76354 4510
rect 76526 4562 76578 4574
rect 76974 4562 77026 4574
rect 76526 4498 76578 4510
rect 76638 4506 76690 4518
rect 13806 4450 13858 4462
rect 16830 4450 16882 4462
rect 15474 4398 15486 4450
rect 15538 4398 15550 4450
rect 13806 4386 13858 4398
rect 16830 4386 16882 4398
rect 18958 4450 19010 4462
rect 23102 4450 23154 4462
rect 21522 4398 21534 4450
rect 21586 4398 21598 4450
rect 18958 4386 19010 4398
rect 23102 4386 23154 4398
rect 23438 4450 23490 4462
rect 23438 4386 23490 4398
rect 23662 4450 23714 4462
rect 23662 4386 23714 4398
rect 24670 4450 24722 4462
rect 37326 4450 37378 4462
rect 39454 4450 39506 4462
rect 47966 4450 48018 4462
rect 29138 4398 29150 4450
rect 29202 4398 29214 4450
rect 32050 4398 32062 4450
rect 32114 4398 32126 4450
rect 34178 4398 34190 4450
rect 34242 4398 34254 4450
rect 38322 4398 38334 4450
rect 38386 4398 38398 4450
rect 46274 4398 46286 4450
rect 46338 4398 46350 4450
rect 24670 4386 24722 4398
rect 37326 4386 37378 4398
rect 39454 4386 39506 4398
rect 47966 4386 48018 4398
rect 49310 4450 49362 4462
rect 56590 4450 56642 4462
rect 49634 4398 49646 4450
rect 49698 4398 49710 4450
rect 53442 4398 53454 4450
rect 53506 4398 53518 4450
rect 53890 4398 53902 4450
rect 53954 4398 53966 4450
rect 49310 4386 49362 4398
rect 56590 4386 56642 4398
rect 56702 4450 56754 4462
rect 56702 4386 56754 4398
rect 56926 4450 56978 4462
rect 65102 4450 65154 4462
rect 57362 4398 57374 4450
rect 57426 4398 57438 4450
rect 61058 4398 61070 4450
rect 61122 4398 61134 4450
rect 63746 4398 63758 4450
rect 63810 4398 63822 4450
rect 56926 4386 56978 4398
rect 65102 4386 65154 4398
rect 67678 4450 67730 4462
rect 76974 4498 77026 4510
rect 86494 4562 86546 4574
rect 86494 4498 86546 4510
rect 87278 4562 87330 4574
rect 87278 4498 87330 4510
rect 87838 4562 87890 4574
rect 87838 4498 87890 4510
rect 90638 4562 90690 4574
rect 110798 4562 110850 4574
rect 105858 4510 105870 4562
rect 105922 4510 105934 4562
rect 90638 4498 90690 4510
rect 110798 4498 110850 4510
rect 113934 4562 113986 4574
rect 113934 4498 113986 4510
rect 115502 4562 115554 4574
rect 132526 4562 132578 4574
rect 122882 4510 122894 4562
rect 122946 4510 122958 4562
rect 115502 4498 115554 4510
rect 132526 4498 132578 4510
rect 142830 4562 142882 4574
rect 142830 4498 142882 4510
rect 149998 4562 150050 4574
rect 149998 4498 150050 4510
rect 69458 4398 69470 4450
rect 69522 4398 69534 4450
rect 73938 4398 73950 4450
rect 74002 4398 74014 4450
rect 76638 4442 76690 4454
rect 101278 4450 101330 4462
rect 110910 4450 110962 4462
rect 79090 4398 79102 4450
rect 79154 4398 79166 4450
rect 82338 4398 82350 4450
rect 82402 4398 82414 4450
rect 83682 4398 83694 4450
rect 83746 4398 83758 4450
rect 89954 4398 89966 4450
rect 90018 4398 90030 4450
rect 92754 4398 92766 4450
rect 92818 4398 92830 4450
rect 94546 4398 94558 4450
rect 94610 4398 94622 4450
rect 99026 4398 99038 4450
rect 99090 4398 99102 4450
rect 101602 4398 101614 4450
rect 101666 4398 101678 4450
rect 104738 4398 104750 4450
rect 104802 4398 104814 4450
rect 67678 4386 67730 4398
rect 101278 4386 101330 4398
rect 110910 4386 110962 4398
rect 113038 4450 113090 4462
rect 113038 4386 113090 4398
rect 115950 4450 116002 4462
rect 121102 4450 121154 4462
rect 119746 4398 119758 4450
rect 119810 4398 119822 4450
rect 115950 4386 116002 4398
rect 121102 4386 121154 4398
rect 121438 4450 121490 4462
rect 126030 4450 126082 4462
rect 122770 4398 122782 4450
rect 122834 4398 122846 4450
rect 121438 4386 121490 4398
rect 126030 4386 126082 4398
rect 127262 4450 127314 4462
rect 135774 4450 135826 4462
rect 141374 4450 141426 4462
rect 129938 4398 129950 4450
rect 130002 4398 130014 4450
rect 131730 4398 131742 4450
rect 131794 4398 131806 4450
rect 136210 4398 136222 4450
rect 136274 4398 136286 4450
rect 137778 4398 137790 4450
rect 137842 4398 137854 4450
rect 144162 4398 144174 4450
rect 144226 4398 144238 4450
rect 148866 4398 148878 4450
rect 148930 4398 148942 4450
rect 149650 4398 149662 4450
rect 149714 4398 149726 4450
rect 127262 4386 127314 4398
rect 135774 4386 135826 4398
rect 141374 4386 141426 4398
rect 13470 4338 13522 4350
rect 24110 4338 24162 4350
rect 25230 4338 25282 4350
rect 15922 4286 15934 4338
rect 15986 4286 15998 4338
rect 16594 4286 16606 4338
rect 16658 4286 16670 4338
rect 17378 4286 17390 4338
rect 17442 4286 17454 4338
rect 22306 4286 22318 4338
rect 22370 4286 22382 4338
rect 22866 4286 22878 4338
rect 22930 4286 22942 4338
rect 24434 4286 24446 4338
rect 24498 4286 24510 4338
rect 13470 4274 13522 4286
rect 24110 4274 24162 4286
rect 25230 4274 25282 4286
rect 25566 4338 25618 4350
rect 25566 4274 25618 4286
rect 25678 4338 25730 4350
rect 33182 4338 33234 4350
rect 41358 4338 41410 4350
rect 29810 4286 29822 4338
rect 29874 4286 29886 4338
rect 34066 4286 34078 4338
rect 34130 4286 34142 4338
rect 36306 4286 36318 4338
rect 36370 4286 36382 4338
rect 38210 4286 38222 4338
rect 38274 4286 38286 4338
rect 40226 4286 40238 4338
rect 40290 4286 40302 4338
rect 41122 4286 41134 4338
rect 41186 4286 41198 4338
rect 25678 4274 25730 4286
rect 33182 4274 33234 4286
rect 41358 4274 41410 4286
rect 41582 4338 41634 4350
rect 48750 4338 48802 4350
rect 43026 4286 43038 4338
rect 43090 4286 43102 4338
rect 41582 4274 41634 4286
rect 48750 4274 48802 4286
rect 51326 4338 51378 4350
rect 64542 4338 64594 4350
rect 51874 4286 51886 4338
rect 51938 4286 51950 4338
rect 55794 4286 55806 4338
rect 55858 4286 55870 4338
rect 61730 4286 61742 4338
rect 61794 4286 61806 4338
rect 51326 4274 51378 4286
rect 64542 4274 64594 4286
rect 66558 4338 66610 4350
rect 72830 4338 72882 4350
rect 86942 4338 86994 4350
rect 68786 4286 68798 4338
rect 68850 4286 68862 4338
rect 73154 4286 73166 4338
rect 73218 4286 73230 4338
rect 82898 4286 82910 4338
rect 82962 4286 82974 4338
rect 86258 4286 86270 4338
rect 86322 4286 86334 4338
rect 66558 4274 66610 4286
rect 72830 4274 72882 4286
rect 86942 4274 86994 4286
rect 87166 4338 87218 4350
rect 87166 4274 87218 4286
rect 87502 4338 87554 4350
rect 109342 4338 109394 4350
rect 110574 4338 110626 4350
rect 98354 4286 98366 4338
rect 98418 4286 98430 4338
rect 105634 4286 105646 4338
rect 105698 4286 105710 4338
rect 106418 4286 106430 4338
rect 106482 4286 106494 4338
rect 109666 4286 109678 4338
rect 109730 4286 109742 4338
rect 87502 4274 87554 4286
rect 109342 4274 109394 4286
rect 110574 4274 110626 4286
rect 112590 4338 112642 4350
rect 117742 4338 117794 4350
rect 124910 4338 124962 4350
rect 115378 4286 115390 4338
rect 115442 4286 115454 4338
rect 117842 4286 117854 4338
rect 117906 4286 117918 4338
rect 124562 4286 124574 4338
rect 124626 4286 124638 4338
rect 112590 4274 112642 4286
rect 117742 4274 117794 4286
rect 124910 4274 124962 4286
rect 127598 4338 127650 4350
rect 127598 4274 127650 4286
rect 127822 4338 127874 4350
rect 141486 4338 141538 4350
rect 132738 4286 132750 4338
rect 132802 4286 132814 4338
rect 135538 4286 135550 4338
rect 135602 4286 135614 4338
rect 137330 4286 137342 4338
rect 137394 4286 137406 4338
rect 127822 4274 127874 4286
rect 141486 4274 141538 4286
rect 141710 4338 141762 4350
rect 141710 4274 141762 4286
rect 141934 4338 141986 4350
rect 141934 4274 141986 4286
rect 142046 4338 142098 4350
rect 143042 4286 143054 4338
rect 143106 4286 143118 4338
rect 142046 4274 142098 4286
rect 13246 4226 13298 4238
rect 13246 4162 13298 4174
rect 15038 4226 15090 4238
rect 26126 4226 26178 4238
rect 30606 4226 30658 4238
rect 33742 4226 33794 4238
rect 41694 4226 41746 4238
rect 71486 4226 71538 4238
rect 112254 4226 112306 4238
rect 18386 4174 18398 4226
rect 18450 4174 18462 4226
rect 19394 4174 19406 4226
rect 19458 4174 19470 4226
rect 27010 4174 27022 4226
rect 27074 4174 27086 4226
rect 31042 4174 31054 4226
rect 31106 4174 31118 4226
rect 35298 4174 35310 4226
rect 35362 4174 35374 4226
rect 39890 4174 39902 4226
rect 39954 4174 39966 4226
rect 42130 4174 42142 4226
rect 42194 4174 42206 4226
rect 43698 4174 43710 4226
rect 43762 4174 43774 4226
rect 45826 4174 45838 4226
rect 45890 4174 45902 4226
rect 47618 4174 47630 4226
rect 47682 4174 47694 4226
rect 55122 4174 55134 4226
rect 55186 4174 55198 4226
rect 58370 4174 58382 4226
rect 58434 4174 58446 4226
rect 58930 4174 58942 4226
rect 58994 4174 59006 4226
rect 62626 4174 62638 4226
rect 62690 4174 62702 4226
rect 76066 4174 76078 4226
rect 76130 4174 76142 4226
rect 80098 4174 80110 4226
rect 80162 4174 80174 4226
rect 85810 4174 85822 4226
rect 85874 4174 85886 4226
rect 93538 4174 93550 4226
rect 93602 4174 93614 4226
rect 102946 4174 102958 4226
rect 103010 4174 103022 4226
rect 103730 4174 103742 4226
rect 103794 4174 103806 4226
rect 109554 4174 109566 4226
rect 109618 4174 109630 4226
rect 15038 4162 15090 4174
rect 26126 4162 26178 4174
rect 30606 4162 30658 4174
rect 33742 4162 33794 4174
rect 41694 4162 41746 4174
rect 71486 4162 71538 4174
rect 112254 4162 112306 4174
rect 115166 4226 115218 4238
rect 121886 4226 121938 4238
rect 117954 4174 117966 4226
rect 118018 4174 118030 4226
rect 120754 4174 120766 4226
rect 120818 4174 120830 4226
rect 115166 4162 115218 4174
rect 121886 4162 121938 4174
rect 122334 4226 122386 4238
rect 135102 4226 135154 4238
rect 139582 4226 139634 4238
rect 130722 4174 130734 4226
rect 130786 4174 130798 4226
rect 138898 4174 138910 4226
rect 138962 4174 138974 4226
rect 122334 4162 122386 4174
rect 135102 4162 135154 4174
rect 139582 4162 139634 4174
rect 143614 4226 143666 4238
rect 146190 4226 146242 4238
rect 145282 4174 145294 4226
rect 145346 4174 145358 4226
rect 143614 4162 143666 4174
rect 146190 4162 146242 4174
rect 147534 4226 147586 4238
rect 147858 4174 147870 4226
rect 147922 4174 147934 4226
rect 147534 4162 147586 4174
rect 15486 4114 15538 4126
rect 15486 4050 15538 4062
rect 96014 4114 96066 4126
rect 96014 4050 96066 4062
rect 107214 4114 107266 4126
rect 109218 4062 109230 4114
rect 109282 4062 109294 4114
rect 118402 4062 118414 4114
rect 118466 4062 118478 4114
rect 107214 4050 107266 4062
rect 1344 3946 158592 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 96638 3946
rect 96690 3894 96742 3946
rect 96794 3894 96846 3946
rect 96898 3894 127358 3946
rect 127410 3894 127462 3946
rect 127514 3894 127566 3946
rect 127618 3894 158078 3946
rect 158130 3894 158182 3946
rect 158234 3894 158286 3946
rect 158338 3894 158592 3946
rect 1344 3860 158592 3894
rect 93214 3778 93266 3790
rect 93214 3714 93266 3726
rect 11342 3666 11394 3678
rect 11342 3602 11394 3614
rect 13358 3666 13410 3678
rect 13358 3602 13410 3614
rect 17054 3666 17106 3678
rect 17054 3602 17106 3614
rect 18510 3666 18562 3678
rect 20974 3666 21026 3678
rect 18722 3614 18734 3666
rect 18786 3614 18798 3666
rect 18510 3602 18562 3614
rect 20974 3602 21026 3614
rect 25454 3666 25506 3678
rect 40798 3666 40850 3678
rect 59054 3666 59106 3678
rect 32162 3614 32174 3666
rect 32226 3614 32238 3666
rect 34290 3614 34302 3666
rect 34354 3614 34366 3666
rect 36754 3614 36766 3666
rect 36818 3614 36830 3666
rect 38882 3614 38894 3666
rect 38946 3614 38958 3666
rect 45490 3614 45502 3666
rect 45554 3614 45566 3666
rect 55010 3614 55022 3666
rect 55074 3614 55086 3666
rect 57138 3614 57150 3666
rect 57202 3614 57214 3666
rect 25454 3602 25506 3614
rect 40798 3602 40850 3614
rect 59054 3602 59106 3614
rect 64878 3666 64930 3678
rect 70478 3666 70530 3678
rect 66434 3614 66446 3666
rect 66498 3614 66510 3666
rect 68562 3614 68574 3666
rect 68626 3614 68638 3666
rect 64878 3602 64930 3614
rect 70478 3602 70530 3614
rect 74846 3666 74898 3678
rect 74846 3602 74898 3614
rect 78990 3666 79042 3678
rect 78990 3602 79042 3614
rect 83022 3666 83074 3678
rect 83022 3602 83074 3614
rect 90190 3666 90242 3678
rect 90190 3602 90242 3614
rect 93102 3666 93154 3678
rect 104750 3666 104802 3678
rect 94098 3614 94110 3666
rect 94162 3614 94174 3666
rect 97906 3614 97918 3666
rect 97970 3614 97982 3666
rect 101938 3614 101950 3666
rect 102002 3614 102014 3666
rect 93102 3602 93154 3614
rect 104750 3602 104802 3614
rect 112926 3666 112978 3678
rect 124574 3666 124626 3678
rect 120978 3614 120990 3666
rect 121042 3614 121054 3666
rect 112926 3602 112978 3614
rect 124574 3602 124626 3614
rect 128382 3666 128434 3678
rect 139806 3666 139858 3678
rect 136098 3614 136110 3666
rect 136162 3614 136174 3666
rect 128382 3602 128434 3614
rect 139806 3602 139858 3614
rect 143614 3666 143666 3678
rect 143614 3602 143666 3614
rect 149774 3666 149826 3678
rect 149774 3602 149826 3614
rect 151566 3666 151618 3678
rect 151566 3602 151618 3614
rect 28702 3554 28754 3566
rect 51214 3554 51266 3566
rect 73502 3554 73554 3566
rect 15250 3502 15262 3554
rect 15314 3502 15326 3554
rect 16258 3502 16270 3554
rect 16322 3502 16334 3554
rect 23314 3502 23326 3554
rect 23378 3502 23390 3554
rect 23762 3502 23774 3554
rect 23826 3502 23838 3554
rect 27794 3502 27806 3554
rect 27858 3502 27870 3554
rect 31154 3502 31166 3554
rect 31218 3502 31230 3554
rect 34962 3502 34974 3554
rect 35026 3502 35038 3554
rect 35970 3502 35982 3554
rect 36034 3502 36046 3554
rect 40002 3502 40014 3554
rect 40066 3502 40078 3554
rect 42914 3502 42926 3554
rect 42978 3502 42990 3554
rect 43698 3502 43710 3554
rect 43762 3502 43774 3554
rect 46834 3502 46846 3554
rect 46898 3502 46910 3554
rect 47618 3502 47630 3554
rect 47682 3502 47694 3554
rect 48514 3502 48526 3554
rect 48578 3502 48590 3554
rect 52098 3502 52110 3554
rect 52162 3502 52174 3554
rect 57810 3502 57822 3554
rect 57874 3502 57886 3554
rect 61394 3502 61406 3554
rect 61458 3502 61470 3554
rect 61954 3502 61966 3554
rect 62018 3502 62030 3554
rect 62850 3502 62862 3554
rect 62914 3502 62926 3554
rect 65874 3502 65886 3554
rect 65938 3502 65950 3554
rect 69234 3502 69246 3554
rect 69298 3502 69310 3554
rect 72370 3502 72382 3554
rect 72434 3502 72446 3554
rect 28702 3490 28754 3502
rect 51214 3490 51266 3502
rect 73502 3490 73554 3502
rect 76526 3554 76578 3566
rect 80782 3554 80834 3566
rect 77186 3502 77198 3554
rect 77250 3502 77262 3554
rect 77970 3502 77982 3554
rect 78034 3502 78046 3554
rect 76526 3490 76578 3502
rect 80782 3490 80834 3502
rect 81118 3554 81170 3566
rect 85486 3554 85538 3566
rect 82002 3502 82014 3554
rect 82066 3502 82078 3554
rect 81118 3490 81170 3502
rect 85486 3490 85538 3502
rect 85822 3554 85874 3566
rect 89630 3554 89682 3566
rect 97246 3554 97298 3566
rect 108670 3554 108722 3566
rect 113262 3554 113314 3566
rect 130398 3554 130450 3566
rect 138238 3554 138290 3566
rect 142046 3554 142098 3566
rect 145854 3554 145906 3566
rect 86034 3502 86046 3554
rect 86098 3502 86110 3554
rect 92306 3502 92318 3554
rect 92370 3502 92382 3554
rect 94994 3502 95006 3554
rect 95058 3502 95070 3554
rect 95218 3502 95230 3554
rect 95282 3502 95294 3554
rect 99698 3502 99710 3554
rect 99762 3502 99774 3554
rect 100930 3502 100942 3554
rect 100994 3502 101006 3554
rect 103954 3502 103966 3554
rect 104018 3502 104030 3554
rect 107538 3502 107550 3554
rect 107602 3502 107614 3554
rect 108994 3502 109006 3554
rect 109058 3502 109070 3554
rect 115266 3502 115278 3554
rect 115330 3502 115342 3554
rect 116162 3502 116174 3554
rect 116226 3502 116238 3554
rect 119074 3502 119086 3554
rect 119138 3502 119150 3554
rect 119746 3502 119758 3554
rect 119810 3502 119822 3554
rect 122882 3502 122894 3554
rect 122946 3502 122958 3554
rect 123554 3502 123566 3554
rect 123618 3502 123630 3554
rect 126690 3502 126702 3554
rect 126754 3502 126766 3554
rect 127362 3502 127374 3554
rect 127426 3502 127438 3554
rect 131170 3502 131182 3554
rect 131234 3502 131246 3554
rect 134306 3502 134318 3554
rect 134370 3502 134382 3554
rect 134978 3502 134990 3554
rect 135042 3502 135054 3554
rect 139234 3502 139246 3554
rect 139298 3502 139310 3554
rect 142594 3502 142606 3554
rect 142658 3502 142670 3554
rect 146514 3502 146526 3554
rect 146578 3502 146590 3554
rect 150546 3502 150558 3554
rect 150610 3502 150622 3554
rect 85822 3490 85874 3502
rect 89630 3490 89682 3502
rect 97246 3490 97298 3502
rect 108670 3490 108722 3502
rect 113262 3490 113314 3502
rect 130398 3490 130450 3502
rect 138238 3490 138290 3502
rect 142046 3490 142098 3502
rect 145854 3490 145906 3502
rect 10558 3442 10610 3454
rect 10558 3378 10610 3390
rect 10782 3442 10834 3454
rect 10782 3378 10834 3390
rect 16046 3442 16098 3454
rect 16046 3378 16098 3390
rect 17502 3442 17554 3454
rect 17502 3378 17554 3390
rect 18062 3442 18114 3454
rect 23998 3442 24050 3454
rect 19730 3390 19742 3442
rect 19794 3390 19806 3442
rect 18062 3378 18114 3390
rect 23998 3378 24050 3390
rect 24558 3442 24610 3454
rect 24558 3378 24610 3390
rect 28366 3442 28418 3454
rect 43934 3442 43986 3454
rect 51550 3442 51602 3454
rect 61742 3442 61794 3454
rect 42690 3390 42702 3442
rect 42754 3390 42766 3442
rect 47394 3390 47406 3442
rect 47458 3390 47470 3442
rect 49634 3390 49646 3442
rect 49698 3390 49710 3442
rect 53554 3390 53566 3442
rect 53618 3390 53630 3442
rect 28366 3378 28418 3390
rect 43934 3378 43986 3390
rect 51550 3378 51602 3390
rect 61742 3378 61794 3390
rect 62638 3442 62690 3454
rect 62638 3378 62690 3390
rect 73166 3442 73218 3454
rect 73166 3378 73218 3390
rect 76078 3442 76130 3454
rect 81006 3442 81058 3454
rect 76962 3390 76974 3442
rect 77026 3390 77038 3442
rect 76078 3378 76130 3390
rect 81006 3378 81058 3390
rect 85598 3442 85650 3454
rect 85598 3378 85650 3390
rect 89294 3442 89346 3454
rect 96910 3442 96962 3454
rect 107326 3442 107378 3454
rect 94322 3390 94334 3442
rect 94386 3390 94398 3442
rect 100706 3390 100718 3442
rect 100770 3390 100782 3442
rect 106866 3390 106878 3442
rect 106930 3390 106942 3442
rect 89294 3378 89346 3390
rect 96910 3378 96962 3390
rect 107326 3378 107378 3390
rect 108334 3442 108386 3454
rect 108334 3378 108386 3390
rect 113710 3442 113762 3454
rect 122670 3442 122722 3454
rect 117618 3390 117630 3442
rect 117682 3390 117694 3442
rect 118850 3390 118862 3442
rect 118914 3390 118926 3442
rect 113710 3378 113762 3390
rect 122670 3378 122722 3390
rect 126478 3442 126530 3454
rect 134094 3442 134146 3454
rect 132738 3390 132750 3442
rect 132802 3390 132814 3442
rect 126478 3378 126530 3390
rect 134094 3378 134146 3390
rect 137902 3442 137954 3454
rect 141698 3390 141710 3442
rect 141762 3390 141774 3442
rect 145506 3390 145518 3442
rect 145570 3390 145582 3442
rect 137902 3378 137954 3390
rect 24894 3330 24946 3342
rect 24894 3266 24946 3278
rect 30606 3330 30658 3342
rect 30606 3266 30658 3278
rect 74286 3330 74338 3342
rect 74286 3266 74338 3278
rect 87054 3330 87106 3342
rect 87054 3266 87106 3278
rect 110014 3330 110066 3342
rect 110014 3266 110066 3278
rect 114606 3330 114658 3342
rect 147534 3330 147586 3342
rect 115042 3278 115054 3330
rect 115106 3278 115118 3330
rect 114606 3266 114658 3278
rect 147534 3266 147586 3278
rect 1344 3162 158592 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 81278 3162
rect 81330 3110 81382 3162
rect 81434 3110 81486 3162
rect 81538 3110 111998 3162
rect 112050 3110 112102 3162
rect 112154 3110 112206 3162
rect 112258 3110 142718 3162
rect 142770 3110 142822 3162
rect 142874 3110 142926 3162
rect 142978 3110 158592 3162
rect 1344 3076 158592 3110
<< via1 >>
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 81278 56422 81330 56474
rect 81382 56422 81434 56474
rect 81486 56422 81538 56474
rect 111998 56422 112050 56474
rect 112102 56422 112154 56474
rect 112206 56422 112258 56474
rect 142718 56422 142770 56474
rect 142822 56422 142874 56474
rect 142926 56422 142978 56474
rect 5070 56254 5122 56306
rect 5854 56254 5906 56306
rect 13470 56254 13522 56306
rect 24894 56254 24946 56306
rect 29710 56254 29762 56306
rect 36318 56254 36370 56306
rect 47742 56254 47794 56306
rect 52558 56254 52610 56306
rect 55358 56254 55410 56306
rect 63982 56254 64034 56306
rect 66782 56254 66834 56306
rect 71598 56254 71650 56306
rect 83022 56254 83074 56306
rect 89630 56254 89682 56306
rect 94446 56254 94498 56306
rect 98254 56254 98306 56306
rect 101054 56254 101106 56306
rect 105870 56254 105922 56306
rect 109678 56254 109730 56306
rect 117294 56254 117346 56306
rect 121102 56254 121154 56306
rect 128718 56254 128770 56306
rect 132526 56254 132578 56306
rect 135326 56254 135378 56306
rect 140142 56254 140194 56306
rect 146750 56254 146802 56306
rect 151566 56254 151618 56306
rect 155374 56254 155426 56306
rect 6190 56142 6242 56194
rect 67118 56142 67170 56194
rect 78206 56142 78258 56194
rect 78542 56142 78594 56194
rect 89966 56142 90018 56194
rect 101390 56142 101442 56194
rect 112478 56142 112530 56194
rect 123902 56142 123954 56194
rect 144510 56142 144562 56194
rect 19854 56030 19906 56082
rect 28702 56030 28754 56082
rect 42702 56030 42754 56082
rect 51550 56030 51602 56082
rect 61742 56030 61794 56082
rect 62974 56030 63026 56082
rect 70590 56030 70642 56082
rect 76974 56030 77026 56082
rect 82014 56030 82066 56082
rect 88398 56030 88450 56082
rect 93438 56030 93490 56082
rect 97582 56030 97634 56082
rect 104862 56030 104914 56082
rect 108670 56030 108722 56082
rect 112702 56030 112754 56082
rect 116286 56030 116338 56082
rect 120094 56030 120146 56082
rect 124126 56030 124178 56082
rect 127710 56030 127762 56082
rect 131518 56030 131570 56082
rect 139246 56030 139298 56082
rect 142942 56030 142994 56082
rect 150782 56030 150834 56082
rect 154590 56030 154642 56082
rect 17502 55918 17554 55970
rect 20974 55918 21026 55970
rect 40350 55918 40402 55970
rect 43822 55918 43874 55970
rect 55918 55918 55970 55970
rect 59390 55918 59442 55970
rect 74622 55918 74674 55970
rect 86046 55918 86098 55970
rect 135774 55918 135826 55970
rect 147198 55918 147250 55970
rect 149774 55918 149826 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 96638 55638 96690 55690
rect 96742 55638 96794 55690
rect 96846 55638 96898 55690
rect 127358 55638 127410 55690
rect 127462 55638 127514 55690
rect 127566 55638 127618 55690
rect 158078 55638 158130 55690
rect 158182 55638 158234 55690
rect 158286 55638 158338 55690
rect 28366 55470 28418 55522
rect 50094 55358 50146 55410
rect 55134 55358 55186 55410
rect 61294 55358 61346 55410
rect 66558 55358 66610 55410
rect 77982 55358 78034 55410
rect 89406 55358 89458 55410
rect 100830 55358 100882 55410
rect 112254 55358 112306 55410
rect 123678 55358 123730 55410
rect 135102 55358 135154 55410
rect 146862 55358 146914 55410
rect 60510 55246 60562 55298
rect 60958 55246 61010 55298
rect 62190 55246 62242 55298
rect 69806 55246 69858 55298
rect 70142 55246 70194 55298
rect 71038 55246 71090 55298
rect 81566 55246 81618 55298
rect 92990 55246 93042 55298
rect 115726 55246 115778 55298
rect 115950 55246 116002 55298
rect 127262 55246 127314 55298
rect 139022 55246 139074 55298
rect 28478 55134 28530 55186
rect 49982 55134 50034 55186
rect 70366 55134 70418 55186
rect 70702 55134 70754 55186
rect 71486 55134 71538 55186
rect 81118 55134 81170 55186
rect 81790 55134 81842 55186
rect 92542 55134 92594 55186
rect 93214 55134 93266 55186
rect 103966 55134 104018 55186
rect 104302 55134 104354 55186
rect 104638 55134 104690 55186
rect 116510 55134 116562 55186
rect 126814 55134 126866 55186
rect 127486 55134 127538 55186
rect 138350 55134 138402 55186
rect 139246 55134 139298 55186
rect 27918 55022 27970 55074
rect 28366 55022 28418 55074
rect 29374 55022 29426 55074
rect 49646 55022 49698 55074
rect 59950 55022 60002 55074
rect 61742 55022 61794 55074
rect 77198 55022 77250 55074
rect 88622 55022 88674 55074
rect 96910 55022 96962 55074
rect 108334 55022 108386 55074
rect 119758 55022 119810 55074
rect 131182 55022 131234 55074
rect 142606 55022 142658 55074
rect 154030 55022 154082 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 81278 54854 81330 54906
rect 81382 54854 81434 54906
rect 81486 54854 81538 54906
rect 111998 54854 112050 54906
rect 112102 54854 112154 54906
rect 112206 54854 112258 54906
rect 142718 54854 142770 54906
rect 142822 54854 142874 54906
rect 142926 54854 142978 54906
rect 116062 54686 116114 54738
rect 115838 54462 115890 54514
rect 116622 54350 116674 54402
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 96638 54070 96690 54122
rect 96742 54070 96794 54122
rect 96846 54070 96898 54122
rect 127358 54070 127410 54122
rect 127462 54070 127514 54122
rect 127566 54070 127618 54122
rect 158078 54070 158130 54122
rect 158182 54070 158234 54122
rect 158286 54070 158338 54122
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 81278 53286 81330 53338
rect 81382 53286 81434 53338
rect 81486 53286 81538 53338
rect 111998 53286 112050 53338
rect 112102 53286 112154 53338
rect 112206 53286 112258 53338
rect 142718 53286 142770 53338
rect 142822 53286 142874 53338
rect 142926 53286 142978 53338
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 96638 52502 96690 52554
rect 96742 52502 96794 52554
rect 96846 52502 96898 52554
rect 127358 52502 127410 52554
rect 127462 52502 127514 52554
rect 127566 52502 127618 52554
rect 158078 52502 158130 52554
rect 158182 52502 158234 52554
rect 158286 52502 158338 52554
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 81278 51718 81330 51770
rect 81382 51718 81434 51770
rect 81486 51718 81538 51770
rect 111998 51718 112050 51770
rect 112102 51718 112154 51770
rect 112206 51718 112258 51770
rect 142718 51718 142770 51770
rect 142822 51718 142874 51770
rect 142926 51718 142978 51770
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 96638 50934 96690 50986
rect 96742 50934 96794 50986
rect 96846 50934 96898 50986
rect 127358 50934 127410 50986
rect 127462 50934 127514 50986
rect 127566 50934 127618 50986
rect 158078 50934 158130 50986
rect 158182 50934 158234 50986
rect 158286 50934 158338 50986
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 81278 50150 81330 50202
rect 81382 50150 81434 50202
rect 81486 50150 81538 50202
rect 111998 50150 112050 50202
rect 112102 50150 112154 50202
rect 112206 50150 112258 50202
rect 142718 50150 142770 50202
rect 142822 50150 142874 50202
rect 142926 50150 142978 50202
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 96638 49366 96690 49418
rect 96742 49366 96794 49418
rect 96846 49366 96898 49418
rect 127358 49366 127410 49418
rect 127462 49366 127514 49418
rect 127566 49366 127618 49418
rect 158078 49366 158130 49418
rect 158182 49366 158234 49418
rect 158286 49366 158338 49418
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 81278 48582 81330 48634
rect 81382 48582 81434 48634
rect 81486 48582 81538 48634
rect 111998 48582 112050 48634
rect 112102 48582 112154 48634
rect 112206 48582 112258 48634
rect 142718 48582 142770 48634
rect 142822 48582 142874 48634
rect 142926 48582 142978 48634
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 96638 47798 96690 47850
rect 96742 47798 96794 47850
rect 96846 47798 96898 47850
rect 127358 47798 127410 47850
rect 127462 47798 127514 47850
rect 127566 47798 127618 47850
rect 158078 47798 158130 47850
rect 158182 47798 158234 47850
rect 158286 47798 158338 47850
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 81278 47014 81330 47066
rect 81382 47014 81434 47066
rect 81486 47014 81538 47066
rect 111998 47014 112050 47066
rect 112102 47014 112154 47066
rect 112206 47014 112258 47066
rect 142718 47014 142770 47066
rect 142822 47014 142874 47066
rect 142926 47014 142978 47066
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 96638 46230 96690 46282
rect 96742 46230 96794 46282
rect 96846 46230 96898 46282
rect 127358 46230 127410 46282
rect 127462 46230 127514 46282
rect 127566 46230 127618 46282
rect 158078 46230 158130 46282
rect 158182 46230 158234 46282
rect 158286 46230 158338 46282
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 81278 45446 81330 45498
rect 81382 45446 81434 45498
rect 81486 45446 81538 45498
rect 111998 45446 112050 45498
rect 112102 45446 112154 45498
rect 112206 45446 112258 45498
rect 142718 45446 142770 45498
rect 142822 45446 142874 45498
rect 142926 45446 142978 45498
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 96638 44662 96690 44714
rect 96742 44662 96794 44714
rect 96846 44662 96898 44714
rect 127358 44662 127410 44714
rect 127462 44662 127514 44714
rect 127566 44662 127618 44714
rect 158078 44662 158130 44714
rect 158182 44662 158234 44714
rect 158286 44662 158338 44714
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 81278 43878 81330 43930
rect 81382 43878 81434 43930
rect 81486 43878 81538 43930
rect 111998 43878 112050 43930
rect 112102 43878 112154 43930
rect 112206 43878 112258 43930
rect 142718 43878 142770 43930
rect 142822 43878 142874 43930
rect 142926 43878 142978 43930
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 96638 43094 96690 43146
rect 96742 43094 96794 43146
rect 96846 43094 96898 43146
rect 127358 43094 127410 43146
rect 127462 43094 127514 43146
rect 127566 43094 127618 43146
rect 158078 43094 158130 43146
rect 158182 43094 158234 43146
rect 158286 43094 158338 43146
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 81278 42310 81330 42362
rect 81382 42310 81434 42362
rect 81486 42310 81538 42362
rect 111998 42310 112050 42362
rect 112102 42310 112154 42362
rect 112206 42310 112258 42362
rect 142718 42310 142770 42362
rect 142822 42310 142874 42362
rect 142926 42310 142978 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 96638 41526 96690 41578
rect 96742 41526 96794 41578
rect 96846 41526 96898 41578
rect 127358 41526 127410 41578
rect 127462 41526 127514 41578
rect 127566 41526 127618 41578
rect 158078 41526 158130 41578
rect 158182 41526 158234 41578
rect 158286 41526 158338 41578
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 81278 40742 81330 40794
rect 81382 40742 81434 40794
rect 81486 40742 81538 40794
rect 111998 40742 112050 40794
rect 112102 40742 112154 40794
rect 112206 40742 112258 40794
rect 142718 40742 142770 40794
rect 142822 40742 142874 40794
rect 142926 40742 142978 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 96638 39958 96690 40010
rect 96742 39958 96794 40010
rect 96846 39958 96898 40010
rect 127358 39958 127410 40010
rect 127462 39958 127514 40010
rect 127566 39958 127618 40010
rect 158078 39958 158130 40010
rect 158182 39958 158234 40010
rect 158286 39958 158338 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 81278 39174 81330 39226
rect 81382 39174 81434 39226
rect 81486 39174 81538 39226
rect 111998 39174 112050 39226
rect 112102 39174 112154 39226
rect 112206 39174 112258 39226
rect 142718 39174 142770 39226
rect 142822 39174 142874 39226
rect 142926 39174 142978 39226
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 96638 38390 96690 38442
rect 96742 38390 96794 38442
rect 96846 38390 96898 38442
rect 127358 38390 127410 38442
rect 127462 38390 127514 38442
rect 127566 38390 127618 38442
rect 158078 38390 158130 38442
rect 158182 38390 158234 38442
rect 158286 38390 158338 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 81278 37606 81330 37658
rect 81382 37606 81434 37658
rect 81486 37606 81538 37658
rect 111998 37606 112050 37658
rect 112102 37606 112154 37658
rect 112206 37606 112258 37658
rect 142718 37606 142770 37658
rect 142822 37606 142874 37658
rect 142926 37606 142978 37658
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 96638 36822 96690 36874
rect 96742 36822 96794 36874
rect 96846 36822 96898 36874
rect 127358 36822 127410 36874
rect 127462 36822 127514 36874
rect 127566 36822 127618 36874
rect 158078 36822 158130 36874
rect 158182 36822 158234 36874
rect 158286 36822 158338 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 81278 36038 81330 36090
rect 81382 36038 81434 36090
rect 81486 36038 81538 36090
rect 111998 36038 112050 36090
rect 112102 36038 112154 36090
rect 112206 36038 112258 36090
rect 142718 36038 142770 36090
rect 142822 36038 142874 36090
rect 142926 36038 142978 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 96638 35254 96690 35306
rect 96742 35254 96794 35306
rect 96846 35254 96898 35306
rect 127358 35254 127410 35306
rect 127462 35254 127514 35306
rect 127566 35254 127618 35306
rect 158078 35254 158130 35306
rect 158182 35254 158234 35306
rect 158286 35254 158338 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 81278 34470 81330 34522
rect 81382 34470 81434 34522
rect 81486 34470 81538 34522
rect 111998 34470 112050 34522
rect 112102 34470 112154 34522
rect 112206 34470 112258 34522
rect 142718 34470 142770 34522
rect 142822 34470 142874 34522
rect 142926 34470 142978 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 96638 33686 96690 33738
rect 96742 33686 96794 33738
rect 96846 33686 96898 33738
rect 127358 33686 127410 33738
rect 127462 33686 127514 33738
rect 127566 33686 127618 33738
rect 158078 33686 158130 33738
rect 158182 33686 158234 33738
rect 158286 33686 158338 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 81278 32902 81330 32954
rect 81382 32902 81434 32954
rect 81486 32902 81538 32954
rect 111998 32902 112050 32954
rect 112102 32902 112154 32954
rect 112206 32902 112258 32954
rect 142718 32902 142770 32954
rect 142822 32902 142874 32954
rect 142926 32902 142978 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 96638 32118 96690 32170
rect 96742 32118 96794 32170
rect 96846 32118 96898 32170
rect 127358 32118 127410 32170
rect 127462 32118 127514 32170
rect 127566 32118 127618 32170
rect 158078 32118 158130 32170
rect 158182 32118 158234 32170
rect 158286 32118 158338 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 81278 31334 81330 31386
rect 81382 31334 81434 31386
rect 81486 31334 81538 31386
rect 111998 31334 112050 31386
rect 112102 31334 112154 31386
rect 112206 31334 112258 31386
rect 142718 31334 142770 31386
rect 142822 31334 142874 31386
rect 142926 31334 142978 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 96638 30550 96690 30602
rect 96742 30550 96794 30602
rect 96846 30550 96898 30602
rect 127358 30550 127410 30602
rect 127462 30550 127514 30602
rect 127566 30550 127618 30602
rect 158078 30550 158130 30602
rect 158182 30550 158234 30602
rect 158286 30550 158338 30602
rect 48862 30270 48914 30322
rect 52110 30270 52162 30322
rect 46062 30158 46114 30210
rect 49310 30158 49362 30210
rect 54798 30158 54850 30210
rect 55246 30158 55298 30210
rect 55806 30158 55858 30210
rect 61070 30158 61122 30210
rect 46734 30046 46786 30098
rect 49982 30046 50034 30098
rect 56254 30046 56306 30098
rect 52782 29934 52834 29986
rect 54126 29934 54178 29986
rect 60510 29934 60562 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 81278 29766 81330 29818
rect 81382 29766 81434 29818
rect 81486 29766 81538 29818
rect 111998 29766 112050 29818
rect 112102 29766 112154 29818
rect 112206 29766 112258 29818
rect 142718 29766 142770 29818
rect 142822 29766 142874 29818
rect 142926 29766 142978 29818
rect 59502 29598 59554 29650
rect 43710 29486 43762 29538
rect 54574 29486 54626 29538
rect 55022 29486 55074 29538
rect 46174 29374 46226 29426
rect 46958 29374 47010 29426
rect 51102 29374 51154 29426
rect 56590 29374 56642 29426
rect 59390 29374 59442 29426
rect 47294 29262 47346 29314
rect 49086 29262 49138 29314
rect 51774 29262 51826 29314
rect 53902 29262 53954 29314
rect 55582 29262 55634 29314
rect 57038 29262 57090 29314
rect 65326 29262 65378 29314
rect 54462 29150 54514 29202
rect 59502 29150 59554 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 96638 28982 96690 29034
rect 96742 28982 96794 29034
rect 96846 28982 96898 29034
rect 127358 28982 127410 29034
rect 127462 28982 127514 29034
rect 127566 28982 127618 29034
rect 158078 28982 158130 29034
rect 158182 28982 158234 29034
rect 158286 28982 158338 29034
rect 32622 28702 32674 28754
rect 48862 28702 48914 28754
rect 56030 28702 56082 28754
rect 56478 28702 56530 28754
rect 56814 28702 56866 28754
rect 73390 28702 73442 28754
rect 29822 28590 29874 28642
rect 49310 28590 49362 28642
rect 49870 28590 49922 28642
rect 50094 28590 50146 28642
rect 50318 28590 50370 28642
rect 50542 28590 50594 28642
rect 53006 28590 53058 28642
rect 53454 28590 53506 28642
rect 53902 28590 53954 28642
rect 55918 28590 55970 28642
rect 57262 28590 57314 28642
rect 57710 28590 57762 28642
rect 58494 28590 58546 28642
rect 59054 28590 59106 28642
rect 59390 28590 59442 28642
rect 60734 28590 60786 28642
rect 62638 28590 62690 28642
rect 62862 28590 62914 28642
rect 63646 28590 63698 28642
rect 69134 28590 69186 28642
rect 72718 28590 72770 28642
rect 30494 28478 30546 28530
rect 44830 28478 44882 28530
rect 45166 28478 45218 28530
rect 49646 28478 49698 28530
rect 55134 28478 55186 28530
rect 33070 28366 33122 28418
rect 49982 28366 50034 28418
rect 51102 28366 51154 28418
rect 54238 28366 54290 28418
rect 57822 28366 57874 28418
rect 58046 28366 58098 28418
rect 59726 28366 59778 28418
rect 65998 28366 66050 28418
rect 66446 28366 66498 28418
rect 69358 28366 69410 28418
rect 70590 28366 70642 28418
rect 71038 28366 71090 28418
rect 72942 28366 72994 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 81278 28198 81330 28250
rect 81382 28198 81434 28250
rect 81486 28198 81538 28250
rect 111998 28198 112050 28250
rect 112102 28198 112154 28250
rect 112206 28198 112258 28250
rect 142718 28198 142770 28250
rect 142822 28198 142874 28250
rect 142926 28198 142978 28250
rect 44158 28030 44210 28082
rect 44718 28030 44770 28082
rect 50878 28030 50930 28082
rect 63982 28030 64034 28082
rect 64766 28030 64818 28082
rect 66110 28030 66162 28082
rect 78654 28030 78706 28082
rect 30942 27918 30994 27970
rect 33182 27918 33234 27970
rect 33854 27918 33906 27970
rect 50990 27918 51042 27970
rect 54014 27918 54066 27970
rect 55246 27918 55298 27970
rect 55582 27918 55634 27970
rect 58046 27918 58098 27970
rect 63758 27918 63810 27970
rect 64654 27918 64706 27970
rect 65326 27918 65378 27970
rect 70926 27918 70978 27970
rect 73726 27918 73778 27970
rect 78206 27918 78258 27970
rect 26910 27806 26962 27858
rect 30718 27806 30770 27858
rect 33406 27806 33458 27858
rect 34190 27806 34242 27858
rect 44606 27806 44658 27858
rect 45278 27806 45330 27858
rect 49422 27806 49474 27858
rect 49646 27806 49698 27858
rect 50318 27806 50370 27858
rect 50542 27806 50594 27858
rect 51214 27806 51266 27858
rect 53230 27806 53282 27858
rect 53342 27806 53394 27858
rect 54350 27806 54402 27858
rect 56926 27806 56978 27858
rect 57374 27806 57426 27858
rect 57710 27806 57762 27858
rect 59278 27806 59330 27858
rect 59502 27806 59554 27858
rect 59838 27806 59890 27858
rect 60622 27806 60674 27858
rect 60846 27806 60898 27858
rect 61070 27806 61122 27858
rect 63646 27806 63698 27858
rect 64542 27806 64594 27858
rect 65102 27806 65154 27858
rect 65662 27806 65714 27858
rect 65886 27806 65938 27858
rect 66222 27806 66274 27858
rect 67118 27806 67170 27858
rect 69694 27806 69746 27858
rect 70366 27806 70418 27858
rect 70702 27806 70754 27858
rect 71150 27806 71202 27858
rect 71486 27806 71538 27858
rect 72718 27806 72770 27858
rect 73950 27806 74002 27858
rect 77646 27806 77698 27858
rect 27582 27694 27634 27746
rect 29710 27694 29762 27746
rect 30158 27694 30210 27746
rect 40350 27694 40402 27746
rect 45054 27694 45106 27746
rect 45726 27694 45778 27746
rect 48974 27694 49026 27746
rect 51774 27694 51826 27746
rect 57150 27694 57202 27746
rect 62078 27694 62130 27746
rect 63310 27694 63362 27746
rect 70814 27694 70866 27746
rect 72270 27694 72322 27746
rect 73166 27694 73218 27746
rect 74286 27694 74338 27746
rect 74734 27694 74786 27746
rect 77758 27694 77810 27746
rect 34190 27582 34242 27634
rect 44830 27582 44882 27634
rect 48862 27582 48914 27634
rect 50766 27582 50818 27634
rect 57822 27582 57874 27634
rect 65662 27582 65714 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 96638 27414 96690 27466
rect 96742 27414 96794 27466
rect 96846 27414 96898 27466
rect 127358 27414 127410 27466
rect 127462 27414 127514 27466
rect 127566 27414 127618 27466
rect 158078 27414 158130 27466
rect 158182 27414 158234 27466
rect 158286 27414 158338 27466
rect 51774 27246 51826 27298
rect 59950 27246 60002 27298
rect 71598 27246 71650 27298
rect 34414 27134 34466 27186
rect 45054 27134 45106 27186
rect 49870 27134 49922 27186
rect 59390 27134 59442 27186
rect 60846 27134 60898 27186
rect 61630 27134 61682 27186
rect 61966 27134 62018 27186
rect 62750 27134 62802 27186
rect 63198 27134 63250 27186
rect 63646 27134 63698 27186
rect 64318 27134 64370 27186
rect 66446 27134 66498 27186
rect 69134 27134 69186 27186
rect 69582 27134 69634 27186
rect 70030 27134 70082 27186
rect 72830 27134 72882 27186
rect 75182 27134 75234 27186
rect 105758 27134 105810 27186
rect 31166 27022 31218 27074
rect 31726 27022 31778 27074
rect 34750 27022 34802 27074
rect 35870 27022 35922 27074
rect 36318 27022 36370 27074
rect 45950 27022 46002 27074
rect 47742 27022 47794 27074
rect 48638 27022 48690 27074
rect 49758 27022 49810 27074
rect 50094 27022 50146 27074
rect 50430 27022 50482 27074
rect 50654 27022 50706 27074
rect 50878 27022 50930 27074
rect 51438 27022 51490 27074
rect 54686 27022 54738 27074
rect 55022 27022 55074 27074
rect 57150 27022 57202 27074
rect 59614 27022 59666 27074
rect 61294 27022 61346 27074
rect 63982 27022 64034 27074
rect 64654 27022 64706 27074
rect 69246 27022 69298 27074
rect 69806 27022 69858 27074
rect 70254 27022 70306 27074
rect 70366 27022 70418 27074
rect 71710 27022 71762 27074
rect 71934 27022 71986 27074
rect 72270 27022 72322 27074
rect 73278 27022 73330 27074
rect 73614 27022 73666 27074
rect 74174 27022 74226 27074
rect 74958 27022 75010 27074
rect 75294 27022 75346 27074
rect 75518 27022 75570 27074
rect 76190 27022 76242 27074
rect 78542 27022 78594 27074
rect 79102 27022 79154 27074
rect 79662 27022 79714 27074
rect 31838 26910 31890 26962
rect 35310 26910 35362 26962
rect 35646 26910 35698 26962
rect 36430 26910 36482 26962
rect 39678 26910 39730 26962
rect 39902 26910 39954 26962
rect 40238 26910 40290 26962
rect 40574 26910 40626 26962
rect 40798 26910 40850 26962
rect 41022 26910 41074 26962
rect 46174 26910 46226 26962
rect 48750 26910 48802 26962
rect 49646 26910 49698 26962
rect 51102 26910 51154 26962
rect 51662 26910 51714 26962
rect 55134 26910 55186 26962
rect 58718 26910 58770 26962
rect 61854 26910 61906 26962
rect 65662 26910 65714 26962
rect 67566 26910 67618 26962
rect 67678 26910 67730 26962
rect 67902 26910 67954 26962
rect 68462 26910 68514 26962
rect 71262 26910 71314 26962
rect 73726 26910 73778 26962
rect 73950 26910 74002 26962
rect 26350 26798 26402 26850
rect 40014 26798 40066 26850
rect 40686 26798 40738 26850
rect 50542 26798 50594 26850
rect 54350 26798 54402 26850
rect 55582 26798 55634 26850
rect 64206 26798 64258 26850
rect 67006 26798 67058 26850
rect 72158 26798 72210 26850
rect 74286 26798 74338 26850
rect 74510 26798 74562 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 81278 26630 81330 26682
rect 81382 26630 81434 26682
rect 81486 26630 81538 26682
rect 111998 26630 112050 26682
rect 112102 26630 112154 26682
rect 112206 26630 112258 26682
rect 142718 26630 142770 26682
rect 142822 26630 142874 26682
rect 142926 26630 142978 26682
rect 24222 26462 24274 26514
rect 25790 26462 25842 26514
rect 26014 26462 26066 26514
rect 26686 26462 26738 26514
rect 27134 26462 27186 26514
rect 31726 26462 31778 26514
rect 41246 26462 41298 26514
rect 41694 26462 41746 26514
rect 41918 26462 41970 26514
rect 46062 26462 46114 26514
rect 47854 26462 47906 26514
rect 48862 26462 48914 26514
rect 50206 26462 50258 26514
rect 51998 26462 52050 26514
rect 64430 26462 64482 26514
rect 65438 26462 65490 26514
rect 71710 26462 71762 26514
rect 72494 26462 72546 26514
rect 73278 26462 73330 26514
rect 75294 26462 75346 26514
rect 75406 26462 75458 26514
rect 107102 26462 107154 26514
rect 24446 26350 24498 26402
rect 24558 26350 24610 26402
rect 30494 26350 30546 26402
rect 32062 26350 32114 26402
rect 36542 26350 36594 26402
rect 38334 26350 38386 26402
rect 38446 26350 38498 26402
rect 39454 26350 39506 26402
rect 42030 26350 42082 26402
rect 42590 26350 42642 26402
rect 43262 26350 43314 26402
rect 43598 26350 43650 26402
rect 48078 26350 48130 26402
rect 49646 26350 49698 26402
rect 49870 26350 49922 26402
rect 50766 26350 50818 26402
rect 50990 26350 51042 26402
rect 51886 26350 51938 26402
rect 52782 26350 52834 26402
rect 53118 26350 53170 26402
rect 55918 26350 55970 26402
rect 56926 26350 56978 26402
rect 58158 26350 58210 26402
rect 63646 26350 63698 26402
rect 68350 26350 68402 26402
rect 70142 26350 70194 26402
rect 72270 26350 72322 26402
rect 72718 26350 72770 26402
rect 73054 26350 73106 26402
rect 73950 26350 74002 26402
rect 75742 26350 75794 26402
rect 105534 26350 105586 26402
rect 106542 26350 106594 26402
rect 24782 26238 24834 26290
rect 25342 26238 25394 26290
rect 25566 26238 25618 26290
rect 30270 26238 30322 26290
rect 30942 26238 30994 26290
rect 31390 26238 31442 26290
rect 35534 26238 35586 26290
rect 35758 26238 35810 26290
rect 36206 26238 36258 26290
rect 39006 26238 39058 26290
rect 39118 26238 39170 26290
rect 39790 26238 39842 26290
rect 40014 26238 40066 26290
rect 40798 26238 40850 26290
rect 41470 26238 41522 26290
rect 42926 26238 42978 26290
rect 44270 26238 44322 26290
rect 44494 26238 44546 26290
rect 45502 26238 45554 26290
rect 48190 26238 48242 26290
rect 48974 26238 49026 26290
rect 50318 26238 50370 26290
rect 50878 26238 50930 26290
rect 54014 26238 54066 26290
rect 54462 26238 54514 26290
rect 55694 26238 55746 26290
rect 56030 26238 56082 26290
rect 57150 26238 57202 26290
rect 57710 26238 57762 26290
rect 59390 26238 59442 26290
rect 60510 26238 60562 26290
rect 62414 26238 62466 26290
rect 63198 26238 63250 26290
rect 63758 26238 63810 26290
rect 67454 26238 67506 26290
rect 67678 26238 67730 26290
rect 70590 26238 70642 26290
rect 72830 26238 72882 26290
rect 73614 26238 73666 26290
rect 73838 26238 73890 26290
rect 74734 26238 74786 26290
rect 75518 26238 75570 26290
rect 77198 26238 77250 26290
rect 77758 26238 77810 26290
rect 86942 26238 86994 26290
rect 104974 26238 105026 26290
rect 105982 26238 106034 26290
rect 25790 26126 25842 26178
rect 35646 26126 35698 26178
rect 36654 26126 36706 26178
rect 37998 26126 38050 26178
rect 39342 26126 39394 26178
rect 41358 26126 41410 26178
rect 45390 26126 45442 26178
rect 46510 26126 46562 26178
rect 53790 26126 53842 26178
rect 59950 26126 60002 26178
rect 60958 26126 61010 26178
rect 61518 26126 61570 26178
rect 64990 26126 65042 26178
rect 67790 26126 67842 26178
rect 68910 26126 68962 26178
rect 74174 26126 74226 26178
rect 76862 26126 76914 26178
rect 86158 26126 86210 26178
rect 86606 26126 86658 26178
rect 104526 26126 104578 26178
rect 104862 26126 104914 26178
rect 107550 26126 107602 26178
rect 30830 26014 30882 26066
rect 31166 26014 31218 26066
rect 36766 26014 36818 26066
rect 38446 26014 38498 26066
rect 40350 26014 40402 26066
rect 44830 26014 44882 26066
rect 45166 26014 45218 26066
rect 45726 26014 45778 26066
rect 46062 26014 46114 26066
rect 48862 26014 48914 26066
rect 52110 26014 52162 26066
rect 54126 26014 54178 26066
rect 73390 26014 73442 26066
rect 106430 26014 106482 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 96638 25846 96690 25898
rect 96742 25846 96794 25898
rect 96846 25846 96898 25898
rect 127358 25846 127410 25898
rect 127462 25846 127514 25898
rect 127566 25846 127618 25898
rect 158078 25846 158130 25898
rect 158182 25846 158234 25898
rect 158286 25846 158338 25898
rect 35198 25678 35250 25730
rect 35534 25678 35586 25730
rect 36318 25678 36370 25730
rect 37438 25678 37490 25730
rect 37550 25678 37602 25730
rect 37774 25678 37826 25730
rect 62190 25678 62242 25730
rect 31054 25566 31106 25618
rect 34638 25566 34690 25618
rect 39006 25566 39058 25618
rect 43486 25566 43538 25618
rect 45838 25566 45890 25618
rect 48078 25566 48130 25618
rect 48638 25566 48690 25618
rect 48974 25566 49026 25618
rect 50878 25566 50930 25618
rect 53118 25566 53170 25618
rect 55918 25566 55970 25618
rect 61182 25566 61234 25618
rect 62638 25566 62690 25618
rect 69918 25566 69970 25618
rect 71598 25566 71650 25618
rect 87278 25566 87330 25618
rect 90302 25566 90354 25618
rect 101838 25566 101890 25618
rect 105534 25566 105586 25618
rect 106766 25566 106818 25618
rect 108670 25566 108722 25618
rect 23438 25454 23490 25506
rect 25790 25454 25842 25506
rect 26574 25454 26626 25506
rect 31502 25454 31554 25506
rect 31950 25454 32002 25506
rect 34862 25454 34914 25506
rect 35758 25454 35810 25506
rect 36094 25454 36146 25506
rect 38894 25454 38946 25506
rect 39566 25454 39618 25506
rect 40014 25454 40066 25506
rect 41246 25454 41298 25506
rect 41694 25454 41746 25506
rect 43934 25454 43986 25506
rect 44718 25454 44770 25506
rect 45390 25454 45442 25506
rect 47294 25454 47346 25506
rect 47742 25454 47794 25506
rect 48862 25454 48914 25506
rect 49086 25454 49138 25506
rect 49422 25454 49474 25506
rect 50094 25454 50146 25506
rect 50542 25454 50594 25506
rect 50766 25454 50818 25506
rect 51774 25454 51826 25506
rect 53006 25454 53058 25506
rect 53342 25454 53394 25506
rect 53790 25454 53842 25506
rect 57598 25454 57650 25506
rect 58046 25454 58098 25506
rect 58494 25454 58546 25506
rect 59054 25454 59106 25506
rect 59502 25454 59554 25506
rect 61854 25454 61906 25506
rect 65550 25454 65602 25506
rect 68910 25454 68962 25506
rect 69470 25454 69522 25506
rect 70478 25454 70530 25506
rect 70702 25454 70754 25506
rect 70814 25454 70866 25506
rect 71150 25454 71202 25506
rect 72046 25454 72098 25506
rect 72718 25454 72770 25506
rect 74734 25454 74786 25506
rect 77310 25454 77362 25506
rect 78094 25454 78146 25506
rect 87614 25454 87666 25506
rect 88174 25454 88226 25506
rect 88958 25454 89010 25506
rect 89742 25454 89794 25506
rect 100494 25454 100546 25506
rect 100942 25454 100994 25506
rect 106094 25454 106146 25506
rect 106542 25454 106594 25506
rect 107662 25454 107714 25506
rect 33966 25342 34018 25394
rect 34302 25342 34354 25394
rect 38558 25342 38610 25394
rect 39342 25342 39394 25394
rect 40462 25342 40514 25394
rect 43598 25342 43650 25394
rect 43822 25342 43874 25394
rect 45166 25342 45218 25394
rect 50318 25342 50370 25394
rect 53902 25342 53954 25394
rect 54462 25342 54514 25394
rect 57150 25342 57202 25394
rect 58830 25342 58882 25394
rect 61630 25342 61682 25394
rect 64766 25342 64818 25394
rect 69918 25342 69970 25394
rect 72606 25342 72658 25394
rect 74846 25342 74898 25394
rect 89854 25342 89906 25394
rect 101390 25342 101442 25394
rect 106990 25342 107042 25394
rect 108222 25342 108274 25394
rect 26910 25230 26962 25282
rect 33630 25230 33682 25282
rect 36430 25230 36482 25282
rect 37438 25230 37490 25282
rect 38222 25230 38274 25282
rect 38446 25230 38498 25282
rect 40126 25230 40178 25282
rect 40238 25230 40290 25282
rect 41022 25230 41074 25282
rect 41134 25230 41186 25282
rect 45054 25230 45106 25282
rect 46398 25230 46450 25282
rect 51326 25230 51378 25282
rect 54238 25230 54290 25282
rect 56254 25230 56306 25282
rect 60734 25230 60786 25282
rect 70590 25230 70642 25282
rect 80446 25230 80498 25282
rect 80894 25230 80946 25282
rect 89518 25230 89570 25282
rect 100830 25230 100882 25282
rect 107886 25230 107938 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 81278 25062 81330 25114
rect 81382 25062 81434 25114
rect 81486 25062 81538 25114
rect 111998 25062 112050 25114
rect 112102 25062 112154 25114
rect 112206 25062 112258 25114
rect 142718 25062 142770 25114
rect 142822 25062 142874 25114
rect 142926 25062 142978 25114
rect 23438 24894 23490 24946
rect 31390 24894 31442 24946
rect 36766 24894 36818 24946
rect 37438 24894 37490 24946
rect 39006 24894 39058 24946
rect 43262 24894 43314 24946
rect 46398 24894 46450 24946
rect 46622 24894 46674 24946
rect 49198 24894 49250 24946
rect 52222 24894 52274 24946
rect 55806 24894 55858 24946
rect 56814 24894 56866 24946
rect 62862 24894 62914 24946
rect 68910 24894 68962 24946
rect 69470 24894 69522 24946
rect 69582 24894 69634 24946
rect 69806 24894 69858 24946
rect 70590 24894 70642 24946
rect 70926 24894 70978 24946
rect 76526 24894 76578 24946
rect 78430 24894 78482 24946
rect 80782 24894 80834 24946
rect 107326 24894 107378 24946
rect 24558 24782 24610 24834
rect 31278 24782 31330 24834
rect 35310 24782 35362 24834
rect 43374 24782 43426 24834
rect 50654 24782 50706 24834
rect 55246 24782 55298 24834
rect 55918 24782 55970 24834
rect 56030 24782 56082 24834
rect 57038 24782 57090 24834
rect 57934 24782 57986 24834
rect 58270 24782 58322 24834
rect 64766 24782 64818 24834
rect 68686 24782 68738 24834
rect 70030 24782 70082 24834
rect 71150 24782 71202 24834
rect 71262 24782 71314 24834
rect 71710 24782 71762 24834
rect 74846 24782 74898 24834
rect 76862 24782 76914 24834
rect 81118 24782 81170 24834
rect 24446 24670 24498 24722
rect 27246 24670 27298 24722
rect 31950 24670 32002 24722
rect 32622 24670 32674 24722
rect 34750 24670 34802 24722
rect 35534 24670 35586 24722
rect 35870 24670 35922 24722
rect 36094 24670 36146 24722
rect 43038 24670 43090 24722
rect 44046 24670 44098 24722
rect 44494 24670 44546 24722
rect 45054 24670 45106 24722
rect 46958 24670 47010 24722
rect 49422 24670 49474 24722
rect 50430 24670 50482 24722
rect 51102 24670 51154 24722
rect 55022 24670 55074 24722
rect 55358 24670 55410 24722
rect 56478 24670 56530 24722
rect 57710 24670 57762 24722
rect 58494 24670 58546 24722
rect 59502 24670 59554 24722
rect 64430 24670 64482 24722
rect 67566 24670 67618 24722
rect 68014 24670 68066 24722
rect 68350 24670 68402 24722
rect 70366 24670 70418 24722
rect 72718 24670 72770 24722
rect 73838 24670 73890 24722
rect 74734 24670 74786 24722
rect 75630 24670 75682 24722
rect 78206 24670 78258 24722
rect 78766 24670 78818 24722
rect 83806 24670 83858 24722
rect 84366 24670 84418 24722
rect 27918 24558 27970 24610
rect 30046 24558 30098 24610
rect 30494 24558 30546 24610
rect 31726 24558 31778 24610
rect 35422 24558 35474 24610
rect 46510 24558 46562 24610
rect 49870 24558 49922 24610
rect 50542 24558 50594 24610
rect 51662 24558 51714 24610
rect 51998 24558 52050 24610
rect 52782 24558 52834 24610
rect 57038 24558 57090 24610
rect 59166 24558 59218 24610
rect 62414 24558 62466 24610
rect 69470 24558 69522 24610
rect 70702 24558 70754 24610
rect 72382 24558 72434 24610
rect 74286 24558 74338 24610
rect 75294 24558 75346 24610
rect 78318 24558 78370 24610
rect 81454 24558 81506 24610
rect 84926 24558 84978 24610
rect 23774 24446 23826 24498
rect 32174 24446 32226 24498
rect 34974 24446 35026 24498
rect 36318 24446 36370 24498
rect 37102 24446 37154 24498
rect 37326 24446 37378 24498
rect 37438 24446 37490 24498
rect 43822 24446 43874 24498
rect 44494 24446 44546 24498
rect 44606 24446 44658 24498
rect 49086 24446 49138 24498
rect 50878 24446 50930 24498
rect 51550 24446 51602 24498
rect 52558 24446 52610 24498
rect 57374 24446 57426 24498
rect 62414 24446 62466 24498
rect 62974 24446 63026 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 96638 24278 96690 24330
rect 96742 24278 96794 24330
rect 96846 24278 96898 24330
rect 127358 24278 127410 24330
rect 127462 24278 127514 24330
rect 127566 24278 127618 24330
rect 158078 24278 158130 24330
rect 158182 24278 158234 24330
rect 158286 24278 158338 24330
rect 27358 24110 27410 24162
rect 46958 24110 47010 24162
rect 50430 24110 50482 24162
rect 53566 24110 53618 24162
rect 27806 23998 27858 24050
rect 33966 23998 34018 24050
rect 43598 23998 43650 24050
rect 48638 23998 48690 24050
rect 50878 23998 50930 24050
rect 52782 23998 52834 24050
rect 58606 23998 58658 24050
rect 64430 23998 64482 24050
rect 67790 23998 67842 24050
rect 69246 23998 69298 24050
rect 73054 23998 73106 24050
rect 31166 23886 31218 23938
rect 34862 23886 34914 23938
rect 35310 23886 35362 23938
rect 35534 23886 35586 23938
rect 39342 23886 39394 23938
rect 39566 23886 39618 23938
rect 40014 23886 40066 23938
rect 43150 23886 43202 23938
rect 45950 23886 46002 23938
rect 46734 23886 46786 23938
rect 47182 23886 47234 23938
rect 47294 23886 47346 23938
rect 47854 23886 47906 23938
rect 50206 23886 50258 23938
rect 50766 23886 50818 23938
rect 51102 23886 51154 23938
rect 51550 23886 51602 23938
rect 51774 23886 51826 23938
rect 52222 23886 52274 23938
rect 54238 23886 54290 23938
rect 54686 23886 54738 23938
rect 57598 23886 57650 23938
rect 58158 23886 58210 23938
rect 64654 23886 64706 23938
rect 65438 23886 65490 23938
rect 68910 23886 68962 23938
rect 73614 23886 73666 23938
rect 74510 23886 74562 23938
rect 74958 23886 75010 23938
rect 75630 23886 75682 23938
rect 76750 23886 76802 23938
rect 78542 23886 78594 23938
rect 86830 23886 86882 23938
rect 27470 23774 27522 23826
rect 28142 23774 28194 23826
rect 28254 23774 28306 23826
rect 28366 23774 28418 23826
rect 31838 23774 31890 23826
rect 40462 23774 40514 23826
rect 45390 23774 45442 23826
rect 45502 23774 45554 23826
rect 46062 23774 46114 23826
rect 46286 23774 46338 23826
rect 54798 23774 54850 23826
rect 60958 23774 61010 23826
rect 68798 23774 68850 23826
rect 69358 23774 69410 23826
rect 74174 23774 74226 23826
rect 80334 23774 80386 23826
rect 27022 23662 27074 23714
rect 27246 23662 27298 23714
rect 28590 23662 28642 23714
rect 34414 23662 34466 23714
rect 35086 23662 35138 23714
rect 39454 23662 39506 23714
rect 42814 23662 42866 23714
rect 45726 23662 45778 23714
rect 47406 23662 47458 23714
rect 48190 23662 48242 23714
rect 50878 23662 50930 23714
rect 51662 23662 51714 23714
rect 53678 23662 53730 23714
rect 53902 23662 53954 23714
rect 54910 23662 54962 23714
rect 59390 23662 59442 23714
rect 61070 23662 61122 23714
rect 61294 23662 61346 23714
rect 68574 23662 68626 23714
rect 75070 23662 75122 23714
rect 76526 23662 76578 23714
rect 86606 23662 86658 23714
rect 92654 23662 92706 23714
rect 93214 23662 93266 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 81278 23494 81330 23546
rect 81382 23494 81434 23546
rect 81486 23494 81538 23546
rect 111998 23494 112050 23546
rect 112102 23494 112154 23546
rect 112206 23494 112258 23546
rect 142718 23494 142770 23546
rect 142822 23494 142874 23546
rect 142926 23494 142978 23546
rect 25342 23326 25394 23378
rect 27806 23326 27858 23378
rect 38334 23326 38386 23378
rect 42030 23326 42082 23378
rect 43374 23326 43426 23378
rect 43710 23326 43762 23378
rect 44606 23326 44658 23378
rect 45054 23326 45106 23378
rect 45166 23326 45218 23378
rect 50878 23326 50930 23378
rect 51326 23326 51378 23378
rect 51550 23326 51602 23378
rect 78654 23326 78706 23378
rect 81566 23326 81618 23378
rect 82574 23326 82626 23378
rect 33518 23214 33570 23266
rect 34078 23214 34130 23266
rect 41022 23214 41074 23266
rect 42142 23214 42194 23266
rect 42366 23214 42418 23266
rect 44158 23214 44210 23266
rect 46398 23214 46450 23266
rect 46958 23214 47010 23266
rect 53678 23214 53730 23266
rect 53790 23214 53842 23266
rect 54686 23214 54738 23266
rect 57822 23214 57874 23266
rect 58382 23214 58434 23266
rect 59054 23214 59106 23266
rect 64654 23214 64706 23266
rect 65550 23214 65602 23266
rect 65774 23214 65826 23266
rect 80222 23214 80274 23266
rect 80894 23214 80946 23266
rect 81790 23214 81842 23266
rect 86382 23214 86434 23266
rect 93326 23214 93378 23266
rect 21870 23102 21922 23154
rect 25454 23102 25506 23154
rect 27694 23102 27746 23154
rect 33294 23102 33346 23154
rect 33630 23102 33682 23154
rect 33966 23102 34018 23154
rect 38558 23102 38610 23154
rect 40798 23102 40850 23154
rect 41134 23102 41186 23154
rect 41470 23102 41522 23154
rect 41806 23102 41858 23154
rect 43486 23102 43538 23154
rect 43934 23102 43986 23154
rect 45278 23102 45330 23154
rect 45614 23102 45666 23154
rect 46286 23102 46338 23154
rect 46622 23102 46674 23154
rect 47182 23102 47234 23154
rect 47742 23102 47794 23154
rect 49870 23102 49922 23154
rect 50094 23102 50146 23154
rect 50318 23102 50370 23154
rect 50766 23102 50818 23154
rect 50990 23102 51042 23154
rect 52782 23102 52834 23154
rect 52894 23102 52946 23154
rect 53118 23102 53170 23154
rect 53342 23102 53394 23154
rect 54014 23102 54066 23154
rect 55022 23102 55074 23154
rect 55694 23102 55746 23154
rect 56814 23102 56866 23154
rect 56926 23102 56978 23154
rect 58606 23102 58658 23154
rect 58830 23102 58882 23154
rect 59838 23102 59890 23154
rect 60286 23102 60338 23154
rect 72494 23102 72546 23154
rect 73054 23102 73106 23154
rect 75742 23102 75794 23154
rect 76078 23102 76130 23154
rect 76302 23102 76354 23154
rect 78430 23102 78482 23154
rect 78878 23102 78930 23154
rect 78990 23102 79042 23154
rect 80670 23102 80722 23154
rect 81118 23102 81170 23154
rect 82126 23102 82178 23154
rect 82462 23102 82514 23154
rect 82686 23102 82738 23154
rect 82910 23102 82962 23154
rect 83358 23102 83410 23154
rect 83582 23102 83634 23154
rect 86718 23102 86770 23154
rect 86942 23102 86994 23154
rect 89742 23102 89794 23154
rect 90302 23102 90354 23154
rect 92878 23102 92930 23154
rect 93550 23102 93602 23154
rect 22542 22990 22594 23042
rect 24670 22990 24722 23042
rect 25902 22990 25954 23042
rect 42590 22990 42642 23042
rect 49086 22990 49138 23042
rect 49534 22990 49586 23042
rect 50542 22990 50594 23042
rect 52334 22990 52386 23042
rect 53006 22990 53058 23042
rect 54350 22990 54402 23042
rect 55358 22990 55410 23042
rect 56590 22990 56642 23042
rect 59166 22990 59218 23042
rect 60958 22990 61010 23042
rect 63086 22990 63138 23042
rect 63870 22990 63922 23042
rect 64766 22990 64818 23042
rect 65438 22990 65490 23042
rect 75406 22990 75458 23042
rect 76190 22990 76242 23042
rect 79550 22990 79602 23042
rect 81678 22990 81730 23042
rect 83134 22990 83186 23042
rect 84030 22990 84082 23042
rect 84478 22990 84530 23042
rect 86494 22990 86546 23042
rect 87390 22990 87442 23042
rect 92654 22990 92706 23042
rect 93102 22990 93154 23042
rect 25342 22878 25394 22930
rect 27806 22878 27858 22930
rect 34078 22878 34130 22930
rect 51662 22878 51714 22930
rect 64430 22878 64482 22930
rect 80110 22878 80162 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 96638 22710 96690 22762
rect 96742 22710 96794 22762
rect 96846 22710 96898 22762
rect 127358 22710 127410 22762
rect 127462 22710 127514 22762
rect 127566 22710 127618 22762
rect 158078 22710 158130 22762
rect 158182 22710 158234 22762
rect 158286 22710 158338 22762
rect 51326 22542 51378 22594
rect 23326 22430 23378 22482
rect 32734 22430 32786 22482
rect 36430 22430 36482 22482
rect 36990 22430 37042 22482
rect 40350 22430 40402 22482
rect 42702 22430 42754 22482
rect 47070 22430 47122 22482
rect 51438 22430 51490 22482
rect 52222 22430 52274 22482
rect 57038 22430 57090 22482
rect 60622 22430 60674 22482
rect 68350 22430 68402 22482
rect 74622 22430 74674 22482
rect 75630 22430 75682 22482
rect 79102 22430 79154 22482
rect 84142 22430 84194 22482
rect 85262 22430 85314 22482
rect 90750 22430 90802 22482
rect 91982 22430 92034 22482
rect 29374 22318 29426 22370
rect 32510 22318 32562 22370
rect 32958 22318 33010 22370
rect 33630 22318 33682 22370
rect 39790 22318 39842 22370
rect 42590 22318 42642 22370
rect 43710 22318 43762 22370
rect 45054 22318 45106 22370
rect 50990 22318 51042 22370
rect 52670 22318 52722 22370
rect 60062 22318 60114 22370
rect 60398 22318 60450 22370
rect 60846 22318 60898 22370
rect 60958 22318 61010 22370
rect 71262 22318 71314 22370
rect 74734 22318 74786 22370
rect 75182 22318 75234 22370
rect 82910 22318 82962 22370
rect 83470 22318 83522 22370
rect 85486 22318 85538 22370
rect 86270 22318 86322 22370
rect 90526 22318 90578 22370
rect 91198 22318 91250 22370
rect 92542 22318 92594 22370
rect 95342 22318 95394 22370
rect 96126 22318 96178 22370
rect 99822 22318 99874 22370
rect 23662 22206 23714 22258
rect 23774 22206 23826 22258
rect 23886 22206 23938 22258
rect 28030 22206 28082 22258
rect 28142 22206 28194 22258
rect 29038 22206 29090 22258
rect 33182 22206 33234 22258
rect 34302 22206 34354 22258
rect 39118 22206 39170 22258
rect 43150 22206 43202 22258
rect 43486 22206 43538 22258
rect 51550 22206 51602 22258
rect 58270 22206 58322 22258
rect 59726 22206 59778 22258
rect 59838 22206 59890 22258
rect 70478 22206 70530 22258
rect 90302 22206 90354 22258
rect 90974 22206 91026 22258
rect 103518 22206 103570 22258
rect 24110 22094 24162 22146
rect 27694 22094 27746 22146
rect 27806 22094 27858 22146
rect 27918 22094 27970 22146
rect 29262 22094 29314 22146
rect 29822 22094 29874 22146
rect 42366 22094 42418 22146
rect 42814 22094 42866 22146
rect 43374 22094 43426 22146
rect 45390 22094 45442 22146
rect 58606 22094 58658 22146
rect 59390 22094 59442 22146
rect 65102 22094 65154 22146
rect 71710 22094 71762 22146
rect 74510 22094 74562 22146
rect 78990 22094 79042 22146
rect 80446 22094 80498 22146
rect 88622 22094 88674 22146
rect 91870 22094 91922 22146
rect 92094 22094 92146 22146
rect 92990 22094 93042 22146
rect 96462 22094 96514 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 81278 21926 81330 21978
rect 81382 21926 81434 21978
rect 81486 21926 81538 21978
rect 111998 21926 112050 21978
rect 112102 21926 112154 21978
rect 112206 21926 112258 21978
rect 142718 21926 142770 21978
rect 142822 21926 142874 21978
rect 142926 21926 142978 21978
rect 26014 21758 26066 21810
rect 43486 21758 43538 21810
rect 47406 21758 47458 21810
rect 47742 21758 47794 21810
rect 47966 21758 48018 21810
rect 49310 21758 49362 21810
rect 50318 21758 50370 21810
rect 52894 21758 52946 21810
rect 53118 21758 53170 21810
rect 55134 21758 55186 21810
rect 57150 21758 57202 21810
rect 59614 21758 59666 21810
rect 60846 21758 60898 21810
rect 80222 21758 80274 21810
rect 82014 21758 82066 21810
rect 82126 21758 82178 21810
rect 86494 21758 86546 21810
rect 86830 21758 86882 21810
rect 88398 21758 88450 21810
rect 93886 21758 93938 21810
rect 98030 21758 98082 21810
rect 24446 21646 24498 21698
rect 27470 21646 27522 21698
rect 31614 21646 31666 21698
rect 33406 21646 33458 21698
rect 34414 21646 34466 21698
rect 42702 21646 42754 21698
rect 42926 21646 42978 21698
rect 46622 21646 46674 21698
rect 47294 21646 47346 21698
rect 47630 21646 47682 21698
rect 51102 21646 51154 21698
rect 55806 21646 55858 21698
rect 60062 21646 60114 21698
rect 21086 21534 21138 21586
rect 24222 21534 24274 21586
rect 24558 21534 24610 21586
rect 26350 21534 26402 21586
rect 26686 21534 26738 21586
rect 31390 21534 31442 21586
rect 31726 21534 31778 21586
rect 33742 21534 33794 21586
rect 34078 21534 34130 21586
rect 41694 21534 41746 21586
rect 42030 21534 42082 21586
rect 46286 21534 46338 21586
rect 50542 21534 50594 21586
rect 50990 21534 51042 21586
rect 52782 21590 52834 21642
rect 73838 21646 73890 21698
rect 86158 21646 86210 21698
rect 87166 21646 87218 21698
rect 88510 21646 88562 21698
rect 93774 21646 93826 21698
rect 97470 21646 97522 21698
rect 98142 21646 98194 21698
rect 109006 21646 109058 21698
rect 51214 21534 51266 21586
rect 51662 21534 51714 21586
rect 52334 21534 52386 21586
rect 54014 21534 54066 21586
rect 54238 21534 54290 21586
rect 54910 21534 54962 21586
rect 55470 21534 55522 21586
rect 56590 21534 56642 21586
rect 59054 21534 59106 21586
rect 59502 21534 59554 21586
rect 59726 21534 59778 21586
rect 60286 21534 60338 21586
rect 60510 21534 60562 21586
rect 60734 21534 60786 21586
rect 67342 21534 67394 21586
rect 69470 21534 69522 21586
rect 74174 21534 74226 21586
rect 74398 21534 74450 21586
rect 74958 21534 75010 21586
rect 76414 21534 76466 21586
rect 77198 21534 77250 21586
rect 81566 21534 81618 21586
rect 82238 21534 82290 21586
rect 87838 21534 87890 21586
rect 88286 21534 88338 21586
rect 90526 21534 90578 21586
rect 91086 21534 91138 21586
rect 93998 21534 94050 21586
rect 94446 21534 94498 21586
rect 97694 21534 97746 21586
rect 98254 21534 98306 21586
rect 104414 21534 104466 21586
rect 108670 21534 108722 21586
rect 21870 21422 21922 21474
rect 23998 21422 24050 21474
rect 29598 21422 29650 21474
rect 30046 21422 30098 21474
rect 32286 21422 32338 21474
rect 33966 21422 34018 21474
rect 34862 21422 34914 21474
rect 36654 21422 36706 21474
rect 41470 21422 41522 21474
rect 43038 21422 43090 21474
rect 44046 21422 44098 21474
rect 47070 21422 47122 21474
rect 48862 21422 48914 21474
rect 49982 21422 50034 21474
rect 51774 21422 51826 21474
rect 52782 21422 52834 21474
rect 64430 21422 64482 21474
rect 66558 21422 66610 21474
rect 67790 21422 67842 21474
rect 68910 21422 68962 21474
rect 73950 21422 74002 21474
rect 75406 21422 75458 21474
rect 79550 21422 79602 21474
rect 93438 21422 93490 21474
rect 103070 21422 103122 21474
rect 103966 21422 104018 21474
rect 108334 21422 108386 21474
rect 42702 21310 42754 21362
rect 43150 21310 43202 21362
rect 46846 21310 46898 21362
rect 48974 21310 49026 21362
rect 49646 21310 49698 21362
rect 49870 21310 49922 21362
rect 51998 21310 52050 21362
rect 53678 21310 53730 21362
rect 74846 21310 74898 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 96638 21142 96690 21194
rect 96742 21142 96794 21194
rect 96846 21142 96898 21194
rect 127358 21142 127410 21194
rect 127462 21142 127514 21194
rect 127566 21142 127618 21194
rect 158078 21142 158130 21194
rect 158182 21142 158234 21194
rect 158286 21142 158338 21194
rect 27582 20974 27634 21026
rect 46398 20974 46450 21026
rect 50206 20974 50258 21026
rect 50654 20974 50706 21026
rect 23326 20862 23378 20914
rect 24558 20862 24610 20914
rect 25006 20862 25058 20914
rect 38558 20862 38610 20914
rect 42030 20862 42082 20914
rect 52110 20862 52162 20914
rect 53678 20862 53730 20914
rect 57374 20862 57426 20914
rect 58270 20862 58322 20914
rect 59838 20862 59890 20914
rect 59950 20862 60002 20914
rect 60510 20862 60562 20914
rect 77534 20862 77586 20914
rect 78430 20862 78482 20914
rect 79326 20862 79378 20914
rect 81454 20862 81506 20914
rect 88734 20862 88786 20914
rect 91310 20862 91362 20914
rect 91982 20862 92034 20914
rect 24110 20750 24162 20802
rect 26686 20750 26738 20802
rect 28590 20750 28642 20802
rect 29374 20750 29426 20802
rect 30046 20750 30098 20802
rect 31838 20750 31890 20802
rect 36878 20750 36930 20802
rect 37326 20750 37378 20802
rect 37774 20750 37826 20802
rect 41806 20750 41858 20802
rect 42702 20750 42754 20802
rect 45054 20750 45106 20802
rect 45390 20750 45442 20802
rect 45614 20750 45666 20802
rect 45950 20750 46002 20802
rect 47406 20750 47458 20802
rect 47742 20750 47794 20802
rect 48974 20750 49026 20802
rect 49310 20750 49362 20802
rect 49534 20750 49586 20802
rect 49870 20750 49922 20802
rect 51326 20750 51378 20802
rect 52558 20750 52610 20802
rect 54350 20750 54402 20802
rect 54798 20750 54850 20802
rect 55918 20750 55970 20802
rect 56366 20750 56418 20802
rect 59054 20750 59106 20802
rect 59390 20750 59442 20802
rect 59614 20750 59666 20802
rect 60622 20750 60674 20802
rect 60958 20750 61010 20802
rect 63310 20750 63362 20802
rect 63646 20750 63698 20802
rect 63870 20750 63922 20802
rect 64094 20750 64146 20802
rect 64766 20750 64818 20802
rect 65214 20750 65266 20802
rect 65550 20750 65602 20802
rect 67006 20750 67058 20802
rect 72046 20750 72098 20802
rect 72830 20750 72882 20802
rect 77086 20750 77138 20802
rect 77758 20750 77810 20802
rect 77982 20750 78034 20802
rect 78542 20750 78594 20802
rect 87614 20750 87666 20802
rect 88398 20750 88450 20802
rect 91870 20750 91922 20802
rect 92094 20750 92146 20802
rect 92430 20750 92482 20802
rect 92878 20750 92930 20802
rect 93438 20750 93490 20802
rect 95566 20750 95618 20802
rect 96350 20750 96402 20802
rect 103518 20750 103570 20802
rect 104302 20750 104354 20802
rect 108222 20750 108274 20802
rect 109006 20750 109058 20802
rect 111694 20750 111746 20802
rect 112366 20750 112418 20802
rect 23662 20638 23714 20690
rect 23774 20638 23826 20690
rect 29150 20638 29202 20690
rect 34750 20638 34802 20690
rect 37550 20638 37602 20690
rect 37998 20638 38050 20690
rect 38110 20638 38162 20690
rect 45838 20638 45890 20690
rect 46846 20638 46898 20690
rect 48190 20638 48242 20690
rect 48526 20638 48578 20690
rect 50094 20638 50146 20690
rect 51662 20638 51714 20690
rect 51774 20638 51826 20690
rect 53006 20638 53058 20690
rect 53230 20638 53282 20690
rect 55134 20638 55186 20690
rect 64318 20638 64370 20690
rect 65774 20638 65826 20690
rect 66222 20638 66274 20690
rect 66558 20638 66610 20690
rect 77422 20638 77474 20690
rect 78766 20638 78818 20690
rect 23886 20526 23938 20578
rect 26462 20526 26514 20578
rect 30606 20526 30658 20578
rect 37214 20526 37266 20578
rect 47070 20526 47122 20578
rect 47294 20526 47346 20578
rect 50766 20526 50818 20578
rect 50878 20526 50930 20578
rect 51550 20526 51602 20578
rect 52894 20526 52946 20578
rect 54126 20526 54178 20578
rect 56814 20526 56866 20578
rect 58830 20526 58882 20578
rect 59166 20526 59218 20578
rect 64430 20526 64482 20578
rect 75182 20526 75234 20578
rect 75630 20526 75682 20578
rect 76526 20526 76578 20578
rect 78318 20526 78370 20578
rect 81566 20526 81618 20578
rect 85262 20526 85314 20578
rect 92766 20526 92818 20578
rect 92990 20526 93042 20578
rect 93774 20526 93826 20578
rect 98702 20526 98754 20578
rect 99150 20526 99202 20578
rect 103294 20526 103346 20578
rect 106654 20526 106706 20578
rect 107998 20526 108050 20578
rect 111358 20526 111410 20578
rect 114830 20526 114882 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 81278 20358 81330 20410
rect 81382 20358 81434 20410
rect 81486 20358 81538 20410
rect 111998 20358 112050 20410
rect 112102 20358 112154 20410
rect 112206 20358 112258 20410
rect 142718 20358 142770 20410
rect 142822 20358 142874 20410
rect 142926 20358 142978 20410
rect 52558 20190 52610 20242
rect 52782 20190 52834 20242
rect 56478 20190 56530 20242
rect 59390 20190 59442 20242
rect 64430 20190 64482 20242
rect 69694 20190 69746 20242
rect 74734 20190 74786 20242
rect 86270 20190 86322 20242
rect 86942 20190 86994 20242
rect 93662 20190 93714 20242
rect 96574 20190 96626 20242
rect 97582 20190 97634 20242
rect 104750 20190 104802 20242
rect 109006 20190 109058 20242
rect 111582 20190 111634 20242
rect 23326 20078 23378 20130
rect 26462 20078 26514 20130
rect 26798 20078 26850 20130
rect 26910 20078 26962 20130
rect 31390 20078 31442 20130
rect 32286 20078 32338 20130
rect 34078 20078 34130 20130
rect 34190 20078 34242 20130
rect 38334 20078 38386 20130
rect 38446 20078 38498 20130
rect 44270 20078 44322 20130
rect 52894 20078 52946 20130
rect 53006 20078 53058 20130
rect 56702 20078 56754 20130
rect 60174 20078 60226 20130
rect 60958 20078 61010 20130
rect 70366 20078 70418 20130
rect 74062 20078 74114 20130
rect 74622 20078 74674 20130
rect 78094 20078 78146 20130
rect 81790 20078 81842 20130
rect 82238 20078 82290 20130
rect 82574 20078 82626 20130
rect 86046 20078 86098 20130
rect 87278 20078 87330 20130
rect 95230 20078 95282 20130
rect 96126 20078 96178 20130
rect 96798 20078 96850 20130
rect 97806 20078 97858 20130
rect 101838 20078 101890 20130
rect 105870 20078 105922 20130
rect 106094 20078 106146 20130
rect 106766 20078 106818 20130
rect 107774 20078 107826 20130
rect 108558 20078 108610 20130
rect 109454 20078 109506 20130
rect 109902 20078 109954 20130
rect 110238 20078 110290 20130
rect 113374 20078 113426 20130
rect 19182 19966 19234 20018
rect 23102 19966 23154 20018
rect 23438 19966 23490 20018
rect 26238 19966 26290 20018
rect 27806 19966 27858 20018
rect 30942 19966 30994 20018
rect 31614 19966 31666 20018
rect 31950 19966 32002 20018
rect 32958 19966 33010 20018
rect 33406 19966 33458 20018
rect 33630 19966 33682 20018
rect 33854 19966 33906 20018
rect 34750 19966 34802 20018
rect 35198 19966 35250 20018
rect 41022 19966 41074 20018
rect 43710 19966 43762 20018
rect 51998 19966 52050 20018
rect 56814 19966 56866 20018
rect 59726 19966 59778 20018
rect 61182 19966 61234 20018
rect 67902 19966 67954 20018
rect 69134 19966 69186 20018
rect 70142 19966 70194 20018
rect 74510 19966 74562 20018
rect 75182 19966 75234 20018
rect 75406 19966 75458 20018
rect 75966 19966 76018 20018
rect 76302 19966 76354 20018
rect 77310 19966 77362 20018
rect 80894 19966 80946 20018
rect 81230 19966 81282 20018
rect 81566 19966 81618 20018
rect 82126 19966 82178 20018
rect 82350 19966 82402 20018
rect 86382 19966 86434 20018
rect 86606 19966 86658 20018
rect 90302 19966 90354 20018
rect 90862 19966 90914 20018
rect 95790 19966 95842 20018
rect 96462 19966 96514 20018
rect 97022 19966 97074 20018
rect 97358 19966 97410 20018
rect 97470 19966 97522 20018
rect 100830 19966 100882 20018
rect 101278 19966 101330 20018
rect 104638 19966 104690 20018
rect 104974 19966 105026 20018
rect 105198 19966 105250 20018
rect 105422 19966 105474 20018
rect 105982 19966 106034 20018
rect 106430 19966 106482 20018
rect 107214 19966 107266 20018
rect 108222 19966 108274 20018
rect 108782 19966 108834 20018
rect 109118 19966 109170 20018
rect 109790 19966 109842 20018
rect 110014 19966 110066 20018
rect 111918 19966 111970 20018
rect 112366 19966 112418 20018
rect 112590 19966 112642 20018
rect 112926 19966 112978 20018
rect 113262 19966 113314 20018
rect 113486 19966 113538 20018
rect 113934 19966 113986 20018
rect 19854 19854 19906 19906
rect 21982 19854 22034 19906
rect 22430 19854 22482 19906
rect 28590 19854 28642 19906
rect 30718 19854 30770 19906
rect 31166 19854 31218 19906
rect 33182 19854 33234 19906
rect 35870 19854 35922 19906
rect 37998 19854 38050 19906
rect 39006 19854 39058 19906
rect 41582 19854 41634 19906
rect 43374 19854 43426 19906
rect 50990 19854 51042 19906
rect 53342 19854 53394 19906
rect 53902 19854 53954 19906
rect 59838 19854 59890 19906
rect 64542 19854 64594 19906
rect 64990 19854 65042 19906
rect 67118 19854 67170 19906
rect 68350 19854 68402 19906
rect 73166 19854 73218 19906
rect 73614 19854 73666 19906
rect 76750 19854 76802 19906
rect 77646 19854 77698 19906
rect 81342 19854 81394 19906
rect 85374 19854 85426 19906
rect 85710 19854 85762 19906
rect 93214 19854 93266 19906
rect 94894 19854 94946 19906
rect 98366 19854 98418 19906
rect 110910 19854 110962 19906
rect 112478 19854 112530 19906
rect 26910 19742 26962 19794
rect 38446 19742 38498 19794
rect 74174 19742 74226 19794
rect 78206 19742 78258 19794
rect 107886 19742 107938 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 96638 19574 96690 19626
rect 96742 19574 96794 19626
rect 96846 19574 96898 19626
rect 127358 19574 127410 19626
rect 127462 19574 127514 19626
rect 127566 19574 127618 19626
rect 158078 19574 158130 19626
rect 158182 19574 158234 19626
rect 158286 19574 158338 19626
rect 22766 19406 22818 19458
rect 43262 19406 43314 19458
rect 52110 19406 52162 19458
rect 53118 19406 53170 19458
rect 85710 19406 85762 19458
rect 86382 19406 86434 19458
rect 94334 19406 94386 19458
rect 94894 19406 94946 19458
rect 28478 19294 28530 19346
rect 37102 19294 37154 19346
rect 40798 19294 40850 19346
rect 49870 19294 49922 19346
rect 52894 19294 52946 19346
rect 55246 19294 55298 19346
rect 58606 19294 58658 19346
rect 66782 19294 66834 19346
rect 68462 19294 68514 19346
rect 70590 19294 70642 19346
rect 71934 19294 71986 19346
rect 73726 19294 73778 19346
rect 74286 19294 74338 19346
rect 82014 19294 82066 19346
rect 86270 19294 86322 19346
rect 86718 19294 86770 19346
rect 90862 19294 90914 19346
rect 94334 19294 94386 19346
rect 95230 19294 95282 19346
rect 95790 19294 95842 19346
rect 98142 19294 98194 19346
rect 105422 19294 105474 19346
rect 108670 19294 108722 19346
rect 112366 19294 112418 19346
rect 114046 19294 114098 19346
rect 23102 19182 23154 19234
rect 23886 19182 23938 19234
rect 25454 19182 25506 19234
rect 33854 19182 33906 19234
rect 37326 19182 37378 19234
rect 37550 19182 37602 19234
rect 37998 19182 38050 19234
rect 39118 19182 39170 19234
rect 41358 19182 41410 19234
rect 43598 19182 43650 19234
rect 47630 19182 47682 19234
rect 48414 19182 48466 19234
rect 48974 19182 49026 19234
rect 51102 19182 51154 19234
rect 51326 19182 51378 19234
rect 51438 19182 51490 19234
rect 51998 19182 52050 19234
rect 53342 19182 53394 19234
rect 55134 19182 55186 19234
rect 56030 19182 56082 19234
rect 58718 19182 58770 19234
rect 60734 19182 60786 19234
rect 61182 19182 61234 19234
rect 63870 19182 63922 19234
rect 64206 19182 64258 19234
rect 66334 19182 66386 19234
rect 67006 19182 67058 19234
rect 67566 19182 67618 19234
rect 71374 19182 71426 19234
rect 77198 19182 77250 19234
rect 86830 19182 86882 19234
rect 87278 19182 87330 19234
rect 90638 19182 90690 19234
rect 96014 19182 96066 19234
rect 97246 19182 97298 19234
rect 106094 19182 106146 19234
rect 109454 19182 109506 19234
rect 112702 19182 112754 19234
rect 23326 19070 23378 19122
rect 23774 19070 23826 19122
rect 26238 19070 26290 19122
rect 30270 19070 30322 19122
rect 36990 19070 37042 19122
rect 39790 19070 39842 19122
rect 42814 19070 42866 19122
rect 46734 19070 46786 19122
rect 46846 19070 46898 19122
rect 47518 19070 47570 19122
rect 48302 19070 48354 19122
rect 50206 19070 50258 19122
rect 52670 19070 52722 19122
rect 53566 19070 53618 19122
rect 54014 19070 54066 19122
rect 55358 19070 55410 19122
rect 55694 19070 55746 19122
rect 58270 19070 58322 19122
rect 62302 19070 62354 19122
rect 64766 19070 64818 19122
rect 66558 19070 66610 19122
rect 72942 19070 72994 19122
rect 75294 19070 75346 19122
rect 75518 19070 75570 19122
rect 78990 19070 79042 19122
rect 87614 19070 87666 19122
rect 91086 19070 91138 19122
rect 91310 19070 91362 19122
rect 97806 19070 97858 19122
rect 99934 19070 99986 19122
rect 104974 19070 105026 19122
rect 105870 19070 105922 19122
rect 107886 19070 107938 19122
rect 113150 19070 113202 19122
rect 22878 18958 22930 19010
rect 23550 18958 23602 19010
rect 24446 18958 24498 19010
rect 29262 18958 29314 19010
rect 43374 18958 43426 19010
rect 46510 18958 46562 19010
rect 49534 18958 49586 19010
rect 49758 18958 49810 19010
rect 49982 18958 50034 19010
rect 50878 18958 50930 19010
rect 51662 18958 51714 19010
rect 52558 18958 52610 19010
rect 54686 18958 54738 19010
rect 54910 18958 54962 19010
rect 55918 18958 55970 19010
rect 61294 18958 61346 19010
rect 62414 18958 62466 19010
rect 67118 18958 67170 19010
rect 73278 18958 73330 19010
rect 74846 18958 74898 19010
rect 75070 18958 75122 19010
rect 75182 18958 75234 19010
rect 85038 18958 85090 19010
rect 85486 18958 85538 19010
rect 85822 18958 85874 19010
rect 86606 18958 86658 19010
rect 87838 18958 87890 19010
rect 87950 18958 88002 19010
rect 88062 18958 88114 19010
rect 88622 18958 88674 19010
rect 91982 18958 92034 19010
rect 92430 18958 92482 19010
rect 93550 18958 93602 19010
rect 94782 18958 94834 19010
rect 96350 18958 96402 19010
rect 96686 18958 96738 19010
rect 96798 18958 96850 19010
rect 96910 18958 96962 19010
rect 98030 18958 98082 19010
rect 98254 18958 98306 19010
rect 98814 18958 98866 19010
rect 99262 18958 99314 19010
rect 100270 18958 100322 19010
rect 112814 18958 112866 19010
rect 112926 18958 112978 19010
rect 114158 18958 114210 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 81278 18790 81330 18842
rect 81382 18790 81434 18842
rect 81486 18790 81538 18842
rect 111998 18790 112050 18842
rect 112102 18790 112154 18842
rect 112206 18790 112258 18842
rect 142718 18790 142770 18842
rect 142822 18790 142874 18842
rect 142926 18790 142978 18842
rect 26350 18622 26402 18674
rect 26686 18622 26738 18674
rect 32174 18622 32226 18674
rect 34302 18622 34354 18674
rect 34862 18622 34914 18674
rect 49534 18622 49586 18674
rect 53454 18622 53506 18674
rect 56702 18622 56754 18674
rect 60062 18622 60114 18674
rect 66782 18622 66834 18674
rect 70142 18622 70194 18674
rect 86158 18622 86210 18674
rect 91534 18622 91586 18674
rect 91646 18622 91698 18674
rect 91758 18622 91810 18674
rect 25342 18510 25394 18562
rect 26462 18510 26514 18562
rect 52446 18510 52498 18562
rect 58606 18510 58658 18562
rect 58718 18510 58770 18562
rect 61966 18510 62018 18562
rect 62526 18510 62578 18562
rect 62638 18510 62690 18562
rect 65102 18510 65154 18562
rect 67678 18510 67730 18562
rect 74622 18510 74674 18562
rect 93550 18510 93602 18562
rect 95790 18510 95842 18562
rect 96350 18510 96402 18562
rect 100382 18510 100434 18562
rect 106430 18510 106482 18562
rect 114942 18510 114994 18562
rect 21534 18398 21586 18450
rect 26910 18398 26962 18450
rect 28814 18398 28866 18450
rect 29822 18398 29874 18450
rect 30046 18398 30098 18450
rect 30270 18398 30322 18450
rect 30494 18398 30546 18450
rect 31838 18398 31890 18450
rect 32510 18398 32562 18450
rect 34638 18398 34690 18450
rect 34750 18398 34802 18450
rect 35310 18398 35362 18450
rect 37326 18398 37378 18450
rect 42142 18398 42194 18450
rect 42590 18398 42642 18450
rect 43598 18398 43650 18450
rect 45390 18398 45442 18450
rect 46286 18398 46338 18450
rect 47518 18398 47570 18450
rect 47630 18398 47682 18450
rect 47742 18398 47794 18450
rect 48190 18398 48242 18450
rect 48862 18398 48914 18450
rect 49310 18398 49362 18450
rect 49982 18398 50034 18450
rect 50318 18398 50370 18450
rect 51214 18398 51266 18450
rect 51886 18398 51938 18450
rect 52110 18398 52162 18450
rect 52670 18398 52722 18450
rect 53118 18398 53170 18450
rect 53342 18398 53394 18450
rect 56926 18398 56978 18450
rect 58382 18398 58434 18450
rect 59502 18398 59554 18450
rect 60734 18398 60786 18450
rect 61630 18398 61682 18450
rect 62862 18398 62914 18450
rect 63422 18398 63474 18450
rect 64430 18398 64482 18450
rect 66558 18398 66610 18450
rect 69022 18398 69074 18450
rect 69470 18398 69522 18450
rect 69582 18398 69634 18450
rect 69694 18398 69746 18450
rect 70702 18398 70754 18450
rect 73278 18398 73330 18450
rect 74062 18398 74114 18450
rect 74174 18398 74226 18450
rect 74286 18398 74338 18450
rect 76078 18398 76130 18450
rect 77758 18398 77810 18450
rect 79550 18398 79602 18450
rect 80446 18398 80498 18450
rect 81118 18398 81170 18450
rect 83470 18398 83522 18450
rect 85822 18398 85874 18450
rect 86382 18398 86434 18450
rect 86830 18398 86882 18450
rect 90302 18398 90354 18450
rect 91086 18398 91138 18450
rect 92206 18398 92258 18450
rect 92542 18398 92594 18450
rect 93102 18398 93154 18450
rect 95342 18398 95394 18450
rect 96126 18398 96178 18450
rect 96686 18398 96738 18450
rect 99710 18398 99762 18450
rect 100046 18398 100098 18450
rect 101390 18398 101442 18450
rect 101726 18398 101778 18450
rect 101950 18398 102002 18450
rect 102510 18398 102562 18450
rect 106094 18398 106146 18450
rect 106990 18398 107042 18450
rect 108670 18398 108722 18450
rect 108894 18398 108946 18450
rect 109342 18398 109394 18450
rect 109566 18398 109618 18450
rect 111694 18398 111746 18450
rect 112142 18398 112194 18450
rect 112366 18398 112418 18450
rect 22206 18286 22258 18338
rect 24334 18286 24386 18338
rect 27358 18286 27410 18338
rect 33742 18286 33794 18338
rect 35646 18286 35698 18338
rect 36206 18286 36258 18338
rect 36990 18286 37042 18338
rect 38110 18286 38162 18338
rect 40238 18286 40290 18338
rect 42702 18286 42754 18338
rect 43150 18286 43202 18338
rect 45726 18286 45778 18338
rect 51774 18286 51826 18338
rect 57374 18286 57426 18338
rect 57822 18286 57874 18338
rect 61070 18286 61122 18338
rect 63086 18286 63138 18338
rect 63758 18286 63810 18338
rect 71598 18286 71650 18338
rect 75630 18286 75682 18338
rect 76638 18286 76690 18338
rect 84030 18286 84082 18338
rect 84478 18286 84530 18338
rect 85038 18286 85090 18338
rect 85486 18286 85538 18338
rect 86270 18286 86322 18338
rect 87166 18286 87218 18338
rect 87950 18286 88002 18338
rect 94446 18286 94498 18338
rect 94782 18286 94834 18338
rect 95902 18286 95954 18338
rect 98926 18286 98978 18338
rect 100830 18286 100882 18338
rect 101838 18286 101890 18338
rect 105758 18286 105810 18338
rect 109118 18286 109170 18338
rect 111022 18286 111074 18338
rect 111918 18286 111970 18338
rect 33182 18174 33234 18226
rect 33518 18174 33570 18226
rect 35422 18174 35474 18226
rect 35646 18174 35698 18226
rect 52894 18174 52946 18226
rect 56590 18174 56642 18226
rect 57262 18174 57314 18226
rect 59726 18174 59778 18226
rect 62078 18174 62130 18226
rect 72942 18174 72994 18226
rect 115054 18174 115106 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 96638 18006 96690 18058
rect 96742 18006 96794 18058
rect 96846 18006 96898 18058
rect 127358 18006 127410 18058
rect 127462 18006 127514 18058
rect 127566 18006 127618 18058
rect 158078 18006 158130 18058
rect 158182 18006 158234 18058
rect 158286 18006 158338 18058
rect 22654 17838 22706 17890
rect 23214 17838 23266 17890
rect 41918 17838 41970 17890
rect 42142 17838 42194 17890
rect 42254 17838 42306 17890
rect 50990 17838 51042 17890
rect 64430 17838 64482 17890
rect 24558 17726 24610 17778
rect 32062 17726 32114 17778
rect 34190 17726 34242 17778
rect 35422 17726 35474 17778
rect 45390 17726 45442 17778
rect 56142 17726 56194 17778
rect 58382 17726 58434 17778
rect 60622 17726 60674 17778
rect 64318 17726 64370 17778
rect 71374 17726 71426 17778
rect 72270 17726 72322 17778
rect 73054 17726 73106 17778
rect 77198 17726 77250 17778
rect 84254 17726 84306 17778
rect 86942 17726 86994 17778
rect 88174 17726 88226 17778
rect 89630 17726 89682 17778
rect 93214 17726 93266 17778
rect 97246 17726 97298 17778
rect 97694 17726 97746 17778
rect 98142 17726 98194 17778
rect 22766 17614 22818 17666
rect 22990 17614 23042 17666
rect 23326 17614 23378 17666
rect 23774 17614 23826 17666
rect 24110 17614 24162 17666
rect 31054 17614 31106 17666
rect 31390 17614 31442 17666
rect 34526 17614 34578 17666
rect 41694 17614 41746 17666
rect 45838 17614 45890 17666
rect 46510 17614 46562 17666
rect 47294 17614 47346 17666
rect 47966 17614 48018 17666
rect 48862 17614 48914 17666
rect 49534 17614 49586 17666
rect 55470 17614 55522 17666
rect 62190 17614 62242 17666
rect 63422 17614 63474 17666
rect 63870 17614 63922 17666
rect 65662 17614 65714 17666
rect 68910 17614 68962 17666
rect 69582 17614 69634 17666
rect 70030 17614 70082 17666
rect 70478 17614 70530 17666
rect 70926 17614 70978 17666
rect 71822 17614 71874 17666
rect 76862 17614 76914 17666
rect 79998 17614 80050 17666
rect 80782 17614 80834 17666
rect 85374 17614 85426 17666
rect 85598 17614 85650 17666
rect 86046 17614 86098 17666
rect 87278 17614 87330 17666
rect 87838 17614 87890 17666
rect 87950 17614 88002 17666
rect 88286 17614 88338 17666
rect 94334 17614 94386 17666
rect 94894 17614 94946 17666
rect 99822 17614 99874 17666
rect 106206 17614 106258 17666
rect 106542 17614 106594 17666
rect 107550 17614 107602 17666
rect 109118 17614 109170 17666
rect 109790 17614 109842 17666
rect 23550 17502 23602 17554
rect 23998 17502 24050 17554
rect 29598 17502 29650 17554
rect 30718 17502 30770 17554
rect 39454 17502 39506 17554
rect 39566 17502 39618 17554
rect 41022 17502 41074 17554
rect 41134 17502 41186 17554
rect 46286 17502 46338 17554
rect 48078 17502 48130 17554
rect 49198 17502 49250 17554
rect 49870 17502 49922 17554
rect 50542 17502 50594 17554
rect 50990 17502 51042 17554
rect 51102 17502 51154 17554
rect 58830 17502 58882 17554
rect 58942 17502 58994 17554
rect 59502 17502 59554 17554
rect 61966 17502 62018 17554
rect 65438 17502 65490 17554
rect 67006 17502 67058 17554
rect 68686 17502 68738 17554
rect 69358 17502 69410 17554
rect 72718 17502 72770 17554
rect 88734 17502 88786 17554
rect 92206 17502 92258 17554
rect 101726 17502 101778 17554
rect 106766 17502 106818 17554
rect 107662 17502 107714 17554
rect 107998 17502 108050 17554
rect 22318 17390 22370 17442
rect 22654 17390 22706 17442
rect 29934 17390 29986 17442
rect 30830 17390 30882 17442
rect 34862 17390 34914 17442
rect 39230 17390 39282 17442
rect 41358 17390 41410 17442
rect 46958 17390 47010 17442
rect 48302 17390 48354 17442
rect 50206 17390 50258 17442
rect 52782 17390 52834 17442
rect 59166 17390 59218 17442
rect 59950 17390 60002 17442
rect 61070 17390 61122 17442
rect 67790 17390 67842 17442
rect 73726 17390 73778 17442
rect 74174 17390 74226 17442
rect 79326 17390 79378 17442
rect 79774 17390 79826 17442
rect 83134 17390 83186 17442
rect 84366 17390 84418 17442
rect 85150 17390 85202 17442
rect 85822 17390 85874 17442
rect 86382 17390 86434 17442
rect 89294 17390 89346 17442
rect 90078 17390 90130 17442
rect 90862 17390 90914 17442
rect 91198 17390 91250 17442
rect 92766 17390 92818 17442
rect 93662 17390 93714 17442
rect 97806 17390 97858 17442
rect 98254 17390 98306 17442
rect 98702 17390 98754 17442
rect 99262 17390 99314 17442
rect 106318 17390 106370 17442
rect 107774 17390 107826 17442
rect 108894 17390 108946 17442
rect 112254 17390 112306 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 81278 17222 81330 17274
rect 81382 17222 81434 17274
rect 81486 17222 81538 17274
rect 111998 17222 112050 17274
rect 112102 17222 112154 17274
rect 112206 17222 112258 17274
rect 142718 17222 142770 17274
rect 142822 17222 142874 17274
rect 142926 17222 142978 17274
rect 19630 17054 19682 17106
rect 23550 17054 23602 17106
rect 25342 17054 25394 17106
rect 28254 17054 28306 17106
rect 30046 17054 30098 17106
rect 36094 17054 36146 17106
rect 38110 17054 38162 17106
rect 44270 17054 44322 17106
rect 49870 17054 49922 17106
rect 51102 17054 51154 17106
rect 51214 17054 51266 17106
rect 51326 17054 51378 17106
rect 51886 17054 51938 17106
rect 52334 17054 52386 17106
rect 56702 17054 56754 17106
rect 58718 17054 58770 17106
rect 60398 17054 60450 17106
rect 63086 17054 63138 17106
rect 64542 17054 64594 17106
rect 75742 17054 75794 17106
rect 79214 17054 79266 17106
rect 80110 17054 80162 17106
rect 80894 17054 80946 17106
rect 81230 17054 81282 17106
rect 82126 17054 82178 17106
rect 83246 17054 83298 17106
rect 83918 17054 83970 17106
rect 87390 17054 87442 17106
rect 89070 17054 89122 17106
rect 89630 17054 89682 17106
rect 90862 17054 90914 17106
rect 92318 17054 92370 17106
rect 92542 17054 92594 17106
rect 93662 17054 93714 17106
rect 93886 17054 93938 17106
rect 95006 17054 95058 17106
rect 96238 17054 96290 17106
rect 97358 17054 97410 17106
rect 99598 17054 99650 17106
rect 99822 17054 99874 17106
rect 100942 17054 100994 17106
rect 102510 17054 102562 17106
rect 105422 17054 105474 17106
rect 109790 17054 109842 17106
rect 109902 17054 109954 17106
rect 115278 17054 115330 17106
rect 21646 16942 21698 16994
rect 28030 16942 28082 16994
rect 30270 16942 30322 16994
rect 31054 16942 31106 16994
rect 31502 16942 31554 16994
rect 32174 16942 32226 16994
rect 33854 16942 33906 16994
rect 38222 16942 38274 16994
rect 38894 16942 38946 16994
rect 39006 16942 39058 16994
rect 45950 16942 46002 16994
rect 47406 16942 47458 16994
rect 47630 16942 47682 16994
rect 48750 16942 48802 16994
rect 53566 16942 53618 16994
rect 57598 16942 57650 16994
rect 63758 16942 63810 16994
rect 68910 16942 68962 16994
rect 79550 16942 79602 16994
rect 80446 16942 80498 16994
rect 81118 16942 81170 16994
rect 81678 16942 81730 16994
rect 81902 16942 81954 16994
rect 82238 16942 82290 16994
rect 82686 16942 82738 16994
rect 94446 16942 94498 16994
rect 98254 16942 98306 16994
rect 100158 16942 100210 16994
rect 101726 16942 101778 16994
rect 104974 16942 105026 16994
rect 105310 16942 105362 16994
rect 115614 16942 115666 16994
rect 19294 16830 19346 16882
rect 20190 16830 20242 16882
rect 26462 16830 26514 16882
rect 26686 16830 26738 16882
rect 27134 16830 27186 16882
rect 27918 16830 27970 16882
rect 30382 16830 30434 16882
rect 30718 16830 30770 16882
rect 31838 16830 31890 16882
rect 32398 16830 32450 16882
rect 35646 16830 35698 16882
rect 37774 16830 37826 16882
rect 38334 16830 38386 16882
rect 38670 16830 38722 16882
rect 40910 16830 40962 16882
rect 47854 16830 47906 16882
rect 48078 16830 48130 16882
rect 49086 16830 49138 16882
rect 50878 16830 50930 16882
rect 52894 16830 52946 16882
rect 57038 16830 57090 16882
rect 60734 16830 60786 16882
rect 60958 16830 61010 16882
rect 62190 16830 62242 16882
rect 62414 16830 62466 16882
rect 63422 16830 63474 16882
rect 66222 16830 66274 16882
rect 66446 16830 66498 16882
rect 72494 16830 72546 16882
rect 76190 16830 76242 16882
rect 76414 16830 76466 16882
rect 76862 16830 76914 16882
rect 81342 16830 81394 16882
rect 83582 16830 83634 16882
rect 86270 16830 86322 16882
rect 87054 16830 87106 16882
rect 89294 16830 89346 16882
rect 89742 16830 89794 16882
rect 89966 16830 90018 16882
rect 93102 16830 93154 16882
rect 96350 16830 96402 16882
rect 96686 16830 96738 16882
rect 97022 16830 97074 16882
rect 97582 16830 97634 16882
rect 97918 16830 97970 16882
rect 100382 16830 100434 16882
rect 100830 16830 100882 16882
rect 101054 16830 101106 16882
rect 101390 16830 101442 16882
rect 101950 16830 102002 16882
rect 105646 16830 105698 16882
rect 106318 16830 106370 16882
rect 108782 16830 108834 16882
rect 109230 16830 109282 16882
rect 109678 16830 109730 16882
rect 111918 16830 111970 16882
rect 112142 16830 112194 16882
rect 112814 16830 112866 16882
rect 20302 16718 20354 16770
rect 26574 16718 26626 16770
rect 41694 16718 41746 16770
rect 43822 16718 43874 16770
rect 55694 16718 55746 16770
rect 61518 16718 61570 16770
rect 62078 16718 62130 16770
rect 73166 16718 73218 16770
rect 75294 16718 75346 16770
rect 76302 16718 76354 16770
rect 77198 16718 77250 16770
rect 77646 16718 77698 16770
rect 78206 16718 78258 16770
rect 78990 16718 79042 16770
rect 88398 16718 88450 16770
rect 90414 16718 90466 16770
rect 91646 16718 91698 16770
rect 96574 16718 96626 16770
rect 97470 16718 97522 16770
rect 98814 16718 98866 16770
rect 101502 16718 101554 16770
rect 102958 16718 103010 16770
rect 103854 16718 103906 16770
rect 104190 16718 104242 16770
rect 50654 16606 50706 16658
rect 82574 16606 82626 16658
rect 98366 16606 98418 16658
rect 115726 16606 115778 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 96638 16438 96690 16490
rect 96742 16438 96794 16490
rect 96846 16438 96898 16490
rect 127358 16438 127410 16490
rect 127462 16438 127514 16490
rect 127566 16438 127618 16490
rect 158078 16438 158130 16490
rect 158182 16438 158234 16490
rect 158286 16438 158338 16490
rect 31166 16270 31218 16322
rect 31950 16270 32002 16322
rect 32622 16270 32674 16322
rect 33406 16270 33458 16322
rect 33742 16270 33794 16322
rect 48414 16270 48466 16322
rect 62078 16270 62130 16322
rect 78542 16270 78594 16322
rect 79326 16270 79378 16322
rect 84142 16270 84194 16322
rect 84926 16270 84978 16322
rect 87390 16270 87442 16322
rect 20750 16158 20802 16210
rect 24558 16158 24610 16210
rect 28478 16158 28530 16210
rect 34974 16158 35026 16210
rect 36430 16158 36482 16210
rect 39902 16158 39954 16210
rect 40910 16158 40962 16210
rect 47518 16158 47570 16210
rect 53006 16158 53058 16210
rect 53566 16158 53618 16210
rect 55918 16158 55970 16210
rect 61070 16158 61122 16210
rect 64318 16158 64370 16210
rect 71262 16158 71314 16210
rect 72046 16158 72098 16210
rect 72494 16158 72546 16210
rect 73166 16158 73218 16210
rect 74286 16158 74338 16210
rect 77982 16158 78034 16210
rect 78430 16158 78482 16210
rect 79998 16158 80050 16210
rect 82126 16158 82178 16210
rect 84142 16158 84194 16210
rect 87166 16158 87218 16210
rect 88958 16158 89010 16210
rect 90750 16158 90802 16210
rect 91982 16158 92034 16210
rect 92878 16158 92930 16210
rect 93998 16158 94050 16210
rect 17950 16046 18002 16098
rect 21646 16046 21698 16098
rect 24894 16046 24946 16098
rect 25566 16046 25618 16098
rect 29822 16046 29874 16098
rect 30046 16046 30098 16098
rect 30494 16046 30546 16098
rect 30830 16046 30882 16098
rect 31838 16046 31890 16098
rect 32510 16046 32562 16098
rect 34078 16046 34130 16098
rect 36990 16046 37042 16098
rect 40238 16046 40290 16098
rect 40574 16046 40626 16098
rect 41134 16046 41186 16098
rect 41358 16046 41410 16098
rect 42030 16046 42082 16098
rect 42142 16046 42194 16098
rect 46846 16046 46898 16098
rect 48078 16046 48130 16098
rect 48638 16046 48690 16098
rect 49198 16046 49250 16098
rect 49534 16046 49586 16098
rect 49870 16046 49922 16098
rect 52894 16046 52946 16098
rect 57486 16046 57538 16098
rect 61406 16046 61458 16098
rect 61966 16046 62018 16098
rect 64542 16046 64594 16098
rect 68462 16046 68514 16098
rect 73278 16046 73330 16098
rect 73614 16046 73666 16098
rect 74846 16046 74898 16098
rect 75070 16046 75122 16098
rect 75294 16046 75346 16098
rect 77086 16046 77138 16098
rect 77646 16046 77698 16098
rect 80558 16046 80610 16098
rect 80782 16046 80834 16098
rect 81342 16046 81394 16098
rect 86942 16046 86994 16098
rect 88846 16046 88898 16098
rect 90638 16046 90690 16098
rect 93550 16046 93602 16098
rect 18622 15934 18674 15986
rect 22430 15934 22482 15986
rect 25230 15934 25282 15986
rect 26350 15934 26402 15986
rect 33630 15934 33682 15986
rect 35758 15934 35810 15986
rect 37774 15934 37826 15986
rect 40798 15934 40850 15986
rect 41694 15934 41746 15986
rect 42814 15934 42866 15986
rect 43150 15934 43202 15986
rect 43598 15934 43650 15986
rect 47294 15934 47346 15986
rect 49758 15934 49810 15986
rect 53118 15934 53170 15986
rect 56590 15934 56642 15986
rect 56926 15934 56978 15986
rect 62078 15934 62130 15986
rect 65102 15934 65154 15986
rect 69134 15934 69186 15986
rect 73054 15934 73106 15986
rect 75630 15934 75682 15986
rect 80334 15934 80386 15986
rect 95342 16270 95394 16322
rect 104638 16270 104690 16322
rect 105310 16270 105362 16322
rect 95342 16158 95394 16210
rect 98814 16158 98866 16210
rect 100270 16158 100322 16210
rect 104414 16158 104466 16210
rect 104862 16158 104914 16210
rect 105310 16158 105362 16210
rect 95790 16046 95842 16098
rect 96462 16046 96514 16098
rect 101502 16046 101554 16098
rect 101950 16046 102002 16098
rect 107886 16046 107938 16098
rect 108558 16046 108610 16098
rect 110238 16046 110290 16098
rect 112366 16046 112418 16098
rect 91086 15934 91138 15986
rect 94782 15934 94834 15986
rect 25118 15822 25170 15874
rect 29598 15822 29650 15874
rect 30270 15822 30322 15874
rect 30382 15822 30434 15874
rect 31054 15822 31106 15874
rect 31950 15822 32002 15874
rect 32622 15822 32674 15874
rect 34414 15822 34466 15874
rect 35534 15822 35586 15874
rect 35870 15822 35922 15874
rect 36094 15822 36146 15874
rect 40350 15822 40402 15874
rect 41806 15822 41858 15874
rect 47406 15822 47458 15874
rect 47630 15822 47682 15874
rect 51774 15822 51826 15874
rect 52222 15822 52274 15874
rect 52670 15822 52722 15874
rect 54126 15822 54178 15874
rect 56254 15822 56306 15874
rect 61518 15822 61570 15874
rect 62638 15822 62690 15874
rect 64094 15822 64146 15874
rect 75182 15822 75234 15874
rect 76302 15822 76354 15874
rect 76974 15822 77026 15874
rect 77198 15822 77250 15874
rect 78990 15822 79042 15874
rect 79438 15822 79490 15874
rect 80558 15822 80610 15874
rect 81678 15822 81730 15874
rect 82686 15822 82738 15874
rect 83134 15822 83186 15874
rect 83582 15822 83634 15874
rect 84590 15822 84642 15874
rect 85150 15822 85202 15874
rect 85598 15822 85650 15874
rect 85934 15822 85986 15874
rect 86494 15822 86546 15874
rect 90862 15822 90914 15874
rect 92430 15822 92482 15874
rect 94558 15822 94610 15874
rect 94894 15822 94946 15874
rect 99822 15822 99874 15874
rect 100830 15822 100882 15874
rect 105758 15822 105810 15874
rect 106318 15822 106370 15874
rect 106990 15822 107042 15874
rect 107998 15822 108050 15874
rect 108110 15822 108162 15874
rect 108894 15822 108946 15874
rect 110350 15822 110402 15874
rect 112478 15822 112530 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 81278 15654 81330 15706
rect 81382 15654 81434 15706
rect 81486 15654 81538 15706
rect 111998 15654 112050 15706
rect 112102 15654 112154 15706
rect 112206 15654 112258 15706
rect 142718 15654 142770 15706
rect 142822 15654 142874 15706
rect 142926 15654 142978 15706
rect 20414 15486 20466 15538
rect 20750 15486 20802 15538
rect 22318 15486 22370 15538
rect 22766 15486 22818 15538
rect 26014 15486 26066 15538
rect 27582 15486 27634 15538
rect 27918 15486 27970 15538
rect 28814 15486 28866 15538
rect 34078 15486 34130 15538
rect 35982 15486 36034 15538
rect 36542 15486 36594 15538
rect 37326 15486 37378 15538
rect 38334 15486 38386 15538
rect 44270 15486 44322 15538
rect 48862 15486 48914 15538
rect 49422 15486 49474 15538
rect 54126 15486 54178 15538
rect 54350 15486 54402 15538
rect 55134 15486 55186 15538
rect 57150 15486 57202 15538
rect 57374 15486 57426 15538
rect 60510 15486 60562 15538
rect 68350 15486 68402 15538
rect 69694 15486 69746 15538
rect 70142 15486 70194 15538
rect 71486 15486 71538 15538
rect 73838 15486 73890 15538
rect 78430 15486 78482 15538
rect 79550 15486 79602 15538
rect 87278 15486 87330 15538
rect 87950 15486 88002 15538
rect 92094 15486 92146 15538
rect 94334 15486 94386 15538
rect 100270 15486 100322 15538
rect 101726 15486 101778 15538
rect 102062 15486 102114 15538
rect 102174 15486 102226 15538
rect 102510 15486 102562 15538
rect 107550 15486 107602 15538
rect 108222 15486 108274 15538
rect 108782 15486 108834 15538
rect 109230 15486 109282 15538
rect 20862 15374 20914 15426
rect 21982 15374 22034 15426
rect 22206 15374 22258 15426
rect 22878 15374 22930 15426
rect 23326 15374 23378 15426
rect 25230 15374 25282 15426
rect 26126 15374 26178 15426
rect 35758 15374 35810 15426
rect 36318 15374 36370 15426
rect 37662 15374 37714 15426
rect 38110 15374 38162 15426
rect 41694 15374 41746 15426
rect 46062 15374 46114 15426
rect 48974 15374 49026 15426
rect 57710 15374 57762 15426
rect 70926 15374 70978 15426
rect 72494 15374 72546 15426
rect 74286 15374 74338 15426
rect 75854 15374 75906 15426
rect 80894 15374 80946 15426
rect 83470 15374 83522 15426
rect 89406 15374 89458 15426
rect 100382 15374 100434 15426
rect 101614 15374 101666 15426
rect 108446 15374 108498 15426
rect 108894 15374 108946 15426
rect 20638 15262 20690 15314
rect 21198 15262 21250 15314
rect 22430 15262 22482 15314
rect 25342 15262 25394 15314
rect 25790 15262 25842 15314
rect 27470 15262 27522 15314
rect 27694 15262 27746 15314
rect 35646 15262 35698 15314
rect 36206 15262 36258 15314
rect 36990 15262 37042 15314
rect 37326 15262 37378 15314
rect 37998 15262 38050 15314
rect 41022 15262 41074 15314
rect 45278 15262 45330 15314
rect 53790 15262 53842 15314
rect 54798 15262 54850 15314
rect 61406 15262 61458 15314
rect 63198 15262 63250 15314
rect 63758 15262 63810 15314
rect 64430 15262 64482 15314
rect 68014 15262 68066 15314
rect 68462 15262 68514 15314
rect 68686 15262 68738 15314
rect 70702 15262 70754 15314
rect 71038 15262 71090 15314
rect 75182 15262 75234 15314
rect 80110 15262 80162 15314
rect 86830 15262 86882 15314
rect 88174 15262 88226 15314
rect 88734 15262 88786 15314
rect 93326 15262 93378 15314
rect 96014 15262 96066 15314
rect 97582 15262 97634 15314
rect 97918 15262 97970 15314
rect 100046 15262 100098 15314
rect 100606 15262 100658 15314
rect 101054 15262 101106 15314
rect 101502 15262 101554 15314
rect 102286 15262 102338 15314
rect 103518 15262 103570 15314
rect 104190 15262 104242 15314
rect 106654 15262 106706 15314
rect 107998 15262 108050 15314
rect 108110 15262 108162 15314
rect 109006 15262 109058 15314
rect 24670 15150 24722 15202
rect 39006 15150 39058 15202
rect 39454 15150 39506 15202
rect 43822 15150 43874 15202
rect 48190 15150 48242 15202
rect 50878 15150 50930 15202
rect 53006 15150 53058 15202
rect 54238 15150 54290 15202
rect 58270 15150 58322 15202
rect 58718 15150 58770 15202
rect 59502 15150 59554 15202
rect 60286 15150 60338 15202
rect 61070 15150 61122 15202
rect 62190 15150 62242 15202
rect 65214 15150 65266 15202
rect 67342 15150 67394 15202
rect 69134 15150 69186 15202
rect 70590 15150 70642 15202
rect 73166 15150 73218 15202
rect 74734 15150 74786 15202
rect 77982 15150 78034 15202
rect 79102 15150 79154 15202
rect 83022 15150 83074 15202
rect 83918 15150 83970 15202
rect 86046 15150 86098 15202
rect 91534 15150 91586 15202
rect 93998 15150 94050 15202
rect 95118 15150 95170 15202
rect 95902 15150 95954 15202
rect 103070 15150 103122 15202
rect 107102 15150 107154 15202
rect 109790 15150 109842 15202
rect 48862 15038 48914 15090
rect 92878 15038 92930 15090
rect 98814 15038 98866 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 96638 14870 96690 14922
rect 96742 14870 96794 14922
rect 96846 14870 96898 14922
rect 127358 14870 127410 14922
rect 127462 14870 127514 14922
rect 127566 14870 127618 14922
rect 158078 14870 158130 14922
rect 158182 14870 158234 14922
rect 158286 14870 158338 14922
rect 37550 14702 37602 14754
rect 37886 14702 37938 14754
rect 38334 14702 38386 14754
rect 39006 14702 39058 14754
rect 39342 14702 39394 14754
rect 39790 14702 39842 14754
rect 44942 14702 44994 14754
rect 57710 14702 57762 14754
rect 19966 14590 20018 14642
rect 33966 14590 34018 14642
rect 37550 14590 37602 14642
rect 39006 14590 39058 14642
rect 42142 14590 42194 14642
rect 48638 14590 48690 14642
rect 57822 14590 57874 14642
rect 62526 14702 62578 14754
rect 63422 14702 63474 14754
rect 58382 14590 58434 14642
rect 59390 14590 59442 14642
rect 62526 14590 62578 14642
rect 62862 14590 62914 14642
rect 63310 14590 63362 14642
rect 71822 14590 71874 14642
rect 72382 14590 72434 14642
rect 17166 14478 17218 14530
rect 31054 14478 31106 14530
rect 37102 14478 37154 14530
rect 47966 14478 48018 14530
rect 52670 14478 52722 14530
rect 52894 14478 52946 14530
rect 53230 14478 53282 14530
rect 58382 14478 58434 14530
rect 61406 14478 61458 14530
rect 61630 14478 61682 14530
rect 73502 14702 73554 14754
rect 74398 14702 74450 14754
rect 81454 14702 81506 14754
rect 89070 14702 89122 14754
rect 94446 14702 94498 14754
rect 72942 14590 72994 14642
rect 76750 14590 76802 14642
rect 83134 14590 83186 14642
rect 85262 14590 85314 14642
rect 92094 14590 92146 14642
rect 95230 14590 95282 14642
rect 98254 14590 98306 14642
rect 98702 14590 98754 14642
rect 99038 14590 99090 14642
rect 106094 14590 106146 14642
rect 110574 14590 110626 14642
rect 62078 14478 62130 14530
rect 69022 14478 69074 14530
rect 72494 14478 72546 14530
rect 77086 14478 77138 14530
rect 79214 14478 79266 14530
rect 80782 14478 80834 14530
rect 82686 14478 82738 14530
rect 84702 14478 84754 14530
rect 86830 14478 86882 14530
rect 88174 14478 88226 14530
rect 88846 14478 88898 14530
rect 90078 14478 90130 14530
rect 92878 14478 92930 14530
rect 93102 14478 93154 14530
rect 94894 14478 94946 14530
rect 99598 14478 99650 14530
rect 100270 14478 100322 14530
rect 103182 14478 103234 14530
rect 103742 14478 103794 14530
rect 106430 14478 106482 14530
rect 106654 14478 106706 14530
rect 106990 14478 107042 14530
rect 107662 14478 107714 14530
rect 108110 14478 108162 14530
rect 17838 14366 17890 14418
rect 29150 14366 29202 14418
rect 29262 14366 29314 14418
rect 31838 14366 31890 14418
rect 38446 14366 38498 14418
rect 44830 14366 44882 14418
rect 64990 14366 65042 14418
rect 65326 14366 65378 14418
rect 65550 14366 65602 14418
rect 65886 14366 65938 14418
rect 66446 14366 66498 14418
rect 66670 14366 66722 14418
rect 66782 14366 66834 14418
rect 69694 14366 69746 14418
rect 75182 14366 75234 14418
rect 77870 14366 77922 14418
rect 81118 14366 81170 14418
rect 81566 14366 81618 14418
rect 20414 14254 20466 14306
rect 25230 14254 25282 14306
rect 29710 14254 29762 14306
rect 34414 14254 34466 14306
rect 34862 14254 34914 14306
rect 35310 14254 35362 14306
rect 35758 14254 35810 14306
rect 38110 14254 38162 14306
rect 39454 14254 39506 14306
rect 39902 14254 39954 14306
rect 41806 14254 41858 14306
rect 42702 14254 42754 14306
rect 46062 14254 46114 14306
rect 47742 14254 47794 14306
rect 48078 14254 48130 14306
rect 49422 14254 49474 14306
rect 49758 14254 49810 14306
rect 53006 14254 53058 14306
rect 54014 14254 54066 14306
rect 54574 14254 54626 14306
rect 57038 14254 57090 14306
rect 57486 14254 57538 14306
rect 60734 14254 60786 14306
rect 61070 14254 61122 14306
rect 61518 14254 61570 14306
rect 64094 14254 64146 14306
rect 64542 14254 64594 14306
rect 65214 14254 65266 14306
rect 66222 14254 66274 14306
rect 68574 14254 68626 14306
rect 73390 14254 73442 14306
rect 73950 14254 74002 14306
rect 74286 14254 74338 14306
rect 74846 14254 74898 14306
rect 75294 14254 75346 14306
rect 81230 14254 81282 14306
rect 81902 14254 81954 14306
rect 84030 14254 84082 14306
rect 85822 14254 85874 14306
rect 86270 14254 86322 14306
rect 90750 14254 90802 14306
rect 91086 14254 91138 14306
rect 92430 14254 92482 14306
rect 96910 14254 96962 14306
rect 97470 14254 97522 14306
rect 97806 14254 97858 14306
rect 99150 14254 99202 14306
rect 102734 14254 102786 14306
rect 106654 14254 106706 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 81278 14086 81330 14138
rect 81382 14086 81434 14138
rect 81486 14086 81538 14138
rect 111998 14086 112050 14138
rect 112102 14086 112154 14138
rect 112206 14086 112258 14138
rect 142718 14086 142770 14138
rect 142822 14086 142874 14138
rect 142926 14086 142978 14138
rect 24558 13918 24610 13970
rect 25678 13918 25730 13970
rect 30158 13918 30210 13970
rect 32510 13918 32562 13970
rect 34190 13918 34242 13970
rect 37102 13918 37154 13970
rect 41694 13918 41746 13970
rect 42142 13918 42194 13970
rect 42590 13918 42642 13970
rect 44494 13918 44546 13970
rect 44942 13918 44994 13970
rect 46398 13918 46450 13970
rect 49198 13918 49250 13970
rect 50206 13918 50258 13970
rect 50766 13918 50818 13970
rect 62862 13918 62914 13970
rect 63758 13918 63810 13970
rect 64542 13918 64594 13970
rect 66670 13918 66722 13970
rect 68910 13918 68962 13970
rect 69470 13918 69522 13970
rect 70814 13918 70866 13970
rect 71262 13918 71314 13970
rect 72382 13918 72434 13970
rect 73502 13918 73554 13970
rect 78654 13918 78706 13970
rect 79214 13918 79266 13970
rect 80334 13918 80386 13970
rect 85934 13918 85986 13970
rect 86942 13918 86994 13970
rect 87390 13918 87442 13970
rect 93102 13918 93154 13970
rect 93886 13918 93938 13970
rect 103742 13918 103794 13970
rect 107214 13918 107266 13970
rect 110574 13918 110626 13970
rect 31166 13806 31218 13858
rect 62526 13806 62578 13858
rect 65662 13806 65714 13858
rect 65774 13806 65826 13858
rect 75518 13806 75570 13858
rect 84590 13806 84642 13858
rect 93550 13806 93602 13858
rect 103630 13806 103682 13858
rect 103966 13806 104018 13858
rect 104190 13806 104242 13858
rect 104638 13806 104690 13858
rect 105198 13806 105250 13858
rect 105534 13806 105586 13858
rect 106094 13806 106146 13858
rect 106654 13806 106706 13858
rect 111470 13806 111522 13858
rect 20078 13694 20130 13746
rect 26686 13694 26738 13746
rect 29710 13694 29762 13746
rect 30382 13694 30434 13746
rect 33854 13694 33906 13746
rect 34302 13694 34354 13746
rect 34638 13694 34690 13746
rect 35310 13694 35362 13746
rect 37438 13694 37490 13746
rect 41022 13694 41074 13746
rect 45838 13694 45890 13746
rect 52670 13694 52722 13746
rect 55134 13694 55186 13746
rect 56590 13694 56642 13746
rect 56814 13694 56866 13746
rect 57150 13694 57202 13746
rect 59390 13694 59442 13746
rect 64430 13694 64482 13746
rect 64654 13694 64706 13746
rect 64990 13694 65042 13746
rect 65438 13694 65490 13746
rect 66222 13694 66274 13746
rect 69134 13694 69186 13746
rect 69582 13694 69634 13746
rect 69806 13694 69858 13746
rect 71038 13694 71090 13746
rect 71374 13694 71426 13746
rect 72494 13694 72546 13746
rect 74958 13694 75010 13746
rect 76414 13694 76466 13746
rect 77422 13694 77474 13746
rect 78206 13694 78258 13746
rect 81118 13694 81170 13746
rect 82574 13694 82626 13746
rect 82910 13694 82962 13746
rect 83918 13694 83970 13746
rect 85710 13694 85762 13746
rect 89070 13694 89122 13746
rect 90750 13694 90802 13746
rect 96014 13694 96066 13746
rect 97806 13694 97858 13746
rect 100270 13694 100322 13746
rect 102734 13694 102786 13746
rect 104526 13694 104578 13746
rect 104862 13694 104914 13746
rect 106206 13694 106258 13746
rect 107662 13694 107714 13746
rect 108222 13694 108274 13746
rect 19742 13582 19794 13634
rect 20190 13582 20242 13634
rect 20974 13582 21026 13634
rect 21422 13582 21474 13634
rect 24670 13582 24722 13634
rect 27358 13582 27410 13634
rect 29486 13582 29538 13634
rect 30270 13582 30322 13634
rect 31614 13582 31666 13634
rect 32174 13582 32226 13634
rect 33518 13582 33570 13634
rect 35086 13582 35138 13634
rect 35758 13582 35810 13634
rect 36206 13582 36258 13634
rect 36766 13582 36818 13634
rect 38222 13582 38274 13634
rect 40350 13582 40402 13634
rect 43150 13582 43202 13634
rect 43710 13582 43762 13634
rect 44158 13582 44210 13634
rect 45614 13582 45666 13634
rect 46846 13582 46898 13634
rect 47406 13582 47458 13634
rect 47742 13582 47794 13634
rect 48190 13582 48242 13634
rect 49646 13582 49698 13634
rect 50878 13582 50930 13634
rect 51886 13582 51938 13634
rect 54462 13582 54514 13634
rect 55918 13582 55970 13634
rect 56702 13582 56754 13634
rect 57598 13582 57650 13634
rect 58046 13582 58098 13634
rect 58606 13582 58658 13634
rect 58942 13582 58994 13634
rect 60062 13582 60114 13634
rect 62190 13582 62242 13634
rect 63310 13582 63362 13634
rect 64990 13582 65042 13634
rect 20414 13470 20466 13522
rect 31278 13470 31330 13522
rect 31614 13470 31666 13522
rect 34190 13470 34242 13522
rect 67230 13582 67282 13634
rect 67678 13582 67730 13634
rect 68126 13582 68178 13634
rect 70366 13582 70418 13634
rect 72942 13582 72994 13634
rect 73950 13582 74002 13634
rect 74398 13582 74450 13634
rect 79326 13582 79378 13634
rect 80782 13582 80834 13634
rect 86494 13582 86546 13634
rect 88062 13582 88114 13634
rect 88846 13582 88898 13634
rect 90526 13582 90578 13634
rect 92654 13582 92706 13634
rect 95230 13582 95282 13634
rect 95902 13582 95954 13634
rect 98030 13582 98082 13634
rect 102062 13582 102114 13634
rect 105086 13582 105138 13634
rect 112030 13582 112082 13634
rect 34974 13470 35026 13522
rect 35534 13470 35586 13522
rect 36318 13470 36370 13522
rect 41806 13470 41858 13522
rect 43150 13470 43202 13522
rect 43934 13470 43986 13522
rect 44830 13470 44882 13522
rect 45502 13470 45554 13522
rect 46062 13470 46114 13522
rect 47070 13470 47122 13522
rect 47742 13470 47794 13522
rect 48078 13470 48130 13522
rect 49310 13470 49362 13522
rect 49758 13470 49810 13522
rect 63086 13470 63138 13522
rect 63310 13470 63362 13522
rect 65214 13470 65266 13522
rect 72382 13470 72434 13522
rect 73390 13470 73442 13522
rect 73838 13470 73890 13522
rect 89182 13470 89234 13522
rect 92654 13470 92706 13522
rect 93438 13470 93490 13522
rect 94670 13470 94722 13522
rect 98814 13470 98866 13522
rect 102622 13470 102674 13522
rect 103182 13470 103234 13522
rect 105646 13470 105698 13522
rect 106094 13470 106146 13522
rect 111582 13470 111634 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 96638 13302 96690 13354
rect 96742 13302 96794 13354
rect 96846 13302 96898 13354
rect 127358 13302 127410 13354
rect 127462 13302 127514 13354
rect 127566 13302 127618 13354
rect 158078 13302 158130 13354
rect 158182 13302 158234 13354
rect 158286 13302 158338 13354
rect 20190 13134 20242 13186
rect 27022 13134 27074 13186
rect 31950 13134 32002 13186
rect 32510 13134 32562 13186
rect 39118 13134 39170 13186
rect 39678 13134 39730 13186
rect 61742 13134 61794 13186
rect 97358 13134 97410 13186
rect 100158 13134 100210 13186
rect 19854 13022 19906 13074
rect 21870 13022 21922 13074
rect 25454 13022 25506 13074
rect 26126 13022 26178 13074
rect 26574 13022 26626 13074
rect 34302 13022 34354 13074
rect 36430 13022 36482 13074
rect 38222 13022 38274 13074
rect 38782 13022 38834 13074
rect 39678 13022 39730 13074
rect 40686 13022 40738 13074
rect 43934 13022 43986 13074
rect 44830 13022 44882 13074
rect 48862 13022 48914 13074
rect 50430 13022 50482 13074
rect 58718 13022 58770 13074
rect 59502 13022 59554 13074
rect 60622 13022 60674 13074
rect 62302 13022 62354 13074
rect 62750 13022 62802 13074
rect 63422 13022 63474 13074
rect 66670 13022 66722 13074
rect 68798 13022 68850 13074
rect 72718 13022 72770 13074
rect 74174 13022 74226 13074
rect 92318 13022 92370 13074
rect 100718 13022 100770 13074
rect 103518 13022 103570 13074
rect 108222 13022 108274 13074
rect 108670 13022 108722 13074
rect 109118 13022 109170 13074
rect 19742 12910 19794 12962
rect 20078 12910 20130 12962
rect 20302 12910 20354 12962
rect 22654 12910 22706 12962
rect 26686 12910 26738 12962
rect 27134 12910 27186 12962
rect 29374 12910 29426 12962
rect 29822 12910 29874 12962
rect 30382 12910 30434 12962
rect 30830 12910 30882 12962
rect 31390 12910 31442 12962
rect 31614 12910 31666 12962
rect 31950 12910 32002 12962
rect 32510 12910 32562 12962
rect 33630 12910 33682 12962
rect 37214 12910 37266 12962
rect 37774 12910 37826 12962
rect 38110 12910 38162 12962
rect 38334 12910 38386 12962
rect 41022 12910 41074 12962
rect 47742 12910 47794 12962
rect 48302 12910 48354 12962
rect 48750 12910 48802 12962
rect 49758 12910 49810 12962
rect 49982 12910 50034 12962
rect 53006 12910 53058 12962
rect 53790 12910 53842 12962
rect 54350 12910 54402 12962
rect 58382 12910 58434 12962
rect 60510 12910 60562 12962
rect 60846 12910 60898 12962
rect 61070 12910 61122 12962
rect 63870 12910 63922 12962
rect 69918 12910 69970 12962
rect 77198 12910 77250 12962
rect 78542 12910 78594 12962
rect 79886 12910 79938 12962
rect 80222 12910 80274 12962
rect 81566 12910 81618 12962
rect 83134 12910 83186 12962
rect 84814 12910 84866 12962
rect 86046 12910 86098 12962
rect 88286 12910 88338 12962
rect 88734 12910 88786 12962
rect 88958 12910 89010 12962
rect 90526 12910 90578 12962
rect 92542 12910 92594 12962
rect 93998 12910 94050 12962
rect 94558 12910 94610 12962
rect 95902 12910 95954 12962
rect 96238 12910 96290 12962
rect 96350 12910 96402 12962
rect 100606 12910 100658 12962
rect 100830 12910 100882 12962
rect 102398 12910 102450 12962
rect 107550 12910 107602 12962
rect 109566 12910 109618 12962
rect 110014 12910 110066 12962
rect 110686 12910 110738 12962
rect 112142 12910 112194 12962
rect 19406 12798 19458 12850
rect 23326 12798 23378 12850
rect 26462 12798 26514 12850
rect 29934 12798 29986 12850
rect 30942 12798 30994 12850
rect 32846 12798 32898 12850
rect 36990 12798 37042 12850
rect 41806 12798 41858 12850
rect 46958 12798 47010 12850
rect 49310 12798 49362 12850
rect 55022 12798 55074 12850
rect 57710 12798 57762 12850
rect 57934 12798 57986 12850
rect 61630 12798 61682 12850
rect 64542 12798 64594 12850
rect 70590 12798 70642 12850
rect 74958 12798 75010 12850
rect 76190 12798 76242 12850
rect 78094 12798 78146 12850
rect 82798 12798 82850 12850
rect 84254 12798 84306 12850
rect 87726 12798 87778 12850
rect 90078 12798 90130 12850
rect 91086 12798 91138 12850
rect 93102 12798 93154 12850
rect 100158 12798 100210 12850
rect 100270 12798 100322 12850
rect 101054 12798 101106 12850
rect 111694 12798 111746 12850
rect 112702 12798 112754 12850
rect 19070 12686 19122 12738
rect 29598 12686 29650 12738
rect 29710 12686 29762 12738
rect 30606 12686 30658 12738
rect 30718 12686 30770 12738
rect 31838 12686 31890 12738
rect 39342 12686 39394 12738
rect 40350 12686 40402 12738
rect 48526 12686 48578 12738
rect 48862 12686 48914 12738
rect 49534 12686 49586 12738
rect 49646 12686 49698 12738
rect 51102 12686 51154 12738
rect 51662 12686 51714 12738
rect 52222 12686 52274 12738
rect 53454 12686 53506 12738
rect 53678 12686 53730 12738
rect 53902 12686 53954 12738
rect 57262 12686 57314 12738
rect 58046 12686 58098 12738
rect 60062 12686 60114 12738
rect 61742 12686 61794 12738
rect 67566 12686 67618 12738
rect 69134 12686 69186 12738
rect 73278 12686 73330 12738
rect 73726 12686 73778 12738
rect 74622 12686 74674 12738
rect 75294 12686 75346 12738
rect 76302 12686 76354 12738
rect 83470 12686 83522 12738
rect 87950 12686 88002 12738
rect 89294 12686 89346 12738
rect 89742 12686 89794 12738
rect 90526 12686 90578 12738
rect 91982 12686 92034 12738
rect 92766 12686 92818 12738
rect 92990 12686 93042 12738
rect 93550 12686 93602 12738
rect 98366 12686 98418 12738
rect 98814 12686 98866 12738
rect 107662 12686 107714 12738
rect 107886 12686 107938 12738
rect 110798 12686 110850 12738
rect 111246 12686 111298 12738
rect 113038 12686 113090 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 81278 12518 81330 12570
rect 81382 12518 81434 12570
rect 81486 12518 81538 12570
rect 111998 12518 112050 12570
rect 112102 12518 112154 12570
rect 112206 12518 112258 12570
rect 142718 12518 142770 12570
rect 142822 12518 142874 12570
rect 142926 12518 142978 12570
rect 18174 12350 18226 12402
rect 18622 12350 18674 12402
rect 18958 12350 19010 12402
rect 21198 12350 21250 12402
rect 21982 12350 22034 12402
rect 23998 12350 24050 12402
rect 24110 12350 24162 12402
rect 27246 12350 27298 12402
rect 27358 12350 27410 12402
rect 29486 12350 29538 12402
rect 36654 12350 36706 12402
rect 37774 12350 37826 12402
rect 39902 12350 39954 12402
rect 40798 12350 40850 12402
rect 43822 12350 43874 12402
rect 45614 12350 45666 12402
rect 46398 12350 46450 12402
rect 47182 12350 47234 12402
rect 47518 12350 47570 12402
rect 47966 12350 48018 12402
rect 49646 12350 49698 12402
rect 54462 12350 54514 12402
rect 19518 12238 19570 12290
rect 19742 12238 19794 12290
rect 21310 12238 21362 12290
rect 21534 12238 21586 12290
rect 22430 12238 22482 12290
rect 25790 12238 25842 12290
rect 26238 12238 26290 12290
rect 29150 12238 29202 12290
rect 29710 12238 29762 12290
rect 31726 12238 31778 12290
rect 32398 12238 32450 12290
rect 37326 12238 37378 12290
rect 37886 12238 37938 12290
rect 42366 12238 42418 12290
rect 42702 12238 42754 12290
rect 45950 12238 46002 12290
rect 48750 12238 48802 12290
rect 19630 12126 19682 12178
rect 20190 12126 20242 12178
rect 20974 12126 21026 12178
rect 21758 12126 21810 12178
rect 22206 12126 22258 12178
rect 22878 12126 22930 12178
rect 23886 12126 23938 12178
rect 24558 12126 24610 12178
rect 25230 12126 25282 12178
rect 25342 12126 25394 12178
rect 25566 12126 25618 12178
rect 29374 12126 29426 12178
rect 30270 12126 30322 12178
rect 31390 12126 31442 12178
rect 32174 12126 32226 12178
rect 35982 12126 36034 12178
rect 36990 12126 37042 12178
rect 37662 12126 37714 12178
rect 40910 12126 40962 12178
rect 41918 12126 41970 12178
rect 42814 12126 42866 12178
rect 43598 12126 43650 12178
rect 44046 12126 44098 12178
rect 44270 12126 44322 12178
rect 44830 12126 44882 12178
rect 45166 12126 45218 12178
rect 45614 12126 45666 12178
rect 46174 12126 46226 12178
rect 46622 12126 46674 12178
rect 49086 12126 49138 12178
rect 49310 12126 49362 12178
rect 18958 12014 19010 12066
rect 19966 12014 20018 12066
rect 28702 12014 28754 12066
rect 32510 12014 32562 12066
rect 34414 12014 34466 12066
rect 38782 12014 38834 12066
rect 39454 12014 39506 12066
rect 40238 12014 40290 12066
rect 46286 12014 46338 12066
rect 19182 11902 19234 11954
rect 27134 11902 27186 11954
rect 40350 11902 40402 11954
rect 43710 11902 43762 11954
rect 45390 11902 45442 11954
rect 54910 12350 54962 12402
rect 56030 12350 56082 12402
rect 59838 12350 59890 12402
rect 60510 12350 60562 12402
rect 60846 12350 60898 12402
rect 64878 12350 64930 12402
rect 70366 12350 70418 12402
rect 73726 12350 73778 12402
rect 78430 12350 78482 12402
rect 84926 12350 84978 12402
rect 85710 12350 85762 12402
rect 88062 12350 88114 12402
rect 90302 12350 90354 12402
rect 90974 12350 91026 12402
rect 104862 12350 104914 12402
rect 105982 12350 106034 12402
rect 109342 12350 109394 12402
rect 110350 12350 110402 12402
rect 110798 12350 110850 12402
rect 113822 12350 113874 12402
rect 49758 12238 49810 12290
rect 50206 12238 50258 12290
rect 50542 12238 50594 12290
rect 54686 12238 54738 12290
rect 55246 12238 55298 12290
rect 57598 12238 57650 12290
rect 61294 12238 61346 12290
rect 65102 12238 65154 12290
rect 75406 12238 75458 12290
rect 77870 12238 77922 12290
rect 79438 12238 79490 12290
rect 83246 12238 83298 12290
rect 84366 12238 84418 12290
rect 85822 12238 85874 12290
rect 88510 12238 88562 12290
rect 89406 12238 89458 12290
rect 90414 12238 90466 12290
rect 93998 12238 94050 12290
rect 104078 12238 104130 12290
rect 105646 12238 105698 12290
rect 106318 12238 106370 12290
rect 106654 12238 106706 12290
rect 106990 12238 107042 12290
rect 107438 12238 107490 12290
rect 107998 12238 108050 12290
rect 108558 12238 108610 12290
rect 51102 12126 51154 12178
rect 54910 12126 54962 12178
rect 56926 12126 56978 12178
rect 64654 12126 64706 12178
rect 65214 12126 65266 12178
rect 68910 12126 68962 12178
rect 69918 12126 69970 12178
rect 70254 12126 70306 12178
rect 70478 12126 70530 12178
rect 74510 12126 74562 12178
rect 76302 12126 76354 12178
rect 78206 12126 78258 12178
rect 79214 12126 79266 12178
rect 79550 12126 79602 12178
rect 80110 12126 80162 12178
rect 81454 12126 81506 12178
rect 83022 12126 83074 12178
rect 84702 12126 84754 12178
rect 86158 12126 86210 12178
rect 89182 12126 89234 12178
rect 90638 12126 90690 12178
rect 91310 12126 91362 12178
rect 91534 12126 91586 12178
rect 94782 12126 94834 12178
rect 96126 12126 96178 12178
rect 97806 12126 97858 12178
rect 102622 12126 102674 12178
rect 102958 12126 103010 12178
rect 103966 12126 104018 12178
rect 104302 12126 104354 12178
rect 104638 12126 104690 12178
rect 105310 12126 105362 12178
rect 107326 12126 107378 12178
rect 107662 12126 107714 12178
rect 108110 12126 108162 12178
rect 108446 12126 108498 12178
rect 109454 12126 109506 12178
rect 51774 12014 51826 12066
rect 53902 12014 53954 12066
rect 61742 12014 61794 12066
rect 62638 12014 62690 12066
rect 62974 12014 63026 12066
rect 63422 12014 63474 12066
rect 63870 12014 63922 12066
rect 65998 12014 66050 12066
rect 68126 12014 68178 12066
rect 69582 12014 69634 12066
rect 71262 12014 71314 12066
rect 71710 12014 71762 12066
rect 72382 12014 72434 12066
rect 72830 12014 72882 12066
rect 73390 12014 73442 12066
rect 74286 12014 74338 12066
rect 87278 12014 87330 12066
rect 91870 12014 91922 12066
rect 95230 12014 95282 12066
rect 95902 12014 95954 12066
rect 98142 12014 98194 12066
rect 99710 12014 99762 12066
rect 101838 12014 101890 12066
rect 103070 12014 103122 12066
rect 109902 12014 109954 12066
rect 111582 12014 111634 12066
rect 112030 12014 112082 12066
rect 112478 12014 112530 12066
rect 112926 12014 112978 12066
rect 113374 12014 113426 12066
rect 49758 11902 49810 11954
rect 61182 11902 61234 11954
rect 61742 11902 61794 11954
rect 64318 11902 64370 11954
rect 64542 11902 64594 11954
rect 72382 11902 72434 11954
rect 72942 11902 72994 11954
rect 85710 11902 85762 11954
rect 98814 11902 98866 11954
rect 107998 11902 108050 11954
rect 108558 11902 108610 11954
rect 109342 11902 109394 11954
rect 111582 11902 111634 11954
rect 112590 11902 112642 11954
rect 113374 11902 113426 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 96638 11734 96690 11786
rect 96742 11734 96794 11786
rect 96846 11734 96898 11786
rect 127358 11734 127410 11786
rect 127462 11734 127514 11786
rect 127566 11734 127618 11786
rect 158078 11734 158130 11786
rect 158182 11734 158234 11786
rect 158286 11734 158338 11786
rect 20302 11566 20354 11618
rect 27582 11566 27634 11618
rect 42926 11566 42978 11618
rect 45950 11566 46002 11618
rect 46398 11566 46450 11618
rect 60622 11566 60674 11618
rect 62974 11566 63026 11618
rect 63310 11566 63362 11618
rect 63534 11566 63586 11618
rect 63982 11566 64034 11618
rect 64654 11566 64706 11618
rect 67006 11566 67058 11618
rect 68910 11566 68962 11618
rect 69134 11566 69186 11618
rect 73278 11566 73330 11618
rect 93550 11566 93602 11618
rect 112702 11566 112754 11618
rect 113486 11566 113538 11618
rect 114382 11566 114434 11618
rect 114830 11566 114882 11618
rect 15598 11454 15650 11506
rect 17726 11454 17778 11506
rect 21310 11454 21362 11506
rect 22542 11454 22594 11506
rect 28702 11454 28754 11506
rect 33518 11454 33570 11506
rect 41806 11454 41858 11506
rect 47854 11454 47906 11506
rect 50766 11454 50818 11506
rect 51662 11454 51714 11506
rect 52110 11454 52162 11506
rect 52782 11454 52834 11506
rect 58718 11454 58770 11506
rect 63534 11454 63586 11506
rect 64878 11454 64930 11506
rect 71038 11454 71090 11506
rect 18510 11342 18562 11394
rect 19742 11342 19794 11394
rect 20078 11342 20130 11394
rect 20526 11342 20578 11394
rect 24782 11342 24834 11394
rect 34414 11342 34466 11394
rect 41134 11342 41186 11394
rect 42254 11342 42306 11394
rect 42926 11342 42978 11394
rect 48526 11342 48578 11394
rect 50094 11342 50146 11394
rect 52670 11342 52722 11394
rect 53006 11342 53058 11394
rect 53230 11342 53282 11394
rect 53566 11342 53618 11394
rect 53790 11342 53842 11394
rect 54574 11342 54626 11394
rect 61406 11342 61458 11394
rect 65438 11342 65490 11394
rect 65886 11342 65938 11394
rect 66334 11342 66386 11394
rect 66446 11342 66498 11394
rect 70142 11342 70194 11394
rect 71598 11342 71650 11394
rect 77086 11454 77138 11506
rect 89070 11454 89122 11506
rect 95230 11454 95282 11506
rect 99150 11454 99202 11506
rect 100606 11454 100658 11506
rect 102958 11454 103010 11506
rect 112590 11454 112642 11506
rect 113486 11454 113538 11506
rect 114382 11454 114434 11506
rect 114830 11454 114882 11506
rect 73054 11342 73106 11394
rect 73278 11342 73330 11394
rect 74398 11342 74450 11394
rect 74846 11342 74898 11394
rect 74958 11342 75010 11394
rect 76078 11342 76130 11394
rect 76750 11342 76802 11394
rect 76974 11342 77026 11394
rect 77198 11342 77250 11394
rect 77422 11342 77474 11394
rect 81902 11342 81954 11394
rect 84142 11342 84194 11394
rect 84814 11342 84866 11394
rect 86270 11342 86322 11394
rect 88510 11342 88562 11394
rect 89182 11342 89234 11394
rect 89854 11342 89906 11394
rect 91982 11342 92034 11394
rect 92318 11342 92370 11394
rect 92654 11342 92706 11394
rect 94110 11342 94162 11394
rect 94558 11342 94610 11394
rect 95566 11342 95618 11394
rect 96910 11342 96962 11394
rect 100270 11342 100322 11394
rect 100382 11342 100434 11394
rect 101278 11342 101330 11394
rect 105870 11342 105922 11394
rect 106430 11342 106482 11394
rect 107774 11342 107826 11394
rect 108558 11342 108610 11394
rect 109230 11342 109282 11394
rect 109902 11342 109954 11394
rect 111022 11342 111074 11394
rect 19070 11230 19122 11282
rect 19406 11230 19458 11282
rect 21422 11230 21474 11282
rect 21646 11230 21698 11282
rect 36318 11230 36370 11282
rect 36430 11230 36482 11282
rect 37326 11230 37378 11282
rect 37662 11230 37714 11282
rect 39006 11230 39058 11282
rect 39118 11230 39170 11282
rect 39342 11230 39394 11282
rect 40686 11230 40738 11282
rect 41246 11230 41298 11282
rect 42590 11230 42642 11282
rect 48190 11230 48242 11282
rect 48750 11230 48802 11282
rect 49534 11230 49586 11282
rect 54126 11230 54178 11282
rect 60510 11230 60562 11282
rect 61630 11230 61682 11282
rect 66894 11230 66946 11282
rect 67006 11230 67058 11282
rect 71934 11230 71986 11282
rect 72718 11230 72770 11282
rect 76302 11230 76354 11282
rect 76414 11230 76466 11282
rect 78990 11230 79042 11282
rect 84030 11230 84082 11282
rect 84478 11230 84530 11282
rect 86942 11230 86994 11282
rect 87726 11230 87778 11282
rect 89406 11230 89458 11282
rect 90974 11230 91026 11282
rect 93102 11230 93154 11282
rect 93662 11230 93714 11282
rect 97246 11230 97298 11282
rect 100718 11230 100770 11282
rect 102510 11230 102562 11282
rect 102622 11286 102674 11338
rect 112142 11342 112194 11394
rect 105086 11230 105138 11282
rect 106206 11230 106258 11282
rect 107550 11230 107602 11282
rect 108110 11230 108162 11282
rect 108782 11230 108834 11282
rect 110686 11230 110738 11282
rect 111470 11230 111522 11282
rect 20190 11118 20242 11170
rect 22094 11118 22146 11170
rect 24446 11118 24498 11170
rect 25342 11118 25394 11170
rect 26014 11118 26066 11170
rect 27694 11118 27746 11170
rect 27806 11118 27858 11170
rect 29262 11118 29314 11170
rect 29934 11118 29986 11170
rect 30270 11118 30322 11170
rect 36094 11118 36146 11170
rect 36990 11118 37042 11170
rect 37998 11118 38050 11170
rect 38334 11118 38386 11170
rect 38670 11118 38722 11170
rect 39790 11118 39842 11170
rect 40126 11118 40178 11170
rect 40350 11118 40402 11170
rect 40574 11118 40626 11170
rect 43822 11118 43874 11170
rect 44270 11118 44322 11170
rect 45054 11118 45106 11170
rect 45502 11118 45554 11170
rect 45838 11118 45890 11170
rect 46286 11118 46338 11170
rect 46958 11118 47010 11170
rect 47406 11118 47458 11170
rect 49086 11118 49138 11170
rect 50318 11118 50370 11170
rect 51214 11118 51266 11170
rect 53678 11118 53730 11170
rect 61966 11118 62018 11170
rect 62078 11118 62130 11170
rect 62190 11118 62242 11170
rect 62414 11118 62466 11170
rect 62974 11118 63026 11170
rect 63982 11118 64034 11170
rect 64318 11118 64370 11170
rect 65102 11118 65154 11170
rect 66222 11118 66274 11170
rect 67902 11118 67954 11170
rect 68574 11118 68626 11170
rect 69022 11118 69074 11170
rect 69358 11118 69410 11170
rect 69806 11118 69858 11170
rect 70478 11118 70530 11170
rect 71262 11118 71314 11170
rect 71486 11118 71538 11170
rect 72046 11118 72098 11170
rect 72270 11118 72322 11170
rect 72830 11118 72882 11170
rect 73614 11118 73666 11170
rect 73950 11118 74002 11170
rect 74622 11118 74674 11170
rect 75630 11118 75682 11170
rect 90190 11118 90242 11170
rect 90638 11118 90690 11170
rect 90862 11118 90914 11170
rect 92430 11118 92482 11170
rect 92766 11118 92818 11170
rect 92990 11118 93042 11170
rect 93550 11118 93602 11170
rect 96350 11118 96402 11170
rect 96574 11118 96626 11170
rect 96798 11118 96850 11170
rect 97358 11118 97410 11170
rect 97806 11118 97858 11170
rect 98254 11118 98306 11170
rect 98702 11118 98754 11170
rect 99822 11118 99874 11170
rect 100942 11118 100994 11170
rect 101166 11118 101218 11170
rect 101614 11118 101666 11170
rect 101950 11118 102002 11170
rect 102286 11118 102338 11170
rect 106990 11118 107042 11170
rect 107998 11118 108050 11170
rect 109454 11118 109506 11170
rect 110126 11118 110178 11170
rect 110798 11118 110850 11170
rect 111582 11118 111634 11170
rect 111806 11118 111858 11170
rect 113038 11118 113090 11170
rect 114046 11118 114098 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 81278 10950 81330 11002
rect 81382 10950 81434 11002
rect 81486 10950 81538 11002
rect 111998 10950 112050 11002
rect 112102 10950 112154 11002
rect 112206 10950 112258 11002
rect 142718 10950 142770 11002
rect 142822 10950 142874 11002
rect 142926 10950 142978 11002
rect 21646 10782 21698 10834
rect 22878 10782 22930 10834
rect 23886 10782 23938 10834
rect 28366 10782 28418 10834
rect 31502 10782 31554 10834
rect 33966 10782 34018 10834
rect 35198 10782 35250 10834
rect 35422 10782 35474 10834
rect 35534 10782 35586 10834
rect 37550 10782 37602 10834
rect 41358 10782 41410 10834
rect 42590 10782 42642 10834
rect 43038 10782 43090 10834
rect 46846 10782 46898 10834
rect 54126 10782 54178 10834
rect 54462 10782 54514 10834
rect 54798 10782 54850 10834
rect 55470 10782 55522 10834
rect 55582 10782 55634 10834
rect 56702 10782 56754 10834
rect 56814 10782 56866 10834
rect 56926 10782 56978 10834
rect 58046 10782 58098 10834
rect 58158 10782 58210 10834
rect 59278 10782 59330 10834
rect 66334 10782 66386 10834
rect 76974 10782 77026 10834
rect 18174 10670 18226 10722
rect 20638 10670 20690 10722
rect 20974 10670 21026 10722
rect 24670 10670 24722 10722
rect 25342 10670 25394 10722
rect 26910 10670 26962 10722
rect 31614 10670 31666 10722
rect 32398 10670 32450 10722
rect 33406 10670 33458 10722
rect 34974 10670 35026 10722
rect 38782 10670 38834 10722
rect 38894 10670 38946 10722
rect 39678 10670 39730 10722
rect 40350 10670 40402 10722
rect 41918 10670 41970 10722
rect 42142 10670 42194 10722
rect 46174 10670 46226 10722
rect 53790 10670 53842 10722
rect 57598 10670 57650 10722
rect 58718 10670 58770 10722
rect 58830 10670 58882 10722
rect 63422 10726 63474 10778
rect 77198 10782 77250 10834
rect 77310 10782 77362 10834
rect 77870 10782 77922 10834
rect 78206 10782 78258 10834
rect 78766 10782 78818 10834
rect 80446 10782 80498 10834
rect 83918 10782 83970 10834
rect 85038 10782 85090 10834
rect 85822 10782 85874 10834
rect 86382 10782 86434 10834
rect 88286 10782 88338 10834
rect 93662 10782 93714 10834
rect 95678 10782 95730 10834
rect 102846 10782 102898 10834
rect 109790 10782 109842 10834
rect 110910 10782 110962 10834
rect 64878 10670 64930 10722
rect 64990 10670 65042 10722
rect 67230 10670 67282 10722
rect 74398 10670 74450 10722
rect 79214 10670 79266 10722
rect 84478 10670 84530 10722
rect 84590 10670 84642 10722
rect 91310 10670 91362 10722
rect 92654 10670 92706 10722
rect 95790 10670 95842 10722
rect 99822 10670 99874 10722
rect 101502 10670 101554 10722
rect 102174 10670 102226 10722
rect 109454 10670 109506 10722
rect 109678 10670 109730 10722
rect 110014 10670 110066 10722
rect 17502 10558 17554 10610
rect 21422 10558 21474 10610
rect 22094 10558 22146 10610
rect 23550 10558 23602 10610
rect 24110 10558 24162 10610
rect 24446 10558 24498 10610
rect 26574 10558 26626 10610
rect 27246 10558 27298 10610
rect 27582 10558 27634 10610
rect 28030 10558 28082 10610
rect 30382 10558 30434 10610
rect 31390 10558 31442 10610
rect 32062 10558 32114 10610
rect 33070 10558 33122 10610
rect 34190 10558 34242 10610
rect 35982 10558 36034 10610
rect 36542 10558 36594 10610
rect 39118 10558 39170 10610
rect 39454 10558 39506 10610
rect 40014 10558 40066 10610
rect 41358 10558 41410 10610
rect 44270 10558 44322 10610
rect 44606 10558 44658 10610
rect 44830 10558 44882 10610
rect 46062 10558 46114 10610
rect 46734 10558 46786 10610
rect 47630 10558 47682 10610
rect 48190 10558 48242 10610
rect 48974 10558 49026 10610
rect 49198 10558 49250 10610
rect 49982 10558 50034 10610
rect 50206 10558 50258 10610
rect 55694 10558 55746 10610
rect 56142 10558 56194 10610
rect 57262 10558 57314 10610
rect 57822 10558 57874 10610
rect 59390 10558 59442 10610
rect 60062 10558 60114 10610
rect 63310 10558 63362 10610
rect 64654 10558 64706 10610
rect 65438 10558 65490 10610
rect 66558 10558 66610 10610
rect 67566 10558 67618 10610
rect 68910 10558 68962 10610
rect 72494 10558 72546 10610
rect 72718 10558 72770 10610
rect 73726 10558 73778 10610
rect 77086 10558 77138 10610
rect 77534 10558 77586 10610
rect 79102 10558 79154 10610
rect 79662 10558 79714 10610
rect 80110 10558 80162 10610
rect 82910 10558 82962 10610
rect 83806 10558 83858 10610
rect 85486 10558 85538 10610
rect 85710 10558 85762 10610
rect 86046 10558 86098 10610
rect 86942 10558 86994 10610
rect 88734 10558 88786 10610
rect 89518 10558 89570 10610
rect 90078 10558 90130 10610
rect 92206 10558 92258 10610
rect 92430 10558 92482 10610
rect 92766 10558 92818 10610
rect 94334 10558 94386 10610
rect 94558 10558 94610 10610
rect 95342 10558 95394 10610
rect 96126 10558 96178 10610
rect 97470 10558 97522 10610
rect 99262 10558 99314 10610
rect 100382 10558 100434 10610
rect 100606 10558 100658 10610
rect 100942 10558 100994 10610
rect 101166 10558 101218 10610
rect 101838 10558 101890 10610
rect 102622 10558 102674 10610
rect 103630 10558 103682 10610
rect 111582 10558 111634 10610
rect 112702 10558 112754 10610
rect 20302 10446 20354 10498
rect 26126 10446 26178 10498
rect 27022 10446 27074 10498
rect 29150 10446 29202 10498
rect 29598 10446 29650 10498
rect 30046 10446 30098 10498
rect 34638 10446 34690 10498
rect 35310 10446 35362 10498
rect 36990 10446 37042 10498
rect 38446 10446 38498 10498
rect 40238 10446 40290 10498
rect 41134 10446 41186 10498
rect 43486 10446 43538 10498
rect 43822 10446 43874 10498
rect 44382 10446 44434 10498
rect 45614 10446 45666 10498
rect 48862 10446 48914 10498
rect 51550 10446 51602 10498
rect 51886 10446 51938 10498
rect 52334 10446 52386 10498
rect 52894 10446 52946 10498
rect 53342 10446 53394 10498
rect 57934 10446 57986 10498
rect 60846 10446 60898 10498
rect 62974 10446 63026 10498
rect 65886 10446 65938 10498
rect 67006 10446 67058 10498
rect 68574 10446 68626 10498
rect 69582 10446 69634 10498
rect 71710 10446 71762 10498
rect 73278 10446 73330 10498
rect 76526 10446 76578 10498
rect 79438 10446 79490 10498
rect 81902 10446 81954 10498
rect 84926 10446 84978 10498
rect 87278 10446 87330 10498
rect 93102 10446 93154 10498
rect 94222 10446 94274 10498
rect 100718 10446 100770 10498
rect 105982 10446 106034 10498
rect 110350 10446 110402 10498
rect 112142 10446 112194 10498
rect 113374 10446 113426 10498
rect 115502 10446 115554 10498
rect 115950 10446 116002 10498
rect 116398 10446 116450 10498
rect 24222 10334 24274 10386
rect 25230 10334 25282 10386
rect 25566 10334 25618 10386
rect 27470 10334 27522 10386
rect 29262 10334 29314 10386
rect 29822 10334 29874 10386
rect 37886 10334 37938 10386
rect 38222 10334 38274 10386
rect 41582 10334 41634 10386
rect 42366 10334 42418 10386
rect 43150 10334 43202 10386
rect 43934 10334 43986 10386
rect 44830 10334 44882 10386
rect 50654 10334 50706 10386
rect 58718 10334 58770 10386
rect 59278 10334 59330 10386
rect 63422 10334 63474 10386
rect 83918 10334 83970 10386
rect 84478 10334 84530 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 96638 10166 96690 10218
rect 96742 10166 96794 10218
rect 96846 10166 96898 10218
rect 127358 10166 127410 10218
rect 127462 10166 127514 10218
rect 127566 10166 127618 10218
rect 158078 10166 158130 10218
rect 158182 10166 158234 10218
rect 158286 10166 158338 10218
rect 19406 9998 19458 10050
rect 19630 9998 19682 10050
rect 45054 9998 45106 10050
rect 45950 9998 46002 10050
rect 59838 9998 59890 10050
rect 64094 9998 64146 10050
rect 66110 9998 66162 10050
rect 67902 9998 67954 10050
rect 116062 9998 116114 10050
rect 117070 9998 117122 10050
rect 18846 9886 18898 9938
rect 19630 9886 19682 9938
rect 20302 9886 20354 9938
rect 21534 9886 21586 9938
rect 22990 9886 23042 9938
rect 25118 9886 25170 9938
rect 26238 9886 26290 9938
rect 30494 9886 30546 9938
rect 31166 9886 31218 9938
rect 40798 9886 40850 9938
rect 42590 9886 42642 9938
rect 43150 9886 43202 9938
rect 45166 9886 45218 9938
rect 47742 9886 47794 9938
rect 50206 9886 50258 9938
rect 53566 9886 53618 9938
rect 55694 9886 55746 9938
rect 56702 9886 56754 9938
rect 58270 9886 58322 9938
rect 59054 9886 59106 9938
rect 60846 9886 60898 9938
rect 66110 9886 66162 9938
rect 67790 9886 67842 9938
rect 70254 9886 70306 9938
rect 75182 9886 75234 9938
rect 78542 9886 78594 9938
rect 80670 9886 80722 9938
rect 81902 9886 81954 9938
rect 85486 9886 85538 9938
rect 94222 9886 94274 9938
rect 97582 9886 97634 9938
rect 99710 9886 99762 9938
rect 101838 9886 101890 9938
rect 104862 9886 104914 9938
rect 109230 9886 109282 9938
rect 116062 9886 116114 9938
rect 22318 9774 22370 9826
rect 25454 9774 25506 9826
rect 29934 9774 29986 9826
rect 30270 9774 30322 9826
rect 30830 9774 30882 9826
rect 31838 9774 31890 9826
rect 32398 9774 32450 9826
rect 33518 9774 33570 9826
rect 34078 9774 34130 9826
rect 35534 9774 35586 9826
rect 36318 9774 36370 9826
rect 37326 9774 37378 9826
rect 37662 9774 37714 9826
rect 38110 9774 38162 9826
rect 43598 9774 43650 9826
rect 45390 9774 45442 9826
rect 46734 9774 46786 9826
rect 48526 9774 48578 9826
rect 48638 9774 48690 9826
rect 49198 9774 49250 9826
rect 49758 9774 49810 9826
rect 50542 9774 50594 9826
rect 52782 9774 52834 9826
rect 56814 9774 56866 9826
rect 57038 9774 57090 9826
rect 57934 9774 57986 9826
rect 58158 9774 58210 9826
rect 59950 9774 60002 9826
rect 61294 9774 61346 9826
rect 62526 9774 62578 9826
rect 63422 9774 63474 9826
rect 63758 9774 63810 9826
rect 67454 9774 67506 9826
rect 70590 9774 70642 9826
rect 72942 9774 72994 9826
rect 73390 9774 73442 9826
rect 73726 9774 73778 9826
rect 74846 9774 74898 9826
rect 75294 9774 75346 9826
rect 75406 9774 75458 9826
rect 76190 9774 76242 9826
rect 81454 9774 81506 9826
rect 82350 9774 82402 9826
rect 83246 9774 83298 9826
rect 83582 9774 83634 9826
rect 84590 9774 84642 9826
rect 86158 9774 86210 9826
rect 86830 9774 86882 9826
rect 87838 9774 87890 9826
rect 89630 9774 89682 9826
rect 91198 9774 91250 9826
rect 91870 9774 91922 9826
rect 92206 9774 92258 9826
rect 92542 9774 92594 9826
rect 92654 9774 92706 9826
rect 93774 9774 93826 9826
rect 93998 9774 94050 9826
rect 95230 9774 95282 9826
rect 96686 9774 96738 9826
rect 99150 9774 99202 9826
rect 102622 9774 102674 9826
rect 103070 9774 103122 9826
rect 103742 9774 103794 9826
rect 104526 9774 104578 9826
rect 104638 9774 104690 9826
rect 105870 9774 105922 9826
rect 106766 9774 106818 9826
rect 107102 9774 107154 9826
rect 107662 9774 107714 9826
rect 107998 9774 108050 9826
rect 108222 9774 108274 9826
rect 112142 9774 112194 9826
rect 113150 9774 113202 9826
rect 113710 9774 113762 9826
rect 114158 9774 114210 9826
rect 114494 9774 114546 9826
rect 115614 9774 115666 9826
rect 29262 9662 29314 9714
rect 31278 9662 31330 9714
rect 32734 9662 32786 9714
rect 33294 9662 33346 9714
rect 35310 9662 35362 9714
rect 38670 9662 38722 9714
rect 41694 9662 41746 9714
rect 44046 9662 44098 9714
rect 44158 9662 44210 9714
rect 45838 9662 45890 9714
rect 45950 9662 46002 9714
rect 46622 9662 46674 9714
rect 48750 9662 48802 9714
rect 51662 9662 51714 9714
rect 56030 9662 56082 9714
rect 56366 9662 56418 9714
rect 56590 9662 56642 9714
rect 57710 9662 57762 9714
rect 59390 9662 59442 9714
rect 59838 9662 59890 9714
rect 60734 9662 60786 9714
rect 61070 9662 61122 9714
rect 61966 9662 62018 9714
rect 62638 9662 62690 9714
rect 63534 9662 63586 9714
rect 64206 9662 64258 9714
rect 65214 9662 65266 9714
rect 69358 9662 69410 9714
rect 69470 9662 69522 9714
rect 70142 9662 70194 9714
rect 70478 9662 70530 9714
rect 70926 9662 70978 9714
rect 71150 9662 71202 9714
rect 71262 9662 71314 9714
rect 72046 9662 72098 9714
rect 72606 9662 72658 9714
rect 73166 9662 73218 9714
rect 73278 9662 73330 9714
rect 74174 9662 74226 9714
rect 82910 9662 82962 9714
rect 85038 9662 85090 9714
rect 85934 9662 85986 9714
rect 86606 9662 86658 9714
rect 87950 9662 88002 9714
rect 88958 9662 89010 9714
rect 90414 9662 90466 9714
rect 92990 9662 93042 9714
rect 95790 9662 95842 9714
rect 99038 9662 99090 9714
rect 103294 9662 103346 9714
rect 103966 9662 104018 9714
rect 104974 9662 105026 9714
rect 106430 9662 106482 9714
rect 111358 9662 111410 9714
rect 112478 9662 112530 9714
rect 112702 9662 112754 9714
rect 113374 9662 113426 9714
rect 113934 9662 113986 9714
rect 114382 9662 114434 9714
rect 20750 9550 20802 9602
rect 21982 9550 22034 9602
rect 28478 9550 28530 9602
rect 29374 9550 29426 9602
rect 33406 9550 33458 9602
rect 36206 9550 36258 9602
rect 36990 9550 37042 9602
rect 44382 9550 44434 9602
rect 46398 9550 46450 9602
rect 47182 9550 47234 9602
rect 48190 9550 48242 9602
rect 50878 9550 50930 9602
rect 52222 9550 52274 9602
rect 56142 9550 56194 9602
rect 58270 9550 58322 9602
rect 61630 9550 61682 9602
rect 62862 9550 62914 9602
rect 64094 9550 64146 9602
rect 64878 9550 64930 9602
rect 65326 9550 65378 9602
rect 65550 9550 65602 9602
rect 66446 9550 66498 9602
rect 67006 9550 67058 9602
rect 68462 9550 68514 9602
rect 69022 9550 69074 9602
rect 69134 9550 69186 9602
rect 71710 9550 71762 9602
rect 72158 9550 72210 9602
rect 72382 9550 72434 9602
rect 72718 9550 72770 9602
rect 74510 9550 74562 9602
rect 75070 9550 75122 9602
rect 76750 9550 76802 9602
rect 77086 9550 77138 9602
rect 77422 9550 77474 9602
rect 77870 9550 77922 9602
rect 78206 9550 78258 9602
rect 82574 9550 82626 9602
rect 83358 9550 83410 9602
rect 84478 9550 84530 9602
rect 84702 9550 84754 9602
rect 84814 9550 84866 9602
rect 86494 9550 86546 9602
rect 92318 9550 92370 9602
rect 92878 9550 92930 9602
rect 93774 9550 93826 9602
rect 105310 9550 105362 9602
rect 106766 9550 106818 9602
rect 108894 9550 108946 9602
rect 112926 9550 112978 9602
rect 113710 9550 113762 9602
rect 115278 9550 115330 9602
rect 115502 9550 115554 9602
rect 116510 9550 116562 9602
rect 116958 9550 117010 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 81278 9382 81330 9434
rect 81382 9382 81434 9434
rect 81486 9382 81538 9434
rect 111998 9382 112050 9434
rect 112102 9382 112154 9434
rect 112206 9382 112258 9434
rect 142718 9382 142770 9434
rect 142822 9382 142874 9434
rect 142926 9382 142978 9434
rect 20974 9214 21026 9266
rect 22878 9214 22930 9266
rect 26798 9214 26850 9266
rect 27470 9214 27522 9266
rect 39678 9214 39730 9266
rect 40798 9214 40850 9266
rect 48302 9214 48354 9266
rect 48974 9214 49026 9266
rect 49310 9214 49362 9266
rect 49758 9214 49810 9266
rect 50318 9214 50370 9266
rect 51998 9214 52050 9266
rect 52558 9214 52610 9266
rect 60398 9214 60450 9266
rect 60846 9214 60898 9266
rect 61182 9214 61234 9266
rect 62414 9214 62466 9266
rect 63086 9214 63138 9266
rect 65886 9214 65938 9266
rect 66110 9214 66162 9266
rect 66670 9214 66722 9266
rect 71710 9214 71762 9266
rect 72494 9214 72546 9266
rect 73390 9214 73442 9266
rect 75854 9214 75906 9266
rect 80446 9214 80498 9266
rect 81230 9214 81282 9266
rect 21422 9102 21474 9154
rect 21758 9102 21810 9154
rect 22430 9102 22482 9154
rect 23998 9102 24050 9154
rect 28366 9102 28418 9154
rect 32174 9102 32226 9154
rect 35646 9102 35698 9154
rect 38670 9102 38722 9154
rect 40910 9102 40962 9154
rect 41918 9102 41970 9154
rect 44494 9102 44546 9154
rect 47518 9102 47570 9154
rect 47630 9102 47682 9154
rect 51326 9102 51378 9154
rect 52894 9102 52946 9154
rect 54350 9102 54402 9154
rect 55358 9102 55410 9154
rect 21870 8990 21922 9042
rect 27134 8990 27186 9042
rect 27806 8990 27858 9042
rect 28926 8990 28978 9042
rect 29486 8990 29538 9042
rect 30046 8990 30098 9042
rect 30382 8990 30434 9042
rect 31502 8990 31554 9042
rect 32510 8990 32562 9042
rect 34414 8990 34466 9042
rect 39790 8990 39842 9042
rect 40014 8990 40066 9042
rect 41134 8990 41186 9042
rect 41358 8990 41410 9042
rect 43822 8990 43874 9042
rect 47294 8990 47346 9042
rect 51214 8990 51266 9042
rect 20414 8878 20466 8930
rect 21534 8878 21586 8930
rect 23438 8878 23490 8930
rect 23662 8878 23714 8930
rect 24670 8878 24722 8930
rect 25566 8878 25618 8930
rect 26126 8878 26178 8930
rect 26574 8878 26626 8930
rect 30830 8878 30882 8930
rect 31838 8878 31890 8930
rect 39230 8878 39282 8930
rect 43038 8878 43090 8930
rect 46622 8878 46674 8930
rect 47182 8878 47234 8930
rect 50654 8878 50706 8930
rect 22318 8766 22370 8818
rect 23326 8766 23378 8818
rect 25566 8766 25618 8818
rect 26462 8766 26514 8818
rect 28142 8766 28194 8818
rect 28478 8766 28530 8818
rect 29038 8766 29090 8818
rect 39006 8766 39058 8818
rect 39678 8766 39730 8818
rect 50990 8766 51042 8818
rect 55806 9102 55858 9154
rect 55918 9102 55970 9154
rect 56926 9102 56978 9154
rect 58270 9102 58322 9154
rect 59166 9102 59218 9154
rect 61742 9102 61794 9154
rect 62078 9102 62130 9154
rect 66446 9102 66498 9154
rect 85822 9158 85874 9210
rect 86158 9214 86210 9266
rect 94446 9214 94498 9266
rect 105534 9214 105586 9266
rect 114830 9214 114882 9266
rect 115390 9214 115442 9266
rect 115950 9214 116002 9266
rect 117182 9214 117234 9266
rect 67342 9102 67394 9154
rect 67902 9102 67954 9154
rect 70590 9102 70642 9154
rect 73726 9102 73778 9154
rect 75406 9102 75458 9154
rect 76190 9102 76242 9154
rect 80110 9102 80162 9154
rect 83358 9102 83410 9154
rect 85934 9102 85986 9154
rect 86494 9102 86546 9154
rect 87278 9102 87330 9154
rect 87390 9102 87442 9154
rect 88734 9102 88786 9154
rect 93326 9102 93378 9154
rect 96350 9102 96402 9154
rect 98142 9102 98194 9154
rect 100382 9102 100434 9154
rect 102286 9102 102338 9154
rect 102846 9102 102898 9154
rect 105422 9102 105474 9154
rect 105758 9102 105810 9154
rect 108334 9102 108386 9154
rect 113150 9102 113202 9154
rect 114158 9102 114210 9154
rect 115614 9102 115666 9154
rect 115726 9102 115778 9154
rect 116174 9102 116226 9154
rect 52782 8990 52834 9042
rect 53118 8990 53170 9042
rect 55246 8990 55298 9042
rect 55582 8990 55634 9042
rect 56142 8990 56194 9042
rect 56590 8990 56642 9042
rect 59054 8990 59106 9042
rect 60398 8990 60450 9042
rect 62750 8990 62802 9042
rect 63422 8990 63474 9042
rect 64318 8990 64370 9042
rect 64654 8990 64706 9042
rect 64990 8990 65042 9042
rect 65774 8990 65826 9042
rect 66334 8990 66386 9042
rect 67230 8990 67282 9042
rect 71374 8990 71426 9042
rect 72718 8990 72770 9042
rect 73054 8990 73106 9042
rect 73390 8990 73442 9042
rect 77534 8990 77586 9042
rect 78430 8990 78482 9042
rect 78766 8990 78818 9042
rect 80334 8990 80386 9042
rect 80782 8990 80834 9042
rect 81902 8990 81954 9042
rect 82686 8990 82738 9042
rect 86270 8990 86322 9042
rect 86606 8990 86658 9042
rect 87950 8990 88002 9042
rect 94110 8990 94162 9042
rect 96574 8990 96626 9042
rect 97918 8990 97970 9042
rect 99710 8990 99762 9042
rect 101054 8990 101106 9042
rect 101278 8990 101330 9042
rect 102510 8990 102562 9042
rect 103630 8990 103682 9042
rect 105198 8990 105250 9042
rect 109006 8990 109058 9042
rect 109678 8990 109730 9042
rect 111582 8990 111634 9042
rect 112926 8990 112978 9042
rect 113262 8990 113314 9042
rect 113486 8990 113538 9042
rect 113934 8990 113986 9042
rect 114606 8990 114658 9042
rect 115166 8990 115218 9042
rect 116286 8990 116338 9042
rect 51550 8878 51602 8930
rect 53566 8878 53618 8930
rect 57486 8878 57538 8930
rect 59278 8878 59330 8930
rect 63982 8878 64034 8930
rect 64542 8878 64594 8930
rect 65438 8878 65490 8930
rect 69246 8878 69298 8930
rect 69582 8878 69634 8930
rect 74062 8878 74114 8930
rect 76638 8878 76690 8930
rect 78318 8878 78370 8930
rect 81454 8878 81506 8930
rect 85486 8878 85538 8930
rect 90862 8878 90914 8930
rect 91198 8878 91250 8930
rect 94894 8878 94946 8930
rect 95790 8878 95842 8930
rect 101614 8878 101666 8930
rect 102398 8878 102450 8930
rect 104526 8878 104578 8930
rect 106206 8878 106258 8930
rect 110574 8878 110626 8930
rect 112142 8878 112194 8930
rect 114382 8878 114434 8930
rect 116734 8878 116786 8930
rect 117630 8878 117682 8930
rect 118078 8878 118130 8930
rect 118638 8878 118690 8930
rect 52222 8766 52274 8818
rect 52558 8766 52610 8818
rect 67342 8766 67394 8818
rect 78654 8766 78706 8818
rect 87278 8766 87330 8818
rect 95902 8766 95954 8818
rect 100830 8766 100882 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 96638 8598 96690 8650
rect 96742 8598 96794 8650
rect 96846 8598 96898 8650
rect 127358 8598 127410 8650
rect 127462 8598 127514 8650
rect 127566 8598 127618 8650
rect 158078 8598 158130 8650
rect 158182 8598 158234 8650
rect 158286 8598 158338 8650
rect 29934 8430 29986 8482
rect 94110 8430 94162 8482
rect 117630 8430 117682 8482
rect 118190 8430 118242 8482
rect 20190 8318 20242 8370
rect 23438 8318 23490 8370
rect 27134 8318 27186 8370
rect 28142 8318 28194 8370
rect 29486 8318 29538 8370
rect 32958 8318 33010 8370
rect 34862 8318 34914 8370
rect 37102 8318 37154 8370
rect 37662 8318 37714 8370
rect 37774 8318 37826 8370
rect 38558 8318 38610 8370
rect 40686 8318 40738 8370
rect 41918 8318 41970 8370
rect 47518 8318 47570 8370
rect 48862 8318 48914 8370
rect 50878 8318 50930 8370
rect 55022 8318 55074 8370
rect 57150 8318 57202 8370
rect 57710 8318 57762 8370
rect 60622 8318 60674 8370
rect 62862 8318 62914 8370
rect 63982 8318 64034 8370
rect 66110 8318 66162 8370
rect 17390 8206 17442 8258
rect 20750 8206 20802 8258
rect 21870 8206 21922 8258
rect 22094 8206 22146 8258
rect 22542 8206 22594 8258
rect 23886 8206 23938 8258
rect 25566 8206 25618 8258
rect 29262 8206 29314 8258
rect 29934 8206 29986 8258
rect 30718 8206 30770 8258
rect 32622 8206 32674 8258
rect 33070 8206 33122 8258
rect 33854 8206 33906 8258
rect 37214 8206 37266 8258
rect 37438 8206 37490 8258
rect 41358 8206 41410 8258
rect 45054 8206 45106 8258
rect 45502 8206 45554 8258
rect 45726 8206 45778 8258
rect 49422 8206 49474 8258
rect 66558 8318 66610 8370
rect 71710 8318 71762 8370
rect 72942 8318 72994 8370
rect 75070 8318 75122 8370
rect 76974 8318 77026 8370
rect 78094 8318 78146 8370
rect 80222 8318 80274 8370
rect 85150 8318 85202 8370
rect 86270 8318 86322 8370
rect 90750 8318 90802 8370
rect 90974 8318 91026 8370
rect 91422 8318 91474 8370
rect 93326 8318 93378 8370
rect 96238 8318 96290 8370
rect 100606 8318 100658 8370
rect 101390 8318 101442 8370
rect 104638 8318 104690 8370
rect 106206 8318 106258 8370
rect 111358 8318 111410 8370
rect 113486 8318 113538 8370
rect 115390 8318 115442 8370
rect 53566 8206 53618 8258
rect 54350 8206 54402 8258
rect 60734 8206 60786 8258
rect 63198 8206 63250 8258
rect 66334 8206 66386 8258
rect 66670 8206 66722 8258
rect 67006 8206 67058 8258
rect 67230 8206 67282 8258
rect 67454 8206 67506 8258
rect 67790 8206 67842 8258
rect 72270 8206 72322 8258
rect 75406 8206 75458 8258
rect 75742 8206 75794 8258
rect 77086 8206 77138 8258
rect 77534 8206 77586 8258
rect 81006 8206 81058 8258
rect 81454 8206 81506 8258
rect 81902 8206 81954 8258
rect 82238 8206 82290 8258
rect 82910 8206 82962 8258
rect 84030 8206 84082 8258
rect 84254 8206 84306 8258
rect 84702 8206 84754 8258
rect 85038 8206 85090 8258
rect 85486 8206 85538 8258
rect 86158 8206 86210 8258
rect 88286 8206 88338 8258
rect 88846 8206 88898 8258
rect 88958 8206 89010 8258
rect 89294 8206 89346 8258
rect 89966 8206 90018 8258
rect 90526 8206 90578 8258
rect 93886 8206 93938 8258
rect 94334 8206 94386 8258
rect 95230 8206 95282 8258
rect 95566 8206 95618 8258
rect 99150 8206 99202 8258
rect 100046 8206 100098 8258
rect 100270 8206 100322 8258
rect 101726 8206 101778 8258
rect 105198 8206 105250 8258
rect 106094 8206 106146 8258
rect 106542 8206 106594 8258
rect 110686 8206 110738 8258
rect 114270 8206 114322 8258
rect 117182 8206 117234 8258
rect 117518 8206 117570 8258
rect 118302 8206 118354 8258
rect 118750 8206 118802 8258
rect 18062 8094 18114 8146
rect 20414 8094 20466 8146
rect 21422 8094 21474 8146
rect 21534 8094 21586 8146
rect 22766 8094 22818 8146
rect 22878 8094 22930 8146
rect 25230 8094 25282 8146
rect 25342 8094 25394 8146
rect 25790 8094 25842 8146
rect 25902 8094 25954 8146
rect 27022 8094 27074 8146
rect 27246 8094 27298 8146
rect 28702 8094 28754 8146
rect 30046 8094 30098 8146
rect 30382 8094 30434 8146
rect 36206 8094 36258 8146
rect 38110 8094 38162 8146
rect 43822 8094 43874 8146
rect 46286 8094 46338 8146
rect 47854 8094 47906 8146
rect 47966 8094 48018 8146
rect 49758 8094 49810 8146
rect 51886 8094 51938 8146
rect 52670 8094 52722 8146
rect 53006 8094 53058 8146
rect 53230 8094 53282 8146
rect 59502 8094 59554 8146
rect 60510 8094 60562 8146
rect 61070 8094 61122 8146
rect 61518 8094 61570 8146
rect 70366 8094 70418 8146
rect 83246 8094 83298 8146
rect 85710 8094 85762 8146
rect 86270 8094 86322 8146
rect 86494 8094 86546 8146
rect 86718 8094 86770 8146
rect 87502 8094 87554 8146
rect 88398 8094 88450 8146
rect 89182 8094 89234 8146
rect 91982 8094 92034 8146
rect 93662 8094 93714 8146
rect 95678 8094 95730 8146
rect 95790 8094 95842 8146
rect 98366 8094 98418 8146
rect 102510 8094 102562 8146
rect 110238 8094 110290 8146
rect 110910 8094 110962 8146
rect 111022 8094 111074 8146
rect 114606 8094 114658 8146
rect 114942 8094 114994 8146
rect 116622 8094 116674 8146
rect 20638 7982 20690 8034
rect 21198 7982 21250 8034
rect 22318 7982 22370 8034
rect 23102 7982 23154 8034
rect 24334 7982 24386 8034
rect 24782 7982 24834 8034
rect 25006 7982 25058 8034
rect 26238 7982 26290 8034
rect 26574 7982 26626 8034
rect 27582 7982 27634 8034
rect 38222 7982 38274 8034
rect 45278 7982 45330 8034
rect 48190 7982 48242 8034
rect 51550 7982 51602 8034
rect 51998 7982 52050 8034
rect 52222 7982 52274 8034
rect 52782 7982 52834 8034
rect 53902 7982 53954 8034
rect 67118 7982 67170 8034
rect 67678 7982 67730 8034
rect 68238 7982 68290 8034
rect 71150 7982 71202 8034
rect 75518 7982 75570 8034
rect 77422 7982 77474 8034
rect 82126 7982 82178 8034
rect 84366 7982 84418 8034
rect 84478 7982 84530 8034
rect 85262 7982 85314 8034
rect 87166 7982 87218 8034
rect 87390 7982 87442 8034
rect 88622 7982 88674 8034
rect 90190 7982 90242 8034
rect 94782 7982 94834 8034
rect 99598 7982 99650 8034
rect 104862 7982 104914 8034
rect 105086 7982 105138 8034
rect 106430 7982 106482 8034
rect 107662 7982 107714 8034
rect 107886 7982 107938 8034
rect 114718 7982 114770 8034
rect 117294 7982 117346 8034
rect 117854 7982 117906 8034
rect 119198 7982 119250 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 81278 7814 81330 7866
rect 81382 7814 81434 7866
rect 81486 7814 81538 7866
rect 111998 7814 112050 7866
rect 112102 7814 112154 7866
rect 112206 7814 112258 7866
rect 142718 7814 142770 7866
rect 142822 7814 142874 7866
rect 142926 7814 142978 7866
rect 23102 7646 23154 7698
rect 24558 7646 24610 7698
rect 26014 7646 26066 7698
rect 28030 7646 28082 7698
rect 29486 7646 29538 7698
rect 32174 7646 32226 7698
rect 35646 7646 35698 7698
rect 40238 7646 40290 7698
rect 41022 7646 41074 7698
rect 49534 7646 49586 7698
rect 50654 7646 50706 7698
rect 51438 7646 51490 7698
rect 56702 7646 56754 7698
rect 57262 7646 57314 7698
rect 64430 7646 64482 7698
rect 65326 7646 65378 7698
rect 65662 7646 65714 7698
rect 66558 7646 66610 7698
rect 85934 7646 85986 7698
rect 87390 7646 87442 7698
rect 94670 7646 94722 7698
rect 95902 7646 95954 7698
rect 110574 7646 110626 7698
rect 110910 7646 110962 7698
rect 111470 7646 111522 7698
rect 118750 7646 118802 7698
rect 119870 7646 119922 7698
rect 23998 7534 24050 7586
rect 24334 7534 24386 7586
rect 24670 7534 24722 7586
rect 27246 7534 27298 7586
rect 28702 7534 28754 7586
rect 31054 7534 31106 7586
rect 34302 7534 34354 7586
rect 34750 7534 34802 7586
rect 37214 7534 37266 7586
rect 39230 7534 39282 7586
rect 39566 7534 39618 7586
rect 42814 7534 42866 7586
rect 49198 7534 49250 7586
rect 49310 7534 49362 7586
rect 54462 7534 54514 7586
rect 56590 7534 56642 7586
rect 57374 7534 57426 7586
rect 58718 7534 58770 7586
rect 63534 7534 63586 7586
rect 67790 7534 67842 7586
rect 71486 7534 71538 7586
rect 72270 7534 72322 7586
rect 72606 7534 72658 7586
rect 73166 7534 73218 7586
rect 74622 7534 74674 7586
rect 78430 7534 78482 7586
rect 82686 7534 82738 7586
rect 88734 7534 88786 7586
rect 92094 7534 92146 7586
rect 92766 7534 92818 7586
rect 94894 7534 94946 7586
rect 95790 7534 95842 7586
rect 96350 7534 96402 7586
rect 98030 7534 98082 7586
rect 100382 7534 100434 7586
rect 102062 7534 102114 7586
rect 106318 7534 106370 7586
rect 108894 7534 108946 7586
rect 114606 7534 114658 7586
rect 116398 7534 116450 7586
rect 120318 7534 120370 7586
rect 19854 7422 19906 7474
rect 22878 7422 22930 7474
rect 23214 7422 23266 7474
rect 23886 7422 23938 7474
rect 28366 7422 28418 7474
rect 28926 7422 28978 7474
rect 29150 7422 29202 7474
rect 29262 7422 29314 7474
rect 32622 7422 32674 7474
rect 33182 7422 33234 7474
rect 33742 7422 33794 7474
rect 34638 7422 34690 7474
rect 38446 7422 38498 7474
rect 39902 7422 39954 7474
rect 41358 7422 41410 7474
rect 42030 7422 42082 7474
rect 45390 7422 45442 7474
rect 50206 7422 50258 7474
rect 52110 7422 52162 7474
rect 52558 7422 52610 7474
rect 53566 7422 53618 7474
rect 54014 7422 54066 7474
rect 54686 7422 54738 7474
rect 55134 7422 55186 7474
rect 55694 7422 55746 7474
rect 56926 7422 56978 7474
rect 57598 7422 57650 7474
rect 58046 7422 58098 7474
rect 66446 7422 66498 7474
rect 67118 7422 67170 7474
rect 72942 7422 72994 7474
rect 73614 7422 73666 7474
rect 73950 7422 74002 7474
rect 78990 7422 79042 7474
rect 81566 7422 81618 7474
rect 86718 7422 86770 7474
rect 87054 7422 87106 7474
rect 87950 7422 88002 7474
rect 91422 7422 91474 7474
rect 91646 7422 91698 7474
rect 93998 7422 94050 7474
rect 94558 7422 94610 7474
rect 95006 7422 95058 7474
rect 96238 7422 96290 7474
rect 97918 7422 97970 7474
rect 99710 7422 99762 7474
rect 102510 7422 102562 7474
rect 103070 7422 103122 7474
rect 103966 7422 104018 7474
rect 104302 7422 104354 7474
rect 105534 7422 105586 7474
rect 115278 7422 115330 7474
rect 117742 7422 117794 7474
rect 20526 7310 20578 7362
rect 22654 7310 22706 7362
rect 25454 7310 25506 7362
rect 26238 7310 26290 7362
rect 29822 7310 29874 7362
rect 33630 7310 33682 7362
rect 44942 7310 44994 7362
rect 46062 7310 46114 7362
rect 48190 7310 48242 7362
rect 48750 7310 48802 7362
rect 49870 7310 49922 7362
rect 54238 7310 54290 7362
rect 60846 7310 60898 7362
rect 61518 7310 61570 7362
rect 64990 7310 65042 7362
rect 66222 7310 66274 7362
rect 69918 7310 69970 7362
rect 70478 7310 70530 7362
rect 73390 7310 73442 7362
rect 76750 7310 76802 7362
rect 77086 7310 77138 7362
rect 79438 7310 79490 7362
rect 86158 7310 86210 7362
rect 90862 7310 90914 7362
rect 91198 7310 91250 7362
rect 92990 7310 93042 7362
rect 100718 7310 100770 7362
rect 104750 7310 104802 7362
rect 108446 7310 108498 7362
rect 110238 7310 110290 7362
rect 112030 7310 112082 7362
rect 112478 7310 112530 7362
rect 117406 7310 117458 7362
rect 118190 7310 118242 7362
rect 119422 7310 119474 7362
rect 23998 7198 24050 7250
rect 41022 7198 41074 7250
rect 41134 7198 41186 7250
rect 48862 7198 48914 7250
rect 66558 7198 66610 7250
rect 94334 7198 94386 7250
rect 103966 7198 104018 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 96638 7030 96690 7082
rect 96742 7030 96794 7082
rect 96846 7030 96898 7082
rect 127358 7030 127410 7082
rect 127462 7030 127514 7082
rect 127566 7030 127618 7082
rect 158078 7030 158130 7082
rect 158182 7030 158234 7082
rect 158286 7030 158338 7082
rect 21982 6862 22034 6914
rect 29486 6862 29538 6914
rect 29598 6862 29650 6914
rect 30382 6862 30434 6914
rect 30606 6862 30658 6914
rect 61070 6862 61122 6914
rect 61294 6862 61346 6914
rect 75742 6862 75794 6914
rect 117294 6862 117346 6914
rect 18622 6750 18674 6802
rect 21646 6750 21698 6802
rect 22318 6750 22370 6802
rect 25118 6750 25170 6802
rect 27246 6750 27298 6802
rect 28590 6750 28642 6802
rect 29262 6750 29314 6802
rect 30830 6750 30882 6802
rect 34974 6750 35026 6802
rect 38446 6750 38498 6802
rect 39006 6750 39058 6802
rect 45614 6750 45666 6802
rect 48638 6750 48690 6802
rect 52110 6750 52162 6802
rect 57710 6750 57762 6802
rect 59950 6750 60002 6802
rect 61630 6750 61682 6802
rect 61854 6750 61906 6802
rect 68910 6750 68962 6802
rect 69918 6750 69970 6802
rect 78206 6750 78258 6802
rect 80110 6750 80162 6802
rect 82350 6750 82402 6802
rect 84702 6750 84754 6802
rect 89406 6750 89458 6802
rect 91982 6750 92034 6802
rect 96014 6750 96066 6802
rect 100270 6750 100322 6802
rect 104862 6750 104914 6802
rect 107550 6750 107602 6802
rect 116846 6750 116898 6802
rect 118190 6750 118242 6802
rect 19854 6638 19906 6690
rect 20302 6638 20354 6690
rect 24334 6638 24386 6690
rect 28142 6638 28194 6690
rect 31390 6638 31442 6690
rect 31726 6638 31778 6690
rect 33182 6638 33234 6690
rect 33518 6638 33570 6690
rect 33854 6638 33906 6690
rect 34078 6638 34130 6690
rect 39566 6638 39618 6690
rect 41582 6638 41634 6690
rect 45054 6638 45106 6690
rect 45390 6638 45442 6690
rect 45838 6638 45890 6690
rect 45950 6638 46002 6690
rect 49198 6638 49250 6690
rect 53678 6638 53730 6690
rect 60734 6638 60786 6690
rect 61742 6638 61794 6690
rect 62302 6638 62354 6690
rect 64318 6638 64370 6690
rect 66558 6638 66610 6690
rect 67230 6638 67282 6690
rect 67790 6638 67842 6690
rect 69358 6638 69410 6690
rect 76414 6638 76466 6690
rect 79550 6638 79602 6690
rect 82238 6638 82290 6690
rect 82462 6638 82514 6690
rect 84142 6638 84194 6690
rect 91310 6638 91362 6690
rect 95454 6638 95506 6690
rect 98142 6638 98194 6690
rect 98926 6638 98978 6690
rect 99710 6638 99762 6690
rect 102398 6638 102450 6690
rect 103070 6638 103122 6690
rect 103742 6638 103794 6690
rect 106654 6638 106706 6690
rect 109678 6638 109730 6690
rect 110350 6638 110402 6690
rect 110910 6638 110962 6690
rect 117182 6638 117234 6690
rect 21758 6526 21810 6578
rect 23550 6526 23602 6578
rect 27694 6526 27746 6578
rect 29150 6526 29202 6578
rect 29934 6526 29986 6578
rect 34638 6526 34690 6578
rect 36094 6526 36146 6578
rect 37438 6526 37490 6578
rect 38894 6526 38946 6578
rect 39118 6526 39170 6578
rect 40686 6526 40738 6578
rect 43374 6526 43426 6578
rect 44046 6526 44098 6578
rect 44158 6526 44210 6578
rect 44382 6526 44434 6578
rect 46510 6526 46562 6578
rect 49982 6526 50034 6578
rect 58606 6526 58658 6578
rect 63422 6526 63474 6578
rect 64878 6526 64930 6578
rect 66334 6526 66386 6578
rect 66894 6526 66946 6578
rect 71710 6526 71762 6578
rect 72494 6526 72546 6578
rect 72830 6526 72882 6578
rect 73390 6526 73442 6578
rect 76974 6526 77026 6578
rect 81118 6526 81170 6578
rect 84366 6526 84418 6578
rect 85934 6526 85986 6578
rect 86606 6526 86658 6578
rect 90638 6526 90690 6578
rect 91198 6526 91250 6578
rect 94222 6526 94274 6578
rect 95230 6526 95282 6578
rect 99822 6526 99874 6578
rect 103406 6526 103458 6578
rect 106094 6526 106146 6578
rect 111358 6526 111410 6578
rect 112366 6526 112418 6578
rect 114718 6526 114770 6578
rect 115502 6526 115554 6578
rect 120318 6526 120370 6578
rect 17838 6414 17890 6466
rect 19070 6414 19122 6466
rect 19630 6414 19682 6466
rect 27582 6414 27634 6466
rect 39790 6414 39842 6466
rect 44830 6414 44882 6466
rect 64990 6414 65042 6466
rect 66782 6414 66834 6466
rect 68462 6414 68514 6466
rect 77982 6414 78034 6466
rect 79774 6414 79826 6466
rect 81790 6414 81842 6466
rect 89070 6414 89122 6466
rect 94894 6414 94946 6466
rect 100046 6414 100098 6466
rect 103630 6414 103682 6466
rect 106542 6414 106594 6466
rect 111806 6414 111858 6466
rect 117294 6414 117346 6466
rect 120878 6414 120930 6466
rect 121662 6414 121714 6466
rect 122558 6414 122610 6466
rect 123790 6414 123842 6466
rect 125806 6414 125858 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 81278 6246 81330 6298
rect 81382 6246 81434 6298
rect 81486 6246 81538 6298
rect 111998 6246 112050 6298
rect 112102 6246 112154 6298
rect 112206 6246 112258 6298
rect 142718 6246 142770 6298
rect 142822 6246 142874 6298
rect 142926 6246 142978 6298
rect 20078 6078 20130 6130
rect 21086 6078 21138 6130
rect 22878 6078 22930 6130
rect 30270 6078 30322 6130
rect 35198 6078 35250 6130
rect 39902 6078 39954 6130
rect 42366 6078 42418 6130
rect 43262 6078 43314 6130
rect 71822 6078 71874 6130
rect 79438 6078 79490 6130
rect 88062 6078 88114 6130
rect 94222 6078 94274 6130
rect 95230 6078 95282 6130
rect 102622 6078 102674 6130
rect 108782 6078 108834 6130
rect 109006 6078 109058 6130
rect 114382 6078 114434 6130
rect 18174 5966 18226 6018
rect 21310 5966 21362 6018
rect 24558 5966 24610 6018
rect 25118 5966 25170 6018
rect 27246 5966 27298 6018
rect 29374 5966 29426 6018
rect 32062 5966 32114 6018
rect 34078 5966 34130 6018
rect 37550 5966 37602 6018
rect 39342 5966 39394 6018
rect 47854 5966 47906 6018
rect 51886 5966 51938 6018
rect 53006 5966 53058 6018
rect 53118 5966 53170 6018
rect 53342 5966 53394 6018
rect 55582 5966 55634 6018
rect 56814 5966 56866 6018
rect 60622 5966 60674 6018
rect 61518 5966 61570 6018
rect 64990 5966 65042 6018
rect 68014 5966 68066 6018
rect 73390 5966 73442 6018
rect 76974 5966 77026 6018
rect 80334 5966 80386 6018
rect 87166 5966 87218 6018
rect 87278 5966 87330 6018
rect 88174 5966 88226 6018
rect 91870 5966 91922 6018
rect 95118 5966 95170 6018
rect 96238 5966 96290 6018
rect 98702 5966 98754 6018
rect 99038 5966 99090 6018
rect 101726 5966 101778 6018
rect 102510 5966 102562 6018
rect 102846 5966 102898 6018
rect 105422 5966 105474 6018
rect 105758 5966 105810 6018
rect 107886 5966 107938 6018
rect 109118 5966 109170 6018
rect 110686 5966 110738 6018
rect 111358 5966 111410 6018
rect 113486 5966 113538 6018
rect 115166 5966 115218 6018
rect 121214 5966 121266 6018
rect 123230 5966 123282 6018
rect 124350 5966 124402 6018
rect 125582 5966 125634 6018
rect 21870 5854 21922 5906
rect 22654 5854 22706 5906
rect 30270 5854 30322 5906
rect 30606 5854 30658 5906
rect 34974 5854 35026 5906
rect 36430 5854 36482 5906
rect 37886 5854 37938 5906
rect 38446 5854 38498 5906
rect 39006 5854 39058 5906
rect 39566 5854 39618 5906
rect 39790 5854 39842 5906
rect 39902 5854 39954 5906
rect 40238 5854 40290 5906
rect 40910 5854 40962 5906
rect 41022 5854 41074 5906
rect 41470 5854 41522 5906
rect 41806 5854 41858 5906
rect 43710 5854 43762 5906
rect 48862 5854 48914 5906
rect 52670 5854 52722 5906
rect 57038 5854 57090 5906
rect 57262 5854 57314 5906
rect 58270 5854 58322 5906
rect 64430 5854 64482 5906
rect 66782 5854 66834 5906
rect 67342 5854 67394 5906
rect 67566 5854 67618 5906
rect 67678 5854 67730 5906
rect 68462 5854 68514 5906
rect 69134 5854 69186 5906
rect 72270 5854 72322 5906
rect 76414 5854 76466 5906
rect 82126 5854 82178 5906
rect 85262 5854 85314 5906
rect 85822 5854 85874 5906
rect 86046 5854 86098 5906
rect 86494 5854 86546 5906
rect 86718 5854 86770 5906
rect 86942 5854 86994 5906
rect 87838 5854 87890 5906
rect 89070 5854 89122 5906
rect 89854 5854 89906 5906
rect 90526 5854 90578 5906
rect 102958 5854 103010 5906
rect 117854 5854 117906 5906
rect 118078 5854 118130 5906
rect 119646 5854 119698 5906
rect 119982 5854 120034 5906
rect 120654 5854 120706 5906
rect 120990 5854 121042 5906
rect 124014 5854 124066 5906
rect 17838 5742 17890 5794
rect 19294 5742 19346 5794
rect 20638 5742 20690 5794
rect 23214 5742 23266 5794
rect 28478 5742 28530 5794
rect 31278 5742 31330 5794
rect 33294 5742 33346 5794
rect 37998 5742 38050 5794
rect 42814 5742 42866 5794
rect 46510 5742 46562 5794
rect 49198 5742 49250 5794
rect 49758 5742 49810 5794
rect 53566 5742 53618 5794
rect 56926 5742 56978 5794
rect 57710 5742 57762 5794
rect 58606 5742 58658 5794
rect 63758 5742 63810 5794
rect 65550 5742 65602 5794
rect 71262 5742 71314 5794
rect 81678 5742 81730 5794
rect 82798 5742 82850 5794
rect 84926 5742 84978 5794
rect 86270 5742 86322 5794
rect 89742 5742 89794 5794
rect 93886 5742 93938 5794
rect 94670 5742 94722 5794
rect 100382 5742 100434 5794
rect 100718 5742 100770 5794
rect 103742 5742 103794 5794
rect 104302 5742 104354 5794
rect 109454 5742 109506 5794
rect 116958 5742 117010 5794
rect 117630 5742 117682 5794
rect 119422 5742 119474 5794
rect 121662 5742 121714 5794
rect 122222 5742 122274 5794
rect 126590 5742 126642 5794
rect 127710 5742 127762 5794
rect 138910 5742 138962 5794
rect 143838 5742 143890 5794
rect 144174 5742 144226 5794
rect 30382 5630 30434 5682
rect 41246 5630 41298 5682
rect 44606 5630 44658 5682
rect 74174 5630 74226 5682
rect 118638 5630 118690 5682
rect 139022 5630 139074 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 96638 5462 96690 5514
rect 96742 5462 96794 5514
rect 96846 5462 96898 5514
rect 127358 5462 127410 5514
rect 127462 5462 127514 5514
rect 127566 5462 127618 5514
rect 158078 5462 158130 5514
rect 158182 5462 158234 5514
rect 158286 5462 158338 5514
rect 15934 5294 15986 5346
rect 21646 5294 21698 5346
rect 32286 5294 32338 5346
rect 36878 5294 36930 5346
rect 40462 5294 40514 5346
rect 45278 5294 45330 5346
rect 45390 5294 45442 5346
rect 45614 5294 45666 5346
rect 52782 5294 52834 5346
rect 60622 5294 60674 5346
rect 68462 5294 68514 5346
rect 98702 5294 98754 5346
rect 99038 5294 99090 5346
rect 102510 5294 102562 5346
rect 125918 5294 125970 5346
rect 16382 5182 16434 5234
rect 17502 5182 17554 5234
rect 19070 5182 19122 5234
rect 19294 5182 19346 5234
rect 23662 5182 23714 5234
rect 25790 5182 25842 5234
rect 26350 5182 26402 5234
rect 27134 5182 27186 5234
rect 32958 5182 33010 5234
rect 34750 5182 34802 5234
rect 39902 5182 39954 5234
rect 43262 5182 43314 5234
rect 46286 5182 46338 5234
rect 48750 5182 48802 5234
rect 57038 5182 57090 5234
rect 61630 5182 61682 5234
rect 64430 5182 64482 5234
rect 69470 5182 69522 5234
rect 74174 5182 74226 5234
rect 76974 5182 77026 5234
rect 79214 5182 79266 5234
rect 80334 5182 80386 5234
rect 85374 5182 85426 5234
rect 89518 5182 89570 5234
rect 89966 5182 90018 5234
rect 92430 5182 92482 5234
rect 102846 5182 102898 5234
rect 108782 5182 108834 5234
rect 110126 5182 110178 5234
rect 113038 5182 113090 5234
rect 116174 5182 116226 5234
rect 120542 5182 120594 5234
rect 121102 5182 121154 5234
rect 123230 5182 123282 5234
rect 134990 5182 135042 5234
rect 140142 5182 140194 5234
rect 142942 5182 142994 5234
rect 150670 5182 150722 5234
rect 15374 5070 15426 5122
rect 15598 5070 15650 5122
rect 16830 5070 16882 5122
rect 21310 5070 21362 5122
rect 21870 5070 21922 5122
rect 22878 5070 22930 5122
rect 26798 5070 26850 5122
rect 29486 5070 29538 5122
rect 33182 5070 33234 5122
rect 35758 5070 35810 5122
rect 40350 5070 40402 5122
rect 42254 5070 42306 5122
rect 43710 5070 43762 5122
rect 45726 5070 45778 5122
rect 50430 5070 50482 5122
rect 51774 5070 51826 5122
rect 52670 5070 52722 5122
rect 53342 5070 53394 5122
rect 53454 5070 53506 5122
rect 53678 5070 53730 5122
rect 53790 5070 53842 5122
rect 54238 5070 54290 5122
rect 54910 5070 54962 5122
rect 60734 5070 60786 5122
rect 63646 5070 63698 5122
rect 65774 5070 65826 5122
rect 67790 5070 67842 5122
rect 68686 5070 68738 5122
rect 69022 5070 69074 5122
rect 71598 5070 71650 5122
rect 72046 5070 72098 5122
rect 77198 5070 77250 5122
rect 79662 5070 79714 5122
rect 82910 5070 82962 5122
rect 83246 5070 83298 5122
rect 83582 5070 83634 5122
rect 84142 5070 84194 5122
rect 85262 5070 85314 5122
rect 85598 5070 85650 5122
rect 86718 5070 86770 5122
rect 94222 5070 94274 5122
rect 95566 5070 95618 5122
rect 98926 5070 98978 5122
rect 103182 5070 103234 5122
rect 103518 5070 103570 5122
rect 103854 5070 103906 5122
rect 111918 5070 111970 5122
rect 113262 5070 113314 5122
rect 116398 5070 116450 5122
rect 129166 5070 129218 5122
rect 132302 5070 132354 5122
rect 137454 5070 137506 5122
rect 138238 5070 138290 5122
rect 142718 5070 142770 5122
rect 147646 5070 147698 5122
rect 148094 5070 148146 5122
rect 149214 5070 149266 5122
rect 17054 4958 17106 5010
rect 20302 4958 20354 5010
rect 22094 4958 22146 5010
rect 28142 4958 28194 5010
rect 29822 4958 29874 5010
rect 34750 4958 34802 5010
rect 35534 4958 35586 5010
rect 39006 4958 39058 5010
rect 48078 4958 48130 5010
rect 50318 4958 50370 5010
rect 51550 4958 51602 5010
rect 52782 4958 52834 5010
rect 59726 4958 59778 5010
rect 60622 4958 60674 5010
rect 64654 4958 64706 5010
rect 67678 4958 67730 5010
rect 71150 4958 71202 5010
rect 72606 4958 72658 5010
rect 75518 4958 75570 5010
rect 77758 4958 77810 5010
rect 82462 4958 82514 5010
rect 84366 4958 84418 5010
rect 87390 4958 87442 5010
rect 90862 4958 90914 5010
rect 91982 4958 92034 5010
rect 92094 4958 92146 5010
rect 93998 4958 94050 5010
rect 95230 4958 95282 5010
rect 96238 4958 96290 5010
rect 99038 4958 99090 5010
rect 100046 4958 100098 5010
rect 103742 4958 103794 5010
rect 104638 4958 104690 5010
rect 106766 4958 106818 5010
rect 107662 4958 107714 5010
rect 111358 4958 111410 5010
rect 113822 4958 113874 5010
rect 116958 4958 117010 5010
rect 118750 4958 118802 5010
rect 122110 4958 122162 5010
rect 125246 4958 125298 5010
rect 128046 4958 128098 5010
rect 128830 4958 128882 5010
rect 133870 4958 133922 5010
rect 141374 4958 141426 5010
rect 143950 4958 144002 5010
rect 144734 4958 144786 5010
rect 145070 4958 145122 5010
rect 149550 4958 149602 5010
rect 17950 4846 18002 4898
rect 18622 4846 18674 4898
rect 21758 4846 21810 4898
rect 22542 4846 22594 4898
rect 57374 4846 57426 4898
rect 70702 4846 70754 4898
rect 76414 4846 76466 4898
rect 83358 4846 83410 4898
rect 85598 4846 85650 4898
rect 91758 4846 91810 4898
rect 111806 4846 111858 4898
rect 113374 4846 113426 4898
rect 117854 4846 117906 4898
rect 133534 4846 133586 4898
rect 135998 4846 136050 4898
rect 138350 4846 138402 4898
rect 147870 4846 147922 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 81278 4678 81330 4730
rect 81382 4678 81434 4730
rect 81486 4678 81538 4730
rect 111998 4678 112050 4730
rect 112102 4678 112154 4730
rect 112206 4678 112258 4730
rect 142718 4678 142770 4730
rect 142822 4678 142874 4730
rect 142926 4678 142978 4730
rect 19070 4510 19122 4562
rect 23886 4510 23938 4562
rect 25342 4510 25394 4562
rect 26686 4510 26738 4562
rect 30718 4510 30770 4562
rect 38670 4510 38722 4562
rect 39118 4510 39170 4562
rect 39342 4510 39394 4562
rect 42590 4510 42642 4562
rect 48078 4510 48130 4562
rect 48302 4510 48354 4562
rect 50430 4510 50482 4562
rect 56030 4510 56082 4562
rect 64542 4510 64594 4562
rect 68574 4510 68626 4562
rect 72494 4510 72546 4562
rect 72718 4510 72770 4562
rect 76302 4510 76354 4562
rect 76526 4510 76578 4562
rect 13806 4398 13858 4450
rect 15486 4398 15538 4450
rect 16830 4398 16882 4450
rect 18958 4398 19010 4450
rect 21534 4398 21586 4450
rect 23102 4398 23154 4450
rect 23438 4398 23490 4450
rect 23662 4398 23714 4450
rect 24670 4398 24722 4450
rect 29150 4398 29202 4450
rect 32062 4398 32114 4450
rect 34190 4398 34242 4450
rect 37326 4398 37378 4450
rect 38334 4398 38386 4450
rect 39454 4398 39506 4450
rect 46286 4398 46338 4450
rect 47966 4398 48018 4450
rect 49310 4398 49362 4450
rect 49646 4398 49698 4450
rect 53454 4398 53506 4450
rect 53902 4398 53954 4450
rect 56590 4398 56642 4450
rect 56702 4398 56754 4450
rect 56926 4398 56978 4450
rect 57374 4398 57426 4450
rect 61070 4398 61122 4450
rect 63758 4398 63810 4450
rect 65102 4398 65154 4450
rect 76638 4454 76690 4506
rect 76974 4510 77026 4562
rect 86494 4510 86546 4562
rect 87278 4510 87330 4562
rect 87838 4510 87890 4562
rect 90638 4510 90690 4562
rect 105870 4510 105922 4562
rect 110798 4510 110850 4562
rect 113934 4510 113986 4562
rect 115502 4510 115554 4562
rect 122894 4510 122946 4562
rect 132526 4510 132578 4562
rect 142830 4510 142882 4562
rect 149998 4510 150050 4562
rect 67678 4398 67730 4450
rect 69470 4398 69522 4450
rect 73950 4398 74002 4450
rect 79102 4398 79154 4450
rect 82350 4398 82402 4450
rect 83694 4398 83746 4450
rect 89966 4398 90018 4450
rect 92766 4398 92818 4450
rect 94558 4398 94610 4450
rect 99038 4398 99090 4450
rect 101278 4398 101330 4450
rect 101614 4398 101666 4450
rect 104750 4398 104802 4450
rect 110910 4398 110962 4450
rect 113038 4398 113090 4450
rect 115950 4398 116002 4450
rect 119758 4398 119810 4450
rect 121102 4398 121154 4450
rect 121438 4398 121490 4450
rect 122782 4398 122834 4450
rect 126030 4398 126082 4450
rect 127262 4398 127314 4450
rect 129950 4398 130002 4450
rect 131742 4398 131794 4450
rect 135774 4398 135826 4450
rect 136222 4398 136274 4450
rect 137790 4398 137842 4450
rect 141374 4398 141426 4450
rect 144174 4398 144226 4450
rect 148878 4398 148930 4450
rect 149662 4398 149714 4450
rect 13470 4286 13522 4338
rect 15934 4286 15986 4338
rect 16606 4286 16658 4338
rect 17390 4286 17442 4338
rect 22318 4286 22370 4338
rect 22878 4286 22930 4338
rect 24110 4286 24162 4338
rect 24446 4286 24498 4338
rect 25230 4286 25282 4338
rect 25566 4286 25618 4338
rect 25678 4286 25730 4338
rect 29822 4286 29874 4338
rect 33182 4286 33234 4338
rect 34078 4286 34130 4338
rect 36318 4286 36370 4338
rect 38222 4286 38274 4338
rect 40238 4286 40290 4338
rect 41134 4286 41186 4338
rect 41358 4286 41410 4338
rect 41582 4286 41634 4338
rect 43038 4286 43090 4338
rect 48750 4286 48802 4338
rect 51326 4286 51378 4338
rect 51886 4286 51938 4338
rect 55806 4286 55858 4338
rect 61742 4286 61794 4338
rect 64542 4286 64594 4338
rect 66558 4286 66610 4338
rect 68798 4286 68850 4338
rect 72830 4286 72882 4338
rect 73166 4286 73218 4338
rect 82910 4286 82962 4338
rect 86270 4286 86322 4338
rect 86942 4286 86994 4338
rect 87166 4286 87218 4338
rect 87502 4286 87554 4338
rect 98366 4286 98418 4338
rect 105646 4286 105698 4338
rect 106430 4286 106482 4338
rect 109342 4286 109394 4338
rect 109678 4286 109730 4338
rect 110574 4286 110626 4338
rect 112590 4286 112642 4338
rect 115390 4286 115442 4338
rect 117742 4286 117794 4338
rect 117854 4286 117906 4338
rect 124574 4286 124626 4338
rect 124910 4286 124962 4338
rect 127598 4286 127650 4338
rect 127822 4286 127874 4338
rect 132750 4286 132802 4338
rect 135550 4286 135602 4338
rect 137342 4286 137394 4338
rect 141486 4286 141538 4338
rect 141710 4286 141762 4338
rect 141934 4286 141986 4338
rect 142046 4286 142098 4338
rect 143054 4286 143106 4338
rect 13246 4174 13298 4226
rect 15038 4174 15090 4226
rect 18398 4174 18450 4226
rect 19406 4174 19458 4226
rect 26126 4174 26178 4226
rect 27022 4174 27074 4226
rect 30606 4174 30658 4226
rect 31054 4174 31106 4226
rect 33742 4174 33794 4226
rect 35310 4174 35362 4226
rect 39902 4174 39954 4226
rect 41694 4174 41746 4226
rect 42142 4174 42194 4226
rect 43710 4174 43762 4226
rect 45838 4174 45890 4226
rect 47630 4174 47682 4226
rect 55134 4174 55186 4226
rect 58382 4174 58434 4226
rect 58942 4174 58994 4226
rect 62638 4174 62690 4226
rect 71486 4174 71538 4226
rect 76078 4174 76130 4226
rect 80110 4174 80162 4226
rect 85822 4174 85874 4226
rect 93550 4174 93602 4226
rect 102958 4174 103010 4226
rect 103742 4174 103794 4226
rect 109566 4174 109618 4226
rect 112254 4174 112306 4226
rect 115166 4174 115218 4226
rect 117966 4174 118018 4226
rect 120766 4174 120818 4226
rect 121886 4174 121938 4226
rect 122334 4174 122386 4226
rect 130734 4174 130786 4226
rect 135102 4174 135154 4226
rect 138910 4174 138962 4226
rect 139582 4174 139634 4226
rect 143614 4174 143666 4226
rect 145294 4174 145346 4226
rect 146190 4174 146242 4226
rect 147534 4174 147586 4226
rect 147870 4174 147922 4226
rect 15486 4062 15538 4114
rect 96014 4062 96066 4114
rect 107214 4062 107266 4114
rect 109230 4062 109282 4114
rect 118414 4062 118466 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 96638 3894 96690 3946
rect 96742 3894 96794 3946
rect 96846 3894 96898 3946
rect 127358 3894 127410 3946
rect 127462 3894 127514 3946
rect 127566 3894 127618 3946
rect 158078 3894 158130 3946
rect 158182 3894 158234 3946
rect 158286 3894 158338 3946
rect 93214 3726 93266 3778
rect 11342 3614 11394 3666
rect 13358 3614 13410 3666
rect 17054 3614 17106 3666
rect 18510 3614 18562 3666
rect 18734 3614 18786 3666
rect 20974 3614 21026 3666
rect 25454 3614 25506 3666
rect 32174 3614 32226 3666
rect 34302 3614 34354 3666
rect 36766 3614 36818 3666
rect 38894 3614 38946 3666
rect 40798 3614 40850 3666
rect 45502 3614 45554 3666
rect 55022 3614 55074 3666
rect 57150 3614 57202 3666
rect 59054 3614 59106 3666
rect 64878 3614 64930 3666
rect 66446 3614 66498 3666
rect 68574 3614 68626 3666
rect 70478 3614 70530 3666
rect 74846 3614 74898 3666
rect 78990 3614 79042 3666
rect 83022 3614 83074 3666
rect 90190 3614 90242 3666
rect 93102 3614 93154 3666
rect 94110 3614 94162 3666
rect 97918 3614 97970 3666
rect 101950 3614 102002 3666
rect 104750 3614 104802 3666
rect 112926 3614 112978 3666
rect 120990 3614 121042 3666
rect 124574 3614 124626 3666
rect 128382 3614 128434 3666
rect 136110 3614 136162 3666
rect 139806 3614 139858 3666
rect 143614 3614 143666 3666
rect 149774 3614 149826 3666
rect 151566 3614 151618 3666
rect 15262 3502 15314 3554
rect 16270 3502 16322 3554
rect 23326 3502 23378 3554
rect 23774 3502 23826 3554
rect 27806 3502 27858 3554
rect 28702 3502 28754 3554
rect 31166 3502 31218 3554
rect 34974 3502 35026 3554
rect 35982 3502 36034 3554
rect 40014 3502 40066 3554
rect 42926 3502 42978 3554
rect 43710 3502 43762 3554
rect 46846 3502 46898 3554
rect 47630 3502 47682 3554
rect 48526 3502 48578 3554
rect 51214 3502 51266 3554
rect 52110 3502 52162 3554
rect 57822 3502 57874 3554
rect 61406 3502 61458 3554
rect 61966 3502 62018 3554
rect 62862 3502 62914 3554
rect 65886 3502 65938 3554
rect 69246 3502 69298 3554
rect 72382 3502 72434 3554
rect 73502 3502 73554 3554
rect 76526 3502 76578 3554
rect 77198 3502 77250 3554
rect 77982 3502 78034 3554
rect 80782 3502 80834 3554
rect 81118 3502 81170 3554
rect 82014 3502 82066 3554
rect 85486 3502 85538 3554
rect 85822 3502 85874 3554
rect 86046 3502 86098 3554
rect 89630 3502 89682 3554
rect 92318 3502 92370 3554
rect 95006 3502 95058 3554
rect 95230 3502 95282 3554
rect 97246 3502 97298 3554
rect 99710 3502 99762 3554
rect 100942 3502 100994 3554
rect 103966 3502 104018 3554
rect 107550 3502 107602 3554
rect 108670 3502 108722 3554
rect 109006 3502 109058 3554
rect 113262 3502 113314 3554
rect 115278 3502 115330 3554
rect 116174 3502 116226 3554
rect 119086 3502 119138 3554
rect 119758 3502 119810 3554
rect 122894 3502 122946 3554
rect 123566 3502 123618 3554
rect 126702 3502 126754 3554
rect 127374 3502 127426 3554
rect 130398 3502 130450 3554
rect 131182 3502 131234 3554
rect 134318 3502 134370 3554
rect 134990 3502 135042 3554
rect 138238 3502 138290 3554
rect 139246 3502 139298 3554
rect 142046 3502 142098 3554
rect 142606 3502 142658 3554
rect 145854 3502 145906 3554
rect 146526 3502 146578 3554
rect 150558 3502 150610 3554
rect 10558 3390 10610 3442
rect 10782 3390 10834 3442
rect 16046 3390 16098 3442
rect 17502 3390 17554 3442
rect 18062 3390 18114 3442
rect 19742 3390 19794 3442
rect 23998 3390 24050 3442
rect 24558 3390 24610 3442
rect 28366 3390 28418 3442
rect 42702 3390 42754 3442
rect 43934 3390 43986 3442
rect 47406 3390 47458 3442
rect 49646 3390 49698 3442
rect 51550 3390 51602 3442
rect 53566 3390 53618 3442
rect 61742 3390 61794 3442
rect 62638 3390 62690 3442
rect 73166 3390 73218 3442
rect 76078 3390 76130 3442
rect 76974 3390 77026 3442
rect 81006 3390 81058 3442
rect 85598 3390 85650 3442
rect 89294 3390 89346 3442
rect 94334 3390 94386 3442
rect 96910 3390 96962 3442
rect 100718 3390 100770 3442
rect 106878 3390 106930 3442
rect 107326 3390 107378 3442
rect 108334 3390 108386 3442
rect 113710 3390 113762 3442
rect 117630 3390 117682 3442
rect 118862 3390 118914 3442
rect 122670 3390 122722 3442
rect 126478 3390 126530 3442
rect 132750 3390 132802 3442
rect 134094 3390 134146 3442
rect 137902 3390 137954 3442
rect 141710 3390 141762 3442
rect 145518 3390 145570 3442
rect 24894 3278 24946 3330
rect 30606 3278 30658 3330
rect 74286 3278 74338 3330
rect 87054 3278 87106 3330
rect 110014 3278 110066 3330
rect 114606 3278 114658 3330
rect 115054 3278 115106 3330
rect 147534 3278 147586 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 81278 3110 81330 3162
rect 81382 3110 81434 3162
rect 81486 3110 81538 3162
rect 111998 3110 112050 3162
rect 112102 3110 112154 3162
rect 112206 3110 112258 3162
rect 142718 3110 142770 3162
rect 142822 3110 142874 3162
rect 142926 3110 142978 3162
<< metal2 >>
rect 5600 59200 5712 60000
rect 9408 59200 9520 60000
rect 13216 59200 13328 60000
rect 17024 59200 17136 60000
rect 20832 59200 20944 60000
rect 24640 59200 24752 60000
rect 28448 59200 28560 60000
rect 32256 59200 32368 60000
rect 36064 59200 36176 60000
rect 39872 59200 39984 60000
rect 43680 59200 43792 60000
rect 47488 59200 47600 60000
rect 51296 59200 51408 60000
rect 55104 59200 55216 60000
rect 58912 59200 59024 60000
rect 62720 59200 62832 60000
rect 66528 59200 66640 60000
rect 70336 59200 70448 60000
rect 74144 59200 74256 60000
rect 77952 59200 78064 60000
rect 81760 59200 81872 60000
rect 85568 59200 85680 60000
rect 89376 59200 89488 60000
rect 93184 59200 93296 60000
rect 96992 59200 97104 60000
rect 100800 59200 100912 60000
rect 104608 59200 104720 60000
rect 108416 59200 108528 60000
rect 112224 59200 112336 60000
rect 116032 59200 116144 60000
rect 119840 59200 119952 60000
rect 123648 59200 123760 60000
rect 127456 59200 127568 60000
rect 131264 59200 131376 60000
rect 135072 59200 135184 60000
rect 138880 59200 138992 60000
rect 142688 59200 142800 60000
rect 146496 59200 146608 60000
rect 150304 59200 150416 60000
rect 154112 59200 154224 60000
rect 5068 56308 5124 56318
rect 5628 56308 5684 59200
rect 5852 56308 5908 56318
rect 5068 56306 5908 56308
rect 5068 56254 5070 56306
rect 5122 56254 5854 56306
rect 5906 56254 5908 56306
rect 5068 56252 5908 56254
rect 13244 56308 13300 59200
rect 13468 56308 13524 56318
rect 13244 56306 13524 56308
rect 13244 56254 13470 56306
rect 13522 56254 13524 56306
rect 13244 56252 13524 56254
rect 5068 56242 5124 56252
rect 5852 56242 5908 56252
rect 13468 56242 13524 56252
rect 6188 56196 6244 56206
rect 6188 56102 6244 56140
rect 9212 56196 9268 56206
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 9212 17108 9268 56140
rect 17052 55972 17108 59200
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 24668 56308 24724 59200
rect 24892 56308 24948 56318
rect 24668 56306 24948 56308
rect 24668 56254 24894 56306
rect 24946 56254 24948 56306
rect 24668 56252 24948 56254
rect 24892 56242 24948 56252
rect 28476 56308 28532 59200
rect 28476 56242 28532 56252
rect 29708 56308 29764 56318
rect 36092 56308 36148 59200
rect 36316 56308 36372 56318
rect 36092 56306 36372 56308
rect 36092 56254 36318 56306
rect 36370 56254 36372 56306
rect 36092 56252 36372 56254
rect 29708 56214 29764 56252
rect 36316 56242 36372 56252
rect 19852 56082 19908 56094
rect 28700 56084 28756 56094
rect 19852 56030 19854 56082
rect 19906 56030 19908 56082
rect 17500 55972 17556 55982
rect 17052 55970 17556 55972
rect 17052 55918 17502 55970
rect 17554 55918 17556 55970
rect 17052 55916 17556 55918
rect 17500 55906 17556 55916
rect 19852 55972 19908 56030
rect 28364 56082 28756 56084
rect 28364 56030 28702 56082
rect 28754 56030 28756 56082
rect 28364 56028 28756 56030
rect 19852 55906 19908 55916
rect 20972 55972 21028 55982
rect 20972 55878 21028 55916
rect 27916 55972 27972 55982
rect 27916 55076 27972 55916
rect 28364 55522 28420 56028
rect 28700 56018 28756 56028
rect 39900 55972 39956 59200
rect 47516 56308 47572 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 47740 56308 47796 56318
rect 47516 56306 47796 56308
rect 47516 56254 47742 56306
rect 47794 56254 47796 56306
rect 47516 56252 47796 56254
rect 47740 56242 47796 56252
rect 51324 56308 51380 59200
rect 51324 56242 51380 56252
rect 52556 56308 52612 56318
rect 52556 56214 52612 56252
rect 55132 56308 55188 59200
rect 55356 56308 55412 56318
rect 55132 56306 55412 56308
rect 55132 56254 55358 56306
rect 55410 56254 55412 56306
rect 55132 56252 55412 56254
rect 42700 56082 42756 56094
rect 42700 56030 42702 56082
rect 42754 56030 42756 56082
rect 40348 55972 40404 55982
rect 39900 55970 40404 55972
rect 39900 55918 40350 55970
rect 40402 55918 40404 55970
rect 39900 55916 40404 55918
rect 40348 55906 40404 55916
rect 42700 55972 42756 56030
rect 50092 56084 50148 56094
rect 42700 55906 42756 55916
rect 43820 55972 43876 55982
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 28364 55470 28366 55522
rect 28418 55470 28420 55522
rect 28364 55458 28420 55470
rect 43820 55468 43876 55916
rect 43708 55412 43876 55468
rect 28476 55186 28532 55198
rect 28476 55134 28478 55186
rect 28530 55134 28532 55186
rect 28364 55076 28420 55086
rect 27916 55074 28420 55076
rect 27916 55022 27918 55074
rect 27970 55022 28366 55074
rect 28418 55022 28420 55074
rect 27916 55020 28420 55022
rect 27916 55010 27972 55020
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 26908 27858 26964 27870
rect 26908 27806 26910 27858
rect 26962 27806 26964 27858
rect 26908 27748 26964 27806
rect 24444 26852 24500 26862
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 24220 26516 24276 26526
rect 24444 26516 24500 26796
rect 25788 26852 25844 26862
rect 24220 26514 24500 26516
rect 24220 26462 24222 26514
rect 24274 26462 24500 26514
rect 24220 26460 24500 26462
rect 24220 26450 24276 26460
rect 24444 26402 24500 26460
rect 25340 26628 25396 26638
rect 24444 26350 24446 26402
rect 24498 26350 24500 26402
rect 24444 26338 24500 26350
rect 24556 26402 24612 26414
rect 24556 26350 24558 26402
rect 24610 26350 24612 26402
rect 23436 25508 23492 25518
rect 23436 25414 23492 25452
rect 24556 25508 24612 26350
rect 24780 26292 24836 26302
rect 24780 26198 24836 26236
rect 25340 26290 25396 26572
rect 25788 26514 25844 26796
rect 26348 26852 26404 26862
rect 26348 26758 26404 26796
rect 26684 26628 26740 26638
rect 25788 26462 25790 26514
rect 25842 26462 25844 26514
rect 25788 26450 25844 26462
rect 26012 26516 26068 26526
rect 26012 26422 26068 26460
rect 26684 26514 26740 26572
rect 26684 26462 26686 26514
rect 26738 26462 26740 26514
rect 26684 26450 26740 26462
rect 25340 26238 25342 26290
rect 25394 26238 25396 26290
rect 25340 26226 25396 26238
rect 25564 26292 25620 26302
rect 25564 26198 25620 26236
rect 23436 25284 23492 25294
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 23436 24946 23492 25228
rect 23436 24894 23438 24946
rect 23490 24894 23492 24946
rect 23436 24882 23492 24894
rect 24556 24834 24612 25452
rect 25788 26178 25844 26190
rect 25788 26126 25790 26178
rect 25842 26126 25844 26178
rect 25788 25506 25844 26126
rect 25788 25454 25790 25506
rect 25842 25454 25844 25506
rect 25788 25442 25844 25454
rect 26572 25506 26628 25518
rect 26572 25454 26574 25506
rect 26626 25454 26628 25506
rect 26572 25284 26628 25454
rect 26908 25284 26964 27692
rect 27580 27746 27636 27758
rect 27580 27694 27582 27746
rect 27634 27694 27636 27746
rect 27580 26908 27636 27694
rect 27356 26852 27636 26908
rect 27020 26628 27076 26638
rect 27020 26292 27076 26572
rect 27132 26516 27188 26526
rect 27132 26422 27188 26460
rect 27020 26236 27188 26292
rect 26572 25282 26964 25284
rect 26572 25230 26910 25282
rect 26962 25230 26964 25282
rect 26572 25228 26964 25230
rect 24556 24782 24558 24834
rect 24610 24782 24612 24834
rect 24556 24770 24612 24782
rect 24444 24722 24500 24734
rect 24444 24670 24446 24722
rect 24498 24670 24500 24722
rect 23772 24500 23828 24510
rect 23548 24498 23828 24500
rect 23548 24446 23774 24498
rect 23826 24446 23828 24498
rect 23548 24444 23828 24446
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 21868 23154 21924 23166
rect 21868 23102 21870 23154
rect 21922 23102 21924 23154
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 21084 21812 21140 21822
rect 21084 21586 21140 21756
rect 21868 21812 21924 23102
rect 22540 23044 22596 23054
rect 22540 22950 22596 22988
rect 23324 23044 23380 23054
rect 23324 22482 23380 22988
rect 23324 22430 23326 22482
rect 23378 22430 23380 22482
rect 23324 22418 23380 22430
rect 21924 21756 22036 21812
rect 21868 21746 21924 21756
rect 21084 21534 21086 21586
rect 21138 21534 21140 21586
rect 21084 21522 21140 21534
rect 21868 21476 21924 21486
rect 21868 21382 21924 21420
rect 21980 20916 22036 21756
rect 21980 20850 22036 20860
rect 23324 21476 23380 21486
rect 23324 20914 23380 21420
rect 23324 20862 23326 20914
rect 23378 20862 23380 20914
rect 23324 20850 23380 20862
rect 23548 20692 23604 24444
rect 23772 24434 23828 24444
rect 23772 22932 23828 22942
rect 23660 22260 23716 22270
rect 23660 22166 23716 22204
rect 23772 22258 23828 22876
rect 23772 22206 23774 22258
rect 23826 22206 23828 22258
rect 23772 22194 23828 22206
rect 23884 22260 23940 22270
rect 23884 22166 23940 22204
rect 24108 22146 24164 22158
rect 24108 22094 24110 22146
rect 24162 22094 24164 22146
rect 23996 21700 24052 21710
rect 24108 21700 24164 22094
rect 24444 21924 24500 24670
rect 26908 24612 26964 25228
rect 26908 24546 26964 24556
rect 27020 23714 27076 23726
rect 27020 23662 27022 23714
rect 27074 23662 27076 23714
rect 24668 23380 24724 23390
rect 24668 23042 24724 23324
rect 25340 23380 25396 23390
rect 25340 23286 25396 23324
rect 24668 22990 24670 23042
rect 24722 22990 24724 23042
rect 24668 22978 24724 22990
rect 25452 23154 25508 23166
rect 25452 23102 25454 23154
rect 25506 23102 25508 23154
rect 25340 22932 25396 22942
rect 25340 22838 25396 22876
rect 25452 22372 25508 23102
rect 25452 22306 25508 22316
rect 25900 23042 25956 23054
rect 25900 22990 25902 23042
rect 25954 22990 25956 23042
rect 24780 22260 24836 22270
rect 24836 22204 24948 22260
rect 24780 22194 24836 22204
rect 24444 21868 24724 21924
rect 23884 21644 23996 21700
rect 24052 21644 24164 21700
rect 24444 21698 24500 21710
rect 24444 21646 24446 21698
rect 24498 21646 24500 21698
rect 23884 21252 23940 21644
rect 23996 21634 24052 21644
rect 24220 21588 24276 21598
rect 24108 21586 24276 21588
rect 24108 21534 24222 21586
rect 24274 21534 24276 21586
rect 24108 21532 24276 21534
rect 23996 21474 24052 21486
rect 23996 21422 23998 21474
rect 24050 21422 24052 21474
rect 23996 21364 24052 21422
rect 23996 21298 24052 21308
rect 23884 21186 23940 21196
rect 23324 20636 23604 20692
rect 23660 21028 23716 21038
rect 24108 21028 24164 21532
rect 24220 21522 24276 21532
rect 24444 21364 24500 21646
rect 24444 21298 24500 21308
rect 24556 21586 24612 21598
rect 24556 21534 24558 21586
rect 24610 21534 24612 21586
rect 23660 20690 23716 20972
rect 23660 20638 23662 20690
rect 23714 20638 23716 20690
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 21980 20244 22036 20254
rect 19180 20018 19236 20030
rect 19180 19966 19182 20018
rect 19234 19966 19236 20018
rect 19180 18564 19236 19966
rect 19852 19908 19908 19918
rect 19852 19814 19908 19852
rect 21980 19906 22036 20188
rect 23324 20244 23380 20636
rect 23660 20626 23716 20638
rect 23772 20972 24164 21028
rect 24220 21252 24276 21262
rect 23772 20690 23828 20972
rect 24108 20804 24164 20814
rect 24220 20804 24276 21196
rect 24556 21140 24612 21534
rect 24108 20802 24276 20804
rect 24108 20750 24110 20802
rect 24162 20750 24276 20802
rect 24108 20748 24276 20750
rect 24332 21084 24612 21140
rect 24108 20738 24164 20748
rect 23772 20638 23774 20690
rect 23826 20638 23828 20690
rect 23772 20626 23828 20638
rect 23884 20580 23940 20590
rect 23884 20578 24276 20580
rect 23884 20526 23886 20578
rect 23938 20526 24276 20578
rect 23884 20524 24276 20526
rect 23884 20514 23940 20524
rect 23884 20356 23940 20366
rect 23324 20130 23380 20188
rect 23324 20078 23326 20130
rect 23378 20078 23380 20130
rect 23324 20066 23380 20078
rect 23772 20300 23884 20356
rect 23100 20018 23156 20030
rect 23100 19966 23102 20018
rect 23154 19966 23156 20018
rect 21980 19854 21982 19906
rect 22034 19854 22036 19906
rect 21980 19842 22036 19854
rect 22428 19906 22484 19918
rect 22428 19854 22430 19906
rect 22482 19854 22484 19906
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19180 18498 19236 18508
rect 21532 18564 21588 18574
rect 21532 18450 21588 18508
rect 22428 18564 22484 19854
rect 22764 19908 22820 19918
rect 22764 19458 22820 19852
rect 22764 19406 22766 19458
rect 22818 19406 22820 19458
rect 22764 19394 22820 19406
rect 23100 19234 23156 19966
rect 23100 19182 23102 19234
rect 23154 19182 23156 19234
rect 23100 19170 23156 19182
rect 23436 20018 23492 20030
rect 23436 19966 23438 20018
rect 23490 19966 23492 20018
rect 23436 19236 23492 19966
rect 23436 19170 23492 19180
rect 23324 19122 23380 19134
rect 23324 19070 23326 19122
rect 23378 19070 23380 19122
rect 22876 19010 22932 19022
rect 22876 18958 22878 19010
rect 22930 18958 22932 19010
rect 22876 18676 22932 18958
rect 22876 18610 22932 18620
rect 22428 18498 22484 18508
rect 21532 18398 21534 18450
rect 21586 18398 21588 18450
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 9212 17042 9268 17052
rect 19628 17108 19684 17118
rect 19628 17014 19684 17052
rect 20188 17108 20244 17118
rect 19292 16882 19348 16894
rect 19292 16830 19294 16882
rect 19346 16830 19348 16882
rect 19292 16772 19348 16830
rect 20188 16882 20244 17052
rect 20188 16830 20190 16882
rect 20242 16830 20244 16882
rect 20188 16818 20244 16830
rect 19292 16706 19348 16716
rect 20300 16772 20356 16782
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 17948 16100 18004 16110
rect 17948 16006 18004 16044
rect 9212 15988 9268 15998
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 9212 800 9268 15932
rect 18620 15986 18676 15998
rect 18620 15934 18622 15986
rect 18674 15934 18676 15986
rect 18620 15540 18676 15934
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 18620 15474 18676 15484
rect 19628 15316 19684 15326
rect 17164 14530 17220 14542
rect 17164 14478 17166 14530
rect 17218 14478 17220 14530
rect 17164 14308 17220 14478
rect 17164 14242 17220 14252
rect 17836 14418 17892 14430
rect 17836 14366 17838 14418
rect 17890 14366 17892 14418
rect 17836 13076 17892 14366
rect 17836 13010 17892 13020
rect 19068 13524 19124 13534
rect 18620 12740 18676 12750
rect 15596 12404 15652 12414
rect 15596 11506 15652 12348
rect 18172 12404 18228 12414
rect 18172 12310 18228 12348
rect 18620 12402 18676 12684
rect 19068 12738 19124 13468
rect 19628 12964 19684 15260
rect 20300 15148 20356 16716
rect 20748 16212 20804 16222
rect 20748 16118 20804 16156
rect 20412 16100 20468 16110
rect 21532 16100 21588 18398
rect 22204 18340 22260 18350
rect 22204 18338 23268 18340
rect 22204 18286 22206 18338
rect 22258 18286 23268 18338
rect 22204 18284 23268 18286
rect 22204 18274 22260 18284
rect 22652 17892 22708 17902
rect 22652 17890 22932 17892
rect 22652 17838 22654 17890
rect 22706 17838 22932 17890
rect 22652 17836 22932 17838
rect 22652 17826 22708 17836
rect 22764 17668 22820 17678
rect 22876 17668 22932 17836
rect 23212 17890 23268 18284
rect 23212 17838 23214 17890
rect 23266 17838 23268 17890
rect 23212 17826 23268 17838
rect 23324 17892 23380 19070
rect 23772 19122 23828 20300
rect 23884 20290 23940 20300
rect 23996 20244 24052 20254
rect 23884 19236 23940 19246
rect 23884 19142 23940 19180
rect 23772 19070 23774 19122
rect 23826 19070 23828 19122
rect 23772 19058 23828 19070
rect 23548 19012 23604 19022
rect 23324 17826 23380 17836
rect 23436 19010 23604 19012
rect 23436 18958 23550 19010
rect 23602 18958 23604 19010
rect 23436 18956 23604 18958
rect 22988 17668 23044 17678
rect 22876 17666 23044 17668
rect 22876 17614 22990 17666
rect 23042 17614 23044 17666
rect 22876 17612 23044 17614
rect 22764 17574 22820 17612
rect 22988 17602 23044 17612
rect 23324 17668 23380 17678
rect 23436 17668 23492 18956
rect 23548 18946 23604 18956
rect 23996 18452 24052 20188
rect 23884 18396 24052 18452
rect 23772 17892 23828 17902
rect 23324 17666 23492 17668
rect 23324 17614 23326 17666
rect 23378 17614 23492 17666
rect 23324 17612 23492 17614
rect 23548 17780 23604 17790
rect 23324 17602 23380 17612
rect 23548 17554 23604 17724
rect 23772 17666 23828 17836
rect 23772 17614 23774 17666
rect 23826 17614 23828 17666
rect 23772 17602 23828 17614
rect 23548 17502 23550 17554
rect 23602 17502 23604 17554
rect 23548 17490 23604 17502
rect 23884 17556 23940 18396
rect 24108 17668 24164 17678
rect 24108 17574 24164 17612
rect 23996 17556 24052 17566
rect 23884 17554 24052 17556
rect 23884 17502 23998 17554
rect 24050 17502 24052 17554
rect 23884 17500 24052 17502
rect 22316 17444 22372 17454
rect 22652 17444 22708 17454
rect 22316 17442 22708 17444
rect 22316 17390 22318 17442
rect 22370 17390 22654 17442
rect 22706 17390 22708 17442
rect 22316 17388 22708 17390
rect 22316 17378 22372 17388
rect 22652 17220 22708 17388
rect 23884 17332 23940 17500
rect 23996 17490 24052 17500
rect 21644 16996 21700 17006
rect 21644 16902 21700 16940
rect 21644 16100 21700 16110
rect 21532 16044 21644 16100
rect 20412 15538 20468 16044
rect 21644 16006 21700 16044
rect 22428 15986 22484 15998
rect 22428 15934 22430 15986
rect 22482 15934 22484 15986
rect 20412 15486 20414 15538
rect 20466 15486 20468 15538
rect 20412 15474 20468 15486
rect 20748 15540 20804 15550
rect 20972 15540 21028 15550
rect 20748 15446 20804 15484
rect 20860 15484 20972 15540
rect 20860 15426 20916 15484
rect 20972 15474 21028 15484
rect 22316 15540 22372 15550
rect 22428 15540 22484 15934
rect 22316 15538 22484 15540
rect 22316 15486 22318 15538
rect 22370 15486 22484 15538
rect 22316 15484 22484 15486
rect 22316 15474 22372 15484
rect 20860 15374 20862 15426
rect 20914 15374 20916 15426
rect 20860 15362 20916 15374
rect 21980 15426 22036 15438
rect 21980 15374 21982 15426
rect 22034 15374 22036 15426
rect 20636 15316 20692 15326
rect 20636 15222 20692 15260
rect 21196 15314 21252 15326
rect 21196 15262 21198 15314
rect 21250 15262 21252 15314
rect 20300 15092 20692 15148
rect 19964 14642 20020 14654
rect 19964 14590 19966 14642
rect 20018 14590 20020 14642
rect 19964 14308 20020 14590
rect 20412 14308 20468 14318
rect 19964 14252 20244 14308
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20076 13972 20132 13982
rect 20188 13972 20244 14252
rect 20412 14214 20468 14252
rect 20132 13916 20244 13972
rect 20076 13746 20132 13916
rect 20076 13694 20078 13746
rect 20130 13694 20132 13746
rect 20076 13682 20132 13694
rect 19740 13634 19796 13646
rect 19740 13582 19742 13634
rect 19794 13582 19796 13634
rect 19740 13524 19796 13582
rect 19740 13458 19796 13468
rect 20188 13634 20244 13646
rect 20188 13582 20190 13634
rect 20242 13582 20244 13634
rect 20076 13300 20132 13310
rect 19852 13076 19908 13086
rect 19852 12982 19908 13020
rect 19740 12964 19796 12974
rect 19404 12962 19796 12964
rect 19404 12910 19742 12962
rect 19794 12910 19796 12962
rect 19404 12908 19796 12910
rect 19404 12850 19460 12908
rect 19404 12798 19406 12850
rect 19458 12798 19460 12850
rect 19404 12786 19460 12798
rect 19068 12686 19070 12738
rect 19122 12686 19124 12738
rect 19068 12628 19124 12686
rect 18620 12350 18622 12402
rect 18674 12350 18676 12402
rect 18620 12338 18676 12350
rect 18844 12572 19124 12628
rect 15596 11454 15598 11506
rect 15650 11454 15652 11506
rect 15596 11442 15652 11454
rect 17724 12180 17780 12190
rect 17724 11506 17780 12124
rect 17724 11454 17726 11506
rect 17778 11454 17780 11506
rect 17724 11442 17780 11454
rect 18508 11394 18564 11406
rect 18508 11342 18510 11394
rect 18562 11342 18564 11394
rect 18172 11172 18228 11182
rect 16940 10724 16996 10734
rect 15932 7812 15988 7822
rect 15932 5346 15988 7756
rect 16940 7812 16996 10668
rect 18172 10722 18228 11116
rect 18172 10670 18174 10722
rect 18226 10670 18228 10722
rect 18172 10658 18228 10670
rect 17500 10612 17556 10622
rect 17500 10518 17556 10556
rect 18508 10612 18564 11342
rect 18844 11284 18900 12572
rect 18956 12404 19012 12414
rect 18956 12310 19012 12348
rect 19516 12290 19572 12908
rect 19740 12898 19796 12908
rect 20076 12962 20132 13244
rect 20188 13186 20244 13582
rect 20412 13524 20468 13534
rect 20412 13430 20468 13468
rect 20188 13134 20190 13186
rect 20242 13134 20244 13186
rect 20188 13122 20244 13134
rect 20076 12910 20078 12962
rect 20130 12910 20132 12962
rect 20076 12898 20132 12910
rect 20300 12962 20356 12974
rect 20300 12910 20302 12962
rect 20354 12910 20356 12962
rect 19628 12740 19684 12750
rect 19628 12404 19684 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19628 12348 19796 12404
rect 19516 12238 19518 12290
rect 19570 12238 19572 12290
rect 19516 12226 19572 12238
rect 19740 12292 19796 12348
rect 19740 12290 19908 12292
rect 19740 12238 19742 12290
rect 19794 12238 19908 12290
rect 19740 12236 19908 12238
rect 19740 12226 19796 12236
rect 19628 12180 19684 12190
rect 19628 12086 19684 12124
rect 18956 12068 19012 12078
rect 18956 11974 19012 12012
rect 19180 11956 19236 11966
rect 19068 11900 19180 11956
rect 18956 11284 19012 11294
rect 18844 11228 18956 11284
rect 18956 11218 19012 11228
rect 19068 11282 19124 11900
rect 19180 11862 19236 11900
rect 19740 11732 19796 11742
rect 19740 11394 19796 11676
rect 19740 11342 19742 11394
rect 19794 11342 19796 11394
rect 19740 11330 19796 11342
rect 19068 11230 19070 11282
rect 19122 11230 19124 11282
rect 19068 11218 19124 11230
rect 19404 11284 19460 11294
rect 18508 9940 18564 10556
rect 19404 10050 19460 11228
rect 19852 11172 19908 12236
rect 20188 12180 20244 12190
rect 20300 12180 20356 12910
rect 20188 12178 20356 12180
rect 20188 12126 20190 12178
rect 20242 12126 20356 12178
rect 20188 12124 20356 12126
rect 19964 12068 20020 12078
rect 19964 11974 20020 12012
rect 20076 11508 20132 11518
rect 20076 11394 20132 11452
rect 20076 11342 20078 11394
rect 20130 11342 20132 11394
rect 20076 11330 20132 11342
rect 20188 11396 20244 12124
rect 20300 11620 20356 11630
rect 20300 11526 20356 11564
rect 20524 11396 20580 11406
rect 20188 11340 20524 11396
rect 20524 11302 20580 11340
rect 19404 9998 19406 10050
rect 19458 9998 19460 10050
rect 19404 9986 19460 9998
rect 19516 11116 19908 11172
rect 20188 11172 20244 11182
rect 18844 9940 18900 9950
rect 18508 9884 18844 9940
rect 18844 9846 18900 9884
rect 16940 7746 16996 7756
rect 17388 8258 17444 8270
rect 17388 8206 17390 8258
rect 17442 8206 17444 8258
rect 17388 7028 17444 8206
rect 18060 8148 18116 8158
rect 18060 8054 18116 8092
rect 19516 7252 19572 11116
rect 20188 11078 20244 11116
rect 20300 11060 20356 11070
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20300 10498 20356 11004
rect 20636 10724 20692 15092
rect 20972 13634 21028 13646
rect 20972 13582 20974 13634
rect 21026 13582 21028 13634
rect 20972 13524 21028 13582
rect 20972 13458 21028 13468
rect 21196 12402 21252 15262
rect 21420 13634 21476 13646
rect 21420 13582 21422 13634
rect 21474 13582 21476 13634
rect 21420 13300 21476 13582
rect 21420 13234 21476 13244
rect 21868 13524 21924 13534
rect 21868 13076 21924 13468
rect 21196 12350 21198 12402
rect 21250 12350 21252 12402
rect 21196 12338 21252 12350
rect 21308 13074 21924 13076
rect 21308 13022 21870 13074
rect 21922 13022 21924 13074
rect 21308 13020 21924 13022
rect 21308 12290 21364 13020
rect 21868 13010 21924 13020
rect 21980 12402 22036 15374
rect 22204 15428 22260 15438
rect 22204 15334 22260 15372
rect 22428 15316 22484 15326
rect 22428 15222 22484 15260
rect 22652 15148 22708 17164
rect 23548 17276 23940 17332
rect 23548 17106 23604 17276
rect 23548 17054 23550 17106
rect 23602 17054 23604 17106
rect 23548 17042 23604 17054
rect 22764 16772 22820 16782
rect 22764 15540 22820 16716
rect 22764 15446 22820 15484
rect 22876 16212 22932 16222
rect 22876 15428 22932 16156
rect 23324 15540 23380 15550
rect 23324 15428 23380 15484
rect 22876 15426 23380 15428
rect 22876 15374 22878 15426
rect 22930 15374 23326 15426
rect 23378 15374 23380 15426
rect 22876 15372 23380 15374
rect 22876 15362 22932 15372
rect 23324 15362 23380 15372
rect 22652 15092 23156 15148
rect 22652 14308 22708 14318
rect 22652 12964 22708 14252
rect 21980 12350 21982 12402
rect 22034 12350 22036 12402
rect 21980 12338 22036 12350
rect 22092 12962 22708 12964
rect 22092 12910 22654 12962
rect 22706 12910 22708 12962
rect 22092 12908 22708 12910
rect 21308 12238 21310 12290
rect 21362 12238 21364 12290
rect 20972 12180 21028 12190
rect 20972 12086 21028 12124
rect 21308 11844 21364 12238
rect 21308 11778 21364 11788
rect 21532 12292 21588 12302
rect 21420 11732 21476 11742
rect 21196 11620 21252 11630
rect 21252 11564 21364 11620
rect 21196 11554 21252 11564
rect 20300 10446 20302 10498
rect 20354 10446 20356 10498
rect 20300 10434 20356 10446
rect 20412 10722 20692 10724
rect 20412 10670 20638 10722
rect 20690 10670 20692 10722
rect 20412 10668 20692 10670
rect 19628 10050 19684 10062
rect 19628 9998 19630 10050
rect 19682 9998 19684 10050
rect 19628 9938 19684 9998
rect 19628 9886 19630 9938
rect 19682 9886 19684 9938
rect 19628 9874 19684 9886
rect 20300 9940 20356 9950
rect 20412 9940 20468 10668
rect 20636 10658 20692 10668
rect 20748 11508 20804 11518
rect 20300 9938 20468 9940
rect 20300 9886 20302 9938
rect 20354 9886 20468 9938
rect 20300 9884 20468 9886
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9268 20244 9278
rect 20188 8484 20244 9212
rect 20188 8370 20244 8428
rect 20188 8318 20190 8370
rect 20242 8318 20244 8370
rect 20188 8306 20244 8318
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19852 7476 19908 7486
rect 19852 7474 20020 7476
rect 19852 7422 19854 7474
rect 19906 7422 20020 7474
rect 19852 7420 20020 7422
rect 19852 7410 19908 7420
rect 19516 7196 19908 7252
rect 17388 6962 17444 6972
rect 18508 7028 18564 7038
rect 16828 6580 16884 6590
rect 16828 5460 16884 6524
rect 17836 6466 17892 6478
rect 17836 6414 17838 6466
rect 17890 6414 17892 6466
rect 17836 6020 17892 6414
rect 18396 6132 18452 6142
rect 18172 6020 18228 6030
rect 17836 6018 18228 6020
rect 17836 5966 18174 6018
rect 18226 5966 18228 6018
rect 17836 5964 18228 5966
rect 17836 5794 17892 5806
rect 17836 5742 17838 5794
rect 17890 5742 17892 5794
rect 15932 5294 15934 5346
rect 15986 5294 15988 5346
rect 15932 5282 15988 5294
rect 16380 5404 16884 5460
rect 16380 5236 16436 5404
rect 16380 5142 16436 5180
rect 16604 5236 16660 5246
rect 11340 5124 11396 5134
rect 11340 3666 11396 5068
rect 15372 5124 15428 5134
rect 15372 5122 15540 5124
rect 15372 5070 15374 5122
rect 15426 5070 15540 5122
rect 15372 5068 15540 5070
rect 15372 5058 15428 5068
rect 13804 4452 13860 4462
rect 13804 4358 13860 4396
rect 15484 4452 15540 5068
rect 15484 4358 15540 4396
rect 15596 5122 15652 5134
rect 15596 5070 15598 5122
rect 15650 5070 15652 5122
rect 13468 4338 13524 4350
rect 13468 4286 13470 4338
rect 13522 4286 13524 4338
rect 13244 4228 13300 4238
rect 13468 4228 13524 4286
rect 15596 4340 15652 5070
rect 15932 4340 15988 4350
rect 15596 4338 16100 4340
rect 15596 4286 15934 4338
rect 15986 4286 16100 4338
rect 15596 4284 16100 4286
rect 15932 4274 15988 4284
rect 13244 4226 13524 4228
rect 13244 4174 13246 4226
rect 13298 4174 13524 4226
rect 13244 4172 13524 4174
rect 15036 4226 15092 4238
rect 15036 4174 15038 4226
rect 15090 4174 15092 4226
rect 11340 3614 11342 3666
rect 11394 3614 11396 3666
rect 11340 3602 11396 3614
rect 11900 3668 11956 3678
rect 10556 3444 10612 3454
rect 10780 3444 10836 3454
rect 10556 3442 10836 3444
rect 10556 3390 10558 3442
rect 10610 3390 10782 3442
rect 10834 3390 10836 3442
rect 10556 3388 10836 3390
rect 10556 800 10612 3388
rect 10780 3378 10836 3388
rect 11900 800 11956 3612
rect 13244 800 13300 4172
rect 13356 3668 13412 3678
rect 13356 3574 13412 3612
rect 15036 3556 15092 4174
rect 15484 4116 15540 4126
rect 15484 4022 15540 4060
rect 15260 3556 15316 3566
rect 15036 3554 15316 3556
rect 15036 3502 15262 3554
rect 15314 3502 15316 3554
rect 15036 3500 15316 3502
rect 14588 3444 14644 3454
rect 14588 800 14644 3388
rect 15260 3388 15316 3500
rect 16044 3442 16100 4284
rect 16604 4338 16660 5180
rect 16828 5122 16884 5404
rect 17500 5572 17556 5582
rect 17500 5234 17556 5516
rect 17500 5182 17502 5234
rect 17554 5182 17556 5234
rect 17500 5170 17556 5182
rect 16828 5070 16830 5122
rect 16882 5070 16884 5122
rect 16828 5058 16884 5070
rect 17052 5124 17108 5134
rect 17052 5010 17108 5068
rect 17052 4958 17054 5010
rect 17106 4958 17108 5010
rect 17052 4946 17108 4958
rect 17836 5012 17892 5742
rect 17836 4946 17892 4956
rect 17948 4898 18004 4910
rect 17948 4846 17950 4898
rect 18002 4846 18004 4898
rect 16828 4452 16884 4462
rect 16828 4358 16884 4396
rect 17388 4340 17444 4350
rect 16604 4286 16606 4338
rect 16658 4286 16660 4338
rect 16604 4274 16660 4286
rect 17052 4338 17444 4340
rect 17052 4286 17390 4338
rect 17442 4286 17444 4338
rect 17052 4284 17444 4286
rect 16044 3390 16046 3442
rect 16098 3390 16100 3442
rect 15260 3332 15764 3388
rect 16044 3378 16100 3390
rect 16156 3668 16212 3678
rect 15708 2884 15764 3332
rect 15708 2818 15764 2828
rect 16156 2660 16212 3612
rect 17052 3668 17108 4284
rect 17388 4274 17444 4284
rect 17052 3574 17108 3612
rect 17836 4116 17892 4126
rect 16268 3554 16324 3566
rect 16268 3502 16270 3554
rect 16322 3502 16324 3554
rect 16268 3444 16324 3502
rect 16268 3378 16324 3388
rect 17500 3444 17556 3482
rect 17500 3378 17556 3388
rect 15932 2604 16212 2660
rect 15932 800 15988 2604
rect 17836 2548 17892 4060
rect 17948 3668 18004 4846
rect 17948 3602 18004 3612
rect 18060 3444 18116 3482
rect 18060 3378 18116 3388
rect 17836 2482 17892 2492
rect 17276 924 17668 980
rect 17276 800 17332 924
rect 9184 0 9296 800
rect 10528 0 10640 800
rect 11872 0 11984 800
rect 13216 0 13328 800
rect 14560 0 14672 800
rect 15904 0 16016 800
rect 17248 0 17360 800
rect 17612 756 17668 924
rect 18172 756 18228 5964
rect 18396 4226 18452 6076
rect 18396 4174 18398 4226
rect 18450 4174 18452 4226
rect 18396 4162 18452 4174
rect 18508 3666 18564 6972
rect 18620 6802 18676 6814
rect 18620 6750 18622 6802
rect 18674 6750 18676 6802
rect 18620 6692 18676 6750
rect 18620 6626 18676 6636
rect 19852 6690 19908 7196
rect 19964 7028 20020 7420
rect 20076 7028 20132 7038
rect 19964 6972 20076 7028
rect 19852 6638 19854 6690
rect 19906 6638 19908 6690
rect 19852 6626 19908 6638
rect 19068 6468 19124 6478
rect 19628 6468 19684 6478
rect 19068 6466 19348 6468
rect 19068 6414 19070 6466
rect 19122 6414 19348 6466
rect 19068 6412 19348 6414
rect 19068 6402 19124 6412
rect 19292 5794 19348 6412
rect 19292 5742 19294 5794
rect 19346 5742 19348 5794
rect 19292 5730 19348 5742
rect 19404 6412 19628 6468
rect 20076 6468 20132 6972
rect 20300 6916 20356 9884
rect 20748 9604 20804 11452
rect 21308 11506 21364 11564
rect 21308 11454 21310 11506
rect 21362 11454 21364 11506
rect 21308 11442 21364 11454
rect 21420 11282 21476 11676
rect 21420 11230 21422 11282
rect 21474 11230 21476 11282
rect 21420 11060 21476 11230
rect 21420 10994 21476 11004
rect 21532 10836 21588 12236
rect 21756 12180 21812 12190
rect 21756 12086 21812 12124
rect 22092 11844 22148 12908
rect 22652 12898 22708 12908
rect 22428 12292 22484 12302
rect 22428 12198 22484 12236
rect 22204 12180 22260 12190
rect 22204 12086 22260 12124
rect 22876 12180 22932 12190
rect 22876 12086 22932 12124
rect 21868 11788 22148 11844
rect 22204 11844 22260 11854
rect 21644 11284 21700 11294
rect 21644 11060 21700 11228
rect 21644 10994 21700 11004
rect 21644 10836 21700 10846
rect 21532 10834 21700 10836
rect 21532 10782 21646 10834
rect 21698 10782 21700 10834
rect 21532 10780 21700 10782
rect 20972 10722 21028 10734
rect 20972 10670 20974 10722
rect 21026 10670 21028 10722
rect 20972 10612 21028 10670
rect 20972 10546 21028 10556
rect 21420 10612 21476 10622
rect 21420 10518 21476 10556
rect 21532 10164 21588 10780
rect 21644 10770 21700 10780
rect 21420 10108 21588 10164
rect 21420 9716 21476 10108
rect 21868 10052 21924 11788
rect 22092 11170 22148 11182
rect 22092 11118 22094 11170
rect 22146 11118 22148 11170
rect 22092 11060 22148 11118
rect 22092 10994 22148 11004
rect 22092 10612 22148 10622
rect 22092 10518 22148 10556
rect 21532 9996 21924 10052
rect 21532 9940 21588 9996
rect 21532 9846 21588 9884
rect 21420 9660 21924 9716
rect 20748 9510 20804 9548
rect 20972 9268 21028 9278
rect 20972 9174 21028 9212
rect 21420 9156 21476 9166
rect 21756 9156 21812 9166
rect 21420 9154 21700 9156
rect 21420 9102 21422 9154
rect 21474 9102 21700 9154
rect 21420 9100 21700 9102
rect 21420 9090 21476 9100
rect 20412 8932 20468 8942
rect 20412 8838 20468 8876
rect 21532 8930 21588 8942
rect 21532 8878 21534 8930
rect 21586 8878 21588 8930
rect 21532 8484 21588 8878
rect 20748 8428 21588 8484
rect 20748 8258 20804 8428
rect 21644 8372 21700 9100
rect 21756 9062 21812 9100
rect 21868 9042 21924 9660
rect 21868 8990 21870 9042
rect 21922 8990 21924 9042
rect 21756 8372 21812 8382
rect 21644 8316 21756 8372
rect 20748 8206 20750 8258
rect 20802 8206 20804 8258
rect 20748 8194 20804 8206
rect 21420 8260 21476 8270
rect 20412 8148 20468 8158
rect 20412 8054 20468 8092
rect 21420 8146 21476 8204
rect 21420 8094 21422 8146
rect 21474 8094 21476 8146
rect 21420 8082 21476 8094
rect 21532 8146 21588 8158
rect 21532 8094 21534 8146
rect 21586 8094 21588 8146
rect 20636 8034 20692 8046
rect 21196 8036 21252 8046
rect 20636 7982 20638 8034
rect 20690 7982 20692 8034
rect 20636 7924 20692 7982
rect 20860 8034 21252 8036
rect 20860 7982 21198 8034
rect 21250 7982 21252 8034
rect 20860 7980 21252 7982
rect 20860 7924 20916 7980
rect 21196 7970 21252 7980
rect 21532 8036 21588 8094
rect 21756 8036 21812 8316
rect 21868 8258 21924 8990
rect 21868 8206 21870 8258
rect 21922 8206 21924 8258
rect 21868 8194 21924 8206
rect 21980 9602 22036 9614
rect 21980 9550 21982 9602
rect 22034 9550 22036 9602
rect 21980 9380 22036 9550
rect 21980 8260 22036 9324
rect 22204 9156 22260 11788
rect 22540 11732 22596 11742
rect 22540 11506 22596 11676
rect 22540 11454 22542 11506
rect 22594 11454 22596 11506
rect 22540 11442 22596 11454
rect 22876 11172 22932 11182
rect 22876 10836 22932 11116
rect 22204 9090 22260 9100
rect 22316 10834 22932 10836
rect 22316 10782 22878 10834
rect 22930 10782 22932 10834
rect 22316 10780 22932 10782
rect 22316 9826 22372 10780
rect 22876 10770 22932 10780
rect 22988 10836 23044 10846
rect 22988 9938 23044 10780
rect 22988 9886 22990 9938
rect 23042 9886 23044 9938
rect 22988 9874 23044 9886
rect 22316 9774 22318 9826
rect 22370 9774 22372 9826
rect 22316 8932 22372 9774
rect 23100 9716 23156 15092
rect 23324 12850 23380 12862
rect 23324 12798 23326 12850
rect 23378 12798 23380 12850
rect 23324 12404 23380 12798
rect 23324 12338 23380 12348
rect 23548 10610 23604 10622
rect 23548 10558 23550 10610
rect 23602 10558 23604 10610
rect 23548 10500 23604 10558
rect 23660 10500 23716 10510
rect 23548 10444 23660 10500
rect 23660 10434 23716 10444
rect 22876 9660 23156 9716
rect 22876 9266 22932 9660
rect 22876 9214 22878 9266
rect 22930 9214 22932 9266
rect 22428 9156 22484 9166
rect 22428 9062 22484 9100
rect 22316 8818 22372 8876
rect 22316 8766 22318 8818
rect 22370 8766 22372 8818
rect 22316 8754 22372 8766
rect 22540 8372 22596 8382
rect 22092 8260 22148 8270
rect 21980 8258 22148 8260
rect 21980 8206 22094 8258
rect 22146 8206 22148 8258
rect 21980 8204 22148 8206
rect 22092 8194 22148 8204
rect 22540 8258 22596 8316
rect 22540 8206 22542 8258
rect 22594 8206 22596 8258
rect 22540 8194 22596 8206
rect 22764 8146 22820 8158
rect 22764 8094 22766 8146
rect 22818 8094 22820 8146
rect 21756 7980 22036 8036
rect 21532 7970 21588 7980
rect 20636 7868 20916 7924
rect 21644 7924 21700 7934
rect 21700 7868 21812 7924
rect 21644 7858 21700 7868
rect 20524 7364 20580 7374
rect 20524 7270 20580 7308
rect 21308 7252 21364 7262
rect 20300 6860 20468 6916
rect 20300 6690 20356 6702
rect 20300 6638 20302 6690
rect 20354 6638 20356 6690
rect 20076 6412 20244 6468
rect 19068 5684 19124 5694
rect 19068 5234 19124 5628
rect 19068 5182 19070 5234
rect 19122 5182 19124 5234
rect 19068 5170 19124 5182
rect 19180 5348 19236 5358
rect 18844 5012 18900 5022
rect 18620 4900 18676 4910
rect 18620 4806 18676 4844
rect 18508 3614 18510 3666
rect 18562 3614 18564 3666
rect 18508 3602 18564 3614
rect 18732 3668 18788 3678
rect 18732 3574 18788 3612
rect 18844 2772 18900 4956
rect 19068 4564 19124 4574
rect 19180 4564 19236 5292
rect 19292 5236 19348 5246
rect 19292 5142 19348 5180
rect 19068 4562 19236 4564
rect 19068 4510 19070 4562
rect 19122 4510 19236 4562
rect 19068 4508 19236 4510
rect 19068 4498 19124 4508
rect 18956 4452 19012 4462
rect 18956 4358 19012 4396
rect 19404 4226 19460 6412
rect 19628 6374 19684 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20076 6132 20132 6142
rect 20188 6132 20244 6412
rect 20076 6130 20244 6132
rect 20076 6078 20078 6130
rect 20130 6078 20244 6130
rect 20076 6076 20244 6078
rect 20076 6066 20132 6076
rect 20300 5348 20356 6638
rect 20412 6580 20468 6860
rect 20412 6514 20468 6524
rect 21084 6468 21140 6478
rect 21084 6130 21140 6412
rect 21084 6078 21086 6130
rect 21138 6078 21140 6130
rect 21084 6066 21140 6078
rect 21308 6018 21364 7196
rect 21308 5966 21310 6018
rect 21362 5966 21364 6018
rect 21308 5954 21364 5966
rect 21644 6802 21700 6814
rect 21644 6750 21646 6802
rect 21698 6750 21700 6802
rect 20300 5282 20356 5292
rect 20636 5794 20692 5806
rect 20636 5742 20638 5794
rect 20690 5742 20692 5794
rect 20300 5012 20356 5022
rect 20300 4918 20356 4956
rect 20636 4900 20692 5742
rect 21532 5460 21588 5470
rect 21308 5124 21364 5134
rect 21308 5030 21364 5068
rect 20636 4834 20692 4844
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 21532 4450 21588 5404
rect 21644 5346 21700 6750
rect 21756 6580 21812 7868
rect 21980 6914 22036 7980
rect 22316 8034 22372 8046
rect 22316 7982 22318 8034
rect 22370 7982 22372 8034
rect 22316 7476 22372 7982
rect 22764 8036 22820 8094
rect 22764 7970 22820 7980
rect 22876 8146 22932 9214
rect 23772 9268 23828 17276
rect 24220 15148 24276 20524
rect 24332 20132 24388 21084
rect 24556 20916 24612 20926
rect 24556 20822 24612 20860
rect 24668 20356 24724 21868
rect 24332 19236 24388 20076
rect 24332 19170 24388 19180
rect 24556 20300 24668 20356
rect 24444 19010 24500 19022
rect 24444 18958 24446 19010
rect 24498 18958 24500 19010
rect 24444 18676 24500 18958
rect 24444 18610 24500 18620
rect 24332 18338 24388 18350
rect 24332 18286 24334 18338
rect 24386 18286 24388 18338
rect 24332 18228 24388 18286
rect 24556 18228 24612 20300
rect 24668 20290 24724 20300
rect 24332 18172 24612 18228
rect 24780 18676 24836 18686
rect 24556 17780 24612 17790
rect 24780 17780 24836 18620
rect 24612 17724 24836 17780
rect 24556 17686 24612 17724
rect 24892 16772 24948 22204
rect 25900 21588 25956 22990
rect 27020 22484 27076 23662
rect 27020 22418 27076 22428
rect 26684 22372 26740 22382
rect 26740 22316 26852 22372
rect 26684 22306 26740 22316
rect 26236 21924 26292 21934
rect 26124 21868 26236 21924
rect 26012 21812 26068 21822
rect 26124 21812 26180 21868
rect 26236 21858 26292 21868
rect 26012 21810 26180 21812
rect 26012 21758 26014 21810
rect 26066 21758 26180 21810
rect 26012 21756 26180 21758
rect 26012 21700 26068 21756
rect 26012 21634 26068 21644
rect 25004 21028 25060 21038
rect 25004 20914 25060 20972
rect 25004 20862 25006 20914
rect 25058 20862 25060 20914
rect 25004 20850 25060 20862
rect 25900 20916 25956 21532
rect 26348 21588 26404 21598
rect 26684 21588 26740 21598
rect 26348 21586 26628 21588
rect 26348 21534 26350 21586
rect 26402 21534 26628 21586
rect 26348 21532 26628 21534
rect 26348 21522 26404 21532
rect 25900 20850 25956 20860
rect 26572 20804 26628 21532
rect 26684 21494 26740 21532
rect 26684 20804 26740 20814
rect 26236 20802 26740 20804
rect 26236 20750 26686 20802
rect 26738 20750 26740 20802
rect 26236 20748 26740 20750
rect 26236 20020 26292 20748
rect 26684 20738 26740 20748
rect 26460 20580 26516 20590
rect 26796 20580 26852 22316
rect 27132 21028 27188 26236
rect 27244 24722 27300 24734
rect 27244 24670 27246 24722
rect 27298 24670 27300 24722
rect 27244 24612 27300 24670
rect 27244 24546 27300 24556
rect 27356 24162 27412 26852
rect 28364 26628 28420 55020
rect 28476 55076 28532 55134
rect 28476 55010 28532 55020
rect 29372 55076 29428 55086
rect 28364 26562 28420 26572
rect 28364 24948 28420 24958
rect 27916 24612 27972 24622
rect 27356 24110 27358 24162
rect 27410 24110 27412 24162
rect 27356 24098 27412 24110
rect 27804 24610 27972 24612
rect 27804 24558 27918 24610
rect 27970 24558 27972 24610
rect 27804 24556 27972 24558
rect 27804 24050 27860 24556
rect 27916 24546 27972 24556
rect 27804 23998 27806 24050
rect 27858 23998 27860 24050
rect 27804 23986 27860 23998
rect 27468 23828 27524 23838
rect 27356 23826 27524 23828
rect 27356 23774 27470 23826
rect 27522 23774 27524 23826
rect 27356 23772 27524 23774
rect 27244 23714 27300 23726
rect 27244 23662 27246 23714
rect 27298 23662 27300 23714
rect 27244 23156 27300 23662
rect 27244 23090 27300 23100
rect 27132 20962 27188 20972
rect 26460 20578 26852 20580
rect 26460 20526 26462 20578
rect 26514 20526 26852 20578
rect 26460 20524 26852 20526
rect 26460 20514 26516 20524
rect 26460 20132 26516 20142
rect 26796 20132 26852 20142
rect 26516 20130 26852 20132
rect 26516 20078 26798 20130
rect 26850 20078 26852 20130
rect 26516 20076 26852 20078
rect 26460 20038 26516 20076
rect 26796 20066 26852 20076
rect 26908 20132 26964 20142
rect 26908 20130 27076 20132
rect 26908 20078 26910 20130
rect 26962 20078 27076 20130
rect 26908 20076 27076 20078
rect 26908 20066 26964 20076
rect 26236 19926 26292 19964
rect 26908 19796 26964 19806
rect 26684 19794 26964 19796
rect 26684 19742 26910 19794
rect 26962 19742 26964 19794
rect 26684 19740 26964 19742
rect 25452 19236 25508 19246
rect 25340 19234 25508 19236
rect 25340 19182 25454 19234
rect 25506 19182 25508 19234
rect 25340 19180 25508 19182
rect 25340 19124 25396 19180
rect 25452 19170 25508 19180
rect 25340 18564 25396 19068
rect 26236 19122 26292 19134
rect 26236 19070 26238 19122
rect 26290 19070 26292 19122
rect 26236 18676 26292 19070
rect 26348 18676 26404 18686
rect 26236 18674 26404 18676
rect 26236 18622 26350 18674
rect 26402 18622 26404 18674
rect 26236 18620 26404 18622
rect 26348 18610 26404 18620
rect 26684 18674 26740 19740
rect 26908 19730 26964 19740
rect 27020 19460 27076 20076
rect 27356 19460 27412 23772
rect 27468 23762 27524 23772
rect 27804 23828 27860 23838
rect 27804 23378 27860 23772
rect 27804 23326 27806 23378
rect 27858 23326 27860 23378
rect 27804 23314 27860 23326
rect 28140 23826 28196 23838
rect 28140 23774 28142 23826
rect 28194 23774 28196 23826
rect 27692 23154 27748 23166
rect 27692 23102 27694 23154
rect 27746 23102 27748 23154
rect 27692 22146 27748 23102
rect 27804 23156 27860 23166
rect 27804 22930 27860 23100
rect 27804 22878 27806 22930
rect 27858 22878 27860 22930
rect 27804 22866 27860 22878
rect 28140 22484 28196 23774
rect 28028 22260 28084 22270
rect 28028 22166 28084 22204
rect 28140 22258 28196 22428
rect 28140 22206 28142 22258
rect 28194 22206 28196 22258
rect 27692 22094 27694 22146
rect 27746 22094 27748 22146
rect 27692 22036 27748 22094
rect 27692 21970 27748 21980
rect 27804 22146 27860 22158
rect 27804 22094 27806 22146
rect 27858 22094 27860 22146
rect 27804 21812 27860 22094
rect 27468 21756 27860 21812
rect 27916 22146 27972 22158
rect 27916 22094 27918 22146
rect 27970 22094 27972 22146
rect 27468 21698 27524 21756
rect 27468 21646 27470 21698
rect 27522 21646 27524 21698
rect 27468 21634 27524 21646
rect 27580 21028 27636 21038
rect 27580 20934 27636 20972
rect 27916 20356 27972 22094
rect 28140 22148 28196 22206
rect 28140 22082 28196 22092
rect 28252 23826 28308 23838
rect 28252 23774 28254 23826
rect 28306 23774 28308 23826
rect 27916 20290 27972 20300
rect 27804 20018 27860 20030
rect 27804 19966 27806 20018
rect 27858 19966 27860 20018
rect 27356 19404 27636 19460
rect 27020 19394 27076 19404
rect 26684 18622 26686 18674
rect 26738 18622 26740 18674
rect 26684 18610 26740 18622
rect 25340 17108 25396 18508
rect 26460 18564 26516 18574
rect 26460 18470 26516 18508
rect 26908 18452 26964 18462
rect 26572 18450 26964 18452
rect 26572 18398 26910 18450
rect 26962 18398 26964 18450
rect 26572 18396 26964 18398
rect 25340 17106 25620 17108
rect 25340 17054 25342 17106
rect 25394 17054 25620 17106
rect 25340 17052 25620 17054
rect 25340 17042 25396 17052
rect 24892 16706 24948 16716
rect 24556 16210 24612 16222
rect 24556 16158 24558 16210
rect 24610 16158 24612 16210
rect 24556 15316 24612 16158
rect 24892 16100 24948 16110
rect 24892 16006 24948 16044
rect 25564 16098 25620 17052
rect 26460 16884 26516 16894
rect 25564 16046 25566 16098
rect 25618 16046 25620 16098
rect 25564 16034 25620 16046
rect 26012 16882 26516 16884
rect 26012 16830 26462 16882
rect 26514 16830 26516 16882
rect 26012 16828 26516 16830
rect 25228 15986 25284 15998
rect 25228 15934 25230 15986
rect 25282 15934 25284 15986
rect 25116 15874 25172 15886
rect 25116 15822 25118 15874
rect 25170 15822 25172 15874
rect 25116 15428 25172 15822
rect 25228 15876 25284 15934
rect 26012 15876 26068 16828
rect 26460 16818 26516 16828
rect 26572 16770 26628 18396
rect 26908 18386 26964 18396
rect 27356 18338 27412 18350
rect 27356 18286 27358 18338
rect 27410 18286 27412 18338
rect 27356 17892 27412 18286
rect 27356 17826 27412 17836
rect 26572 16718 26574 16770
rect 26626 16718 26628 16770
rect 26572 16706 26628 16718
rect 26684 16882 26740 16894
rect 26684 16830 26686 16882
rect 26738 16830 26740 16882
rect 25228 15820 26068 15876
rect 25788 15540 25844 15550
rect 25228 15428 25284 15438
rect 25116 15372 25228 15428
rect 25228 15334 25284 15372
rect 24556 15250 24612 15260
rect 25340 15316 25396 15326
rect 25340 15222 25396 15260
rect 25788 15314 25844 15484
rect 26012 15538 26068 15820
rect 26348 15986 26404 15998
rect 26348 15934 26350 15986
rect 26402 15934 26404 15986
rect 26012 15486 26014 15538
rect 26066 15486 26068 15538
rect 26012 15474 26068 15486
rect 26124 15540 26180 15550
rect 26124 15426 26180 15484
rect 26124 15374 26126 15426
rect 26178 15374 26180 15426
rect 26124 15362 26180 15374
rect 25788 15262 25790 15314
rect 25842 15262 25844 15314
rect 24668 15202 24724 15214
rect 24668 15150 24670 15202
rect 24722 15150 24724 15202
rect 24668 15148 24724 15150
rect 24220 15092 24612 15148
rect 24668 15092 24948 15148
rect 24556 13972 24612 15092
rect 24108 13970 24612 13972
rect 24108 13918 24558 13970
rect 24610 13918 24612 13970
rect 24108 13916 24612 13918
rect 23996 12404 24052 12414
rect 23996 12310 24052 12348
rect 24108 12402 24164 13916
rect 24556 13906 24612 13916
rect 24668 13634 24724 13646
rect 24668 13582 24670 13634
rect 24722 13582 24724 13634
rect 24108 12350 24110 12402
rect 24162 12350 24164 12402
rect 24108 12338 24164 12350
rect 24220 13300 24276 13310
rect 23884 12178 23940 12190
rect 24220 12180 24276 13244
rect 24668 13076 24724 13582
rect 24668 13010 24724 13020
rect 24780 12404 24836 12414
rect 23884 12126 23886 12178
rect 23938 12126 23940 12178
rect 23884 11844 23940 12126
rect 23884 11778 23940 11788
rect 23996 12124 24276 12180
rect 24556 12180 24612 12190
rect 23884 10836 23940 10846
rect 23884 10742 23940 10780
rect 23772 9202 23828 9212
rect 23996 9154 24052 12124
rect 24556 12086 24612 12124
rect 24668 11844 24724 11854
rect 24332 11396 24388 11406
rect 24332 11172 24388 11340
rect 24444 11172 24500 11182
rect 24332 11170 24500 11172
rect 24332 11118 24446 11170
rect 24498 11118 24500 11170
rect 24332 11116 24500 11118
rect 24108 10612 24164 10622
rect 24332 10612 24388 11116
rect 24444 11106 24500 11116
rect 24668 10722 24724 11788
rect 24780 11394 24836 12348
rect 24892 11732 24948 15092
rect 25228 14306 25284 14318
rect 25228 14254 25230 14306
rect 25282 14254 25284 14306
rect 25228 14196 25284 14254
rect 25228 14130 25284 14140
rect 25676 14308 25732 14318
rect 24892 11666 24948 11676
rect 25004 14084 25060 14094
rect 25004 12740 25060 14028
rect 25676 13970 25732 14252
rect 25788 14196 25844 15262
rect 26348 15148 26404 15934
rect 26684 15316 26740 16830
rect 27132 16882 27188 16894
rect 27132 16830 27134 16882
rect 27186 16830 27188 16882
rect 27132 16660 27188 16830
rect 27132 16594 27188 16604
rect 27580 15538 27636 19404
rect 27804 19124 27860 19966
rect 27804 19058 27860 19068
rect 27580 15486 27582 15538
rect 27634 15486 27636 15538
rect 27580 15474 27636 15486
rect 27804 17444 27860 17454
rect 26684 15250 26740 15260
rect 27468 15314 27524 15326
rect 27468 15262 27470 15314
rect 27522 15262 27524 15314
rect 26348 15092 26628 15148
rect 25788 14130 25844 14140
rect 25676 13918 25678 13970
rect 25730 13918 25732 13970
rect 25676 13906 25732 13918
rect 26124 13300 26180 13310
rect 24780 11342 24782 11394
rect 24834 11342 24836 11394
rect 24780 11330 24836 11342
rect 25004 10836 25060 12684
rect 25452 13076 25508 13086
rect 25228 12178 25284 12190
rect 25228 12126 25230 12178
rect 25282 12126 25284 12178
rect 25228 11956 25284 12126
rect 25340 12180 25396 12190
rect 25340 12086 25396 12124
rect 25452 12068 25508 13020
rect 26124 13074 26180 13244
rect 26124 13022 26126 13074
rect 26178 13022 26180 13074
rect 26124 13010 26180 13022
rect 26572 13074 26628 15092
rect 26684 14308 26740 14318
rect 26684 13746 26740 14252
rect 26684 13694 26686 13746
rect 26738 13694 26740 13746
rect 26684 13682 26740 13694
rect 27356 13636 27412 13646
rect 27356 13542 27412 13580
rect 27356 13412 27412 13422
rect 26572 13022 26574 13074
rect 26626 13022 26628 13074
rect 26572 13010 26628 13022
rect 26684 13300 26740 13310
rect 26684 12962 26740 13244
rect 27020 13188 27076 13198
rect 27020 13186 27300 13188
rect 27020 13134 27022 13186
rect 27074 13134 27300 13186
rect 27020 13132 27300 13134
rect 27020 13122 27076 13132
rect 26684 12910 26686 12962
rect 26738 12910 26740 12962
rect 26684 12898 26740 12910
rect 27132 12962 27188 12974
rect 27132 12910 27134 12962
rect 27186 12910 27188 12962
rect 26460 12850 26516 12862
rect 26460 12798 26462 12850
rect 26514 12798 26516 12850
rect 25788 12404 25844 12414
rect 25564 12292 25620 12302
rect 25564 12180 25620 12236
rect 25788 12290 25844 12348
rect 25788 12238 25790 12290
rect 25842 12238 25844 12290
rect 25788 12226 25844 12238
rect 26236 12292 26292 12302
rect 26236 12198 26292 12236
rect 25564 12178 25732 12180
rect 25564 12126 25566 12178
rect 25618 12126 25732 12178
rect 25564 12124 25732 12126
rect 25564 12114 25620 12124
rect 25452 12002 25508 12012
rect 25228 11890 25284 11900
rect 25340 11172 25396 11182
rect 25396 11116 25508 11172
rect 25340 11078 25396 11116
rect 24668 10670 24670 10722
rect 24722 10670 24724 10722
rect 24668 10658 24724 10670
rect 24780 10780 25060 10836
rect 24108 10610 24388 10612
rect 24108 10558 24110 10610
rect 24162 10558 24388 10610
rect 24108 10556 24388 10558
rect 24444 10610 24500 10622
rect 24444 10558 24446 10610
rect 24498 10558 24500 10610
rect 24108 10546 24164 10556
rect 24444 10500 24500 10558
rect 24780 10500 24836 10780
rect 24500 10444 24836 10500
rect 25340 10722 25396 10734
rect 25340 10670 25342 10722
rect 25394 10670 25396 10722
rect 24444 10406 24500 10444
rect 24220 10388 24276 10398
rect 24220 10294 24276 10332
rect 25228 10388 25284 10398
rect 25228 10294 25284 10332
rect 25116 9940 25172 9950
rect 25340 9940 25396 10670
rect 25172 9884 25396 9940
rect 25116 9846 25172 9884
rect 25452 9826 25508 11116
rect 25564 10388 25620 10398
rect 25564 10294 25620 10332
rect 25452 9774 25454 9826
rect 25506 9774 25508 9826
rect 25452 9762 25508 9774
rect 25676 9604 25732 12124
rect 26460 11844 26516 12798
rect 27132 12740 27188 12910
rect 27132 12674 27188 12684
rect 27244 12402 27300 13132
rect 27244 12350 27246 12402
rect 27298 12350 27300 12402
rect 27244 12338 27300 12350
rect 27356 12402 27412 13356
rect 27356 12350 27358 12402
rect 27410 12350 27412 12402
rect 27356 12338 27412 12350
rect 26460 11778 26516 11788
rect 26796 11956 26852 11966
rect 23996 9102 23998 9154
rect 24050 9102 24052 9154
rect 23996 9090 24052 9102
rect 25452 9548 25732 9604
rect 26012 11170 26068 11182
rect 26012 11118 26014 11170
rect 26066 11118 26068 11170
rect 22876 8094 22878 8146
rect 22930 8094 22932 8146
rect 22876 7812 22932 8094
rect 23212 8988 23492 9044
rect 22316 7410 22372 7420
rect 22652 7756 22932 7812
rect 23100 8034 23156 8046
rect 23100 7982 23102 8034
rect 23154 7982 23156 8034
rect 22652 7362 22708 7756
rect 23100 7698 23156 7982
rect 23100 7646 23102 7698
rect 23154 7646 23156 7698
rect 23100 7634 23156 7646
rect 23212 7700 23268 8988
rect 23436 8930 23492 8988
rect 23660 8932 23716 8942
rect 23436 8878 23438 8930
rect 23490 8878 23492 8930
rect 23436 8866 23492 8878
rect 23548 8930 23716 8932
rect 23548 8878 23662 8930
rect 23714 8878 23716 8930
rect 23548 8876 23716 8878
rect 23324 8818 23380 8830
rect 23324 8766 23326 8818
rect 23378 8766 23380 8818
rect 23324 8372 23380 8766
rect 23436 8372 23492 8382
rect 23324 8370 23492 8372
rect 23324 8318 23438 8370
rect 23490 8318 23492 8370
rect 23324 8316 23492 8318
rect 23436 8260 23492 8316
rect 23212 7644 23380 7700
rect 22652 7310 22654 7362
rect 22706 7310 22708 7362
rect 22652 7298 22708 7310
rect 22876 7474 22932 7486
rect 22876 7422 22878 7474
rect 22930 7422 22932 7474
rect 22876 7364 22932 7422
rect 23212 7476 23268 7486
rect 23212 7382 23268 7420
rect 22876 7298 22932 7308
rect 21980 6862 21982 6914
rect 22034 6862 22036 6914
rect 21980 6850 22036 6862
rect 22540 7140 22596 7150
rect 21756 6486 21812 6524
rect 22316 6802 22372 6814
rect 22316 6750 22318 6802
rect 22370 6750 22372 6802
rect 21868 5908 21924 5918
rect 21868 5814 21924 5852
rect 22316 5460 22372 6750
rect 22316 5394 22372 5404
rect 22540 6692 22596 7084
rect 22764 7028 22820 7038
rect 21644 5294 21646 5346
rect 21698 5294 21700 5346
rect 21644 5282 21700 5294
rect 21868 5348 21924 5358
rect 21756 5236 21812 5246
rect 21756 4898 21812 5180
rect 21868 5122 21924 5292
rect 21868 5070 21870 5122
rect 21922 5070 21924 5122
rect 21868 5058 21924 5070
rect 21756 4846 21758 4898
rect 21810 4846 21812 4898
rect 21756 4834 21812 4846
rect 22092 5010 22148 5022
rect 22092 4958 22094 5010
rect 22146 4958 22148 5010
rect 21532 4398 21534 4450
rect 21586 4398 21588 4450
rect 21532 4386 21588 4398
rect 22092 4340 22148 4958
rect 22540 4898 22596 6636
rect 22652 6804 22708 6814
rect 22652 5906 22708 6748
rect 22652 5854 22654 5906
rect 22706 5854 22708 5906
rect 22652 5842 22708 5854
rect 22764 5124 22820 6972
rect 22876 6580 22932 6590
rect 22876 6130 22932 6524
rect 23324 6132 23380 7644
rect 23436 7028 23492 8204
rect 23436 6962 23492 6972
rect 23548 6804 23604 8876
rect 23660 8866 23716 8876
rect 24444 8932 24500 8942
rect 23884 8260 23940 8270
rect 23884 8166 23940 8204
rect 24332 8034 24388 8046
rect 24332 7982 24334 8034
rect 24386 7982 24388 8034
rect 24332 7924 24388 7982
rect 24332 7858 24388 7868
rect 23996 7588 24052 7598
rect 24332 7588 24388 7598
rect 23996 7586 24388 7588
rect 23996 7534 23998 7586
rect 24050 7534 24334 7586
rect 24386 7534 24388 7586
rect 23996 7532 24388 7534
rect 23996 7522 24052 7532
rect 24332 7522 24388 7532
rect 22876 6078 22878 6130
rect 22930 6078 22932 6130
rect 22876 6066 22932 6078
rect 22988 6076 23324 6132
rect 22876 5124 22932 5134
rect 22540 4846 22542 4898
rect 22594 4846 22596 4898
rect 22540 4834 22596 4846
rect 22652 5122 22932 5124
rect 22652 5070 22878 5122
rect 22930 5070 22932 5122
rect 22652 5068 22932 5070
rect 22092 4274 22148 4284
rect 22316 4340 22372 4350
rect 22652 4340 22708 5068
rect 22876 5058 22932 5068
rect 22316 4338 22708 4340
rect 22316 4286 22318 4338
rect 22370 4286 22708 4338
rect 22316 4284 22708 4286
rect 22876 4452 22932 4462
rect 22876 4338 22932 4396
rect 22876 4286 22878 4338
rect 22930 4286 22932 4338
rect 22316 4274 22372 4284
rect 22876 4274 22932 4286
rect 19404 4174 19406 4226
rect 19458 4174 19460 4226
rect 19404 4162 19460 4174
rect 20188 3668 20244 3678
rect 19740 3444 19796 3482
rect 19740 3378 19796 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 2996 20244 3612
rect 20972 3668 21028 3678
rect 20972 3574 21028 3612
rect 18620 2716 18900 2772
rect 19964 2940 20244 2996
rect 21308 3444 21364 3454
rect 22988 3388 23044 6076
rect 23324 6038 23380 6076
rect 23436 6748 23604 6804
rect 23884 7474 23940 7486
rect 23884 7422 23886 7474
rect 23938 7422 23940 7474
rect 23436 6580 23492 6748
rect 23212 5908 23268 5918
rect 23212 5794 23268 5852
rect 23212 5742 23214 5794
rect 23266 5742 23268 5794
rect 23212 5730 23268 5742
rect 23212 5012 23268 5022
rect 23436 5012 23492 6524
rect 23548 6578 23604 6590
rect 23548 6526 23550 6578
rect 23602 6526 23604 6578
rect 23548 5236 23604 6526
rect 23548 5170 23604 5180
rect 23660 6580 23716 6590
rect 23660 5234 23716 6524
rect 23660 5182 23662 5234
rect 23714 5182 23716 5234
rect 23660 5170 23716 5182
rect 23268 4956 23380 5012
rect 23436 4956 23716 5012
rect 23212 4946 23268 4956
rect 23324 4564 23380 4956
rect 18620 800 18676 2716
rect 19964 800 20020 2940
rect 21308 800 21364 3388
rect 22652 3332 23044 3388
rect 23100 4450 23156 4462
rect 23100 4398 23102 4450
rect 23154 4398 23156 4450
rect 22652 800 22708 3332
rect 23100 2996 23156 4398
rect 23324 4452 23380 4508
rect 23436 4452 23492 4462
rect 23324 4450 23492 4452
rect 23324 4398 23438 4450
rect 23490 4398 23492 4450
rect 23324 4396 23492 4398
rect 23436 4386 23492 4396
rect 23660 4450 23716 4956
rect 23884 4562 23940 7422
rect 24444 7364 24500 8876
rect 24668 8932 24724 8942
rect 24668 8930 24948 8932
rect 24668 8878 24670 8930
rect 24722 8878 24948 8930
rect 24668 8876 24948 8878
rect 24668 8866 24724 8876
rect 24668 8036 24724 8046
rect 24556 7700 24612 7710
rect 24556 7606 24612 7644
rect 24668 7588 24724 7980
rect 24668 7494 24724 7532
rect 24780 8034 24836 8046
rect 24780 7982 24782 8034
rect 24834 7982 24836 8034
rect 24220 7308 24500 7364
rect 24556 7364 24612 7374
rect 23996 7250 24052 7262
rect 23996 7198 23998 7250
rect 24050 7198 24052 7250
rect 23996 6580 24052 7198
rect 23996 6514 24052 6524
rect 24220 6356 24276 7308
rect 24332 7028 24388 7038
rect 24332 6690 24388 6972
rect 24332 6638 24334 6690
rect 24386 6638 24388 6690
rect 24332 6626 24388 6638
rect 24556 6356 24612 7308
rect 24780 7252 24836 7982
rect 24780 7186 24836 7196
rect 24780 6468 24836 6478
rect 24892 6468 24948 8876
rect 25228 8596 25284 8606
rect 25452 8596 25508 9548
rect 26012 9156 26068 11118
rect 26124 10836 26180 10846
rect 26124 10498 26180 10780
rect 26572 10612 26628 10622
rect 26572 10518 26628 10556
rect 26124 10446 26126 10498
rect 26178 10446 26180 10498
rect 26124 9604 26180 10446
rect 26236 10500 26292 10510
rect 26236 9938 26292 10444
rect 26236 9886 26238 9938
rect 26290 9886 26292 9938
rect 26236 9874 26292 9886
rect 26796 10388 26852 11900
rect 27132 11956 27188 11966
rect 27132 11862 27188 11900
rect 26908 11844 26964 11854
rect 26908 10724 26964 11788
rect 27244 10836 27300 10846
rect 26908 10722 27188 10724
rect 26908 10670 26910 10722
rect 26962 10670 27188 10722
rect 26908 10668 27188 10670
rect 26908 10658 26964 10668
rect 27020 10500 27076 10510
rect 27020 10406 27076 10444
rect 26124 9268 26180 9548
rect 26124 9212 26404 9268
rect 25676 9100 26068 9156
rect 25564 8930 25620 8942
rect 25564 8878 25566 8930
rect 25618 8878 25620 8930
rect 25564 8818 25620 8878
rect 25564 8766 25566 8818
rect 25618 8766 25620 8818
rect 25564 8754 25620 8766
rect 25284 8540 25508 8596
rect 25228 8484 25284 8540
rect 25116 8428 25284 8484
rect 25004 8034 25060 8046
rect 25004 7982 25006 8034
rect 25058 7982 25060 8034
rect 25004 6804 25060 7982
rect 25116 7924 25172 8428
rect 25228 8316 25508 8372
rect 25228 8146 25284 8316
rect 25452 8260 25508 8316
rect 25564 8260 25620 8270
rect 25452 8258 25620 8260
rect 25452 8206 25566 8258
rect 25618 8206 25620 8258
rect 25452 8204 25620 8206
rect 25564 8194 25620 8204
rect 25228 8094 25230 8146
rect 25282 8094 25284 8146
rect 25228 8082 25284 8094
rect 25340 8146 25396 8158
rect 25340 8094 25342 8146
rect 25394 8094 25396 8146
rect 25116 7868 25284 7924
rect 25116 6804 25172 6814
rect 25004 6802 25172 6804
rect 25004 6750 25118 6802
rect 25170 6750 25172 6802
rect 25004 6748 25172 6750
rect 25116 6738 25172 6748
rect 24836 6412 24948 6468
rect 24780 6402 24836 6412
rect 23884 4510 23886 4562
rect 23938 4510 23940 4562
rect 23884 4498 23940 4510
rect 23996 6300 24276 6356
rect 24332 6300 24612 6356
rect 23660 4398 23662 4450
rect 23714 4398 23716 4450
rect 23660 4386 23716 4398
rect 23772 3892 23828 3902
rect 23324 3556 23380 3566
rect 23324 3554 23604 3556
rect 23324 3502 23326 3554
rect 23378 3502 23604 3554
rect 23324 3500 23604 3502
rect 23324 3490 23380 3500
rect 23548 3108 23604 3500
rect 23772 3554 23828 3836
rect 23772 3502 23774 3554
rect 23826 3502 23828 3554
rect 23772 3490 23828 3502
rect 23996 3442 24052 6300
rect 24108 4340 24164 4350
rect 24108 4246 24164 4284
rect 23996 3390 23998 3442
rect 24050 3390 24052 3442
rect 23996 3378 24052 3390
rect 24332 3388 24388 6300
rect 24556 6020 24612 6030
rect 25116 6020 25172 6030
rect 24556 6018 25172 6020
rect 24556 5966 24558 6018
rect 24610 5966 25118 6018
rect 25170 5966 25172 6018
rect 24556 5964 25172 5966
rect 24556 5954 24612 5964
rect 25116 5954 25172 5964
rect 25228 5684 25284 7868
rect 25228 5618 25284 5628
rect 25340 4562 25396 8094
rect 25564 7812 25620 7822
rect 25452 7362 25508 7374
rect 25452 7310 25454 7362
rect 25506 7310 25508 7362
rect 25452 7252 25508 7310
rect 25452 7186 25508 7196
rect 25564 4564 25620 7756
rect 25676 7476 25732 9100
rect 26124 8930 26180 8942
rect 26124 8878 26126 8930
rect 26178 8878 26180 8930
rect 26012 8708 26068 8718
rect 25788 8260 25844 8270
rect 25788 8146 25844 8204
rect 25788 8094 25790 8146
rect 25842 8094 25844 8146
rect 25788 8082 25844 8094
rect 25900 8146 25956 8158
rect 25900 8094 25902 8146
rect 25954 8094 25956 8146
rect 25676 7410 25732 7420
rect 25788 7700 25844 7710
rect 25788 5234 25844 7644
rect 25900 7588 25956 8094
rect 26012 7698 26068 8652
rect 26012 7646 26014 7698
rect 26066 7646 26068 7698
rect 26012 7634 26068 7646
rect 25900 6580 25956 7532
rect 25900 6514 25956 6524
rect 25788 5182 25790 5234
rect 25842 5182 25844 5234
rect 25788 5170 25844 5182
rect 25900 5684 25956 5694
rect 25340 4510 25342 4562
rect 25394 4510 25396 4562
rect 25340 4498 25396 4510
rect 25452 4508 25620 4564
rect 25676 5012 25732 5022
rect 25676 4564 25732 4956
rect 24668 4450 24724 4462
rect 24668 4398 24670 4450
rect 24722 4398 24724 4450
rect 24444 4340 24500 4350
rect 24444 4246 24500 4284
rect 24668 4004 24724 4398
rect 25228 4340 25284 4350
rect 25452 4340 25508 4508
rect 25228 4338 25508 4340
rect 25228 4286 25230 4338
rect 25282 4286 25508 4338
rect 25228 4284 25508 4286
rect 25564 4338 25620 4350
rect 25564 4286 25566 4338
rect 25618 4286 25620 4338
rect 25228 4228 25284 4284
rect 25228 4162 25284 4172
rect 25564 4116 25620 4286
rect 25676 4338 25732 4508
rect 25676 4286 25678 4338
rect 25730 4286 25732 4338
rect 25676 4274 25732 4286
rect 25900 4116 25956 5628
rect 26124 4564 26180 8878
rect 26236 8034 26292 8046
rect 26236 7982 26238 8034
rect 26290 7982 26292 8034
rect 26236 7812 26292 7982
rect 26236 7746 26292 7756
rect 26236 7362 26292 7374
rect 26236 7310 26238 7362
rect 26290 7310 26292 7362
rect 26236 6804 26292 7310
rect 26236 6738 26292 6748
rect 26348 6580 26404 9212
rect 26796 9266 26852 10332
rect 27132 9828 27188 10668
rect 27244 10610 27300 10780
rect 27468 10612 27524 15262
rect 27692 15314 27748 15326
rect 27692 15262 27694 15314
rect 27746 15262 27748 15314
rect 27692 12180 27748 15262
rect 27692 12114 27748 12124
rect 27580 11956 27636 11966
rect 27580 11618 27636 11900
rect 27580 11566 27582 11618
rect 27634 11566 27636 11618
rect 27580 11554 27636 11566
rect 27692 11844 27748 11854
rect 27692 11396 27748 11788
rect 27244 10558 27246 10610
rect 27298 10558 27300 10610
rect 27244 10546 27300 10558
rect 27356 10556 27524 10612
rect 27580 11340 27748 11396
rect 27580 10610 27636 11340
rect 27580 10558 27582 10610
rect 27634 10558 27636 10610
rect 27356 10052 27412 10556
rect 27580 10546 27636 10558
rect 27692 11170 27748 11182
rect 27692 11118 27694 11170
rect 27746 11118 27748 11170
rect 27468 10388 27524 10398
rect 27692 10388 27748 11118
rect 27468 10386 27748 10388
rect 27468 10334 27470 10386
rect 27522 10334 27748 10386
rect 27468 10332 27748 10334
rect 27804 11170 27860 17388
rect 28252 17106 28308 23774
rect 28364 23826 28420 24892
rect 28364 23774 28366 23826
rect 28418 23774 28420 23826
rect 28364 23762 28420 23774
rect 28588 23716 28644 23726
rect 28588 23714 28756 23716
rect 28588 23662 28590 23714
rect 28642 23662 28756 23714
rect 28588 23660 28756 23662
rect 28588 23650 28644 23660
rect 28588 20804 28644 20814
rect 28588 20710 28644 20748
rect 28588 19908 28644 19918
rect 28588 19814 28644 19852
rect 28476 19460 28532 19470
rect 28476 19346 28532 19404
rect 28476 19294 28478 19346
rect 28530 19294 28532 19346
rect 28476 19282 28532 19294
rect 28700 18452 28756 23660
rect 29372 22596 29428 55020
rect 43708 55076 43764 55412
rect 50092 55410 50148 56028
rect 51548 56084 51604 56094
rect 51548 55990 51604 56028
rect 50092 55358 50094 55410
rect 50146 55358 50148 55410
rect 50092 55346 50148 55358
rect 55132 55410 55188 56252
rect 55356 56242 55412 56252
rect 55916 55970 55972 55982
rect 55916 55918 55918 55970
rect 55970 55918 55972 55970
rect 55916 55468 55972 55918
rect 58940 55972 58996 59200
rect 62748 56308 62804 59200
rect 62748 56242 62804 56252
rect 63980 56308 64036 56318
rect 63980 56214 64036 56252
rect 66556 56308 66612 59200
rect 66780 56308 66836 56318
rect 66556 56306 66836 56308
rect 66556 56254 66782 56306
rect 66834 56254 66836 56306
rect 66556 56252 66836 56254
rect 61292 56084 61348 56094
rect 59388 55972 59444 55982
rect 58940 55970 59444 55972
rect 58940 55918 59390 55970
rect 59442 55918 59444 55970
rect 58940 55916 59444 55918
rect 59388 55906 59444 55916
rect 55916 55412 56084 55468
rect 55132 55358 55134 55410
rect 55186 55358 55188 55410
rect 55132 55346 55188 55358
rect 49980 55186 50036 55198
rect 49980 55134 49982 55186
rect 50034 55134 50036 55186
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 37884 30884 37940 30894
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 32844 30324 32900 30334
rect 32620 28754 32676 28766
rect 32620 28702 32622 28754
rect 32674 28702 32676 28754
rect 29820 28642 29876 28654
rect 29820 28590 29822 28642
rect 29874 28590 29876 28642
rect 29708 27746 29764 27758
rect 29708 27694 29710 27746
rect 29762 27694 29764 27746
rect 29708 27636 29764 27694
rect 29820 27748 29876 28590
rect 30492 28532 30548 28542
rect 29820 27682 29876 27692
rect 29932 28530 30548 28532
rect 29932 28478 30494 28530
rect 30546 28478 30548 28530
rect 29932 28476 30548 28478
rect 29708 27570 29764 27580
rect 29372 22530 29428 22540
rect 29372 22372 29428 22382
rect 29372 22278 29428 22316
rect 29036 22260 29092 22270
rect 29036 22166 29092 22204
rect 29148 22148 29204 22158
rect 29148 20690 29204 22092
rect 29260 22148 29316 22158
rect 29820 22148 29876 22158
rect 29260 22146 29876 22148
rect 29260 22094 29262 22146
rect 29314 22094 29822 22146
rect 29874 22094 29876 22146
rect 29260 22092 29876 22094
rect 29260 22082 29316 22092
rect 29596 21474 29652 22092
rect 29820 21812 29876 22092
rect 29820 21746 29876 21756
rect 29596 21422 29598 21474
rect 29650 21422 29652 21474
rect 29596 21410 29652 21422
rect 29372 20804 29428 20814
rect 29148 20638 29150 20690
rect 29202 20638 29204 20690
rect 29148 20626 29204 20638
rect 29260 20748 29372 20804
rect 29148 20356 29204 20366
rect 28700 17668 28756 18396
rect 28700 17602 28756 17612
rect 28812 19124 28868 19134
rect 28812 18450 28868 19068
rect 28812 18398 28814 18450
rect 28866 18398 28868 18450
rect 28252 17054 28254 17106
rect 28306 17054 28308 17106
rect 28252 17042 28308 17054
rect 28028 16996 28084 17006
rect 28028 16994 28196 16996
rect 28028 16942 28030 16994
rect 28082 16942 28196 16994
rect 28028 16940 28196 16942
rect 28028 16930 28084 16940
rect 27916 16882 27972 16894
rect 27916 16830 27918 16882
rect 27970 16830 27972 16882
rect 27916 16660 27972 16830
rect 27916 15538 27972 16604
rect 27916 15486 27918 15538
rect 27970 15486 27972 15538
rect 27916 15474 27972 15486
rect 28140 11620 28196 16940
rect 28476 16210 28532 16222
rect 28476 16158 28478 16210
rect 28530 16158 28532 16210
rect 28476 15148 28532 16158
rect 28812 16212 28868 18398
rect 28812 15538 28868 16156
rect 28812 15486 28814 15538
rect 28866 15486 28868 15538
rect 28812 15474 28868 15486
rect 28252 15092 28532 15148
rect 28252 13412 28308 15092
rect 28476 15026 28532 15036
rect 29036 15316 29092 15326
rect 29036 13972 29092 15260
rect 29148 14420 29204 20300
rect 29260 19010 29316 20748
rect 29372 20710 29428 20748
rect 29260 18958 29262 19010
rect 29314 18958 29316 19010
rect 29260 18900 29316 18958
rect 29260 18834 29316 18844
rect 29596 18452 29652 18462
rect 29820 18452 29876 18462
rect 29596 17554 29652 18396
rect 29596 17502 29598 17554
rect 29650 17502 29652 17554
rect 29596 17490 29652 17502
rect 29708 18450 29876 18452
rect 29708 18398 29822 18450
rect 29874 18398 29876 18450
rect 29708 18396 29876 18398
rect 29932 18452 29988 28476
rect 30492 28466 30548 28476
rect 32620 28084 32676 28702
rect 32620 28018 32676 28028
rect 30940 27972 30996 27982
rect 30940 27878 30996 27916
rect 31612 27972 31668 27982
rect 30716 27858 30772 27870
rect 30716 27806 30718 27858
rect 30770 27806 30772 27858
rect 30156 27748 30212 27758
rect 30156 27654 30212 27692
rect 30716 27636 30772 27806
rect 30716 27076 30772 27580
rect 31164 27076 31220 27086
rect 30716 27074 31220 27076
rect 30716 27022 31166 27074
rect 31218 27022 31220 27074
rect 30716 27020 31220 27022
rect 31164 27010 31220 27020
rect 31388 27076 31444 27086
rect 30492 26402 30548 26414
rect 30492 26350 30494 26402
rect 30546 26350 30548 26402
rect 30268 26292 30324 26302
rect 30156 26236 30268 26292
rect 30044 24612 30100 24622
rect 30156 24612 30212 26236
rect 30268 26198 30324 26236
rect 30492 26068 30548 26350
rect 30940 26292 30996 26302
rect 30940 26198 30996 26236
rect 31388 26290 31444 27020
rect 31612 26516 31668 27916
rect 31724 27860 31780 27870
rect 31724 27076 31780 27804
rect 31724 26982 31780 27020
rect 31836 26962 31892 26974
rect 31836 26910 31838 26962
rect 31890 26910 31892 26962
rect 31836 26628 31892 26910
rect 31836 26562 31892 26572
rect 31724 26516 31780 26526
rect 31388 26238 31390 26290
rect 31442 26238 31444 26290
rect 31388 26226 31444 26238
rect 31500 26514 31780 26516
rect 31500 26462 31726 26514
rect 31778 26462 31780 26514
rect 31500 26460 31780 26462
rect 30492 26002 30548 26012
rect 30828 26068 30884 26078
rect 31164 26068 31220 26078
rect 31500 26068 31556 26460
rect 31724 26450 31780 26460
rect 32060 26402 32116 26414
rect 32060 26350 32062 26402
rect 32114 26350 32116 26402
rect 30828 26066 31108 26068
rect 30828 26014 30830 26066
rect 30882 26014 31108 26066
rect 30828 26012 31108 26014
rect 30828 26002 30884 26012
rect 31052 25618 31108 26012
rect 31164 26066 31556 26068
rect 31164 26014 31166 26066
rect 31218 26014 31556 26066
rect 31164 26012 31556 26014
rect 31836 26068 31892 26078
rect 31164 26002 31220 26012
rect 31052 25566 31054 25618
rect 31106 25566 31108 25618
rect 31052 25554 31108 25566
rect 31500 25506 31556 25518
rect 31500 25454 31502 25506
rect 31554 25454 31556 25506
rect 31388 24948 31444 24958
rect 31388 24854 31444 24892
rect 31276 24836 31332 24846
rect 31276 24742 31332 24780
rect 30044 24610 30212 24612
rect 30044 24558 30046 24610
rect 30098 24558 30212 24610
rect 30044 24556 30212 24558
rect 30492 24612 30548 24622
rect 31500 24612 31556 25454
rect 31836 24836 31892 26012
rect 31948 25508 32004 25518
rect 31948 25414 32004 25452
rect 31836 24724 31892 24780
rect 31948 24724 32004 24734
rect 31836 24722 32004 24724
rect 31836 24670 31950 24722
rect 32002 24670 32004 24722
rect 31836 24668 32004 24670
rect 31948 24658 32004 24668
rect 31724 24612 31780 24622
rect 31500 24610 31780 24612
rect 31500 24558 31726 24610
rect 31778 24558 31780 24610
rect 31500 24556 31780 24558
rect 30044 24546 30100 24556
rect 30492 23716 30548 24556
rect 30492 23650 30548 23660
rect 31164 23938 31220 23950
rect 31164 23886 31166 23938
rect 31218 23886 31220 23938
rect 31164 23716 31220 23886
rect 31164 23650 31220 23660
rect 31500 22596 31556 22606
rect 30716 21700 30772 21710
rect 30044 21476 30100 21486
rect 30044 21382 30100 21420
rect 30044 20804 30100 20814
rect 30044 20710 30100 20748
rect 30604 20578 30660 20590
rect 30604 20526 30606 20578
rect 30658 20526 30660 20578
rect 30268 20020 30324 20030
rect 30156 19964 30268 20020
rect 30044 18452 30100 18462
rect 29932 18450 30100 18452
rect 29932 18398 30046 18450
rect 30098 18398 30100 18450
rect 29932 18396 30100 18398
rect 29596 15876 29652 15886
rect 29596 15782 29652 15820
rect 29708 15148 29764 18396
rect 29820 18386 29876 18396
rect 30044 18386 30100 18396
rect 29932 17442 29988 17454
rect 29932 17390 29934 17442
rect 29986 17390 29988 17442
rect 29932 16884 29988 17390
rect 30044 17108 30100 17118
rect 30156 17108 30212 19964
rect 30268 19954 30324 19964
rect 30268 19124 30324 19134
rect 30604 19124 30660 20526
rect 30716 19906 30772 21644
rect 31388 21586 31444 21598
rect 31388 21534 31390 21586
rect 31442 21534 31444 21586
rect 31388 20130 31444 21534
rect 31388 20078 31390 20130
rect 31442 20078 31444 20130
rect 31388 20066 31444 20078
rect 30940 20020 30996 20030
rect 30940 19926 30996 19964
rect 30716 19854 30718 19906
rect 30770 19854 30772 19906
rect 30716 19842 30772 19854
rect 31164 19908 31220 19918
rect 31164 19814 31220 19852
rect 30324 19068 30660 19124
rect 30268 19030 30324 19068
rect 31052 19012 31108 19022
rect 30268 18452 30324 18462
rect 30268 18358 30324 18396
rect 30492 18452 30548 18462
rect 30492 18358 30548 18396
rect 31052 17666 31108 18956
rect 31500 18900 31556 22540
rect 31612 21700 31668 24556
rect 31724 24546 31780 24556
rect 32060 24612 32116 26350
rect 32620 24724 32676 24734
rect 32620 24630 32676 24668
rect 32060 24500 32116 24556
rect 32172 24500 32228 24510
rect 32060 24498 32228 24500
rect 32060 24446 32174 24498
rect 32226 24446 32228 24498
rect 32060 24444 32228 24446
rect 31836 23826 31892 23838
rect 31836 23774 31838 23826
rect 31890 23774 31892 23826
rect 31836 22484 31892 23774
rect 32172 23828 32228 24444
rect 32172 23762 32228 23772
rect 31836 22418 31892 22428
rect 32732 22484 32788 22494
rect 32732 22390 32788 22428
rect 32508 22372 32564 22382
rect 31612 21606 31668 21644
rect 32060 22370 32564 22372
rect 32060 22318 32510 22370
rect 32562 22318 32564 22370
rect 32060 22316 32564 22318
rect 31724 21586 31780 21598
rect 31724 21534 31726 21586
rect 31778 21534 31780 21586
rect 31724 20132 31780 21534
rect 31724 20066 31780 20076
rect 31836 20802 31892 20814
rect 31836 20750 31838 20802
rect 31890 20750 31892 20802
rect 31612 20018 31668 20030
rect 31612 19966 31614 20018
rect 31666 19966 31668 20018
rect 31612 19908 31668 19966
rect 31612 19842 31668 19852
rect 31836 19236 31892 20750
rect 31948 20018 32004 20030
rect 31948 19966 31950 20018
rect 32002 19966 32004 20018
rect 31948 19796 32004 19966
rect 31948 19730 32004 19740
rect 31836 19170 31892 19180
rect 32060 19124 32116 22316
rect 32508 22306 32564 22316
rect 32284 21476 32340 21486
rect 32284 21474 32452 21476
rect 32284 21422 32286 21474
rect 32338 21422 32452 21474
rect 32284 21420 32452 21422
rect 32284 21410 32340 21420
rect 32284 20132 32340 20142
rect 32284 20038 32340 20076
rect 32396 19908 32452 21420
rect 32396 19842 32452 19852
rect 31948 19068 32116 19124
rect 32172 19796 32228 19806
rect 31500 18844 31892 18900
rect 31052 17614 31054 17666
rect 31106 17614 31108 17666
rect 31052 17602 31108 17614
rect 31388 18564 31444 18574
rect 31388 17666 31444 18508
rect 31836 18450 31892 18844
rect 31836 18398 31838 18450
rect 31890 18398 31892 18450
rect 31836 18340 31892 18398
rect 31836 18274 31892 18284
rect 31388 17614 31390 17666
rect 31442 17614 31444 17666
rect 31388 17602 31444 17614
rect 30716 17554 30772 17566
rect 30716 17502 30718 17554
rect 30770 17502 30772 17554
rect 30716 17108 30772 17502
rect 30828 17444 30884 17454
rect 30828 17350 30884 17388
rect 31164 17108 31220 17118
rect 30044 17106 30212 17108
rect 30044 17054 30046 17106
rect 30098 17054 30212 17106
rect 30044 17052 30212 17054
rect 30268 17052 30660 17108
rect 30716 17052 30884 17108
rect 30044 17042 30100 17052
rect 30268 16994 30324 17052
rect 30268 16942 30270 16994
rect 30322 16942 30324 16994
rect 30268 16930 30324 16942
rect 29988 16828 30100 16884
rect 29932 16818 29988 16828
rect 29820 16100 29876 16110
rect 29820 16006 29876 16044
rect 30044 16098 30100 16828
rect 30380 16882 30436 16894
rect 30380 16830 30382 16882
rect 30434 16830 30436 16882
rect 30380 16772 30436 16830
rect 30380 16706 30436 16716
rect 30044 16046 30046 16098
rect 30098 16046 30100 16098
rect 30044 16034 30100 16046
rect 30492 16100 30548 16110
rect 30492 16006 30548 16044
rect 30268 15874 30324 15886
rect 30268 15822 30270 15874
rect 30322 15822 30324 15874
rect 30268 15148 30324 15822
rect 30380 15874 30436 15886
rect 30380 15822 30382 15874
rect 30434 15822 30436 15874
rect 30380 15764 30436 15822
rect 30380 15698 30436 15708
rect 29708 15092 30100 15148
rect 30268 15092 30548 15148
rect 29148 14326 29204 14364
rect 29260 14420 29316 14430
rect 29260 14418 29540 14420
rect 29260 14366 29262 14418
rect 29314 14366 29540 14418
rect 29260 14364 29540 14366
rect 29260 14354 29316 14364
rect 29484 13972 29540 14364
rect 29708 14308 29764 14318
rect 29708 14214 29764 14252
rect 29036 13916 29428 13972
rect 28252 13346 28308 13356
rect 29372 12962 29428 13916
rect 29484 13916 29876 13972
rect 29484 13634 29540 13916
rect 29484 13582 29486 13634
rect 29538 13582 29540 13634
rect 29484 13570 29540 13582
rect 29708 13746 29764 13758
rect 29708 13694 29710 13746
rect 29762 13694 29764 13746
rect 29708 12964 29764 13694
rect 29372 12910 29374 12962
rect 29426 12910 29428 12962
rect 29372 12898 29428 12910
rect 29484 12908 29764 12964
rect 29820 12962 29876 13916
rect 29820 12910 29822 12962
rect 29874 12910 29876 12962
rect 28140 11554 28196 11564
rect 28364 12740 28420 12750
rect 28364 11844 28420 12684
rect 29148 12404 29204 12414
rect 29148 12290 29204 12348
rect 29484 12402 29540 12908
rect 29820 12898 29876 12910
rect 29932 12852 29988 12862
rect 29932 12758 29988 12796
rect 29596 12738 29652 12750
rect 29596 12686 29598 12738
rect 29650 12686 29652 12738
rect 29596 12628 29652 12686
rect 29708 12740 29764 12750
rect 29708 12738 29876 12740
rect 29708 12686 29710 12738
rect 29762 12686 29876 12738
rect 29708 12684 29876 12686
rect 29708 12674 29764 12684
rect 29596 12562 29652 12572
rect 29484 12350 29486 12402
rect 29538 12350 29540 12402
rect 29484 12338 29540 12350
rect 29148 12238 29150 12290
rect 29202 12238 29204 12290
rect 29148 12226 29204 12238
rect 29708 12292 29764 12302
rect 29708 12198 29764 12236
rect 28812 12180 28868 12190
rect 28700 12068 28756 12078
rect 27804 11118 27806 11170
rect 27858 11118 27860 11170
rect 27468 10322 27524 10332
rect 27356 9996 27636 10052
rect 27132 9772 27524 9828
rect 26796 9214 26798 9266
rect 26850 9214 26852 9266
rect 26796 9202 26852 9214
rect 27468 9266 27524 9772
rect 27468 9214 27470 9266
rect 27522 9214 27524 9266
rect 27468 9202 27524 9214
rect 27020 9044 27076 9054
rect 26572 8932 26628 8942
rect 26572 8930 26740 8932
rect 26572 8878 26574 8930
rect 26626 8878 26740 8930
rect 26572 8876 26740 8878
rect 26572 8866 26628 8876
rect 26236 6524 26404 6580
rect 26460 8818 26516 8830
rect 26460 8766 26462 8818
rect 26514 8766 26516 8818
rect 26236 5012 26292 6524
rect 26460 6356 26516 8766
rect 26572 8036 26628 8046
rect 26572 7942 26628 7980
rect 26460 6290 26516 6300
rect 26684 6244 26740 8876
rect 27020 8146 27076 8988
rect 27132 9042 27188 9054
rect 27132 8990 27134 9042
rect 27186 8990 27188 9042
rect 27132 8932 27188 8990
rect 27132 8866 27188 8876
rect 27580 8708 27636 9996
rect 27804 9492 27860 11118
rect 28028 10948 28084 10958
rect 28028 10612 28084 10892
rect 28364 10834 28420 11788
rect 28588 12066 28756 12068
rect 28588 12014 28702 12066
rect 28754 12014 28756 12066
rect 28588 12012 28756 12014
rect 28364 10782 28366 10834
rect 28418 10782 28420 10834
rect 28364 10770 28420 10782
rect 28476 11620 28532 11630
rect 28028 10518 28084 10556
rect 28476 9828 28532 11564
rect 28252 9772 28532 9828
rect 27916 9492 27972 9502
rect 27804 9436 27916 9492
rect 27916 9426 27972 9436
rect 27132 8652 27636 8708
rect 27804 9042 27860 9054
rect 27804 8990 27806 9042
rect 27858 8990 27860 9042
rect 27804 8932 27860 8990
rect 27132 8370 27188 8652
rect 27804 8484 27860 8876
rect 28140 8820 28196 8830
rect 27804 8418 27860 8428
rect 28028 8818 28196 8820
rect 28028 8766 28142 8818
rect 28194 8766 28196 8818
rect 28028 8764 28196 8766
rect 27132 8318 27134 8370
rect 27186 8318 27188 8370
rect 27132 8306 27188 8318
rect 28028 8372 28084 8764
rect 28140 8754 28196 8764
rect 27020 8094 27022 8146
rect 27074 8094 27076 8146
rect 26684 6178 26740 6188
rect 26908 6468 26964 6478
rect 26796 6132 26852 6142
rect 26348 5908 26404 5918
rect 26348 5234 26404 5852
rect 26348 5182 26350 5234
rect 26402 5182 26404 5234
rect 26348 5170 26404 5182
rect 26796 5122 26852 6076
rect 26796 5070 26798 5122
rect 26850 5070 26852 5122
rect 26796 5058 26852 5070
rect 26236 4956 26404 5012
rect 26124 4508 26292 4564
rect 25564 4060 25956 4116
rect 26124 4226 26180 4238
rect 26124 4174 26126 4226
rect 26178 4174 26180 4226
rect 24668 3938 24724 3948
rect 26124 3892 26180 4174
rect 26236 4116 26292 4508
rect 26236 4050 26292 4060
rect 26348 3892 26404 4956
rect 26124 3836 26404 3892
rect 26460 4676 26516 4686
rect 26908 4676 26964 6412
rect 25452 3666 25508 3678
rect 25452 3614 25454 3666
rect 25506 3614 25508 3666
rect 24108 3332 24388 3388
rect 24556 3442 24612 3454
rect 24556 3390 24558 3442
rect 24610 3390 24612 3442
rect 24108 3220 24164 3332
rect 23548 3042 23604 3052
rect 23996 3164 24164 3220
rect 24556 3220 24612 3390
rect 25452 3388 25508 3614
rect 24892 3332 24948 3342
rect 24892 3238 24948 3276
rect 25340 3332 25508 3388
rect 23100 2930 23156 2940
rect 23996 800 24052 3164
rect 24556 3154 24612 3164
rect 25340 800 25396 3332
rect 26460 980 26516 4620
rect 26684 4620 26964 4676
rect 26684 4562 26740 4620
rect 26684 4510 26686 4562
rect 26738 4510 26740 4562
rect 26684 4498 26740 4510
rect 27020 4226 27076 8094
rect 27244 8148 27300 8158
rect 27244 8146 27412 8148
rect 27244 8094 27246 8146
rect 27298 8094 27412 8146
rect 27244 8092 27412 8094
rect 27244 8082 27300 8092
rect 27356 8036 27412 8092
rect 27580 8036 27636 8046
rect 27356 8034 27636 8036
rect 27356 7982 27582 8034
rect 27634 7982 27636 8034
rect 27356 7980 27636 7982
rect 27244 7588 27300 7598
rect 27244 7494 27300 7532
rect 27244 6804 27300 6814
rect 27356 6804 27412 7980
rect 27580 7970 27636 7980
rect 28028 7698 28084 8316
rect 28140 8372 28196 8382
rect 28252 8372 28308 9772
rect 28476 9602 28532 9614
rect 28476 9550 28478 9602
rect 28530 9550 28532 9602
rect 28476 9492 28532 9550
rect 28476 9426 28532 9436
rect 28364 9154 28420 9166
rect 28364 9102 28366 9154
rect 28418 9102 28420 9154
rect 28364 8932 28420 9102
rect 28364 8866 28420 8876
rect 28140 8370 28252 8372
rect 28140 8318 28142 8370
rect 28194 8318 28252 8370
rect 28140 8316 28252 8318
rect 28140 8306 28196 8316
rect 28252 8278 28308 8316
rect 28476 8818 28532 8830
rect 28476 8766 28478 8818
rect 28530 8766 28532 8818
rect 28028 7646 28030 7698
rect 28082 7646 28084 7698
rect 28028 7634 28084 7646
rect 28364 8036 28420 8046
rect 27244 6802 27412 6804
rect 27244 6750 27246 6802
rect 27298 6750 27412 6802
rect 27244 6748 27412 6750
rect 28364 7474 28420 7980
rect 28364 7422 28366 7474
rect 28418 7422 28420 7474
rect 27244 6738 27300 6748
rect 28140 6692 28196 6702
rect 28140 6598 28196 6636
rect 27692 6580 27748 6590
rect 27692 6578 27972 6580
rect 27692 6526 27694 6578
rect 27746 6526 27972 6578
rect 27692 6524 27972 6526
rect 27692 6514 27748 6524
rect 27580 6468 27636 6478
rect 27580 6374 27636 6412
rect 27356 6356 27412 6366
rect 27244 6020 27300 6030
rect 27244 5926 27300 5964
rect 27356 5908 27412 6300
rect 27356 5842 27412 5852
rect 27132 5234 27188 5246
rect 27132 5182 27134 5234
rect 27186 5182 27188 5234
rect 27132 4452 27188 5182
rect 27916 5236 27972 6524
rect 28364 6468 28420 7422
rect 28476 7476 28532 8766
rect 28476 7410 28532 7420
rect 28588 7364 28644 12012
rect 28700 12002 28756 12012
rect 28700 11508 28756 11518
rect 28700 11414 28756 11452
rect 28700 8148 28756 8158
rect 28812 8148 28868 12124
rect 29372 12178 29428 12190
rect 29372 12126 29374 12178
rect 29426 12126 29428 12178
rect 28924 11508 28980 11518
rect 28924 10724 28980 11452
rect 29372 11396 29428 12126
rect 28924 10658 28980 10668
rect 29036 11340 29428 11396
rect 29820 11396 29876 12684
rect 29932 11396 29988 11406
rect 29820 11340 29932 11396
rect 29036 10276 29092 11340
rect 29932 11330 29988 11340
rect 29260 11172 29316 11182
rect 29932 11172 29988 11182
rect 29316 11116 29764 11172
rect 29260 11078 29316 11116
rect 29148 10500 29204 10510
rect 29596 10500 29652 10510
rect 29148 10498 29316 10500
rect 29148 10446 29150 10498
rect 29202 10446 29316 10498
rect 29148 10444 29316 10446
rect 29148 10434 29204 10444
rect 29260 10386 29316 10444
rect 29260 10334 29262 10386
rect 29314 10334 29316 10386
rect 29260 10322 29316 10334
rect 29484 10498 29652 10500
rect 29484 10446 29598 10498
rect 29650 10446 29652 10498
rect 29484 10444 29652 10446
rect 29036 10220 29204 10276
rect 28924 9156 28980 9166
rect 28924 9042 28980 9100
rect 28924 8990 28926 9042
rect 28978 8990 28980 9042
rect 28924 8978 28980 8990
rect 29036 8818 29092 8830
rect 29036 8766 29038 8818
rect 29090 8766 29092 8818
rect 29036 8708 29092 8766
rect 29148 8820 29204 10220
rect 29372 9828 29428 9838
rect 29260 9714 29316 9726
rect 29260 9662 29262 9714
rect 29314 9662 29316 9714
rect 29260 9156 29316 9662
rect 29260 9090 29316 9100
rect 29372 9602 29428 9772
rect 29484 9716 29540 10444
rect 29596 10434 29652 10444
rect 29708 10388 29764 11116
rect 29932 11078 29988 11116
rect 29932 10724 29988 10734
rect 30044 10724 30100 15092
rect 30156 14420 30212 14430
rect 30156 13970 30212 14364
rect 30156 13918 30158 13970
rect 30210 13918 30212 13970
rect 30156 13906 30212 13918
rect 30492 13972 30548 15092
rect 30380 13748 30436 13758
rect 30380 13654 30436 13692
rect 30268 13636 30324 13646
rect 30268 13542 30324 13580
rect 30492 13524 30548 13916
rect 30380 13468 30548 13524
rect 30380 12962 30436 13468
rect 30604 12964 30660 17052
rect 30828 16996 30884 17052
rect 31052 16996 31108 17006
rect 30828 16994 31108 16996
rect 30828 16942 31054 16994
rect 31106 16942 31108 16994
rect 30828 16940 31108 16942
rect 30716 16884 30772 16894
rect 30772 16828 30884 16884
rect 30716 16790 30772 16828
rect 30828 16098 30884 16828
rect 30828 16046 30830 16098
rect 30882 16046 30884 16098
rect 30828 16034 30884 16046
rect 31052 16772 31108 16940
rect 31052 16100 31108 16716
rect 31164 16322 31220 17052
rect 31500 16994 31556 17006
rect 31500 16942 31502 16994
rect 31554 16942 31556 16994
rect 31500 16884 31556 16942
rect 31500 16818 31556 16828
rect 31836 16884 31892 16894
rect 31836 16790 31892 16828
rect 31164 16270 31166 16322
rect 31218 16270 31220 16322
rect 31164 16258 31220 16270
rect 31948 16322 32004 19068
rect 32060 18676 32116 18686
rect 32060 17778 32116 18620
rect 32172 18674 32228 19740
rect 32844 18676 32900 30268
rect 36876 29092 36932 29102
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 33068 28418 33124 28430
rect 33068 28366 33070 28418
rect 33122 28366 33124 28418
rect 33068 23716 33124 28366
rect 33404 28084 33460 28094
rect 33180 27970 33236 27982
rect 33180 27918 33182 27970
rect 33234 27918 33236 27970
rect 33180 27860 33236 27918
rect 33180 27794 33236 27804
rect 33404 27972 33460 28028
rect 33852 27972 33908 27982
rect 33404 27970 33908 27972
rect 33404 27918 33854 27970
rect 33906 27918 33908 27970
rect 33404 27916 33908 27918
rect 33404 27858 33460 27916
rect 33852 27906 33908 27916
rect 34188 27972 34244 27982
rect 33404 27806 33406 27858
rect 33458 27806 33460 27858
rect 33404 27794 33460 27806
rect 34188 27858 34244 27916
rect 34188 27806 34190 27858
rect 34242 27806 34244 27858
rect 34188 27794 34244 27806
rect 35756 27972 35812 27982
rect 34188 27636 34244 27646
rect 34188 27634 34468 27636
rect 34188 27582 34190 27634
rect 34242 27582 34468 27634
rect 34188 27580 34468 27582
rect 34188 27570 34244 27580
rect 34412 27186 34468 27580
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34412 27134 34414 27186
rect 34466 27134 34468 27186
rect 34412 27122 34468 27134
rect 34748 27074 34804 27086
rect 34748 27022 34750 27074
rect 34802 27022 34804 27074
rect 34636 26404 34692 26414
rect 34636 25732 34692 26348
rect 34748 26068 34804 27022
rect 35308 26962 35364 26974
rect 35308 26910 35310 26962
rect 35362 26910 35364 26962
rect 35308 26292 35364 26910
rect 35644 26964 35700 26974
rect 35644 26870 35700 26908
rect 35756 26852 35812 27916
rect 35868 27860 35924 27870
rect 35868 27076 35924 27804
rect 36316 27076 36372 27086
rect 35868 27074 36372 27076
rect 35868 27022 35870 27074
rect 35922 27022 36318 27074
rect 36370 27022 36372 27074
rect 35868 27020 36372 27022
rect 35868 27010 35924 27020
rect 36316 27010 36372 27020
rect 36428 26962 36484 26974
rect 36428 26910 36430 26962
rect 36482 26910 36484 26962
rect 35756 26796 35924 26852
rect 35532 26292 35588 26302
rect 35308 26236 35532 26292
rect 35532 26198 35588 26236
rect 35756 26290 35812 26302
rect 35756 26238 35758 26290
rect 35810 26238 35812 26290
rect 34748 26002 34804 26012
rect 35644 26178 35700 26190
rect 35644 26126 35646 26178
rect 35698 26126 35700 26178
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 25732 35252 25742
rect 34636 25676 35028 25732
rect 34636 25620 34692 25676
rect 34300 25618 34692 25620
rect 34300 25566 34638 25618
rect 34690 25566 34692 25618
rect 34300 25564 34692 25566
rect 33964 25396 34020 25406
rect 33628 25284 33684 25294
rect 33964 25284 34020 25340
rect 34300 25394 34356 25564
rect 34636 25554 34692 25564
rect 34300 25342 34302 25394
rect 34354 25342 34356 25394
rect 34300 25330 34356 25342
rect 34860 25508 34916 25518
rect 33684 25228 34020 25284
rect 33628 25190 33684 25228
rect 34748 24724 34804 24734
rect 34748 24630 34804 24668
rect 33964 24052 34020 24062
rect 33964 24050 34244 24052
rect 33964 23998 33966 24050
rect 34018 23998 34244 24050
rect 33964 23996 34244 23998
rect 33964 23986 34020 23996
rect 33068 23650 33124 23660
rect 33516 23266 33572 23278
rect 33516 23214 33518 23266
rect 33570 23214 33572 23266
rect 33292 23156 33348 23166
rect 32956 23154 33348 23156
rect 32956 23102 33294 23154
rect 33346 23102 33348 23154
rect 32956 23100 33348 23102
rect 32956 22370 33012 23100
rect 33292 23090 33348 23100
rect 33516 23156 33572 23214
rect 34076 23268 34132 23278
rect 34076 23174 34132 23212
rect 33516 23090 33572 23100
rect 33628 23156 33684 23166
rect 33964 23156 34020 23166
rect 33628 23154 34020 23156
rect 33628 23102 33630 23154
rect 33682 23102 33966 23154
rect 34018 23102 34020 23154
rect 33628 23100 34020 23102
rect 33628 23090 33684 23100
rect 32956 22318 32958 22370
rect 33010 22318 33012 22370
rect 32956 22306 33012 22318
rect 33628 22370 33684 22382
rect 33628 22318 33630 22370
rect 33682 22318 33684 22370
rect 33180 22258 33236 22270
rect 33180 22206 33182 22258
rect 33234 22206 33236 22258
rect 33180 21700 33236 22206
rect 33404 21700 33460 21710
rect 33180 21644 33404 21700
rect 33404 21606 33460 21644
rect 33628 21476 33684 22318
rect 33740 22372 33796 23100
rect 33964 23090 34020 23100
rect 34188 23156 34244 23996
rect 34860 23938 34916 25452
rect 34972 24500 35028 25676
rect 35196 25638 35252 25676
rect 35532 25732 35588 25742
rect 35644 25732 35700 26126
rect 35756 26180 35812 26238
rect 35756 26114 35812 26124
rect 35532 25730 35700 25732
rect 35532 25678 35534 25730
rect 35586 25678 35700 25730
rect 35532 25676 35700 25678
rect 35756 25844 35812 25854
rect 35532 25666 35588 25676
rect 35756 25506 35812 25788
rect 35756 25454 35758 25506
rect 35810 25454 35812 25506
rect 35756 25442 35812 25454
rect 35308 24836 35364 24846
rect 35308 24742 35364 24780
rect 35756 24836 35812 24846
rect 35532 24724 35588 24734
rect 35532 24722 35700 24724
rect 35532 24670 35534 24722
rect 35586 24670 35700 24722
rect 35532 24668 35700 24670
rect 35532 24658 35588 24668
rect 35420 24610 35476 24622
rect 35420 24558 35422 24610
rect 35474 24558 35476 24610
rect 35420 24500 35476 24558
rect 34972 24498 35140 24500
rect 34972 24446 34974 24498
rect 35026 24446 35140 24498
rect 34972 24444 35140 24446
rect 35420 24444 35588 24500
rect 34972 24434 35028 24444
rect 34860 23886 34862 23938
rect 34914 23886 34916 23938
rect 34860 23874 34916 23886
rect 34972 24052 35028 24062
rect 34188 23090 34244 23100
rect 34412 23716 34468 23726
rect 34972 23716 35028 23996
rect 35084 23940 35140 24444
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35308 23940 35364 23950
rect 35084 23938 35364 23940
rect 35084 23886 35310 23938
rect 35362 23886 35364 23938
rect 35084 23884 35364 23886
rect 35308 23874 35364 23884
rect 35532 23938 35588 24444
rect 35532 23886 35534 23938
rect 35586 23886 35588 23938
rect 35532 23874 35588 23886
rect 35084 23716 35140 23726
rect 34972 23714 35140 23716
rect 34972 23662 35086 23714
rect 35138 23662 35140 23714
rect 34972 23660 35140 23662
rect 33740 22306 33796 22316
rect 34076 22930 34132 22942
rect 34076 22878 34078 22930
rect 34130 22878 34132 22930
rect 33628 21410 33684 21420
rect 33740 21586 33796 21598
rect 33740 21534 33742 21586
rect 33794 21534 33796 21586
rect 32956 20018 33012 20030
rect 32956 19966 32958 20018
rect 33010 19966 33012 20018
rect 32956 19012 33012 19966
rect 33404 20020 33460 20030
rect 33404 19926 33460 19964
rect 33628 20018 33684 20030
rect 33628 19966 33630 20018
rect 33682 19966 33684 20018
rect 32956 18946 33012 18956
rect 33180 19906 33236 19918
rect 33180 19854 33182 19906
rect 33234 19854 33236 19906
rect 32172 18622 32174 18674
rect 32226 18622 32228 18674
rect 32172 18610 32228 18622
rect 32284 18620 32900 18676
rect 33180 18676 33236 19854
rect 33628 19908 33684 19966
rect 33628 19348 33684 19852
rect 33628 19282 33684 19292
rect 32060 17726 32062 17778
rect 32114 17726 32116 17778
rect 32060 17714 32116 17726
rect 32172 16994 32228 17006
rect 32172 16942 32174 16994
rect 32226 16942 32228 16994
rect 32172 16772 32228 16942
rect 32172 16706 32228 16716
rect 31948 16270 31950 16322
rect 32002 16270 32004 16322
rect 31948 16258 32004 16270
rect 31052 16034 31108 16044
rect 31836 16100 31892 16110
rect 31836 16006 31892 16044
rect 31052 15876 31108 15886
rect 31052 15148 31108 15820
rect 31948 15874 32004 15886
rect 31948 15822 31950 15874
rect 32002 15822 32004 15874
rect 31052 15092 31220 15148
rect 31052 14530 31108 14542
rect 31052 14478 31054 14530
rect 31106 14478 31108 14530
rect 31052 14308 31108 14478
rect 31052 14242 31108 14252
rect 31164 14084 31220 15092
rect 31948 15092 32004 15822
rect 32284 15148 32340 18620
rect 33180 18610 33236 18620
rect 33740 18564 33796 21534
rect 34076 21586 34132 22878
rect 34300 22260 34356 22270
rect 34076 21534 34078 21586
rect 34130 21534 34132 21586
rect 34076 21522 34132 21534
rect 34188 22258 34356 22260
rect 34188 22206 34302 22258
rect 34354 22206 34356 22258
rect 34188 22204 34356 22206
rect 33964 21474 34020 21486
rect 33964 21422 33966 21474
rect 34018 21422 34020 21474
rect 33964 21364 34020 21422
rect 34188 21364 34244 22204
rect 34300 22194 34356 22204
rect 34412 22036 34468 23660
rect 35084 23650 35140 23660
rect 35644 23492 35700 24668
rect 35644 23426 35700 23436
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34300 21980 34468 22036
rect 34300 21476 34356 21980
rect 34412 21756 34916 21812
rect 34412 21700 34468 21756
rect 34412 21606 34468 21644
rect 34636 21588 34692 21598
rect 34412 21476 34468 21486
rect 34300 21420 34412 21476
rect 34412 21410 34468 21420
rect 33964 21308 34244 21364
rect 34076 20130 34132 20142
rect 34076 20078 34078 20130
rect 34130 20078 34132 20130
rect 33852 20020 33908 20030
rect 33852 19926 33908 19964
rect 34076 19796 34132 20078
rect 34188 20132 34244 20142
rect 34188 20038 34244 20076
rect 33628 18508 33796 18564
rect 33852 19236 33908 19246
rect 32508 18450 32564 18462
rect 32508 18398 32510 18450
rect 32562 18398 32564 18450
rect 32508 18228 32564 18398
rect 33180 18228 33236 18238
rect 33516 18228 33572 18238
rect 32508 18226 33236 18228
rect 32508 18174 33182 18226
rect 33234 18174 33236 18226
rect 32508 18172 33236 18174
rect 32620 18004 32676 18014
rect 32396 16884 32452 16894
rect 32396 16790 32452 16828
rect 32620 16322 32676 17948
rect 33180 17668 33236 18172
rect 33180 17602 33236 17612
rect 33404 18172 33516 18228
rect 32620 16270 32622 16322
rect 32674 16270 32676 16322
rect 32620 16258 32676 16270
rect 33404 16324 33460 18172
rect 33516 18134 33572 18172
rect 33628 18004 33684 18508
rect 33628 17938 33684 17948
rect 33740 18340 33796 18350
rect 33740 17780 33796 18284
rect 33404 16230 33460 16268
rect 33628 17724 33796 17780
rect 32508 16100 32564 16110
rect 32508 16006 32564 16044
rect 33628 15988 33684 17724
rect 33852 16994 33908 19180
rect 34076 17780 34132 19740
rect 34300 19236 34356 19246
rect 34300 18674 34356 19180
rect 34300 18622 34302 18674
rect 34354 18622 34356 18674
rect 34300 18610 34356 18622
rect 34636 18676 34692 21532
rect 34860 21474 34916 21756
rect 35644 21588 35700 21598
rect 35756 21588 35812 24780
rect 35868 24722 35924 26796
rect 36204 26292 36260 26302
rect 36204 26290 36372 26292
rect 36204 26238 36206 26290
rect 36258 26238 36372 26290
rect 36204 26236 36372 26238
rect 36204 26226 36260 26236
rect 36316 25732 36372 26236
rect 36428 26180 36484 26910
rect 36540 26404 36596 26414
rect 36540 26310 36596 26348
rect 36652 26180 36708 26190
rect 36428 26124 36596 26180
rect 36316 25638 36372 25676
rect 36092 25506 36148 25518
rect 36540 25508 36596 26124
rect 36652 26086 36708 26124
rect 36764 26068 36820 26078
rect 36764 25974 36820 26012
rect 36092 25454 36094 25506
rect 36146 25454 36148 25506
rect 36092 25284 36148 25454
rect 36092 25218 36148 25228
rect 36204 25452 36596 25508
rect 35868 24670 35870 24722
rect 35922 24670 35924 24722
rect 35868 24658 35924 24670
rect 36092 24724 36148 24734
rect 36204 24724 36260 25452
rect 36428 25284 36484 25294
rect 36876 25284 36932 29036
rect 37436 26292 37492 26302
rect 37436 25730 37492 26236
rect 37772 26180 37828 26190
rect 37436 25678 37438 25730
rect 37490 25678 37492 25730
rect 37436 25666 37492 25678
rect 37548 26068 37604 26078
rect 37548 25730 37604 26012
rect 37548 25678 37550 25730
rect 37602 25678 37604 25730
rect 36428 25282 36932 25284
rect 36428 25230 36430 25282
rect 36482 25230 36932 25282
rect 36428 25228 36932 25230
rect 36988 25284 37044 25294
rect 37436 25284 37492 25294
rect 36428 25218 36484 25228
rect 36988 25172 37044 25228
rect 36764 25116 37044 25172
rect 37324 25282 37492 25284
rect 37324 25230 37438 25282
rect 37490 25230 37492 25282
rect 37324 25228 37492 25230
rect 36764 24946 36820 25116
rect 36764 24894 36766 24946
rect 36818 24894 36820 24946
rect 36764 24882 36820 24894
rect 36092 24722 36204 24724
rect 36092 24670 36094 24722
rect 36146 24670 36204 24722
rect 36092 24668 36204 24670
rect 36092 24658 36148 24668
rect 36204 24630 36260 24668
rect 36988 24836 37044 24846
rect 36988 24612 37044 24780
rect 37100 24724 37156 24734
rect 37324 24724 37380 25228
rect 37436 25218 37492 25228
rect 37436 24948 37492 24958
rect 37548 24948 37604 25678
rect 37772 25730 37828 26124
rect 37772 25678 37774 25730
rect 37826 25678 37828 25730
rect 37772 25666 37828 25678
rect 37436 24946 37604 24948
rect 37436 24894 37438 24946
rect 37490 24894 37604 24946
rect 37436 24892 37604 24894
rect 37436 24882 37492 24892
rect 37156 24668 37268 24724
rect 37324 24668 37604 24724
rect 37100 24658 37156 24668
rect 36316 24500 36372 24510
rect 36988 24500 37044 24556
rect 37100 24500 37156 24510
rect 36988 24498 37156 24500
rect 36988 24446 37102 24498
rect 37154 24446 37156 24498
rect 36988 24444 37156 24446
rect 37212 24500 37268 24668
rect 37324 24500 37380 24510
rect 37212 24498 37380 24500
rect 37212 24446 37326 24498
rect 37378 24446 37380 24498
rect 37212 24444 37380 24446
rect 36316 24406 36372 24444
rect 37100 24434 37156 24444
rect 37324 24434 37380 24444
rect 37436 24500 37492 24510
rect 37436 23604 37492 24444
rect 37548 23940 37604 24668
rect 37548 23874 37604 23884
rect 37436 23538 37492 23548
rect 36428 23268 36484 23278
rect 36428 22484 36484 23212
rect 36428 22390 36484 22428
rect 36988 22820 37044 22830
rect 36988 22482 37044 22764
rect 36988 22430 36990 22482
rect 37042 22430 37044 22482
rect 36988 22418 37044 22430
rect 35700 21532 35812 21588
rect 37212 22260 37268 22270
rect 35644 21522 35700 21532
rect 34860 21422 34862 21474
rect 34914 21422 34916 21474
rect 34748 20690 34804 20702
rect 34748 20638 34750 20690
rect 34802 20638 34804 20690
rect 34748 20020 34804 20638
rect 34860 20356 34916 21422
rect 35532 21476 35588 21486
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34860 20290 34916 20300
rect 35196 20020 35252 20030
rect 35532 20020 35588 21420
rect 36652 21476 36708 21486
rect 36652 21382 36708 21420
rect 36876 20804 36932 20814
rect 36764 20802 36932 20804
rect 36764 20750 36878 20802
rect 36930 20750 36932 20802
rect 36764 20748 36932 20750
rect 34748 20018 35588 20020
rect 34748 19966 34750 20018
rect 34802 19966 35198 20018
rect 35250 19966 35588 20018
rect 34748 19964 35588 19966
rect 34748 19954 34804 19964
rect 35196 19954 35252 19964
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34860 18676 34916 18686
rect 34636 18674 34916 18676
rect 34636 18622 34862 18674
rect 34914 18622 34916 18674
rect 34636 18620 34916 18622
rect 34860 18610 34916 18620
rect 35532 18564 35588 19964
rect 36092 20020 36148 20030
rect 35868 19908 35924 19918
rect 35868 19814 35924 19852
rect 34636 18450 34692 18462
rect 34636 18398 34638 18450
rect 34690 18398 34692 18450
rect 34188 17780 34244 17790
rect 34076 17778 34244 17780
rect 34076 17726 34190 17778
rect 34242 17726 34244 17778
rect 34076 17724 34244 17726
rect 34188 17714 34244 17724
rect 34524 17668 34580 17678
rect 34524 17574 34580 17612
rect 33852 16942 33854 16994
rect 33906 16942 33908 16994
rect 33852 16930 33908 16942
rect 33740 16884 33796 16894
rect 33740 16324 33796 16828
rect 34636 16772 34692 18398
rect 34748 18452 34804 18462
rect 34748 18358 34804 18396
rect 35308 18452 35364 18462
rect 35308 18450 35476 18452
rect 35308 18398 35310 18450
rect 35362 18398 35476 18450
rect 35308 18396 35476 18398
rect 35308 18386 35364 18396
rect 35420 18226 35476 18396
rect 35420 18174 35422 18226
rect 35474 18174 35476 18226
rect 35420 18162 35476 18174
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35420 17780 35476 17790
rect 35532 17780 35588 18508
rect 35420 17778 35588 17780
rect 35420 17726 35422 17778
rect 35474 17726 35588 17778
rect 35420 17724 35588 17726
rect 35644 18338 35700 18350
rect 35644 18286 35646 18338
rect 35698 18286 35700 18338
rect 35644 18226 35700 18286
rect 35644 18174 35646 18226
rect 35698 18174 35700 18226
rect 35644 17780 35700 18174
rect 35420 17714 35476 17724
rect 35644 17714 35700 17724
rect 34860 17444 34916 17454
rect 34860 17350 34916 17388
rect 36092 17108 36148 19964
rect 36204 18338 36260 18350
rect 36204 18286 36206 18338
rect 36258 18286 36260 18338
rect 36204 18228 36260 18286
rect 36204 18004 36260 18172
rect 36204 17938 36260 17948
rect 35644 17106 36372 17108
rect 35644 17054 36094 17106
rect 36146 17054 36372 17106
rect 35644 17052 36372 17054
rect 35644 16882 35700 17052
rect 36092 17042 36148 17052
rect 35644 16830 35646 16882
rect 35698 16830 35700 16882
rect 35644 16818 35700 16830
rect 35980 16884 36036 16894
rect 34636 16706 34692 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34972 16324 35028 16334
rect 33740 16322 34132 16324
rect 33740 16270 33742 16322
rect 33794 16270 34132 16322
rect 33740 16268 34132 16270
rect 33740 16258 33796 16268
rect 34076 16098 34132 16268
rect 34972 16210 35028 16268
rect 34972 16158 34974 16210
rect 35026 16158 35028 16210
rect 34972 16146 35028 16158
rect 34076 16046 34078 16098
rect 34130 16046 34132 16098
rect 34076 16034 34132 16046
rect 35756 15988 35812 15998
rect 33628 15986 34020 15988
rect 33628 15934 33630 15986
rect 33682 15934 34020 15986
rect 33628 15932 34020 15934
rect 33628 15922 33684 15932
rect 32172 15092 32340 15148
rect 32620 15874 32676 15886
rect 32620 15822 32622 15874
rect 32674 15822 32676 15874
rect 32004 15036 32116 15092
rect 31948 15026 32004 15036
rect 31052 14028 31220 14084
rect 31836 14418 31892 14430
rect 31836 14366 31838 14418
rect 31890 14366 31892 14418
rect 30380 12910 30382 12962
rect 30434 12910 30436 12962
rect 30380 12898 30436 12910
rect 30492 12908 30660 12964
rect 30828 12964 30884 12974
rect 30268 12180 30324 12190
rect 30268 12086 30324 12124
rect 30268 11620 30324 11630
rect 30324 11564 30436 11620
rect 30268 11554 30324 11564
rect 30268 11170 30324 11182
rect 30268 11118 30270 11170
rect 30322 11118 30324 11170
rect 30044 10668 30212 10724
rect 29932 10500 29988 10668
rect 30044 10500 30100 10510
rect 29932 10498 30100 10500
rect 29932 10446 30046 10498
rect 30098 10446 30100 10498
rect 29932 10444 30100 10446
rect 30044 10434 30100 10444
rect 29484 9660 29652 9716
rect 29372 9550 29374 9602
rect 29426 9550 29428 9602
rect 29260 8820 29316 8830
rect 29148 8764 29260 8820
rect 29260 8754 29316 8764
rect 29036 8642 29092 8652
rect 29260 8258 29316 8270
rect 29260 8206 29262 8258
rect 29314 8206 29316 8258
rect 29260 8148 29316 8206
rect 28812 8092 29316 8148
rect 28700 8054 28756 8092
rect 28700 7812 28756 7822
rect 28700 7586 28756 7756
rect 28812 7700 28868 7710
rect 28924 7700 28980 8092
rect 29372 8036 29428 9550
rect 29484 9044 29540 9054
rect 29484 8950 29540 8988
rect 29484 8372 29540 8382
rect 29484 8278 29540 8316
rect 28868 7644 28980 7700
rect 29036 7980 29428 8036
rect 28812 7634 28868 7644
rect 28700 7534 28702 7586
rect 28754 7534 28756 7586
rect 28700 7522 28756 7534
rect 28924 7474 28980 7486
rect 28924 7422 28926 7474
rect 28978 7422 28980 7474
rect 28588 7308 28756 7364
rect 28588 6916 28644 6926
rect 28588 6802 28644 6860
rect 28588 6750 28590 6802
rect 28642 6750 28644 6802
rect 28588 6738 28644 6750
rect 28364 6402 28420 6412
rect 28476 5794 28532 5806
rect 28476 5742 28478 5794
rect 28530 5742 28532 5794
rect 27916 5180 28420 5236
rect 28140 5010 28196 5022
rect 28140 4958 28142 5010
rect 28194 4958 28196 5010
rect 27132 4386 27188 4396
rect 28028 4788 28084 4798
rect 27020 4174 27022 4226
rect 27074 4174 27076 4226
rect 27020 4162 27076 4174
rect 27804 4228 27860 4238
rect 27804 3554 27860 4172
rect 27804 3502 27806 3554
rect 27858 3502 27860 3554
rect 27804 3490 27860 3502
rect 26460 924 26740 980
rect 26684 800 26740 924
rect 28028 800 28084 4732
rect 28140 4676 28196 4958
rect 28140 4610 28196 4620
rect 28364 3442 28420 5180
rect 28476 4452 28532 5742
rect 28700 4788 28756 7308
rect 28812 7028 28868 7038
rect 28812 5012 28868 6972
rect 28924 6356 28980 7422
rect 29036 6804 29092 7980
rect 29484 7700 29540 7710
rect 29372 7698 29540 7700
rect 29372 7646 29486 7698
rect 29538 7646 29540 7698
rect 29372 7644 29540 7646
rect 29148 7476 29204 7486
rect 29148 7382 29204 7420
rect 29260 7474 29316 7486
rect 29260 7422 29262 7474
rect 29314 7422 29316 7474
rect 29260 7028 29316 7422
rect 29260 6962 29316 6972
rect 29260 6804 29316 6814
rect 29036 6748 29260 6804
rect 29260 6710 29316 6748
rect 29148 6578 29204 6590
rect 29148 6526 29150 6578
rect 29202 6526 29204 6578
rect 29148 6468 29204 6526
rect 29148 6402 29204 6412
rect 28924 6290 28980 6300
rect 28812 4946 28868 4956
rect 28924 6020 28980 6030
rect 28700 4722 28756 4732
rect 28476 4386 28532 4396
rect 28924 4004 28980 5964
rect 29372 6018 29428 7644
rect 29484 7634 29540 7644
rect 29596 7252 29652 9660
rect 29484 7196 29652 7252
rect 29484 7140 29540 7196
rect 29484 7074 29540 7084
rect 29596 7028 29652 7038
rect 29484 6916 29540 6926
rect 29484 6822 29540 6860
rect 29596 6914 29652 6972
rect 29596 6862 29598 6914
rect 29650 6862 29652 6914
rect 29596 6850 29652 6862
rect 29372 5966 29374 6018
rect 29426 5966 29428 6018
rect 29372 5954 29428 5966
rect 29596 6020 29652 6030
rect 29484 5124 29540 5134
rect 29484 5030 29540 5068
rect 29148 4452 29204 4462
rect 29148 4358 29204 4396
rect 28924 3938 28980 3948
rect 28700 3556 28756 3566
rect 28700 3462 28756 3500
rect 28364 3390 28366 3442
rect 28418 3390 28420 3442
rect 28364 3378 28420 3390
rect 29596 3388 29652 5964
rect 29708 4340 29764 10332
rect 29820 10386 29876 10398
rect 29820 10334 29822 10386
rect 29874 10334 29876 10386
rect 29820 7588 29876 10334
rect 29932 9828 29988 9838
rect 29932 9734 29988 9772
rect 30156 9604 30212 10668
rect 30268 10388 30324 11118
rect 30380 10610 30436 11564
rect 30380 10558 30382 10610
rect 30434 10558 30436 10610
rect 30380 10546 30436 10558
rect 30492 10500 30548 12908
rect 30828 12870 30884 12908
rect 30940 12852 30996 12862
rect 30604 12738 30660 12750
rect 30604 12686 30606 12738
rect 30658 12686 30660 12738
rect 30604 12628 30660 12686
rect 30604 12562 30660 12572
rect 30716 12738 30772 12750
rect 30716 12686 30718 12738
rect 30770 12686 30772 12738
rect 30716 12404 30772 12686
rect 30716 12348 30884 12404
rect 30828 11732 30884 12348
rect 30940 12180 30996 12796
rect 30940 12114 30996 12124
rect 31052 12516 31108 14028
rect 31164 13860 31220 13870
rect 31164 13766 31220 13804
rect 31500 13860 31556 13870
rect 31388 13748 31444 13758
rect 31276 13522 31332 13534
rect 31276 13470 31278 13522
rect 31330 13470 31332 13522
rect 31276 12740 31332 13470
rect 31388 12962 31444 13692
rect 31388 12910 31390 12962
rect 31442 12910 31444 12962
rect 31388 12898 31444 12910
rect 31500 13300 31556 13804
rect 31612 13634 31668 13646
rect 31612 13582 31614 13634
rect 31666 13582 31668 13634
rect 31612 13522 31668 13582
rect 31612 13470 31614 13522
rect 31666 13470 31668 13522
rect 31612 13458 31668 13470
rect 31500 12964 31556 13244
rect 31724 13412 31780 13422
rect 31612 12964 31668 12974
rect 31500 12962 31668 12964
rect 31500 12910 31614 12962
rect 31666 12910 31668 12962
rect 31500 12908 31668 12910
rect 31612 12898 31668 12908
rect 31276 12684 31668 12740
rect 30828 11676 30996 11732
rect 30828 11396 30884 11406
rect 30492 10444 30772 10500
rect 30268 10332 30660 10388
rect 30492 10052 30548 10062
rect 30492 9938 30548 9996
rect 30492 9886 30494 9938
rect 30546 9886 30548 9938
rect 29932 9548 30212 9604
rect 30268 9826 30324 9838
rect 30268 9774 30270 9826
rect 30322 9774 30324 9826
rect 29932 8482 29988 9548
rect 30268 9492 30324 9774
rect 30156 9436 30324 9492
rect 30044 9044 30100 9054
rect 30044 8950 30100 8988
rect 29932 8430 29934 8482
rect 29986 8430 29988 8482
rect 29932 8418 29988 8430
rect 29932 8260 29988 8270
rect 29932 8166 29988 8204
rect 30044 8146 30100 8158
rect 30044 8094 30046 8146
rect 30098 8094 30100 8146
rect 30044 7812 30100 8094
rect 30044 7746 30100 7756
rect 29820 7532 30100 7588
rect 29820 7362 29876 7374
rect 29820 7310 29822 7362
rect 29874 7310 29876 7362
rect 29820 6132 29876 7310
rect 29932 6580 29988 6590
rect 29932 6486 29988 6524
rect 29820 6066 29876 6076
rect 30044 6020 30100 7532
rect 30156 6916 30212 9436
rect 30380 9044 30436 9054
rect 30268 9042 30436 9044
rect 30268 8990 30382 9042
rect 30434 8990 30436 9042
rect 30268 8988 30436 8990
rect 30268 8820 30324 8988
rect 30380 8978 30436 8988
rect 30492 8820 30548 9886
rect 30604 9604 30660 10332
rect 30604 9538 30660 9548
rect 30268 8754 30324 8764
rect 30380 8764 30548 8820
rect 30716 9044 30772 10444
rect 30828 9826 30884 11340
rect 30940 10612 30996 11676
rect 30940 10546 30996 10556
rect 30828 9774 30830 9826
rect 30882 9774 30884 9826
rect 30828 9762 30884 9774
rect 31052 9604 31108 12460
rect 31388 12178 31444 12190
rect 31388 12126 31390 12178
rect 31442 12126 31444 12178
rect 31388 10836 31444 12126
rect 31612 10948 31668 12684
rect 31724 12290 31780 13356
rect 31836 12738 31892 14366
rect 31948 13188 32004 13198
rect 31948 13094 32004 13132
rect 32060 13076 32116 15036
rect 32172 13634 32228 15092
rect 32508 14308 32564 14318
rect 32508 13970 32564 14252
rect 32508 13918 32510 13970
rect 32562 13918 32564 13970
rect 32508 13906 32564 13918
rect 32172 13582 32174 13634
rect 32226 13582 32228 13634
rect 32172 13412 32228 13582
rect 32172 13346 32228 13356
rect 32284 13188 32340 13198
rect 32508 13188 32564 13198
rect 32340 13186 32564 13188
rect 32340 13134 32510 13186
rect 32562 13134 32564 13186
rect 32340 13132 32564 13134
rect 32284 13122 32340 13132
rect 32508 13122 32564 13132
rect 32060 13020 32228 13076
rect 31948 12964 32004 12974
rect 31948 12962 32116 12964
rect 31948 12910 31950 12962
rect 32002 12910 32116 12962
rect 31948 12908 32116 12910
rect 31948 12898 32004 12908
rect 31836 12686 31838 12738
rect 31890 12686 31892 12738
rect 31836 12674 31892 12686
rect 32060 12740 32116 12908
rect 32060 12674 32116 12684
rect 31724 12238 31726 12290
rect 31778 12238 31780 12290
rect 31724 12226 31780 12238
rect 32172 12178 32228 13020
rect 32508 12964 32564 12974
rect 32508 12870 32564 12908
rect 32620 12516 32676 15822
rect 33964 15876 34020 15932
rect 35644 15986 35812 15988
rect 35644 15934 35758 15986
rect 35810 15934 35812 15986
rect 35644 15932 35812 15934
rect 34412 15876 34468 15886
rect 33964 15820 34132 15876
rect 34076 15538 34132 15820
rect 34412 15782 34468 15820
rect 35532 15874 35588 15886
rect 35532 15822 35534 15874
rect 35586 15822 35588 15874
rect 34076 15486 34078 15538
rect 34130 15486 34132 15538
rect 34076 15474 34132 15486
rect 34860 15540 34916 15550
rect 33964 15428 34020 15438
rect 33964 14642 34020 15372
rect 33964 14590 33966 14642
rect 34018 14590 34020 14642
rect 33516 14308 33572 14318
rect 33572 14252 33684 14308
rect 33516 14242 33572 14252
rect 33516 13636 33572 13646
rect 33516 13542 33572 13580
rect 33628 12964 33684 14252
rect 33516 12962 33684 12964
rect 33516 12910 33630 12962
rect 33682 12910 33684 12962
rect 33516 12908 33684 12910
rect 32172 12126 32174 12178
rect 32226 12126 32228 12178
rect 32172 12114 32228 12126
rect 32284 12460 32676 12516
rect 32844 12852 32900 12862
rect 32060 12068 32116 12078
rect 31612 10892 31780 10948
rect 31388 10610 31444 10780
rect 31388 10558 31390 10610
rect 31442 10558 31444 10610
rect 31388 10546 31444 10558
rect 31500 10834 31556 10846
rect 31500 10782 31502 10834
rect 31554 10782 31556 10834
rect 31052 9538 31108 9548
rect 31164 9938 31220 9950
rect 31164 9886 31166 9938
rect 31218 9886 31220 9938
rect 30156 6850 30212 6860
rect 30268 8484 30324 8494
rect 30268 6130 30324 8428
rect 30380 8146 30436 8764
rect 30380 8094 30382 8146
rect 30434 8094 30436 8146
rect 30380 8082 30436 8094
rect 30492 8372 30548 8382
rect 30492 7028 30548 8316
rect 30716 8260 30772 8988
rect 30828 8930 30884 8942
rect 30828 8878 30830 8930
rect 30882 8878 30884 8930
rect 30828 8484 30884 8878
rect 30828 8418 30884 8428
rect 30716 8166 30772 8204
rect 31052 7588 31108 7598
rect 31052 7494 31108 7532
rect 30268 6078 30270 6130
rect 30322 6078 30324 6130
rect 30268 6066 30324 6078
rect 30380 6916 30436 6926
rect 30492 6916 30548 6972
rect 30380 6914 30548 6916
rect 30380 6862 30382 6914
rect 30434 6862 30548 6914
rect 30380 6860 30548 6862
rect 30604 6916 30660 6926
rect 30044 5954 30100 5964
rect 30268 5908 30324 5918
rect 30380 5908 30436 6860
rect 30604 6822 30660 6860
rect 30828 6804 30884 6814
rect 30828 6710 30884 6748
rect 30268 5906 30436 5908
rect 30268 5854 30270 5906
rect 30322 5854 30436 5906
rect 30268 5852 30436 5854
rect 30492 6692 30548 6702
rect 30268 5842 30324 5852
rect 30380 5684 30436 5694
rect 30492 5684 30548 6636
rect 30604 6580 30660 6590
rect 30604 5906 30660 6524
rect 30604 5854 30606 5906
rect 30658 5854 30660 5906
rect 30604 5842 30660 5854
rect 30380 5682 30548 5684
rect 30380 5630 30382 5682
rect 30434 5630 30548 5682
rect 30380 5628 30548 5630
rect 30380 5618 30436 5628
rect 29820 5010 29876 5022
rect 29820 4958 29822 5010
rect 29874 4958 29876 5010
rect 29820 4788 29876 4958
rect 29820 4722 29876 4732
rect 30716 5012 30772 5022
rect 30716 4562 30772 4956
rect 30716 4510 30718 4562
rect 30770 4510 30772 4562
rect 30716 4498 30772 4510
rect 29820 4340 29876 4350
rect 29708 4284 29820 4340
rect 29820 4246 29876 4284
rect 30604 4228 30660 4238
rect 30604 4134 30660 4172
rect 31052 4226 31108 4238
rect 31052 4174 31054 4226
rect 31106 4174 31108 4226
rect 31052 3556 31108 4174
rect 31052 3490 31108 3500
rect 31164 3554 31220 9886
rect 31276 9716 31332 9726
rect 31500 9716 31556 10782
rect 31612 10724 31668 10734
rect 31612 10630 31668 10668
rect 31276 9714 31556 9716
rect 31276 9662 31278 9714
rect 31330 9662 31556 9714
rect 31276 9660 31556 9662
rect 31276 9650 31332 9660
rect 31500 9042 31556 9054
rect 31500 8990 31502 9042
rect 31554 8990 31556 9042
rect 31388 7812 31444 7822
rect 31388 7252 31444 7756
rect 31388 6690 31444 7196
rect 31388 6638 31390 6690
rect 31442 6638 31444 6690
rect 31388 6626 31444 6638
rect 31276 5794 31332 5806
rect 31276 5742 31278 5794
rect 31330 5742 31332 5794
rect 31276 3892 31332 5742
rect 31500 5796 31556 8990
rect 31724 8596 31780 10892
rect 32060 10610 32116 12012
rect 32060 10558 32062 10610
rect 32114 10558 32116 10610
rect 32060 10546 32116 10558
rect 31948 10500 32004 10510
rect 31836 9828 31892 9838
rect 31948 9828 32004 10444
rect 32284 9940 32340 12460
rect 32396 12290 32452 12302
rect 32396 12238 32398 12290
rect 32450 12238 32452 12290
rect 32396 10722 32452 12238
rect 32844 12292 32900 12796
rect 32844 12226 32900 12236
rect 32396 10670 32398 10722
rect 32450 10670 32452 10722
rect 32396 10052 32452 10670
rect 32508 12066 32564 12078
rect 32508 12014 32510 12066
rect 32562 12014 32564 12066
rect 32508 10724 32564 12014
rect 33516 11506 33572 12908
rect 33628 12898 33684 12908
rect 33852 13746 33908 13758
rect 33852 13694 33854 13746
rect 33906 13694 33908 13746
rect 33852 12740 33908 13694
rect 33964 12964 34020 14590
rect 34300 15092 34356 15102
rect 34188 13972 34244 13982
rect 34076 13970 34244 13972
rect 34076 13918 34190 13970
rect 34242 13918 34244 13970
rect 34076 13916 34244 13918
rect 34076 13188 34132 13916
rect 34188 13906 34244 13916
rect 34300 13746 34356 15036
rect 34412 14308 34468 14318
rect 34860 14308 34916 15484
rect 35532 15540 35588 15822
rect 35532 15474 35588 15484
rect 35644 15876 35700 15932
rect 35756 15922 35812 15932
rect 35644 15316 35700 15820
rect 35868 15874 35924 15886
rect 35868 15822 35870 15874
rect 35922 15822 35924 15874
rect 35868 15540 35924 15822
rect 35868 15474 35924 15484
rect 35980 15538 36036 16828
rect 36092 15876 36148 15886
rect 36092 15782 36148 15820
rect 36316 15764 36372 17052
rect 36428 16212 36484 16222
rect 36428 16118 36484 16156
rect 36316 15708 36484 15764
rect 35980 15486 35982 15538
rect 36034 15486 36036 15538
rect 35980 15474 36036 15486
rect 35644 15250 35700 15260
rect 35756 15426 35812 15438
rect 35756 15374 35758 15426
rect 35810 15374 35812 15426
rect 35756 15148 35812 15374
rect 36316 15428 36372 15438
rect 36316 15334 36372 15372
rect 36204 15316 36260 15326
rect 36204 15222 36260 15260
rect 36428 15148 36484 15708
rect 36540 15540 36596 15550
rect 36764 15540 36820 20748
rect 36876 20738 36932 20748
rect 37212 20578 37268 22204
rect 37324 20860 37716 20916
rect 37324 20802 37380 20860
rect 37324 20750 37326 20802
rect 37378 20750 37380 20802
rect 37324 20738 37380 20750
rect 37660 20804 37716 20860
rect 37772 20804 37828 20814
rect 37660 20802 37828 20804
rect 37660 20750 37774 20802
rect 37826 20750 37828 20802
rect 37660 20748 37828 20750
rect 37772 20738 37828 20748
rect 37212 20526 37214 20578
rect 37266 20526 37268 20578
rect 37212 20514 37268 20526
rect 37548 20692 37604 20702
rect 37100 19908 37156 19918
rect 37100 19346 37156 19852
rect 37100 19294 37102 19346
rect 37154 19294 37156 19346
rect 37100 19282 37156 19294
rect 37324 19348 37380 19358
rect 37324 19234 37380 19292
rect 37324 19182 37326 19234
rect 37378 19182 37380 19234
rect 37324 19170 37380 19182
rect 37548 19236 37604 20636
rect 37548 19142 37604 19180
rect 36988 19122 37044 19134
rect 36988 19070 36990 19122
rect 37042 19070 37044 19122
rect 36988 18564 37044 19070
rect 36876 18508 37044 18564
rect 36876 16884 36932 18508
rect 37324 18450 37380 18462
rect 37324 18398 37326 18450
rect 37378 18398 37380 18450
rect 36988 18338 37044 18350
rect 36988 18286 36990 18338
rect 37042 18286 37044 18338
rect 36988 18116 37044 18286
rect 37324 18116 37380 18398
rect 36988 18060 37380 18116
rect 36876 16818 36932 16828
rect 36988 16212 37044 16222
rect 37100 16212 37156 18060
rect 37772 17108 37828 17118
rect 37884 17108 37940 30828
rect 43708 29540 43764 55020
rect 49644 55076 49700 55086
rect 49980 55076 50036 55134
rect 49700 55020 50036 55076
rect 50988 55076 51044 55086
rect 49644 54982 49700 55020
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50988 43708 51044 55020
rect 50988 43652 51268 43708
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 51212 38668 51268 43652
rect 56028 38668 56084 55412
rect 61292 55410 61348 56028
rect 61292 55358 61294 55410
rect 61346 55358 61348 55410
rect 61292 55346 61348 55358
rect 61740 56082 61796 56094
rect 61740 56030 61742 56082
rect 61794 56030 61796 56082
rect 60508 55298 60564 55310
rect 60508 55246 60510 55298
rect 60562 55246 60564 55298
rect 59948 55076 60004 55086
rect 59948 54982 60004 55020
rect 60508 55076 60564 55246
rect 60956 55300 61012 55310
rect 60956 55206 61012 55244
rect 61740 55300 61796 56030
rect 62972 56084 63028 56094
rect 62972 55990 63028 56028
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 66556 55410 66612 56252
rect 66780 56242 66836 56252
rect 70364 56308 70420 59200
rect 70364 56242 70420 56252
rect 71596 56308 71652 56318
rect 71596 56214 71652 56252
rect 67116 56196 67172 56206
rect 67116 56102 67172 56140
rect 68012 56196 68068 56206
rect 66556 55358 66558 55410
rect 66610 55358 66612 55410
rect 66556 55346 66612 55358
rect 60508 55010 60564 55020
rect 61740 55074 61796 55244
rect 62188 55300 62244 55310
rect 62188 55206 62244 55244
rect 62972 55300 63028 55310
rect 61740 55022 61742 55074
rect 61794 55022 61796 55074
rect 61740 38668 61796 55022
rect 51212 38612 51492 38668
rect 56028 38612 56420 38668
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 46844 32004 46900 32014
rect 46060 30210 46116 30222
rect 46060 30158 46062 30210
rect 46114 30158 46116 30210
rect 43708 29538 44212 29540
rect 43708 29486 43710 29538
rect 43762 29486 44212 29538
rect 43708 29484 44212 29486
rect 43708 29474 43764 29484
rect 43372 28868 43428 28878
rect 40348 27746 40404 27758
rect 40348 27694 40350 27746
rect 40402 27694 40404 27746
rect 39676 26962 39732 26974
rect 39676 26910 39678 26962
rect 39730 26910 39732 26962
rect 38556 26740 38612 26750
rect 38332 26628 38388 26638
rect 38332 26404 38388 26572
rect 38556 26516 38612 26684
rect 38332 26310 38388 26348
rect 38444 26460 38836 26516
rect 38444 26402 38500 26460
rect 38444 26350 38446 26402
rect 38498 26350 38500 26402
rect 37996 26292 38052 26302
rect 37996 26178 38052 26236
rect 38444 26292 38500 26350
rect 38444 26226 38500 26236
rect 37996 26126 37998 26178
rect 38050 26126 38052 26178
rect 37996 25396 38052 26126
rect 38444 26068 38500 26078
rect 38444 26066 38612 26068
rect 38444 26014 38446 26066
rect 38498 26014 38612 26066
rect 38444 26012 38612 26014
rect 38444 26002 38500 26012
rect 37996 25330 38052 25340
rect 38556 25394 38612 26012
rect 38556 25342 38558 25394
rect 38610 25342 38612 25394
rect 38556 25330 38612 25342
rect 38780 25508 38836 26460
rect 39452 26404 39508 26414
rect 39452 26310 39508 26348
rect 39004 26290 39060 26302
rect 39004 26238 39006 26290
rect 39058 26238 39060 26290
rect 39004 26180 39060 26238
rect 39116 26292 39172 26302
rect 39116 26290 39284 26292
rect 39116 26238 39118 26290
rect 39170 26238 39284 26290
rect 39116 26236 39284 26238
rect 39116 26226 39172 26236
rect 39004 25844 39060 26124
rect 39004 25788 39172 25844
rect 39004 25618 39060 25630
rect 39004 25566 39006 25618
rect 39058 25566 39060 25618
rect 38220 25284 38276 25294
rect 38220 25190 38276 25228
rect 38444 25282 38500 25294
rect 38444 25230 38446 25282
rect 38498 25230 38500 25282
rect 38444 24948 38500 25230
rect 38780 24948 38836 25452
rect 38892 25506 38948 25518
rect 38892 25454 38894 25506
rect 38946 25454 38948 25506
rect 38892 25396 38948 25454
rect 38892 25330 38948 25340
rect 39004 25172 39060 25566
rect 39116 25396 39172 25788
rect 39228 25620 39284 26236
rect 39340 26178 39396 26190
rect 39340 26126 39342 26178
rect 39394 26126 39396 26178
rect 39340 25732 39396 26126
rect 39676 26180 39732 26910
rect 39900 26964 39956 26974
rect 39900 26516 39956 26908
rect 40124 26964 40180 26974
rect 39900 26450 39956 26460
rect 40012 26850 40068 26862
rect 40012 26798 40014 26850
rect 40066 26798 40068 26850
rect 39788 26292 39844 26302
rect 39788 26198 39844 26236
rect 40012 26290 40068 26798
rect 40012 26238 40014 26290
rect 40066 26238 40068 26290
rect 40012 26226 40068 26238
rect 39676 26114 39732 26124
rect 39340 25676 40068 25732
rect 39228 25564 39508 25620
rect 39340 25396 39396 25406
rect 39116 25394 39396 25396
rect 39116 25342 39342 25394
rect 39394 25342 39396 25394
rect 39116 25340 39396 25342
rect 39340 25330 39396 25340
rect 39004 25116 39172 25172
rect 39004 24948 39060 24958
rect 38780 24946 39060 24948
rect 38780 24894 39006 24946
rect 39058 24894 39060 24946
rect 38780 24892 39060 24894
rect 38444 24882 38500 24892
rect 39004 24882 39060 24892
rect 38556 24500 38612 24510
rect 38444 24444 38556 24500
rect 38332 23492 38388 23502
rect 38332 23378 38388 23436
rect 38332 23326 38334 23378
rect 38386 23326 38388 23378
rect 38332 23314 38388 23326
rect 37996 22820 38052 22830
rect 37996 20690 38052 22764
rect 38444 20916 38500 24444
rect 38556 24434 38612 24444
rect 39116 23940 39172 25116
rect 39452 25060 39508 25564
rect 39564 25508 39620 25518
rect 39564 25414 39620 25452
rect 40012 25506 40068 25676
rect 40124 25620 40180 26908
rect 40236 26962 40292 26974
rect 40236 26910 40238 26962
rect 40290 26910 40292 26962
rect 40236 26404 40292 26910
rect 40348 26964 40404 27694
rect 40572 26964 40628 26974
rect 40348 26962 40628 26964
rect 40348 26910 40574 26962
rect 40626 26910 40628 26962
rect 40348 26908 40628 26910
rect 40572 26740 40628 26908
rect 40796 26964 40852 26974
rect 40796 26870 40852 26908
rect 41020 26962 41076 26974
rect 41020 26910 41022 26962
rect 41074 26910 41076 26962
rect 40572 26674 40628 26684
rect 40684 26850 40740 26862
rect 40684 26798 40686 26850
rect 40738 26798 40740 26850
rect 40236 26338 40292 26348
rect 40684 26292 40740 26798
rect 40796 26292 40852 26302
rect 40684 26290 40852 26292
rect 40684 26238 40798 26290
rect 40850 26238 40852 26290
rect 40684 26236 40852 26238
rect 40796 26226 40852 26236
rect 40348 26066 40404 26078
rect 40348 26014 40350 26066
rect 40402 26014 40404 26066
rect 40124 25564 40292 25620
rect 40012 25454 40014 25506
rect 40066 25454 40068 25506
rect 40012 25442 40068 25454
rect 40124 25284 40180 25294
rect 40124 25190 40180 25228
rect 40236 25282 40292 25564
rect 40348 25508 40404 26014
rect 41020 25956 41076 26910
rect 41244 26516 41300 26526
rect 41692 26516 41748 26526
rect 41244 26514 41748 26516
rect 41244 26462 41246 26514
rect 41298 26462 41694 26514
rect 41746 26462 41748 26514
rect 41244 26460 41748 26462
rect 41244 26450 41300 26460
rect 41692 26450 41748 26460
rect 41916 26516 41972 26526
rect 41916 26422 41972 26460
rect 42028 26404 42084 26414
rect 42028 26310 42084 26348
rect 42588 26404 42644 26414
rect 42588 26310 42644 26348
rect 43260 26404 43316 26414
rect 43260 26310 43316 26348
rect 41468 26292 41524 26302
rect 42812 26292 42868 26302
rect 41468 26198 41524 26236
rect 42700 26236 42812 26292
rect 41356 26180 41412 26190
rect 41356 26086 41412 26124
rect 40348 25442 40404 25452
rect 40796 25900 41076 25956
rect 40460 25396 40516 25406
rect 40460 25302 40516 25340
rect 40236 25230 40238 25282
rect 40290 25230 40292 25282
rect 39452 24994 39508 25004
rect 40236 24724 40292 25230
rect 40236 24658 40292 24668
rect 39340 23940 39396 23950
rect 39116 23938 39396 23940
rect 39116 23886 39342 23938
rect 39394 23886 39396 23938
rect 39116 23884 39396 23886
rect 39340 23874 39396 23884
rect 39564 23940 39620 23950
rect 39564 23846 39620 23884
rect 40012 23938 40068 23950
rect 40012 23886 40014 23938
rect 40066 23886 40068 23938
rect 40012 23828 40068 23886
rect 40012 23762 40068 23772
rect 40460 23828 40516 23838
rect 40460 23734 40516 23772
rect 39452 23716 39508 23726
rect 39452 23622 39508 23660
rect 38556 23604 38612 23614
rect 38556 23154 38612 23548
rect 40796 23492 40852 25900
rect 41244 25508 41300 25518
rect 41244 25414 41300 25452
rect 41692 25506 41748 25518
rect 41692 25454 41694 25506
rect 41746 25454 41748 25506
rect 41020 25284 41076 25294
rect 41020 25190 41076 25228
rect 41132 25282 41188 25294
rect 41132 25230 41134 25282
rect 41186 25230 41188 25282
rect 41132 24724 41188 25230
rect 41132 24658 41188 24668
rect 40796 23426 40852 23436
rect 41132 23380 41188 23390
rect 41020 23268 41076 23278
rect 41020 23174 41076 23212
rect 38556 23102 38558 23154
rect 38610 23102 38612 23154
rect 38556 23090 38612 23102
rect 40796 23154 40852 23166
rect 40796 23102 40798 23154
rect 40850 23102 40852 23154
rect 40796 23044 40852 23102
rect 41132 23154 41188 23324
rect 41132 23102 41134 23154
rect 41186 23102 41188 23154
rect 41132 23090 41188 23102
rect 41468 23154 41524 23166
rect 41468 23102 41470 23154
rect 41522 23102 41524 23154
rect 39788 22484 39844 22494
rect 39788 22370 39844 22428
rect 40348 22484 40404 22494
rect 40348 22390 40404 22428
rect 39788 22318 39790 22370
rect 39842 22318 39844 22370
rect 39788 22306 39844 22318
rect 39116 22260 39172 22270
rect 39116 22166 39172 22204
rect 38556 20916 38612 20926
rect 38444 20914 38612 20916
rect 38444 20862 38558 20914
rect 38610 20862 38612 20914
rect 38444 20860 38612 20862
rect 37996 20638 37998 20690
rect 38050 20638 38052 20690
rect 37996 20626 38052 20638
rect 38108 20690 38164 20702
rect 38108 20638 38110 20690
rect 38162 20638 38164 20690
rect 38108 20132 38164 20638
rect 38444 20692 38500 20860
rect 38556 20850 38612 20860
rect 38444 20626 38500 20636
rect 40012 20244 40068 20254
rect 38332 20132 38388 20142
rect 38164 20130 38388 20132
rect 38164 20078 38334 20130
rect 38386 20078 38388 20130
rect 38164 20076 38388 20078
rect 38108 20066 38164 20076
rect 38332 20066 38388 20076
rect 38444 20132 38500 20142
rect 38444 20038 38500 20076
rect 39004 20132 39060 20142
rect 37996 19908 38052 19918
rect 37996 19814 38052 19852
rect 39004 19908 39060 20076
rect 39004 19814 39060 19852
rect 38444 19794 38500 19806
rect 38444 19742 38446 19794
rect 38498 19742 38500 19794
rect 38220 19348 38276 19358
rect 38444 19348 38500 19742
rect 38276 19292 38500 19348
rect 39116 19460 39172 19470
rect 38220 19282 38276 19292
rect 37996 19236 38052 19246
rect 37996 19142 38052 19180
rect 39116 19234 39172 19404
rect 39900 19236 39956 19246
rect 39116 19182 39118 19234
rect 39170 19182 39172 19234
rect 39116 19170 39172 19182
rect 39788 19180 39900 19236
rect 39788 19122 39844 19180
rect 39788 19070 39790 19122
rect 39842 19070 39844 19122
rect 39788 19058 39844 19070
rect 38108 18338 38164 18350
rect 38108 18286 38110 18338
rect 38162 18286 38164 18338
rect 37884 17052 38052 17108
rect 37044 16156 37156 16212
rect 37212 16884 37268 16894
rect 36988 16098 37044 16156
rect 36988 16046 36990 16098
rect 37042 16046 37044 16098
rect 36988 16034 37044 16046
rect 36540 15538 36820 15540
rect 36540 15486 36542 15538
rect 36594 15486 36820 15538
rect 36540 15484 36820 15486
rect 36988 15876 37044 15886
rect 36540 15474 36596 15484
rect 36988 15314 37044 15820
rect 36988 15262 36990 15314
rect 37042 15262 37044 15314
rect 36988 15250 37044 15262
rect 37212 15316 37268 16828
rect 37772 16882 37828 17052
rect 37772 16830 37774 16882
rect 37826 16830 37828 16882
rect 37772 16818 37828 16830
rect 37996 16660 38052 17052
rect 38108 17106 38164 18286
rect 39452 17668 39508 17678
rect 39004 17556 39060 17566
rect 38108 17054 38110 17106
rect 38162 17054 38164 17106
rect 38108 17042 38164 17054
rect 38220 17444 38276 17454
rect 38220 16994 38276 17388
rect 39004 17332 39060 17500
rect 39452 17554 39508 17612
rect 39452 17502 39454 17554
rect 39506 17502 39508 17554
rect 39452 17490 39508 17502
rect 39564 17556 39620 17566
rect 39564 17462 39620 17500
rect 39228 17444 39284 17454
rect 39228 17350 39284 17388
rect 38220 16942 38222 16994
rect 38274 16942 38276 16994
rect 38220 16930 38276 16942
rect 38892 16994 38948 17006
rect 38892 16942 38894 16994
rect 38946 16942 38948 16994
rect 38332 16882 38388 16894
rect 38332 16830 38334 16882
rect 38386 16830 38388 16882
rect 37884 16604 38052 16660
rect 38220 16660 38276 16670
rect 37772 15988 37828 15998
rect 37324 15986 37828 15988
rect 37324 15934 37774 15986
rect 37826 15934 37828 15986
rect 37324 15932 37828 15934
rect 37324 15538 37380 15932
rect 37772 15922 37828 15932
rect 37324 15486 37326 15538
rect 37378 15486 37380 15538
rect 37324 15474 37380 15486
rect 37660 15764 37716 15774
rect 37660 15426 37716 15708
rect 37660 15374 37662 15426
rect 37714 15374 37716 15426
rect 37660 15362 37716 15374
rect 37324 15316 37380 15326
rect 37212 15314 37380 15316
rect 37212 15262 37326 15314
rect 37378 15262 37380 15314
rect 37212 15260 37380 15262
rect 37324 15250 37380 15260
rect 35532 15092 35812 15148
rect 36204 15092 36484 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34412 14214 34468 14252
rect 34748 14306 34916 14308
rect 34748 14254 34862 14306
rect 34914 14254 34916 14306
rect 34748 14252 34916 14254
rect 34300 13694 34302 13746
rect 34354 13694 34356 13746
rect 34300 13636 34356 13694
rect 34636 13748 34692 13758
rect 34636 13654 34692 13692
rect 34300 13570 34356 13580
rect 34188 13524 34244 13534
rect 34188 13430 34244 13468
rect 34076 13132 34356 13188
rect 34300 13074 34356 13132
rect 34300 13022 34302 13074
rect 34354 13022 34356 13074
rect 34300 13010 34356 13022
rect 33964 12898 34020 12908
rect 33852 12674 33908 12684
rect 33516 11454 33518 11506
rect 33570 11454 33572 11506
rect 33516 11442 33572 11454
rect 34412 12066 34468 12078
rect 34412 12014 34414 12066
rect 34466 12014 34468 12066
rect 34412 11394 34468 12014
rect 34412 11342 34414 11394
rect 34466 11342 34468 11394
rect 34300 11172 34356 11182
rect 33964 10834 34020 10846
rect 33964 10782 33966 10834
rect 34018 10782 34020 10834
rect 32508 10658 32564 10668
rect 33404 10724 33460 10734
rect 33404 10630 33460 10668
rect 33068 10612 33124 10622
rect 33068 10518 33124 10556
rect 32956 10500 33012 10510
rect 32396 9996 32676 10052
rect 32340 9884 32452 9940
rect 32284 9874 32340 9884
rect 31836 9826 32004 9828
rect 31836 9774 31838 9826
rect 31890 9774 32004 9826
rect 31836 9772 32004 9774
rect 32396 9826 32452 9884
rect 32396 9774 32398 9826
rect 32450 9774 32452 9826
rect 31836 9762 31892 9772
rect 32396 9762 32452 9774
rect 32620 9716 32676 9996
rect 32956 9940 33012 10444
rect 33404 9940 33460 9950
rect 32956 9884 33236 9940
rect 32732 9716 32788 9726
rect 32620 9714 32788 9716
rect 32620 9662 32734 9714
rect 32786 9662 32788 9714
rect 32620 9660 32788 9662
rect 32172 9154 32228 9166
rect 32172 9102 32174 9154
rect 32226 9102 32228 9154
rect 31836 8930 31892 8942
rect 31836 8878 31838 8930
rect 31890 8878 31892 8930
rect 31836 8820 31892 8878
rect 31836 8754 31892 8764
rect 31724 8540 31892 8596
rect 31500 5730 31556 5740
rect 31612 8484 31668 8494
rect 31276 3826 31332 3836
rect 31164 3502 31166 3554
rect 31218 3502 31220 3554
rect 31164 3490 31220 3502
rect 29372 3332 29652 3388
rect 30604 3332 30660 3342
rect 29372 800 29428 3332
rect 30604 3330 30772 3332
rect 30604 3278 30606 3330
rect 30658 3278 30772 3330
rect 30604 3276 30772 3278
rect 30604 3266 30660 3276
rect 30716 800 30772 3276
rect 31612 1652 31668 8428
rect 31724 6916 31780 6926
rect 31724 6690 31780 6860
rect 31724 6638 31726 6690
rect 31778 6638 31780 6690
rect 31724 6626 31780 6638
rect 31836 5572 31892 8540
rect 32172 8372 32228 9102
rect 32508 9044 32564 9054
rect 32508 8950 32564 8988
rect 32172 8306 32228 8316
rect 32620 8260 32676 8270
rect 32620 8166 32676 8204
rect 32732 8148 32788 9660
rect 32956 9716 33012 9726
rect 32956 8370 33012 9660
rect 32956 8318 32958 8370
rect 33010 8318 33012 8370
rect 32956 8306 33012 8318
rect 33068 9492 33124 9502
rect 33068 8258 33124 9436
rect 33068 8206 33070 8258
rect 33122 8206 33124 8258
rect 33068 8194 33124 8206
rect 32732 8082 32788 8092
rect 32172 7924 32228 7934
rect 32172 7698 32228 7868
rect 32172 7646 32174 7698
rect 32226 7646 32228 7698
rect 32172 7634 32228 7646
rect 32284 7588 32340 7598
rect 32060 6244 32116 6254
rect 31836 4788 31892 5516
rect 31836 4722 31892 4732
rect 31948 6188 32060 6244
rect 31948 3388 32004 6188
rect 32060 6178 32116 6188
rect 32060 6020 32116 6030
rect 32060 5926 32116 5964
rect 32284 5346 32340 7532
rect 32620 7476 32676 7486
rect 32620 7382 32676 7420
rect 33180 7474 33236 9884
rect 33292 9884 33404 9940
rect 33292 9714 33348 9884
rect 33404 9874 33460 9884
rect 33516 9828 33572 9838
rect 33516 9734 33572 9772
rect 33292 9662 33294 9714
rect 33346 9662 33348 9714
rect 33292 9650 33348 9662
rect 33404 9604 33460 9614
rect 33404 9602 33572 9604
rect 33404 9550 33406 9602
rect 33458 9550 33572 9602
rect 33404 9548 33572 9550
rect 33404 9538 33460 9548
rect 33516 8372 33572 9548
rect 33516 8316 33796 8372
rect 33180 7422 33182 7474
rect 33234 7422 33236 7474
rect 33180 7410 33236 7422
rect 33404 8260 33460 8270
rect 33180 6690 33236 6702
rect 33180 6638 33182 6690
rect 33234 6638 33236 6690
rect 33180 6580 33236 6638
rect 33180 6514 33236 6524
rect 33404 6468 33460 8204
rect 33516 8148 33572 8158
rect 33516 6690 33572 8092
rect 33740 7474 33796 8316
rect 33852 8258 33908 8270
rect 33852 8206 33854 8258
rect 33906 8206 33908 8258
rect 33852 8148 33908 8206
rect 33852 8082 33908 8092
rect 33740 7422 33742 7474
rect 33794 7422 33796 7474
rect 33740 7410 33796 7422
rect 33516 6638 33518 6690
rect 33570 6638 33572 6690
rect 33516 6626 33572 6638
rect 33628 7362 33684 7374
rect 33628 7310 33630 7362
rect 33682 7310 33684 7362
rect 33404 6412 33572 6468
rect 33292 5794 33348 5806
rect 33292 5742 33294 5794
rect 33346 5742 33348 5794
rect 32284 5294 32286 5346
rect 32338 5294 32340 5346
rect 32284 5282 32340 5294
rect 32956 5348 33012 5358
rect 32956 5234 33012 5292
rect 32956 5182 32958 5234
rect 33010 5182 33012 5234
rect 32956 5170 33012 5182
rect 33180 5122 33236 5134
rect 33180 5070 33182 5122
rect 33234 5070 33236 5122
rect 33180 5012 33236 5070
rect 33180 4946 33236 4956
rect 32060 4900 32116 4910
rect 32060 4452 32116 4844
rect 32060 4358 32116 4396
rect 33180 4338 33236 4350
rect 33180 4286 33182 4338
rect 33234 4286 33236 4338
rect 32172 4228 32228 4238
rect 32172 3666 32228 4172
rect 33180 4004 33236 4286
rect 33180 3938 33236 3948
rect 32172 3614 32174 3666
rect 32226 3614 32228 3666
rect 32172 3602 32228 3614
rect 31948 3332 32116 3388
rect 31612 1586 31668 1596
rect 32060 800 32116 3332
rect 33292 3220 33348 5742
rect 33292 3154 33348 3164
rect 33404 4116 33460 4126
rect 33404 800 33460 4060
rect 33516 2660 33572 6412
rect 33628 3108 33684 7310
rect 33852 7028 33908 7038
rect 33852 6690 33908 6972
rect 33852 6638 33854 6690
rect 33906 6638 33908 6690
rect 33852 4340 33908 6638
rect 33964 4564 34020 10782
rect 34188 10610 34244 10622
rect 34188 10558 34190 10610
rect 34242 10558 34244 10610
rect 34188 10500 34244 10558
rect 34188 10434 34244 10444
rect 34076 9826 34132 9838
rect 34076 9774 34078 9826
rect 34130 9774 34132 9826
rect 34076 9604 34132 9774
rect 34076 9538 34132 9548
rect 34076 7812 34132 7822
rect 34076 7140 34132 7756
rect 34300 7586 34356 11116
rect 34412 9042 34468 11342
rect 34636 11620 34692 11630
rect 34636 10498 34692 11564
rect 34748 10724 34804 14252
rect 34860 14242 34916 14252
rect 35308 14306 35364 14318
rect 35308 14254 35310 14306
rect 35362 14254 35364 14306
rect 35308 13972 35364 14254
rect 35308 13906 35364 13916
rect 35308 13746 35364 13758
rect 35308 13694 35310 13746
rect 35362 13694 35364 13746
rect 35084 13634 35140 13646
rect 35084 13582 35086 13634
rect 35138 13582 35140 13634
rect 34972 13522 35028 13534
rect 34972 13470 34974 13522
rect 35026 13470 35028 13522
rect 34972 12852 35028 13470
rect 35084 13524 35140 13582
rect 35308 13524 35364 13694
rect 35532 13524 35588 15092
rect 35756 14420 35812 14430
rect 35756 14308 35812 14364
rect 35308 13522 35588 13524
rect 35308 13470 35534 13522
rect 35586 13470 35588 13522
rect 35308 13468 35588 13470
rect 35084 13458 35140 13468
rect 35532 13458 35588 13468
rect 35644 14306 35812 14308
rect 35644 14254 35758 14306
rect 35810 14254 35812 14306
rect 35644 14252 35812 14254
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 34972 12786 35028 12796
rect 35084 12628 35140 12638
rect 35084 11284 35140 12572
rect 35532 12180 35588 12190
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35532 11620 35588 12124
rect 35084 10836 35140 11228
rect 35420 11396 35476 11406
rect 35196 10836 35252 10846
rect 35084 10834 35252 10836
rect 35084 10782 35198 10834
rect 35250 10782 35252 10834
rect 35084 10780 35252 10782
rect 35196 10770 35252 10780
rect 35420 10834 35476 11340
rect 35420 10782 35422 10834
rect 35474 10782 35476 10834
rect 35420 10770 35476 10782
rect 35532 10834 35588 11564
rect 35532 10782 35534 10834
rect 35586 10782 35588 10834
rect 35532 10770 35588 10782
rect 34972 10724 35028 10734
rect 34748 10722 35028 10724
rect 34748 10670 34974 10722
rect 35026 10670 35028 10722
rect 34748 10668 35028 10670
rect 34972 10658 35028 10668
rect 34636 10446 34638 10498
rect 34690 10446 34692 10498
rect 34636 10164 34692 10446
rect 35084 10612 35140 10622
rect 35084 10164 35140 10556
rect 35308 10498 35364 10510
rect 35308 10446 35310 10498
rect 35362 10446 35364 10498
rect 35308 10388 35364 10446
rect 35644 10388 35700 14252
rect 35756 14242 35812 14252
rect 35868 13972 35924 13982
rect 35756 13634 35812 13646
rect 35756 13582 35758 13634
rect 35810 13582 35812 13634
rect 35756 13524 35812 13582
rect 35756 13458 35812 13468
rect 35308 10332 35588 10388
rect 34636 10108 35140 10164
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35084 10052 35140 10108
rect 35084 9996 35476 10052
rect 35308 9716 35364 9726
rect 35308 9622 35364 9660
rect 35196 9604 35252 9614
rect 35084 9548 35196 9604
rect 35420 9604 35476 9996
rect 35532 9826 35588 10332
rect 35532 9774 35534 9826
rect 35586 9774 35588 9826
rect 35532 9762 35588 9774
rect 35420 9548 35588 9604
rect 34412 8990 34414 9042
rect 34466 8990 34468 9042
rect 34412 8978 34468 8990
rect 34524 9268 34580 9278
rect 34300 7534 34302 7586
rect 34354 7534 34356 7586
rect 34300 7522 34356 7534
rect 34076 6692 34132 7084
rect 34076 6690 34244 6692
rect 34076 6638 34078 6690
rect 34130 6638 34244 6690
rect 34076 6636 34244 6638
rect 34076 6626 34132 6636
rect 34076 6244 34132 6254
rect 34076 6018 34132 6188
rect 34076 5966 34078 6018
rect 34130 5966 34132 6018
rect 34076 5954 34132 5966
rect 33964 4498 34020 4508
rect 34188 4450 34244 6636
rect 34524 6356 34580 9212
rect 34748 9044 34804 9054
rect 34636 8148 34692 8158
rect 34636 7474 34692 8092
rect 34636 7422 34638 7474
rect 34690 7422 34692 7474
rect 34636 6804 34692 7422
rect 34636 6738 34692 6748
rect 34748 7586 34804 8988
rect 34748 7534 34750 7586
rect 34802 7534 34804 7586
rect 34188 4398 34190 4450
rect 34242 4398 34244 4450
rect 34188 4386 34244 4398
rect 34300 6300 34580 6356
rect 34636 6578 34692 6590
rect 34636 6526 34638 6578
rect 34690 6526 34692 6578
rect 34076 4340 34132 4350
rect 33852 4338 34132 4340
rect 33852 4286 34078 4338
rect 34130 4286 34132 4338
rect 33852 4284 34132 4286
rect 34076 4274 34132 4284
rect 33740 4228 33796 4238
rect 33740 4134 33796 4172
rect 34300 3666 34356 6300
rect 34636 6020 34692 6526
rect 34636 5954 34692 5964
rect 34748 5234 34804 7534
rect 34748 5182 34750 5234
rect 34802 5182 34804 5234
rect 34748 5170 34804 5182
rect 34860 8370 34916 8382
rect 34860 8318 34862 8370
rect 34914 8318 34916 8370
rect 34748 5010 34804 5022
rect 34748 4958 34750 5010
rect 34802 4958 34804 5010
rect 34636 4788 34692 4798
rect 34748 4788 34804 4958
rect 34692 4732 34804 4788
rect 34636 4722 34692 4732
rect 34748 4564 34804 4732
rect 34860 4788 34916 8318
rect 34972 6802 35028 6814
rect 34972 6750 34974 6802
rect 35026 6750 35028 6802
rect 34972 5906 35028 6750
rect 35084 6132 35140 9548
rect 35196 9538 35252 9548
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 6132 35252 6142
rect 35084 6130 35252 6132
rect 35084 6078 35198 6130
rect 35250 6078 35252 6130
rect 35084 6076 35252 6078
rect 35196 6066 35252 6076
rect 34972 5854 34974 5906
rect 35026 5854 35028 5906
rect 34972 5842 35028 5854
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34860 4722 34916 4732
rect 35308 5236 35364 5246
rect 34860 4564 34916 4574
rect 34748 4508 34860 4564
rect 34860 4498 34916 4508
rect 34300 3614 34302 3666
rect 34354 3614 34356 3666
rect 34300 3602 34356 3614
rect 34636 4452 34692 4462
rect 34636 3388 34692 4396
rect 34972 4340 35028 4350
rect 34972 3556 35028 4284
rect 35308 4226 35364 5180
rect 35532 5010 35588 9548
rect 35644 9154 35700 10332
rect 35644 9102 35646 9154
rect 35698 9102 35700 9154
rect 35644 8260 35700 9102
rect 35644 8194 35700 8204
rect 35756 11060 35812 11070
rect 35644 7700 35700 7710
rect 35756 7700 35812 11004
rect 35868 8820 35924 13916
rect 36204 13634 36260 15092
rect 37548 14754 37604 14766
rect 37548 14702 37550 14754
rect 37602 14702 37604 14754
rect 37548 14642 37604 14702
rect 37884 14754 37940 16604
rect 38108 15426 38164 15438
rect 38108 15374 38110 15426
rect 38162 15374 38164 15426
rect 37996 15316 38052 15326
rect 37996 15222 38052 15260
rect 38108 15148 38164 15374
rect 37884 14702 37886 14754
rect 37938 14702 37940 14754
rect 37884 14690 37940 14702
rect 37996 15092 38164 15148
rect 37548 14590 37550 14642
rect 37602 14590 37604 14642
rect 37548 14578 37604 14590
rect 37100 14532 37156 14542
rect 37100 14438 37156 14476
rect 37324 14532 37380 14542
rect 37100 14308 37156 14318
rect 37100 13970 37156 14252
rect 37100 13918 37102 13970
rect 37154 13918 37156 13970
rect 37100 13906 37156 13918
rect 36204 13582 36206 13634
rect 36258 13582 36260 13634
rect 35980 12180 36036 12190
rect 36204 12180 36260 13582
rect 36652 13748 36708 13758
rect 35980 12178 36260 12180
rect 35980 12126 35982 12178
rect 36034 12126 36260 12178
rect 35980 12124 36260 12126
rect 36316 13522 36372 13534
rect 36316 13470 36318 13522
rect 36370 13470 36372 13522
rect 36316 13076 36372 13470
rect 36428 13076 36484 13086
rect 36316 13074 36484 13076
rect 36316 13022 36430 13074
rect 36482 13022 36484 13074
rect 36316 13020 36484 13022
rect 35980 12114 36036 12124
rect 35980 11508 36036 11518
rect 35980 10836 36036 11452
rect 36316 11282 36372 13020
rect 36428 13010 36484 13020
rect 36652 12964 36708 13692
rect 37100 13748 37156 13758
rect 36764 13636 36820 13646
rect 36764 13542 36820 13580
rect 36652 12402 36708 12908
rect 37100 13524 37156 13692
rect 36988 12852 37044 12862
rect 36988 12758 37044 12796
rect 36652 12350 36654 12402
rect 36706 12350 36708 12402
rect 36652 12338 36708 12350
rect 36988 12178 37044 12190
rect 36988 12126 36990 12178
rect 37042 12126 37044 12178
rect 36540 12068 36596 12078
rect 36316 11230 36318 11282
rect 36370 11230 36372 11282
rect 36316 11218 36372 11230
rect 36428 11282 36484 11294
rect 36428 11230 36430 11282
rect 36482 11230 36484 11282
rect 36092 11172 36148 11182
rect 36092 11078 36148 11116
rect 35980 10780 36148 10836
rect 35980 10610 36036 10622
rect 35980 10558 35982 10610
rect 36034 10558 36036 10610
rect 35980 10052 36036 10558
rect 35980 9986 36036 9996
rect 35868 8754 35924 8764
rect 35644 7698 35812 7700
rect 35644 7646 35646 7698
rect 35698 7646 35812 7698
rect 35644 7644 35812 7646
rect 35644 7634 35700 7644
rect 36092 6578 36148 10780
rect 36316 10500 36372 10510
rect 36316 9826 36372 10444
rect 36316 9774 36318 9826
rect 36370 9774 36372 9826
rect 36316 9762 36372 9774
rect 36204 9604 36260 9614
rect 36204 9602 36372 9604
rect 36204 9550 36206 9602
rect 36258 9550 36372 9602
rect 36204 9548 36372 9550
rect 36204 9538 36260 9548
rect 36204 8146 36260 8158
rect 36204 8094 36206 8146
rect 36258 8094 36260 8146
rect 36204 7028 36260 8094
rect 36316 7252 36372 9548
rect 36428 9492 36484 11230
rect 36540 10836 36596 12012
rect 36988 11844 37044 12126
rect 36988 11778 37044 11788
rect 36988 11172 37044 11182
rect 37100 11172 37156 13468
rect 37212 12962 37268 12974
rect 37212 12910 37214 12962
rect 37266 12910 37268 12962
rect 37212 11844 37268 12910
rect 37324 12628 37380 14476
rect 37436 14308 37492 14318
rect 37436 13746 37492 14252
rect 37436 13694 37438 13746
rect 37490 13694 37492 13746
rect 37436 13524 37492 13694
rect 37436 13458 37492 13468
rect 37548 13636 37604 13646
rect 37324 12572 37492 12628
rect 37212 11778 37268 11788
rect 37324 12404 37380 12414
rect 37324 12290 37380 12348
rect 37324 12238 37326 12290
rect 37378 12238 37380 12290
rect 37324 11282 37380 12238
rect 37324 11230 37326 11282
rect 37378 11230 37380 11282
rect 37324 11218 37380 11230
rect 36988 11170 37156 11172
rect 36988 11118 36990 11170
rect 37042 11118 37156 11170
rect 36988 11116 37156 11118
rect 36988 10948 37044 11116
rect 36988 10882 37044 10892
rect 36540 10610 36596 10780
rect 36540 10558 36542 10610
rect 36594 10558 36596 10610
rect 36540 10546 36596 10558
rect 36988 10500 37044 10510
rect 37436 10500 37492 12572
rect 37548 11060 37604 13580
rect 37772 12962 37828 12974
rect 37772 12910 37774 12962
rect 37826 12910 37828 12962
rect 37772 12402 37828 12910
rect 37772 12350 37774 12402
rect 37826 12350 37828 12402
rect 37772 12338 37828 12350
rect 37884 12852 37940 12862
rect 37884 12290 37940 12796
rect 37884 12238 37886 12290
rect 37938 12238 37940 12290
rect 37884 12226 37940 12238
rect 37660 12180 37716 12190
rect 37660 12086 37716 12124
rect 37996 11396 38052 15092
rect 38108 14306 38164 14318
rect 38108 14254 38110 14306
rect 38162 14254 38164 14306
rect 38108 13748 38164 14254
rect 38220 13972 38276 16604
rect 38332 16324 38388 16830
rect 38668 16884 38724 16894
rect 38668 16790 38724 16828
rect 38892 16772 38948 16942
rect 39004 16994 39060 17276
rect 39004 16942 39006 16994
rect 39058 16942 39060 16994
rect 39004 16930 39060 16942
rect 39900 16772 39956 19180
rect 38892 16716 39956 16772
rect 38332 15764 38388 16268
rect 39900 16210 39956 16716
rect 39900 16158 39902 16210
rect 39954 16158 39956 16210
rect 39900 16146 39956 16158
rect 38332 15698 38388 15708
rect 38332 15540 38388 15550
rect 38332 15446 38388 15484
rect 39004 15204 39060 15242
rect 39004 15138 39060 15148
rect 39452 15202 39508 15214
rect 39452 15150 39454 15202
rect 39506 15150 39508 15202
rect 38332 14754 38388 14766
rect 38332 14702 38334 14754
rect 38386 14702 38388 14754
rect 38332 14196 38388 14702
rect 39004 14754 39060 14766
rect 39004 14702 39006 14754
rect 39058 14702 39060 14754
rect 39004 14642 39060 14702
rect 39004 14590 39006 14642
rect 39058 14590 39060 14642
rect 39004 14578 39060 14590
rect 39340 14754 39396 14766
rect 39340 14702 39342 14754
rect 39394 14702 39396 14754
rect 38444 14420 38500 14430
rect 38444 14326 38500 14364
rect 39340 14308 39396 14702
rect 39452 14532 39508 15150
rect 39788 14754 39844 14766
rect 39788 14702 39790 14754
rect 39842 14702 39844 14754
rect 39452 14476 39620 14532
rect 39452 14308 39508 14318
rect 39340 14306 39508 14308
rect 39340 14254 39454 14306
rect 39506 14254 39508 14306
rect 39340 14252 39508 14254
rect 39452 14242 39508 14252
rect 39564 14308 39620 14476
rect 38332 14140 38500 14196
rect 38220 13906 38276 13916
rect 38108 13682 38164 13692
rect 38220 13634 38276 13646
rect 38220 13582 38222 13634
rect 38274 13582 38276 13634
rect 38108 13188 38164 13198
rect 38108 12962 38164 13132
rect 38220 13074 38276 13582
rect 38220 13022 38222 13074
rect 38274 13022 38276 13074
rect 38220 13010 38276 13022
rect 38108 12910 38110 12962
rect 38162 12910 38164 12962
rect 38108 12898 38164 12910
rect 38332 12964 38388 12974
rect 38332 12870 38388 12908
rect 37996 11330 38052 11340
rect 37660 11284 37716 11294
rect 37660 11190 37716 11228
rect 37548 10834 37604 11004
rect 37548 10782 37550 10834
rect 37602 10782 37604 10834
rect 37548 10770 37604 10782
rect 37996 11170 38052 11182
rect 37996 11118 37998 11170
rect 38050 11118 38052 11170
rect 37996 10612 38052 11118
rect 38332 11170 38388 11182
rect 38332 11118 38334 11170
rect 38386 11118 38388 11170
rect 38332 10948 38388 11118
rect 38332 10882 38388 10892
rect 36988 10406 37044 10444
rect 37212 10444 37492 10500
rect 37548 10556 37828 10612
rect 37996 10556 38388 10612
rect 37100 10052 37156 10062
rect 36428 9426 36484 9436
rect 36988 9602 37044 9614
rect 36988 9550 36990 9602
rect 37042 9550 37044 9602
rect 36988 9492 37044 9550
rect 36988 9426 37044 9436
rect 37100 9268 37156 9996
rect 36988 9212 37156 9268
rect 36988 8484 37044 9212
rect 37212 8484 37268 10444
rect 37548 10052 37604 10556
rect 37772 10388 37828 10556
rect 37884 10388 37940 10398
rect 37772 10386 38164 10388
rect 37772 10334 37886 10386
rect 37938 10334 38164 10386
rect 37772 10332 38164 10334
rect 37884 10322 37940 10332
rect 37324 9996 37604 10052
rect 37324 9826 37380 9996
rect 37324 9774 37326 9826
rect 37378 9774 37380 9826
rect 37324 9762 37380 9774
rect 37660 9826 37716 9838
rect 37660 9774 37662 9826
rect 37714 9774 37716 9826
rect 37548 9716 37604 9726
rect 37660 9716 37716 9774
rect 38108 9826 38164 10332
rect 38108 9774 38110 9826
rect 38162 9774 38164 9826
rect 38108 9762 38164 9774
rect 38220 10386 38276 10398
rect 38220 10334 38222 10386
rect 38274 10334 38276 10386
rect 37604 9660 37716 9716
rect 37772 9716 37828 9726
rect 37548 9650 37604 9660
rect 37212 8428 37380 8484
rect 36988 7588 37044 8428
rect 37100 8372 37156 8382
rect 37100 8278 37156 8316
rect 37212 8258 37268 8270
rect 37212 8206 37214 8258
rect 37266 8206 37268 8258
rect 37212 8148 37268 8206
rect 37212 8082 37268 8092
rect 37212 7588 37268 7598
rect 36988 7586 37268 7588
rect 36988 7534 37214 7586
rect 37266 7534 37268 7586
rect 36988 7532 37268 7534
rect 37212 7522 37268 7532
rect 36316 7196 36820 7252
rect 36204 6972 36708 7028
rect 36092 6526 36094 6578
rect 36146 6526 36148 6578
rect 35532 4958 35534 5010
rect 35586 4958 35588 5010
rect 35532 4946 35588 4958
rect 35756 5908 35812 5918
rect 35756 5122 35812 5852
rect 35756 5070 35758 5122
rect 35810 5070 35812 5122
rect 35308 4174 35310 4226
rect 35362 4174 35364 4226
rect 35308 4162 35364 4174
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34972 3462 35028 3500
rect 34636 3332 34804 3388
rect 33628 3042 33684 3052
rect 33516 2594 33572 2604
rect 34748 800 34804 3332
rect 35756 1092 35812 5070
rect 36092 5012 36148 6526
rect 36428 6804 36484 6814
rect 36428 5908 36484 6748
rect 36428 5906 36596 5908
rect 36428 5854 36430 5906
rect 36482 5854 36596 5906
rect 36428 5852 36596 5854
rect 36428 5842 36484 5852
rect 36092 4946 36148 4956
rect 36316 4340 36372 4350
rect 36540 4340 36596 5852
rect 36652 5348 36708 6972
rect 36764 5684 36820 7196
rect 37324 6244 37380 8428
rect 37660 8372 37716 8382
rect 37436 8260 37492 8270
rect 37436 8258 37604 8260
rect 37436 8206 37438 8258
rect 37490 8206 37604 8258
rect 37436 8204 37604 8206
rect 37436 8194 37492 8204
rect 37548 6692 37604 8204
rect 37660 6804 37716 8316
rect 37772 8370 37828 9660
rect 37772 8318 37774 8370
rect 37826 8318 37828 8370
rect 37772 8306 37828 8318
rect 37884 8820 37940 8830
rect 37660 6738 37716 6748
rect 37548 6626 37604 6636
rect 37436 6578 37492 6590
rect 37436 6526 37438 6578
rect 37490 6526 37492 6578
rect 37436 6468 37492 6526
rect 37436 6402 37492 6412
rect 36988 5796 37044 5806
rect 37324 5796 37380 6188
rect 37548 6020 37604 6030
rect 37548 5926 37604 5964
rect 37884 5906 37940 8764
rect 38220 8596 38276 10334
rect 38332 9828 38388 10556
rect 38444 10498 38500 14140
rect 39452 14084 39508 14094
rect 38780 13188 38836 13198
rect 38780 13074 38836 13132
rect 38780 13022 38782 13074
rect 38834 13022 38836 13074
rect 38780 13010 38836 13022
rect 39116 13186 39172 13198
rect 39116 13134 39118 13186
rect 39170 13134 39172 13186
rect 38780 12068 38836 12078
rect 38780 12066 38948 12068
rect 38780 12014 38782 12066
rect 38834 12014 38948 12066
rect 38780 12012 38948 12014
rect 38780 12002 38836 12012
rect 38444 10446 38446 10498
rect 38498 10446 38500 10498
rect 38444 10276 38500 10446
rect 38444 10210 38500 10220
rect 38556 11396 38612 11406
rect 38556 10052 38612 11340
rect 38668 11170 38724 11182
rect 38668 11118 38670 11170
rect 38722 11118 38724 11170
rect 38668 10612 38724 11118
rect 38780 10948 38836 10958
rect 38892 10948 38948 12012
rect 39004 11284 39060 11294
rect 39004 11190 39060 11228
rect 39116 11282 39172 13134
rect 39340 12740 39396 12750
rect 39116 11230 39118 11282
rect 39170 11230 39172 11282
rect 39116 11218 39172 11230
rect 39228 12738 39396 12740
rect 39228 12686 39342 12738
rect 39394 12686 39396 12738
rect 39228 12684 39396 12686
rect 39228 12180 39284 12684
rect 39340 12674 39396 12684
rect 38892 10892 39060 10948
rect 38780 10722 38836 10892
rect 38780 10670 38782 10722
rect 38834 10670 38836 10722
rect 38780 10658 38836 10670
rect 38892 10722 38948 10734
rect 38892 10670 38894 10722
rect 38946 10670 38948 10722
rect 38668 10546 38724 10556
rect 38892 10500 38948 10670
rect 38332 9156 38388 9772
rect 38332 9090 38388 9100
rect 38444 9996 38612 10052
rect 38780 10444 38948 10500
rect 38220 8530 38276 8540
rect 38444 8372 38500 9996
rect 38556 9828 38612 9838
rect 38556 9604 38612 9772
rect 38668 9716 38724 9726
rect 38668 9622 38724 9660
rect 38556 9538 38612 9548
rect 38668 9156 38724 9166
rect 38668 9062 38724 9100
rect 38556 8372 38612 8382
rect 38444 8370 38612 8372
rect 38444 8318 38558 8370
rect 38610 8318 38612 8370
rect 38444 8316 38612 8318
rect 38556 8306 38612 8316
rect 37884 5854 37886 5906
rect 37938 5854 37940 5906
rect 37884 5842 37940 5854
rect 38108 8146 38164 8158
rect 38108 8094 38110 8146
rect 38162 8094 38164 8146
rect 38108 6580 38164 8094
rect 38220 8036 38276 8046
rect 38220 8034 38388 8036
rect 38220 7982 38222 8034
rect 38274 7982 38388 8034
rect 38220 7980 38388 7982
rect 38220 7970 38276 7980
rect 37044 5740 37268 5796
rect 36988 5730 37044 5740
rect 36764 5618 36820 5628
rect 36876 5348 36932 5358
rect 36652 5346 36932 5348
rect 36652 5294 36878 5346
rect 36930 5294 36932 5346
rect 36652 5292 36932 5294
rect 36876 5282 36932 5292
rect 37212 5236 37268 5740
rect 37324 5730 37380 5740
rect 37996 5796 38052 5806
rect 38108 5796 38164 6524
rect 37996 5794 38164 5796
rect 37996 5742 37998 5794
rect 38050 5742 38164 5794
rect 37996 5740 38164 5742
rect 38220 6020 38276 6030
rect 37996 5730 38052 5740
rect 36316 4338 36596 4340
rect 36316 4286 36318 4338
rect 36370 4286 36596 4338
rect 36316 4284 36596 4286
rect 36876 4900 36932 4910
rect 36316 4228 36372 4284
rect 36316 4162 36372 4172
rect 36204 3668 36260 3678
rect 35980 3556 36036 3566
rect 35980 3462 36036 3500
rect 36204 1652 36260 3612
rect 36764 3668 36820 3678
rect 36876 3668 36932 4844
rect 37212 4452 37268 5180
rect 37436 5012 37492 5022
rect 37324 4452 37380 4462
rect 37212 4450 37380 4452
rect 37212 4398 37326 4450
rect 37378 4398 37380 4450
rect 37212 4396 37380 4398
rect 37324 4386 37380 4396
rect 36764 3666 36932 3668
rect 36764 3614 36766 3666
rect 36818 3614 36932 3666
rect 36764 3612 36932 3614
rect 36764 3602 36820 3612
rect 35756 1026 35812 1036
rect 36092 1596 36260 1652
rect 36092 800 36148 1596
rect 37436 800 37492 4956
rect 38220 4338 38276 5964
rect 38332 5908 38388 7980
rect 38444 7476 38500 7486
rect 38444 7474 38612 7476
rect 38444 7422 38446 7474
rect 38498 7422 38612 7474
rect 38444 7420 38612 7422
rect 38444 7410 38500 7420
rect 38444 6802 38500 6814
rect 38444 6750 38446 6802
rect 38498 6750 38500 6802
rect 38444 6132 38500 6750
rect 38556 6692 38612 7420
rect 38612 6636 38724 6692
rect 38556 6626 38612 6636
rect 38444 6076 38612 6132
rect 38332 5842 38388 5852
rect 38444 5906 38500 5918
rect 38444 5854 38446 5906
rect 38498 5854 38500 5906
rect 38444 5796 38500 5854
rect 38332 5236 38388 5246
rect 38332 4450 38388 5180
rect 38332 4398 38334 4450
rect 38386 4398 38388 4450
rect 38332 4386 38388 4398
rect 38220 4286 38222 4338
rect 38274 4286 38276 4338
rect 38220 4274 38276 4286
rect 38444 2548 38500 5740
rect 38556 3556 38612 6076
rect 38668 4562 38724 6636
rect 38668 4510 38670 4562
rect 38722 4510 38724 4562
rect 38668 4498 38724 4510
rect 38780 3668 38836 10444
rect 39004 9044 39060 10892
rect 38892 8988 39060 9044
rect 39116 10610 39172 10622
rect 39116 10558 39118 10610
rect 39170 10558 39172 10610
rect 38892 7364 38948 8988
rect 39004 8818 39060 8830
rect 39004 8766 39006 8818
rect 39058 8766 39060 8818
rect 39004 8596 39060 8766
rect 39004 8530 39060 8540
rect 39116 8484 39172 10558
rect 39228 9604 39284 12124
rect 39452 12066 39508 14028
rect 39564 13972 39620 14252
rect 39564 13906 39620 13916
rect 39676 14196 39732 14206
rect 39676 13186 39732 14140
rect 39676 13134 39678 13186
rect 39730 13134 39732 13186
rect 39676 13074 39732 13134
rect 39676 13022 39678 13074
rect 39730 13022 39732 13074
rect 39676 13010 39732 13022
rect 39788 12180 39844 14702
rect 39900 14306 39956 14318
rect 39900 14254 39902 14306
rect 39954 14254 39956 14306
rect 39900 14084 39956 14254
rect 39900 14018 39956 14028
rect 39900 12404 39956 12414
rect 40012 12404 40068 20188
rect 40236 19572 40292 19582
rect 40236 18338 40292 19516
rect 40796 19346 40852 22988
rect 41468 22708 41524 23102
rect 41468 22642 41524 22652
rect 41692 21586 41748 25454
rect 42252 23828 42308 23838
rect 41916 23492 41972 23502
rect 41804 23154 41860 23166
rect 41804 23102 41806 23154
rect 41858 23102 41860 23154
rect 41804 23044 41860 23102
rect 41804 22978 41860 22988
rect 41916 22932 41972 23436
rect 42028 23380 42084 23390
rect 42028 23286 42084 23324
rect 42140 23268 42196 23306
rect 42140 23202 42196 23212
rect 41916 22866 41972 22876
rect 41692 21534 41694 21586
rect 41746 21534 41748 21586
rect 41468 21476 41524 21486
rect 41468 21382 41524 21420
rect 41692 20916 41748 21534
rect 41692 20850 41748 20860
rect 41916 22484 41972 22494
rect 41804 20802 41860 20814
rect 41804 20750 41806 20802
rect 41858 20750 41860 20802
rect 41804 20132 41860 20750
rect 41356 20076 41860 20132
rect 41020 20018 41076 20030
rect 41020 19966 41022 20018
rect 41074 19966 41076 20018
rect 41020 19572 41076 19966
rect 41020 19506 41076 19516
rect 40796 19294 40798 19346
rect 40850 19294 40852 19346
rect 40796 19282 40852 19294
rect 41356 19236 41412 20076
rect 41132 19234 41412 19236
rect 41132 19182 41358 19234
rect 41410 19182 41412 19234
rect 41132 19180 41412 19182
rect 41020 18452 41076 18462
rect 40236 18286 40238 18338
rect 40290 18286 40292 18338
rect 40236 18274 40292 18286
rect 40908 18396 41020 18452
rect 40236 17556 40292 17566
rect 40236 16098 40292 17500
rect 40908 16884 40964 18396
rect 41020 18386 41076 18396
rect 41020 17556 41076 17566
rect 41020 17462 41076 17500
rect 41132 17554 41188 19180
rect 41356 19170 41412 19180
rect 41580 19906 41636 19918
rect 41580 19854 41582 19906
rect 41634 19854 41636 19906
rect 41580 19124 41636 19854
rect 41580 17668 41636 19068
rect 41692 18228 41748 20076
rect 41916 18676 41972 22428
rect 42252 22148 42308 23772
rect 42588 23828 42644 23838
rect 42364 23268 42420 23278
rect 42364 23174 42420 23212
rect 42588 23042 42644 23772
rect 42588 22990 42590 23042
rect 42642 22990 42644 23042
rect 42588 22978 42644 22990
rect 42700 22820 42756 26236
rect 42812 26226 42868 26236
rect 42924 26292 42980 26302
rect 42924 26290 43204 26292
rect 42924 26238 42926 26290
rect 42978 26238 43204 26290
rect 42924 26236 43204 26238
rect 42924 26226 42980 26236
rect 43148 25396 43204 26236
rect 43148 24948 43204 25340
rect 43260 24948 43316 24958
rect 43148 24946 43316 24948
rect 43148 24894 43262 24946
rect 43314 24894 43316 24946
rect 43148 24892 43316 24894
rect 43260 24882 43316 24892
rect 43372 24834 43428 28812
rect 44156 28084 44212 29484
rect 45164 29428 45220 29438
rect 44828 28532 44884 28542
rect 44716 28530 44884 28532
rect 44716 28478 44830 28530
rect 44882 28478 44884 28530
rect 44716 28476 44884 28478
rect 44156 28082 44660 28084
rect 44156 28030 44158 28082
rect 44210 28030 44660 28082
rect 44156 28028 44660 28030
rect 44156 28018 44212 28028
rect 44604 27858 44660 28028
rect 44716 28082 44772 28476
rect 44828 28466 44884 28476
rect 45164 28530 45220 29372
rect 46060 29316 46116 30158
rect 46732 30098 46788 30110
rect 46732 30046 46734 30098
rect 46786 30046 46788 30098
rect 46172 29428 46228 29438
rect 46172 29334 46228 29372
rect 46060 29250 46116 29260
rect 45164 28478 45166 28530
rect 45218 28478 45220 28530
rect 45164 28466 45220 28478
rect 46732 28420 46788 30046
rect 46732 28354 46788 28364
rect 44716 28030 44718 28082
rect 44770 28030 44772 28082
rect 44716 28018 44772 28030
rect 46060 27972 46116 27982
rect 44604 27806 44606 27858
rect 44658 27806 44660 27858
rect 44604 27794 44660 27806
rect 45276 27858 45332 27870
rect 45276 27806 45278 27858
rect 45330 27806 45332 27858
rect 45052 27748 45108 27758
rect 45052 27654 45108 27692
rect 44828 27636 44884 27646
rect 44828 27542 44884 27580
rect 45052 27412 45108 27422
rect 45052 27188 45108 27356
rect 44492 27186 45108 27188
rect 44492 27134 45054 27186
rect 45106 27134 45108 27186
rect 44492 27132 45108 27134
rect 43596 26402 43652 26414
rect 43596 26350 43598 26402
rect 43650 26350 43652 26402
rect 43596 26292 43652 26350
rect 43596 26226 43652 26236
rect 44268 26292 44324 26302
rect 44492 26292 44548 27132
rect 45052 27122 45108 27132
rect 44268 26198 44324 26236
rect 44380 26290 44548 26292
rect 44380 26238 44494 26290
rect 44546 26238 44548 26290
rect 44380 26236 44548 26238
rect 44380 25956 44436 26236
rect 44492 26226 44548 26236
rect 44604 26292 44660 26302
rect 43932 25900 44436 25956
rect 43484 25620 43540 25630
rect 43932 25620 43988 25900
rect 43484 25618 43988 25620
rect 43484 25566 43486 25618
rect 43538 25566 43988 25618
rect 43484 25564 43988 25566
rect 43484 25554 43540 25564
rect 43932 25506 43988 25564
rect 43932 25454 43934 25506
rect 43986 25454 43988 25506
rect 43932 25442 43988 25454
rect 44044 25732 44100 25742
rect 43596 25396 43652 25406
rect 43820 25396 43876 25406
rect 43596 25394 43764 25396
rect 43596 25342 43598 25394
rect 43650 25342 43764 25394
rect 43596 25340 43764 25342
rect 43596 25330 43652 25340
rect 43708 25284 43764 25340
rect 43820 25302 43876 25340
rect 43708 25218 43764 25228
rect 43372 24782 43374 24834
rect 43426 24782 43428 24834
rect 43036 24724 43092 24734
rect 43372 24724 43428 24782
rect 43036 24722 43428 24724
rect 43036 24670 43038 24722
rect 43090 24670 43428 24722
rect 43036 24668 43428 24670
rect 44044 24722 44100 25676
rect 44604 25396 44660 26236
rect 44716 26180 44772 26190
rect 44716 25506 44772 26124
rect 44828 26066 44884 26078
rect 44828 26014 44830 26066
rect 44882 26014 44884 26066
rect 44828 25732 44884 26014
rect 45164 26066 45220 26078
rect 45164 26014 45166 26066
rect 45218 26014 45220 26066
rect 45164 25956 45220 26014
rect 44828 25666 44884 25676
rect 44940 25900 45164 25956
rect 44716 25454 44718 25506
rect 44770 25454 44772 25506
rect 44716 25442 44772 25454
rect 44604 25330 44660 25340
rect 44044 24670 44046 24722
rect 44098 24670 44100 24722
rect 43036 24658 43092 24668
rect 43148 24052 43204 24668
rect 44044 24658 44100 24670
rect 44492 24724 44548 24734
rect 44940 24724 44996 25900
rect 45164 25890 45220 25900
rect 45276 25620 45332 27806
rect 45724 27746 45780 27758
rect 45724 27694 45726 27746
rect 45778 27694 45780 27746
rect 45724 27636 45780 27694
rect 45724 27188 45780 27580
rect 45724 27122 45780 27132
rect 45948 27636 46004 27646
rect 45948 27074 46004 27580
rect 45948 27022 45950 27074
rect 46002 27022 46004 27074
rect 45836 26964 45892 26974
rect 45388 26628 45444 26638
rect 45388 26178 45444 26572
rect 45500 26292 45556 26302
rect 45500 26290 45668 26292
rect 45500 26238 45502 26290
rect 45554 26238 45668 26290
rect 45500 26236 45668 26238
rect 45500 26226 45556 26236
rect 45388 26126 45390 26178
rect 45442 26126 45444 26178
rect 45388 26114 45444 26126
rect 45612 26068 45668 26236
rect 45724 26068 45780 26078
rect 45612 26066 45780 26068
rect 45612 26014 45726 26066
rect 45778 26014 45780 26066
rect 45612 26012 45780 26014
rect 45724 26002 45780 26012
rect 45276 25554 45332 25564
rect 45836 25618 45892 26908
rect 45836 25566 45838 25618
rect 45890 25566 45892 25618
rect 45836 25554 45892 25566
rect 45388 25508 45444 25518
rect 45388 25414 45444 25452
rect 45164 25394 45220 25406
rect 45164 25342 45166 25394
rect 45218 25342 45220 25394
rect 45052 25282 45108 25294
rect 45052 25230 45054 25282
rect 45106 25230 45108 25282
rect 45052 24948 45108 25230
rect 45164 25284 45220 25342
rect 45164 25218 45220 25228
rect 45052 24882 45108 24892
rect 45500 24836 45556 24846
rect 45052 24724 45108 24734
rect 44492 24722 45108 24724
rect 44492 24670 44494 24722
rect 44546 24670 45054 24722
rect 45106 24670 45108 24722
rect 44492 24668 45108 24670
rect 44492 24658 44548 24668
rect 45052 24658 45108 24668
rect 43820 24498 43876 24510
rect 43820 24446 43822 24498
rect 43874 24446 43876 24498
rect 43596 24052 43652 24062
rect 43148 24050 43652 24052
rect 43148 23998 43598 24050
rect 43650 23998 43652 24050
rect 43148 23996 43652 23998
rect 43148 23938 43204 23996
rect 43596 23986 43652 23996
rect 43820 24052 43876 24446
rect 43820 23986 43876 23996
rect 44492 24498 44548 24510
rect 44492 24446 44494 24498
rect 44546 24446 44548 24498
rect 43148 23886 43150 23938
rect 43202 23886 43204 23938
rect 43148 23874 43204 23886
rect 44492 23940 44548 24446
rect 44492 23874 44548 23884
rect 44604 24498 44660 24510
rect 44604 24446 44606 24498
rect 44658 24446 44660 24498
rect 44604 23828 44660 24446
rect 44828 24388 44884 24398
rect 44604 23762 44660 23772
rect 44716 24332 44828 24388
rect 42812 23714 42868 23726
rect 42812 23662 42814 23714
rect 42866 23662 42868 23714
rect 42812 23604 42868 23662
rect 42812 23538 42868 23548
rect 43372 23604 43428 23614
rect 43372 23378 43428 23548
rect 43372 23326 43374 23378
rect 43426 23326 43428 23378
rect 43372 23314 43428 23326
rect 43708 23492 43764 23502
rect 43708 23378 43764 23436
rect 44604 23380 44660 23390
rect 44716 23380 44772 24332
rect 44828 24322 44884 24332
rect 45388 24052 45444 24062
rect 45276 23996 45388 24052
rect 45164 23828 45220 23838
rect 43708 23326 43710 23378
rect 43762 23326 43764 23378
rect 43708 23314 43764 23326
rect 44156 23378 44772 23380
rect 44156 23326 44606 23378
rect 44658 23326 44772 23378
rect 44156 23324 44772 23326
rect 45052 23492 45108 23502
rect 45052 23378 45108 23436
rect 45052 23326 45054 23378
rect 45106 23326 45108 23378
rect 44156 23266 44212 23324
rect 44604 23314 44660 23324
rect 44156 23214 44158 23266
rect 44210 23214 44212 23266
rect 44156 23202 44212 23214
rect 43484 23156 43540 23166
rect 42588 22764 42756 22820
rect 43260 23154 43540 23156
rect 43260 23102 43486 23154
rect 43538 23102 43540 23154
rect 43260 23100 43540 23102
rect 42588 22708 42644 22764
rect 42588 22370 42644 22652
rect 42700 22596 42756 22606
rect 42700 22482 42756 22540
rect 42700 22430 42702 22482
rect 42754 22430 42756 22482
rect 42700 22418 42756 22430
rect 42588 22318 42590 22370
rect 42642 22318 42644 22370
rect 42588 22306 42644 22318
rect 43148 22258 43204 22270
rect 43148 22206 43150 22258
rect 43202 22206 43204 22258
rect 42364 22148 42420 22158
rect 42252 22146 42420 22148
rect 42252 22094 42366 22146
rect 42418 22094 42420 22146
rect 42252 22092 42420 22094
rect 42364 21700 42420 22092
rect 42812 22146 42868 22158
rect 42812 22094 42814 22146
rect 42866 22094 42868 22146
rect 42700 21700 42756 21710
rect 42364 21698 42756 21700
rect 42364 21646 42702 21698
rect 42754 21646 42756 21698
rect 42364 21644 42756 21646
rect 42700 21634 42756 21644
rect 42028 21588 42084 21598
rect 42028 21494 42084 21532
rect 42700 21362 42756 21374
rect 42700 21310 42702 21362
rect 42754 21310 42756 21362
rect 42028 20914 42084 20926
rect 42028 20862 42030 20914
rect 42082 20862 42084 20914
rect 42028 19572 42084 20862
rect 42700 20802 42756 21310
rect 42700 20750 42702 20802
rect 42754 20750 42756 20802
rect 42700 20738 42756 20750
rect 42812 20244 42868 22094
rect 42924 21698 42980 21710
rect 42924 21646 42926 21698
rect 42978 21646 42980 21698
rect 42924 21476 42980 21646
rect 43036 21476 43092 21486
rect 42924 21474 43092 21476
rect 42924 21422 43038 21474
rect 43090 21422 43092 21474
rect 42924 21420 43092 21422
rect 42028 19506 42084 19516
rect 42700 20188 42868 20244
rect 41804 18620 41972 18676
rect 42140 19460 42196 19470
rect 41804 18452 41860 18620
rect 41804 18386 41860 18396
rect 42140 18450 42196 19404
rect 42364 19348 42420 19358
rect 42364 18676 42420 19292
rect 42140 18398 42142 18450
rect 42194 18398 42196 18450
rect 41916 18340 41972 18350
rect 41916 18228 41972 18284
rect 41692 18172 41972 18228
rect 41916 17890 41972 18172
rect 41916 17838 41918 17890
rect 41970 17838 41972 17890
rect 41916 17826 41972 17838
rect 42140 17890 42196 18398
rect 42140 17838 42142 17890
rect 42194 17838 42196 17890
rect 42140 17826 42196 17838
rect 42252 18620 42420 18676
rect 42588 18676 42644 18686
rect 42252 17890 42308 18620
rect 42588 18450 42644 18620
rect 42588 18398 42590 18450
rect 42642 18398 42644 18450
rect 42588 18386 42644 18398
rect 42700 18338 42756 20188
rect 42812 19124 42868 19134
rect 42812 19030 42868 19068
rect 43036 18900 43092 21420
rect 43148 21362 43204 22206
rect 43148 21310 43150 21362
rect 43202 21310 43204 21362
rect 43148 21298 43204 21310
rect 43260 19796 43316 23100
rect 43484 23090 43540 23100
rect 43932 23154 43988 23166
rect 43932 23102 43934 23154
rect 43986 23102 43988 23154
rect 43484 22932 43540 22942
rect 43372 22260 43428 22270
rect 43372 22146 43428 22204
rect 43372 22094 43374 22146
rect 43426 22094 43428 22146
rect 43372 22082 43428 22094
rect 43484 22258 43540 22876
rect 43708 22708 43764 22718
rect 43708 22370 43764 22652
rect 43708 22318 43710 22370
rect 43762 22318 43764 22370
rect 43708 22306 43764 22318
rect 43484 22206 43486 22258
rect 43538 22206 43540 22258
rect 43484 21810 43540 22206
rect 43484 21758 43486 21810
rect 43538 21758 43540 21810
rect 43484 21746 43540 21758
rect 43932 21252 43988 23102
rect 45052 22370 45108 23326
rect 45164 23378 45220 23772
rect 45164 23326 45166 23378
rect 45218 23326 45220 23378
rect 45164 23314 45220 23326
rect 45276 23380 45332 23996
rect 45388 23986 45444 23996
rect 45388 23826 45444 23838
rect 45388 23774 45390 23826
rect 45442 23774 45444 23826
rect 45388 23604 45444 23774
rect 45500 23826 45556 24780
rect 45948 24164 46004 27022
rect 46060 26514 46116 27916
rect 46172 27748 46228 27758
rect 46172 27076 46228 27692
rect 46172 26962 46228 27020
rect 46172 26910 46174 26962
rect 46226 26910 46228 26962
rect 46172 26898 46228 26910
rect 46732 27188 46788 27198
rect 46060 26462 46062 26514
rect 46114 26462 46116 26514
rect 46060 26066 46116 26462
rect 46060 26014 46062 26066
rect 46114 26014 46116 26066
rect 46060 26002 46116 26014
rect 46508 26178 46564 26190
rect 46508 26126 46510 26178
rect 46562 26126 46564 26178
rect 46508 25956 46564 26126
rect 46508 25890 46564 25900
rect 46396 25284 46452 25294
rect 46620 25284 46676 25294
rect 46396 25282 46564 25284
rect 46396 25230 46398 25282
rect 46450 25230 46564 25282
rect 46396 25228 46564 25230
rect 46396 25218 46452 25228
rect 46396 24948 46452 24958
rect 46396 24854 46452 24892
rect 46508 24836 46564 25228
rect 46620 24946 46676 25228
rect 46620 24894 46622 24946
rect 46674 24894 46676 24946
rect 46620 24882 46676 24894
rect 46508 24770 46564 24780
rect 45500 23774 45502 23826
rect 45554 23774 45556 23826
rect 45500 23762 45556 23774
rect 45612 24108 46004 24164
rect 46508 24610 46564 24622
rect 46508 24558 46510 24610
rect 46562 24558 46564 24610
rect 45388 23538 45444 23548
rect 45276 23324 45556 23380
rect 45276 23156 45332 23166
rect 45276 23062 45332 23100
rect 45052 22318 45054 22370
rect 45106 22318 45108 22370
rect 45052 22306 45108 22318
rect 45388 22148 45444 22158
rect 45388 22054 45444 22092
rect 43932 21186 43988 21196
rect 44044 21474 44100 21486
rect 44044 21422 44046 21474
rect 44098 21422 44100 21474
rect 44044 20692 44100 21422
rect 44044 20626 44100 20636
rect 44268 20804 44324 20814
rect 44268 20130 44324 20748
rect 45052 20804 45108 20814
rect 45388 20804 45444 20814
rect 45052 20802 45444 20804
rect 45052 20750 45054 20802
rect 45106 20750 45390 20802
rect 45442 20750 45444 20802
rect 45052 20748 45444 20750
rect 45052 20738 45108 20748
rect 45388 20692 45444 20748
rect 45388 20626 45444 20636
rect 44268 20078 44270 20130
rect 44322 20078 44324 20130
rect 44268 20066 44324 20078
rect 43708 20018 43764 20030
rect 43708 19966 43710 20018
rect 43762 19966 43764 20018
rect 43148 19740 43316 19796
rect 43372 19906 43428 19918
rect 43372 19854 43374 19906
rect 43426 19854 43428 19906
rect 43148 19124 43204 19740
rect 43260 19572 43316 19582
rect 43260 19458 43316 19516
rect 43260 19406 43262 19458
rect 43314 19406 43316 19458
rect 43260 19394 43316 19406
rect 43372 19348 43428 19854
rect 43372 19282 43428 19292
rect 43148 19058 43204 19068
rect 43596 19234 43652 19246
rect 43596 19182 43598 19234
rect 43650 19182 43652 19234
rect 43372 19010 43428 19022
rect 43372 18958 43374 19010
rect 43426 18958 43428 19010
rect 43036 18844 43316 18900
rect 42700 18286 42702 18338
rect 42754 18286 42756 18338
rect 42700 18274 42756 18286
rect 43148 18340 43204 18350
rect 43148 18246 43204 18284
rect 42252 17838 42254 17890
rect 42306 17838 42308 17890
rect 42252 17826 42308 17838
rect 42364 17780 42420 17790
rect 41692 17668 41748 17678
rect 41636 17666 41748 17668
rect 41636 17614 41694 17666
rect 41746 17614 41748 17666
rect 41636 17612 41748 17614
rect 41580 17574 41636 17612
rect 41692 17602 41748 17612
rect 41132 17502 41134 17554
rect 41186 17502 41188 17554
rect 41132 17490 41188 17502
rect 41356 17444 41412 17454
rect 41244 17442 41412 17444
rect 41244 17390 41358 17442
rect 41410 17390 41412 17442
rect 41244 17388 41412 17390
rect 40908 16882 41076 16884
rect 40908 16830 40910 16882
rect 40962 16830 41076 16882
rect 40908 16828 41076 16830
rect 40908 16818 40964 16828
rect 40908 16212 40964 16222
rect 40908 16118 40964 16156
rect 40236 16046 40238 16098
rect 40290 16046 40292 16098
rect 40236 16034 40292 16046
rect 40572 16100 40628 16110
rect 40572 16006 40628 16044
rect 40796 15986 40852 15998
rect 40796 15934 40798 15986
rect 40850 15934 40852 15986
rect 40348 15876 40404 15886
rect 40348 15782 40404 15820
rect 40796 15764 40852 15934
rect 40796 15698 40852 15708
rect 41020 15314 41076 16828
rect 41132 16100 41188 16110
rect 41244 16100 41300 17388
rect 41356 17378 41412 17388
rect 41692 16770 41748 16782
rect 41692 16718 41694 16770
rect 41746 16718 41748 16770
rect 41132 16098 41300 16100
rect 41132 16046 41134 16098
rect 41186 16046 41300 16098
rect 41132 16044 41300 16046
rect 41356 16324 41412 16334
rect 41356 16098 41412 16268
rect 41692 16212 41748 16718
rect 41692 16146 41748 16156
rect 42140 16324 42196 16334
rect 41356 16046 41358 16098
rect 41410 16046 41412 16098
rect 41132 16034 41188 16044
rect 41356 16034 41412 16046
rect 41804 16100 41860 16110
rect 42028 16100 42084 16110
rect 41860 16098 42084 16100
rect 41860 16046 42030 16098
rect 42082 16046 42084 16098
rect 41860 16044 42084 16046
rect 41804 16034 41860 16044
rect 42028 16034 42084 16044
rect 42140 16098 42196 16268
rect 42140 16046 42142 16098
rect 42194 16046 42196 16098
rect 42140 16034 42196 16046
rect 41692 15986 41748 15998
rect 41692 15934 41694 15986
rect 41746 15934 41748 15986
rect 41692 15764 41748 15934
rect 41692 15698 41748 15708
rect 41804 15874 41860 15886
rect 41804 15822 41806 15874
rect 41858 15822 41860 15874
rect 41692 15428 41748 15438
rect 41804 15428 41860 15822
rect 41692 15426 41860 15428
rect 41692 15374 41694 15426
rect 41746 15374 41860 15426
rect 41692 15372 41860 15374
rect 41692 15362 41748 15372
rect 41020 15262 41022 15314
rect 41074 15262 41076 15314
rect 41020 15250 41076 15262
rect 42140 14756 42196 14766
rect 42140 14644 42196 14700
rect 41692 14642 42196 14644
rect 41692 14590 42142 14642
rect 42194 14590 42196 14642
rect 41692 14588 42196 14590
rect 39900 12402 40068 12404
rect 39900 12350 39902 12402
rect 39954 12350 40068 12402
rect 39900 12348 40068 12350
rect 39900 12338 39956 12348
rect 40012 12180 40068 12348
rect 39788 12124 39956 12180
rect 39452 12014 39454 12066
rect 39506 12014 39508 12066
rect 39452 11508 39508 12014
rect 39452 11442 39508 11452
rect 39564 11844 39620 11854
rect 39340 11284 39396 11294
rect 39340 11190 39396 11228
rect 39564 11172 39620 11788
rect 39788 11172 39844 11182
rect 39564 11170 39844 11172
rect 39564 11118 39790 11170
rect 39842 11118 39844 11170
rect 39564 11116 39844 11118
rect 39452 10612 39508 10622
rect 39564 10612 39620 11116
rect 39788 11106 39844 11116
rect 39676 10724 39732 10734
rect 39676 10630 39732 10668
rect 39452 10610 39620 10612
rect 39452 10558 39454 10610
rect 39506 10558 39620 10610
rect 39452 10556 39620 10558
rect 39452 10052 39508 10556
rect 39452 9986 39508 9996
rect 39340 9604 39396 9614
rect 39228 9548 39340 9604
rect 39340 9538 39396 9548
rect 39676 9268 39732 9278
rect 39676 9174 39732 9212
rect 39788 9044 39844 9054
rect 39340 9042 39844 9044
rect 39340 8990 39790 9042
rect 39842 8990 39844 9042
rect 39340 8988 39844 8990
rect 39116 8418 39172 8428
rect 39228 8930 39284 8942
rect 39228 8878 39230 8930
rect 39282 8878 39284 8930
rect 39228 8372 39284 8878
rect 39228 8306 39284 8316
rect 39228 7586 39284 7598
rect 39228 7534 39230 7586
rect 39282 7534 39284 7586
rect 38892 7308 39172 7364
rect 39004 7140 39060 7150
rect 38892 7084 39004 7140
rect 38892 6578 38948 7084
rect 39004 7074 39060 7084
rect 39004 6916 39060 6926
rect 39004 6802 39060 6860
rect 39004 6750 39006 6802
rect 39058 6750 39060 6802
rect 39004 6738 39060 6750
rect 39116 6804 39172 7308
rect 39228 7252 39284 7534
rect 39228 7186 39284 7196
rect 39340 7140 39396 8988
rect 39788 8978 39844 8988
rect 39676 8818 39732 8830
rect 39676 8766 39678 8818
rect 39730 8766 39732 8818
rect 39564 8708 39620 8718
rect 39340 7074 39396 7084
rect 39452 8652 39564 8708
rect 39340 6916 39396 6926
rect 39116 6748 39284 6804
rect 38892 6526 38894 6578
rect 38946 6526 38948 6578
rect 38892 5236 38948 6526
rect 39004 6580 39060 6590
rect 39004 5906 39060 6524
rect 39116 6578 39172 6590
rect 39116 6526 39118 6578
rect 39170 6526 39172 6578
rect 39116 6132 39172 6526
rect 39228 6468 39284 6748
rect 39228 6402 39284 6412
rect 39116 6066 39172 6076
rect 39340 6018 39396 6860
rect 39340 5966 39342 6018
rect 39394 5966 39396 6018
rect 39340 5954 39396 5966
rect 39452 6356 39508 8652
rect 39564 8642 39620 8652
rect 39564 7924 39620 7934
rect 39564 7586 39620 7868
rect 39564 7534 39566 7586
rect 39618 7534 39620 7586
rect 39564 7028 39620 7534
rect 39564 6962 39620 6972
rect 39676 6804 39732 8766
rect 39676 6738 39732 6748
rect 39788 8596 39844 8606
rect 39564 6692 39620 6702
rect 39564 6598 39620 6636
rect 39004 5854 39006 5906
rect 39058 5854 39060 5906
rect 39004 5842 39060 5854
rect 39452 5908 39508 6300
rect 39788 6466 39844 8540
rect 39900 8148 39956 12124
rect 40012 12114 40068 12124
rect 40124 14084 40180 14094
rect 40124 11620 40180 14028
rect 41692 13970 41748 14588
rect 42140 14578 42196 14588
rect 42364 14644 42420 17724
rect 43260 16436 43316 18844
rect 43372 18676 43428 18958
rect 43372 18610 43428 18620
rect 43596 18450 43652 19182
rect 43708 19236 43764 19966
rect 43708 19170 43764 19180
rect 45388 19012 45444 19022
rect 43596 18398 43598 18450
rect 43650 18398 43652 18450
rect 43596 16772 43652 18398
rect 44268 18452 44324 18462
rect 44268 17106 44324 18396
rect 45388 18450 45444 18956
rect 45388 18398 45390 18450
rect 45442 18398 45444 18450
rect 45388 18386 45444 18398
rect 44268 17054 44270 17106
rect 44322 17054 44324 17106
rect 43820 16772 43876 16782
rect 43596 16770 43876 16772
rect 43596 16718 43822 16770
rect 43874 16718 43876 16770
rect 43596 16716 43876 16718
rect 43820 16706 43876 16716
rect 43260 16370 43316 16380
rect 42812 16324 42868 16334
rect 42812 15986 42868 16268
rect 42812 15934 42814 15986
rect 42866 15934 42868 15986
rect 42812 15922 42868 15934
rect 43148 15988 43204 15998
rect 43596 15988 43652 15998
rect 43148 15986 43652 15988
rect 43148 15934 43150 15986
rect 43202 15934 43598 15986
rect 43650 15934 43652 15986
rect 43148 15932 43652 15934
rect 43148 15922 43204 15932
rect 42364 14578 42420 14588
rect 41692 13918 41694 13970
rect 41746 13918 41748 13970
rect 41020 13748 41076 13758
rect 41020 13654 41076 13692
rect 41692 13748 41748 13918
rect 40348 13636 40404 13646
rect 40348 13542 40404 13580
rect 40684 13524 40740 13534
rect 40684 13076 40740 13468
rect 40684 13074 41076 13076
rect 40684 13022 40686 13074
rect 40738 13022 41076 13074
rect 40684 13020 41076 13022
rect 40684 13010 40740 13020
rect 41020 12962 41076 13020
rect 41020 12910 41022 12962
rect 41074 12910 41076 12962
rect 41020 12898 41076 12910
rect 40348 12738 40404 12750
rect 40348 12686 40350 12738
rect 40402 12686 40404 12738
rect 40348 12628 40404 12686
rect 40348 12572 41524 12628
rect 40796 12404 40852 12414
rect 40796 12402 41188 12404
rect 40796 12350 40798 12402
rect 40850 12350 41188 12402
rect 40796 12348 41188 12350
rect 40796 12338 40852 12348
rect 40908 12180 40964 12190
rect 40908 12086 40964 12124
rect 40124 11554 40180 11564
rect 40236 12066 40292 12078
rect 40236 12014 40238 12066
rect 40290 12014 40292 12066
rect 40236 11508 40292 12014
rect 40348 11956 40404 11966
rect 40348 11862 40404 11900
rect 40236 11442 40292 11452
rect 40012 11396 40068 11406
rect 40012 10610 40068 11340
rect 41132 11394 41188 12348
rect 41132 11342 41134 11394
rect 41186 11342 41188 11394
rect 41132 11330 41188 11342
rect 40684 11282 40740 11294
rect 40684 11230 40686 11282
rect 40738 11230 40740 11282
rect 40124 11172 40180 11182
rect 40236 11172 40292 11182
rect 40124 11170 40236 11172
rect 40124 11118 40126 11170
rect 40178 11118 40236 11170
rect 40124 11116 40236 11118
rect 40124 11106 40180 11116
rect 40012 10558 40014 10610
rect 40066 10558 40068 10610
rect 40012 10546 40068 10558
rect 40124 10948 40180 10958
rect 40012 9716 40068 9726
rect 40012 9042 40068 9660
rect 40012 8990 40014 9042
rect 40066 8990 40068 9042
rect 40012 8978 40068 8990
rect 39900 8082 39956 8092
rect 39900 7476 39956 7486
rect 40124 7476 40180 10892
rect 40236 10724 40292 11116
rect 40348 11172 40404 11182
rect 40348 11170 40516 11172
rect 40348 11118 40350 11170
rect 40402 11118 40516 11170
rect 40348 11116 40516 11118
rect 40348 11106 40404 11116
rect 40348 10724 40404 10734
rect 40236 10722 40404 10724
rect 40236 10670 40350 10722
rect 40402 10670 40404 10722
rect 40236 10668 40404 10670
rect 40348 10658 40404 10668
rect 40236 10498 40292 10510
rect 40236 10446 40238 10498
rect 40290 10446 40292 10498
rect 40236 10388 40292 10446
rect 40236 10322 40292 10332
rect 40460 9940 40516 11116
rect 40572 11170 40628 11182
rect 40572 11118 40574 11170
rect 40626 11118 40628 11170
rect 40572 10500 40628 11118
rect 40572 10434 40628 10444
rect 40460 9874 40516 9884
rect 40684 9268 40740 11230
rect 41244 11284 41300 11294
rect 41244 11190 41300 11228
rect 41356 10836 41412 10846
rect 41020 10834 41412 10836
rect 41020 10782 41358 10834
rect 41410 10782 41412 10834
rect 41020 10780 41412 10782
rect 40796 10052 40852 10062
rect 40796 9938 40852 9996
rect 40796 9886 40798 9938
rect 40850 9886 40852 9938
rect 40796 9874 40852 9886
rect 40908 9940 40964 9950
rect 40908 9716 40964 9884
rect 40908 9650 40964 9660
rect 40796 9268 40852 9278
rect 40684 9266 40852 9268
rect 40684 9214 40798 9266
rect 40850 9214 40852 9266
rect 40684 9212 40852 9214
rect 40796 9202 40852 9212
rect 40908 9154 40964 9166
rect 40908 9102 40910 9154
rect 40962 9102 40964 9154
rect 40908 9044 40964 9102
rect 40572 8988 40964 9044
rect 40348 8484 40404 8494
rect 40236 7700 40292 7710
rect 40236 7606 40292 7644
rect 40124 7420 40292 7476
rect 39900 7382 39956 7420
rect 39788 6414 39790 6466
rect 39842 6414 39844 6466
rect 39564 5908 39620 5918
rect 39452 5906 39620 5908
rect 39452 5854 39566 5906
rect 39618 5854 39620 5906
rect 39452 5852 39620 5854
rect 39564 5842 39620 5852
rect 39788 5906 39844 6414
rect 40012 7252 40068 7262
rect 39900 6132 39956 6142
rect 40012 6132 40068 7196
rect 39900 6130 40068 6132
rect 39900 6078 39902 6130
rect 39954 6078 40068 6130
rect 39900 6076 40068 6078
rect 40124 6468 40180 6478
rect 39900 6066 39956 6076
rect 39788 5854 39790 5906
rect 39842 5854 39844 5906
rect 39788 5842 39844 5854
rect 39900 5908 39956 5918
rect 39900 5814 39956 5852
rect 40012 5684 40068 5694
rect 38892 5170 38948 5180
rect 39900 5236 39956 5246
rect 39004 5010 39060 5022
rect 39004 4958 39006 5010
rect 39058 4958 39060 5010
rect 39004 4116 39060 4958
rect 39452 4788 39508 4798
rect 39116 4676 39172 4686
rect 39116 4562 39172 4620
rect 39116 4510 39118 4562
rect 39170 4510 39172 4562
rect 39116 4498 39172 4510
rect 39340 4564 39396 4574
rect 39340 4470 39396 4508
rect 39452 4450 39508 4732
rect 39452 4398 39454 4450
rect 39506 4398 39508 4450
rect 39452 4386 39508 4398
rect 39900 4226 39956 5180
rect 39900 4174 39902 4226
rect 39954 4174 39956 4226
rect 39900 4162 39956 4174
rect 39004 4050 39060 4060
rect 38892 3668 38948 3678
rect 38780 3666 38948 3668
rect 38780 3614 38894 3666
rect 38946 3614 38948 3666
rect 38780 3612 38948 3614
rect 38892 3602 38948 3612
rect 38556 3490 38612 3500
rect 40012 3554 40068 5628
rect 40012 3502 40014 3554
rect 40066 3502 40068 3554
rect 40012 3490 40068 3502
rect 38444 2482 38500 2492
rect 38780 3444 38836 3454
rect 38780 800 38836 3388
rect 40124 800 40180 6412
rect 40236 6132 40292 7420
rect 40236 6066 40292 6076
rect 40236 5908 40292 5918
rect 40236 5814 40292 5852
rect 40236 5684 40292 5694
rect 40236 5124 40292 5628
rect 40236 4338 40292 5068
rect 40348 5122 40404 8428
rect 40572 6916 40628 8988
rect 41020 8932 41076 10780
rect 41356 10770 41412 10780
rect 41356 10612 41412 10622
rect 41356 10518 41412 10556
rect 41132 10500 41188 10510
rect 41132 10406 41188 10444
rect 41356 9940 41412 9950
rect 41244 9884 41356 9940
rect 40684 8876 41076 8932
rect 41132 9042 41188 9054
rect 41132 8990 41134 9042
rect 41186 8990 41188 9042
rect 40684 8370 40740 8876
rect 40684 8318 40686 8370
rect 40738 8318 40740 8370
rect 40684 8306 40740 8318
rect 41020 7700 41076 7710
rect 40572 6850 40628 6860
rect 40796 7698 41076 7700
rect 40796 7646 41022 7698
rect 41074 7646 41076 7698
rect 40796 7644 41076 7646
rect 40684 6578 40740 6590
rect 40684 6526 40686 6578
rect 40738 6526 40740 6578
rect 40684 6132 40740 6526
rect 40684 6066 40740 6076
rect 40348 5070 40350 5122
rect 40402 5070 40404 5122
rect 40348 5058 40404 5070
rect 40460 5346 40516 5358
rect 40460 5294 40462 5346
rect 40514 5294 40516 5346
rect 40236 4286 40238 4338
rect 40290 4286 40292 4338
rect 40236 4274 40292 4286
rect 40460 2884 40516 5294
rect 40796 4900 40852 7644
rect 41020 7634 41076 7644
rect 41132 7700 41188 8990
rect 41132 7634 41188 7644
rect 41244 7476 41300 9884
rect 41356 9874 41412 9884
rect 41468 9716 41524 12572
rect 41580 10388 41636 10398
rect 41580 10294 41636 10332
rect 41692 9940 41748 13692
rect 41804 14306 41860 14318
rect 41804 14254 41806 14306
rect 41858 14254 41860 14306
rect 41804 13522 41860 14254
rect 42700 14308 42756 14318
rect 42700 14306 42980 14308
rect 42700 14254 42702 14306
rect 42754 14254 42980 14306
rect 42700 14252 42980 14254
rect 42700 14242 42756 14252
rect 42588 14084 42644 14094
rect 42140 13972 42196 13982
rect 42140 13878 42196 13916
rect 42588 13970 42644 14028
rect 42588 13918 42590 13970
rect 42642 13918 42644 13970
rect 42588 13906 42644 13918
rect 41804 13470 41806 13522
rect 41858 13470 41860 13522
rect 41804 13458 41860 13470
rect 42812 13076 42868 13086
rect 41804 12850 41860 12862
rect 41804 12798 41806 12850
rect 41858 12798 41860 12850
rect 41804 12404 41860 12798
rect 41804 12338 41860 12348
rect 42364 12292 42420 12302
rect 42364 12198 42420 12236
rect 42700 12290 42756 12302
rect 42700 12238 42702 12290
rect 42754 12238 42756 12290
rect 41916 12180 41972 12190
rect 41916 12086 41972 12124
rect 42700 11788 42756 12238
rect 42476 11732 42756 11788
rect 42812 12178 42868 13020
rect 42812 12126 42814 12178
rect 42866 12126 42868 12178
rect 42812 11844 42868 12126
rect 42924 12180 42980 14252
rect 43148 13634 43204 13646
rect 43148 13582 43150 13634
rect 43202 13582 43204 13634
rect 43148 13522 43204 13582
rect 43148 13470 43150 13522
rect 43202 13470 43204 13522
rect 43148 12516 43204 13470
rect 43204 12460 43316 12516
rect 43148 12450 43204 12460
rect 42924 12124 43204 12180
rect 42812 11778 42868 11788
rect 42924 11956 42980 11966
rect 41692 9874 41748 9884
rect 41804 11506 41860 11518
rect 41804 11454 41806 11506
rect 41858 11454 41860 11506
rect 41692 9716 41748 9726
rect 41468 9714 41748 9716
rect 41468 9662 41694 9714
rect 41746 9662 41748 9714
rect 41468 9660 41748 9662
rect 41356 9042 41412 9054
rect 41356 8990 41358 9042
rect 41410 8990 41412 9042
rect 41356 8708 41412 8990
rect 41356 8642 41412 8652
rect 41356 8260 41412 8270
rect 41356 8166 41412 8204
rect 41356 7476 41412 7486
rect 41244 7474 41412 7476
rect 41244 7422 41358 7474
rect 41410 7422 41412 7474
rect 41244 7420 41412 7422
rect 41020 7252 41076 7262
rect 41020 7158 41076 7196
rect 41132 7250 41188 7262
rect 41132 7198 41134 7250
rect 41186 7198 41188 7250
rect 41020 7028 41076 7038
rect 41020 6020 41076 6972
rect 41132 6692 41188 7198
rect 41132 6626 41188 6636
rect 41356 6468 41412 7420
rect 41580 7476 41636 7486
rect 41580 6692 41636 7420
rect 41580 6598 41636 6636
rect 41356 6412 41636 6468
rect 40908 5908 40964 5918
rect 40908 5814 40964 5852
rect 41020 5906 41076 5964
rect 41020 5854 41022 5906
rect 41074 5854 41076 5906
rect 41020 5842 41076 5854
rect 41468 6132 41524 6142
rect 41468 5906 41524 6076
rect 41468 5854 41470 5906
rect 41522 5854 41524 5906
rect 41244 5682 41300 5694
rect 41244 5630 41246 5682
rect 41298 5630 41300 5682
rect 40796 4834 40852 4844
rect 41132 5348 41188 5358
rect 41132 4338 41188 5292
rect 41244 5236 41300 5630
rect 41244 5170 41300 5180
rect 41132 4286 41134 4338
rect 41186 4286 41188 4338
rect 41132 4274 41188 4286
rect 41356 5124 41412 5134
rect 41356 4338 41412 5068
rect 41468 4900 41524 5854
rect 41468 4834 41524 4844
rect 41356 4286 41358 4338
rect 41410 4286 41412 4338
rect 41356 4274 41412 4286
rect 41468 4452 41524 4462
rect 40796 3668 40852 3678
rect 40796 3574 40852 3612
rect 40460 2818 40516 2828
rect 41468 800 41524 4396
rect 41580 4338 41636 6412
rect 41692 5572 41748 9660
rect 41804 6692 41860 11454
rect 42252 11396 42308 11406
rect 42476 11396 42532 11732
rect 42252 11394 42420 11396
rect 42252 11342 42254 11394
rect 42306 11342 42420 11394
rect 42252 11340 42420 11342
rect 42252 11330 42308 11340
rect 41916 10836 41972 10846
rect 41916 10722 41972 10780
rect 41916 10670 41918 10722
rect 41970 10670 41972 10722
rect 41916 10658 41972 10670
rect 42140 10724 42196 10734
rect 42140 10630 42196 10668
rect 42364 10386 42420 11340
rect 42476 11330 42532 11340
rect 42700 11620 42756 11630
rect 42588 11284 42644 11294
rect 42588 11190 42644 11228
rect 42588 10836 42644 10846
rect 42700 10836 42756 11564
rect 42924 11618 42980 11900
rect 42924 11566 42926 11618
rect 42978 11566 42980 11618
rect 42924 11554 42980 11566
rect 43036 11732 43092 11742
rect 42644 10780 42756 10836
rect 42812 11508 42868 11518
rect 42588 10742 42644 10780
rect 42364 10334 42366 10386
rect 42418 10334 42420 10386
rect 42364 10322 42420 10334
rect 42476 10500 42532 10510
rect 42252 10164 42308 10174
rect 42140 10108 42252 10164
rect 41916 9154 41972 9166
rect 41916 9102 41918 9154
rect 41970 9102 41972 9154
rect 41916 8370 41972 9102
rect 41916 8318 41918 8370
rect 41970 8318 41972 8370
rect 41916 8306 41972 8318
rect 42028 8260 42084 8270
rect 42028 7474 42084 8204
rect 42028 7422 42030 7474
rect 42082 7422 42084 7474
rect 42028 7410 42084 7422
rect 41804 6626 41860 6636
rect 41916 6020 41972 6030
rect 41804 5964 41916 6020
rect 41804 5906 41860 5964
rect 41916 5954 41972 5964
rect 41804 5854 41806 5906
rect 41858 5854 41860 5906
rect 41804 5842 41860 5854
rect 41692 5516 41860 5572
rect 41580 4286 41582 4338
rect 41634 4286 41636 4338
rect 41580 4274 41636 4286
rect 41692 4228 41748 4238
rect 41692 4134 41748 4172
rect 41804 3444 41860 5516
rect 42140 4900 42196 10108
rect 42252 10098 42308 10108
rect 42252 6580 42308 6590
rect 42252 5124 42308 6524
rect 42364 6356 42420 6366
rect 42364 6130 42420 6300
rect 42364 6078 42366 6130
rect 42418 6078 42420 6130
rect 42364 6066 42420 6078
rect 42252 5030 42308 5068
rect 42140 4844 42308 4900
rect 42140 4226 42196 4238
rect 42140 4174 42142 4226
rect 42194 4174 42196 4226
rect 42140 4004 42196 4174
rect 42140 3938 42196 3948
rect 41804 3378 41860 3388
rect 42252 980 42308 4844
rect 42476 2324 42532 10444
rect 42812 10052 42868 11452
rect 42924 11396 42980 11406
rect 43036 11396 43092 11676
rect 42924 11394 43092 11396
rect 42924 11342 42926 11394
rect 42978 11342 43092 11394
rect 42924 11340 43092 11342
rect 42924 11330 42980 11340
rect 43148 11284 43204 12124
rect 43036 11228 43204 11284
rect 43036 11172 43092 11228
rect 42700 9996 42868 10052
rect 42924 11116 43092 11172
rect 42588 9938 42644 9950
rect 42588 9886 42590 9938
rect 42642 9886 42644 9938
rect 42588 5012 42644 9886
rect 42588 4946 42644 4956
rect 42588 4564 42644 4574
rect 42588 4470 42644 4508
rect 42700 3442 42756 9996
rect 42812 8036 42868 8046
rect 42812 7586 42868 7980
rect 42812 7534 42814 7586
rect 42866 7534 42868 7586
rect 42812 7522 42868 7534
rect 42812 5796 42868 5806
rect 42812 5702 42868 5740
rect 42924 5684 42980 11116
rect 43036 10948 43092 10958
rect 43036 10834 43092 10892
rect 43036 10782 43038 10834
rect 43090 10782 43092 10834
rect 43036 10164 43092 10782
rect 43036 10098 43092 10108
rect 43148 10388 43204 10398
rect 43148 9938 43204 10332
rect 43148 9886 43150 9938
rect 43202 9886 43204 9938
rect 43148 9874 43204 9886
rect 43260 9156 43316 12460
rect 43148 9100 43316 9156
rect 43036 8930 43092 8942
rect 43036 8878 43038 8930
rect 43090 8878 43092 8930
rect 43036 8596 43092 8878
rect 43148 8820 43204 9100
rect 43372 9044 43428 15932
rect 43596 15922 43652 15932
rect 43820 15876 43876 15886
rect 43820 15202 43876 15820
rect 44268 15540 44324 17054
rect 45388 17780 45444 17790
rect 45500 17780 45556 23324
rect 45612 23154 45668 24108
rect 46060 24052 46116 24062
rect 46508 24052 46564 24558
rect 46732 24164 46788 27132
rect 46732 24098 46788 24108
rect 45948 23996 46060 24052
rect 45948 23938 46004 23996
rect 46060 23986 46116 23996
rect 46172 23996 46564 24052
rect 45948 23886 45950 23938
rect 46002 23886 46004 23938
rect 45948 23874 46004 23886
rect 46060 23826 46116 23838
rect 46060 23774 46062 23826
rect 46114 23774 46116 23826
rect 45724 23716 45780 23726
rect 46060 23716 46116 23774
rect 45724 23714 46116 23716
rect 45724 23662 45726 23714
rect 45778 23662 46116 23714
rect 45724 23660 46116 23662
rect 45724 23650 45780 23660
rect 46172 23604 46228 23996
rect 46732 23940 46788 23950
rect 46732 23846 46788 23884
rect 46284 23828 46340 23838
rect 46284 23734 46340 23772
rect 46396 23716 46452 23726
rect 45612 23102 45614 23154
rect 45666 23102 45668 23154
rect 45612 21700 45668 23102
rect 45612 21634 45668 21644
rect 46060 23548 46228 23604
rect 46284 23604 46340 23614
rect 45612 20916 45668 20926
rect 45612 20802 45668 20860
rect 45612 20750 45614 20802
rect 45666 20750 45668 20802
rect 45612 20244 45668 20750
rect 45836 20916 45892 20926
rect 45836 20690 45892 20860
rect 45948 20804 46004 20814
rect 45948 20710 46004 20748
rect 45836 20638 45838 20690
rect 45890 20638 45892 20690
rect 45836 20626 45892 20638
rect 45612 20178 45668 20188
rect 46060 19236 46116 23548
rect 46284 23154 46340 23548
rect 46396 23266 46452 23660
rect 46844 23604 46900 31948
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 48300 30996 48356 31006
rect 46956 29428 47012 29438
rect 46956 29426 47124 29428
rect 46956 29374 46958 29426
rect 47010 29374 47124 29426
rect 46956 29372 47124 29374
rect 46956 29362 47012 29372
rect 47068 29316 47124 29372
rect 47292 29316 47348 29326
rect 47068 29260 47292 29316
rect 46956 24722 47012 24734
rect 46956 24670 46958 24722
rect 47010 24670 47012 24722
rect 46956 24162 47012 24670
rect 46956 24110 46958 24162
rect 47010 24110 47012 24162
rect 46956 24098 47012 24110
rect 46396 23214 46398 23266
rect 46450 23214 46452 23266
rect 46396 23202 46452 23214
rect 46508 23548 46900 23604
rect 46284 23102 46286 23154
rect 46338 23102 46340 23154
rect 46284 23090 46340 23102
rect 46284 21586 46340 21598
rect 46284 21534 46286 21586
rect 46338 21534 46340 21586
rect 46284 19684 46340 21534
rect 46396 21028 46452 21038
rect 46508 21028 46564 23548
rect 46956 23268 47012 23278
rect 46956 23174 47012 23212
rect 46620 23156 46676 23166
rect 46620 23154 46788 23156
rect 46620 23102 46622 23154
rect 46674 23102 46788 23154
rect 46620 23100 46788 23102
rect 46620 23090 46676 23100
rect 46620 21700 46676 21710
rect 46620 21606 46676 21644
rect 46396 21026 46564 21028
rect 46396 20974 46398 21026
rect 46450 20974 46564 21026
rect 46396 20972 46564 20974
rect 46396 20962 46452 20972
rect 46732 20804 46788 23100
rect 47068 22484 47124 29260
rect 47292 29222 47348 29260
rect 47740 27074 47796 27086
rect 47740 27022 47742 27074
rect 47794 27022 47796 27074
rect 47292 25732 47348 25742
rect 47740 25732 47796 27022
rect 47964 26964 48020 26974
rect 47852 26852 47908 26862
rect 47852 26514 47908 26796
rect 47852 26462 47854 26514
rect 47906 26462 47908 26514
rect 47852 26450 47908 26462
rect 47348 25676 47796 25732
rect 47292 25506 47348 25676
rect 47292 25454 47294 25506
rect 47346 25454 47348 25506
rect 47292 25442 47348 25454
rect 47740 25506 47796 25518
rect 47740 25454 47742 25506
rect 47794 25454 47796 25506
rect 47740 25284 47796 25454
rect 47740 25218 47796 25228
rect 47180 24164 47236 24174
rect 47964 24164 48020 26908
rect 48076 26402 48132 26414
rect 48076 26350 48078 26402
rect 48130 26350 48132 26402
rect 48076 26292 48132 26350
rect 48076 26226 48132 26236
rect 48188 26290 48244 26302
rect 48188 26238 48190 26290
rect 48242 26238 48244 26290
rect 48188 25844 48244 26238
rect 48188 25778 48244 25788
rect 48076 25732 48132 25742
rect 48076 25618 48132 25676
rect 48076 25566 48078 25618
rect 48130 25566 48132 25618
rect 48076 25554 48132 25566
rect 47180 23938 47236 24108
rect 47740 24108 48020 24164
rect 47628 24052 47684 24062
rect 47180 23886 47182 23938
rect 47234 23886 47236 23938
rect 47180 23492 47236 23886
rect 47292 23940 47348 23950
rect 47292 23846 47348 23884
rect 47180 23426 47236 23436
rect 47404 23714 47460 23726
rect 47404 23662 47406 23714
rect 47458 23662 47460 23714
rect 47180 23154 47236 23166
rect 47180 23102 47182 23154
rect 47234 23102 47236 23154
rect 47180 22596 47236 23102
rect 47404 22820 47460 23662
rect 47628 23156 47684 23996
rect 47628 22932 47684 23100
rect 47740 23154 47796 24108
rect 47852 23940 47908 23950
rect 47852 23938 48244 23940
rect 47852 23886 47854 23938
rect 47906 23886 48244 23938
rect 47852 23884 48244 23886
rect 47852 23874 47908 23884
rect 48188 23714 48244 23884
rect 48188 23662 48190 23714
rect 48242 23662 48244 23714
rect 47852 23268 47908 23278
rect 47908 23212 48020 23268
rect 47852 23202 47908 23212
rect 47740 23102 47742 23154
rect 47794 23102 47796 23154
rect 47740 23044 47796 23102
rect 47740 22988 47908 23044
rect 47628 22876 47796 22932
rect 47404 22754 47460 22764
rect 47180 22530 47236 22540
rect 47068 22390 47124 22428
rect 46844 22148 46900 22158
rect 46900 22092 47012 22148
rect 46844 22082 46900 22092
rect 46844 21700 46900 21710
rect 46844 21362 46900 21644
rect 46844 21310 46846 21362
rect 46898 21310 46900 21362
rect 46844 21298 46900 21310
rect 46732 20738 46788 20748
rect 46844 20692 46900 20702
rect 46844 20598 46900 20636
rect 46956 20468 47012 22092
rect 47404 21812 47460 21822
rect 47404 21810 47684 21812
rect 47404 21758 47406 21810
rect 47458 21758 47684 21810
rect 47404 21756 47684 21758
rect 47404 21746 47460 21756
rect 47292 21698 47348 21710
rect 47292 21646 47294 21698
rect 47346 21646 47348 21698
rect 47292 21644 47348 21646
rect 47628 21698 47684 21756
rect 47740 21810 47796 22876
rect 47740 21758 47742 21810
rect 47794 21758 47796 21810
rect 47740 21746 47796 21758
rect 47628 21646 47630 21698
rect 47682 21646 47684 21698
rect 47292 21588 47572 21644
rect 47628 21634 47684 21646
rect 47852 21588 47908 22988
rect 47964 21810 48020 23212
rect 48188 23044 48244 23662
rect 47964 21758 47966 21810
rect 48018 21758 48020 21810
rect 47964 21746 48020 21758
rect 48076 22820 48132 22830
rect 47068 21476 47124 21486
rect 47516 21476 47572 21588
rect 47068 21382 47124 21420
rect 47292 21420 47572 21476
rect 47740 21532 47908 21588
rect 47068 20580 47124 20590
rect 47292 20580 47348 21420
rect 47404 21140 47460 21150
rect 47404 20804 47460 21084
rect 47740 20916 47796 21532
rect 47404 20802 47572 20804
rect 47404 20750 47406 20802
rect 47458 20750 47572 20802
rect 47404 20748 47572 20750
rect 47404 20738 47460 20748
rect 47068 20486 47124 20524
rect 47180 20578 47348 20580
rect 47180 20526 47294 20578
rect 47346 20526 47348 20578
rect 47180 20524 47348 20526
rect 46284 19618 46340 19628
rect 46732 20412 47012 20468
rect 46060 19170 46116 19180
rect 46732 19122 46788 20412
rect 46732 19070 46734 19122
rect 46786 19070 46788 19122
rect 46732 19058 46788 19070
rect 46844 19122 46900 19134
rect 46844 19070 46846 19122
rect 46898 19070 46900 19122
rect 46284 19012 46340 19022
rect 46284 18452 46340 18956
rect 46508 19010 46564 19022
rect 46508 18958 46510 19010
rect 46562 18958 46564 19010
rect 46508 18452 46564 18958
rect 46844 18788 46900 19070
rect 46844 18722 46900 18732
rect 46284 18450 46452 18452
rect 46284 18398 46286 18450
rect 46338 18398 46452 18450
rect 46284 18396 46452 18398
rect 46284 18386 46340 18396
rect 45724 18338 45780 18350
rect 45724 18286 45726 18338
rect 45778 18286 45780 18338
rect 45724 17892 45780 18286
rect 45724 17826 45780 17836
rect 45388 17778 45556 17780
rect 45388 17726 45390 17778
rect 45442 17726 45556 17778
rect 45388 17724 45556 17726
rect 44268 15446 44324 15484
rect 45276 15540 45332 15550
rect 45276 15314 45332 15484
rect 45276 15262 45278 15314
rect 45330 15262 45332 15314
rect 45276 15250 45332 15262
rect 43820 15150 43822 15202
rect 43874 15150 43876 15202
rect 43820 15138 43876 15150
rect 44940 14756 44996 14766
rect 45388 14756 45444 17724
rect 45836 17668 45892 17678
rect 45836 17574 45892 17612
rect 46284 17668 46340 17678
rect 46284 17554 46340 17612
rect 46284 17502 46286 17554
rect 46338 17502 46340 17554
rect 46284 17490 46340 17502
rect 45724 17220 45780 17230
rect 45724 15148 45780 17164
rect 46172 17220 46228 17230
rect 45948 16996 46004 17006
rect 45948 16902 46004 16940
rect 46060 16884 46116 16894
rect 46060 15426 46116 16828
rect 46060 15374 46062 15426
rect 46114 15374 46116 15426
rect 46060 15362 46116 15374
rect 45724 15092 46004 15148
rect 44940 14754 45220 14756
rect 44940 14702 44942 14754
rect 44994 14702 45220 14754
rect 44940 14700 45220 14702
rect 44940 14690 44996 14700
rect 44940 14532 44996 14542
rect 44996 14476 45108 14532
rect 44940 14466 44996 14476
rect 44828 14418 44884 14430
rect 44828 14366 44830 14418
rect 44882 14366 44884 14418
rect 44492 14084 44548 14094
rect 44492 13970 44548 14028
rect 44492 13918 44494 13970
rect 44546 13918 44548 13970
rect 44492 13906 44548 13918
rect 43708 13634 43764 13646
rect 43708 13582 43710 13634
rect 43762 13582 43764 13634
rect 43596 12178 43652 12190
rect 43596 12126 43598 12178
rect 43650 12126 43652 12178
rect 43596 11844 43652 12126
rect 43708 12180 43764 13582
rect 44156 13634 44212 13646
rect 44156 13582 44158 13634
rect 44210 13582 44212 13634
rect 43932 13522 43988 13534
rect 43932 13470 43934 13522
rect 43986 13470 43988 13522
rect 43932 13076 43988 13470
rect 43932 12982 43988 13020
rect 43820 12404 43876 12414
rect 44156 12404 44212 13582
rect 44828 13522 44884 14366
rect 44940 13972 44996 13982
rect 45052 13972 45108 14476
rect 44940 13970 45108 13972
rect 44940 13918 44942 13970
rect 44994 13918 45108 13970
rect 44940 13916 45108 13918
rect 44940 13906 44996 13916
rect 44828 13470 44830 13522
rect 44882 13470 44884 13522
rect 44828 13458 44884 13470
rect 45164 13412 45220 14700
rect 45388 14690 45444 14700
rect 45836 13746 45892 13758
rect 45836 13694 45838 13746
rect 45890 13694 45892 13746
rect 45612 13634 45668 13646
rect 45612 13582 45614 13634
rect 45666 13582 45668 13634
rect 45500 13524 45556 13534
rect 45164 13346 45220 13356
rect 45388 13522 45556 13524
rect 45388 13470 45502 13522
rect 45554 13470 45556 13522
rect 45388 13468 45556 13470
rect 44828 13074 44884 13086
rect 44828 13022 44830 13074
rect 44882 13022 44884 13074
rect 44828 12852 44884 13022
rect 44828 12786 44884 12796
rect 45388 12404 45444 13468
rect 45500 13458 45556 13468
rect 45612 12628 45668 13582
rect 45836 12852 45892 13694
rect 45836 12786 45892 12796
rect 43820 12310 43876 12348
rect 43932 12348 44212 12404
rect 45052 12348 45444 12404
rect 45500 12572 45668 12628
rect 43708 12124 43876 12180
rect 43708 11956 43764 11966
rect 43708 11862 43764 11900
rect 43596 10612 43652 11788
rect 43820 11396 43876 12124
rect 43596 10546 43652 10556
rect 43708 11340 43876 11396
rect 43372 8978 43428 8988
rect 43484 10498 43540 10510
rect 43484 10446 43486 10498
rect 43538 10446 43540 10498
rect 43148 8764 43428 8820
rect 43036 8540 43316 8596
rect 42924 5236 42980 5628
rect 42924 5170 42980 5180
rect 43036 8372 43092 8382
rect 43036 4338 43092 8316
rect 43036 4286 43038 4338
rect 43090 4286 43092 4338
rect 43036 4274 43092 4286
rect 43148 6580 43204 6590
rect 42924 3556 42980 3566
rect 42924 3462 42980 3500
rect 42700 3390 42702 3442
rect 42754 3390 42756 3442
rect 42700 3378 42756 3390
rect 43148 3332 43204 6524
rect 43260 6130 43316 8540
rect 43260 6078 43262 6130
rect 43314 6078 43316 6130
rect 43260 6066 43316 6078
rect 43372 6578 43428 8764
rect 43372 6526 43374 6578
rect 43426 6526 43428 6578
rect 43372 6020 43428 6526
rect 43372 5954 43428 5964
rect 43484 8148 43540 10446
rect 43596 10164 43652 10174
rect 43596 9826 43652 10108
rect 43596 9774 43598 9826
rect 43650 9774 43652 9826
rect 43596 9762 43652 9774
rect 43708 9828 43764 11340
rect 43820 11170 43876 11182
rect 43820 11118 43822 11170
rect 43874 11118 43876 11170
rect 43820 10724 43876 11118
rect 43932 11060 43988 12348
rect 44044 12178 44100 12190
rect 44268 12180 44324 12190
rect 44828 12180 44884 12190
rect 44044 12126 44046 12178
rect 44098 12126 44100 12178
rect 44044 12068 44100 12126
rect 44044 12002 44100 12012
rect 44156 12178 44884 12180
rect 44156 12126 44270 12178
rect 44322 12126 44830 12178
rect 44882 12126 44884 12178
rect 44156 12124 44884 12126
rect 43932 10994 43988 11004
rect 44156 11060 44212 12124
rect 44268 12114 44324 12124
rect 44828 12114 44884 12124
rect 45052 11396 45108 12348
rect 44940 11340 45108 11396
rect 45164 12178 45220 12190
rect 45164 12126 45166 12178
rect 45218 12126 45220 12178
rect 44940 11284 44996 11340
rect 44268 11172 44324 11182
rect 44268 11170 44548 11172
rect 44268 11118 44270 11170
rect 44322 11118 44548 11170
rect 44268 11116 44548 11118
rect 44268 11106 44324 11116
rect 44156 10994 44212 11004
rect 43820 10668 44212 10724
rect 43820 10498 43876 10510
rect 43820 10446 43822 10498
rect 43874 10446 43876 10498
rect 43820 10052 43876 10446
rect 43932 10386 43988 10398
rect 43932 10334 43934 10386
rect 43986 10334 43988 10386
rect 43932 10164 43988 10334
rect 43932 10098 43988 10108
rect 44156 10276 44212 10668
rect 44268 10612 44324 10622
rect 44268 10518 44324 10556
rect 44156 10052 44212 10220
rect 44380 10498 44436 10510
rect 44380 10446 44382 10498
rect 44434 10446 44436 10498
rect 44156 9996 44324 10052
rect 43820 9986 43876 9996
rect 44156 9828 44212 9838
rect 43708 9772 43988 9828
rect 43820 9042 43876 9054
rect 43820 8990 43822 9042
rect 43874 8990 43876 9042
rect 43820 8372 43876 8990
rect 43820 8306 43876 8316
rect 43820 8148 43876 8158
rect 43484 8146 43876 8148
rect 43484 8094 43822 8146
rect 43874 8094 43876 8146
rect 43484 8092 43876 8094
rect 43260 5236 43316 5246
rect 43260 5142 43316 5180
rect 43148 3266 43204 3276
rect 42476 2258 42532 2268
rect 42252 914 42308 924
rect 42812 924 43092 980
rect 42812 800 42868 924
rect 17612 700 18228 756
rect 18592 0 18704 800
rect 19936 0 20048 800
rect 21280 0 21392 800
rect 22624 0 22736 800
rect 23968 0 24080 800
rect 25312 0 25424 800
rect 26656 0 26768 800
rect 28000 0 28112 800
rect 29344 0 29456 800
rect 30688 0 30800 800
rect 32032 0 32144 800
rect 33376 0 33488 800
rect 34720 0 34832 800
rect 36064 0 36176 800
rect 37408 0 37520 800
rect 38752 0 38864 800
rect 40096 0 40208 800
rect 41440 0 41552 800
rect 42784 0 42896 800
rect 43036 756 43092 924
rect 43484 756 43540 8092
rect 43820 8082 43876 8092
rect 43932 7812 43988 9772
rect 44044 9714 44100 9726
rect 44044 9662 44046 9714
rect 44098 9662 44100 9714
rect 44044 7924 44100 9662
rect 44156 9714 44212 9772
rect 44156 9662 44158 9714
rect 44210 9662 44212 9714
rect 44156 9650 44212 9662
rect 44268 8036 44324 9996
rect 44380 9828 44436 10446
rect 44492 10052 44548 11116
rect 44604 10612 44660 10622
rect 44828 10612 44884 10622
rect 44604 10518 44660 10556
rect 44716 10610 44884 10612
rect 44716 10558 44830 10610
rect 44882 10558 44884 10610
rect 44716 10556 44884 10558
rect 44716 10500 44772 10556
rect 44828 10546 44884 10556
rect 44716 10434 44772 10444
rect 44828 10386 44884 10398
rect 44828 10334 44830 10386
rect 44882 10334 44884 10386
rect 44492 9986 44548 9996
rect 44716 10052 44772 10062
rect 44380 9772 44548 9828
rect 44380 9602 44436 9614
rect 44380 9550 44382 9602
rect 44434 9550 44436 9602
rect 44380 8260 44436 9550
rect 44492 9154 44548 9772
rect 44492 9102 44494 9154
rect 44546 9102 44548 9154
rect 44492 9090 44548 9102
rect 44716 9156 44772 9996
rect 44828 9940 44884 10334
rect 44940 10052 44996 11228
rect 45052 11170 45108 11182
rect 45052 11118 45054 11170
rect 45106 11118 45108 11170
rect 45052 10276 45108 11118
rect 45164 11172 45220 12126
rect 45388 11956 45444 11966
rect 45500 11956 45556 12572
rect 45836 12516 45892 12526
rect 45612 12404 45668 12414
rect 45612 12310 45668 12348
rect 45388 11954 45556 11956
rect 45388 11902 45390 11954
rect 45442 11902 45556 11954
rect 45388 11900 45556 11902
rect 45612 12178 45668 12190
rect 45612 12126 45614 12178
rect 45666 12126 45668 12178
rect 45388 11890 45444 11900
rect 45612 11844 45668 12126
rect 45612 11778 45668 11788
rect 45836 11844 45892 12460
rect 45836 11778 45892 11788
rect 45948 12290 46004 15092
rect 46060 14306 46116 14318
rect 46060 14254 46062 14306
rect 46114 14254 46116 14306
rect 46060 13522 46116 14254
rect 46060 13470 46062 13522
rect 46114 13470 46116 13522
rect 46060 13458 46116 13470
rect 46172 12404 46228 17164
rect 46396 14980 46452 18396
rect 46508 18386 46564 18396
rect 46508 17666 46564 17678
rect 46508 17614 46510 17666
rect 46562 17614 46564 17666
rect 46508 16996 46564 17614
rect 46956 17442 47012 17454
rect 46956 17390 46958 17442
rect 47010 17390 47012 17442
rect 46956 17220 47012 17390
rect 46956 17154 47012 17164
rect 46508 16212 46564 16940
rect 46508 16146 46564 16156
rect 46844 16098 46900 16110
rect 46844 16046 46846 16098
rect 46898 16046 46900 16098
rect 46844 15148 46900 16046
rect 47180 15876 47236 20524
rect 47292 20514 47348 20524
rect 47292 20244 47348 20254
rect 47348 20188 47460 20244
rect 47292 20178 47348 20188
rect 47292 17668 47348 17678
rect 47292 17574 47348 17612
rect 47404 17444 47460 20188
rect 47516 19122 47572 20748
rect 47740 20802 47796 20860
rect 47740 20750 47742 20802
rect 47794 20750 47796 20802
rect 47740 20738 47796 20750
rect 48076 20580 48132 22764
rect 48188 21476 48244 22988
rect 48188 21410 48244 21420
rect 48188 20692 48244 20702
rect 48300 20692 48356 30940
rect 49756 30772 49812 30782
rect 48860 30322 48916 30334
rect 48860 30270 48862 30322
rect 48914 30270 48916 30322
rect 48860 28980 48916 30270
rect 49308 30210 49364 30222
rect 49308 30158 49310 30210
rect 49362 30158 49364 30210
rect 49308 29988 49364 30158
rect 49308 29922 49364 29932
rect 49084 29316 49140 29326
rect 49084 29222 49140 29260
rect 49420 29092 49476 29102
rect 49476 29036 49588 29092
rect 49420 29026 49476 29036
rect 49308 28980 49364 28990
rect 48860 28924 49308 28980
rect 48860 28756 48916 28766
rect 48860 28754 49028 28756
rect 48860 28702 48862 28754
rect 48914 28702 49028 28754
rect 48860 28700 49028 28702
rect 48860 28690 48916 28700
rect 48244 20636 48356 20692
rect 48524 28532 48580 28542
rect 48524 20690 48580 28476
rect 48972 27746 49028 28700
rect 49308 28642 49364 28924
rect 49308 28590 49310 28642
rect 49362 28590 49364 28642
rect 49308 28578 49364 28590
rect 49420 28644 49476 28654
rect 49420 27858 49476 28588
rect 49420 27806 49422 27858
rect 49474 27806 49476 27858
rect 49420 27794 49476 27806
rect 48972 27694 48974 27746
rect 49026 27694 49028 27746
rect 48860 27636 48916 27646
rect 48860 27542 48916 27580
rect 48636 27524 48692 27534
rect 48636 27074 48692 27468
rect 48636 27022 48638 27074
rect 48690 27022 48692 27074
rect 48636 27010 48692 27022
rect 48748 26964 48804 26974
rect 48748 26870 48804 26908
rect 48860 26516 48916 26526
rect 48972 26516 49028 27694
rect 49420 27076 49476 27086
rect 48916 26460 49028 26516
rect 49196 27020 49420 27076
rect 48860 26422 48916 26460
rect 48860 26292 48916 26302
rect 48748 26236 48860 26292
rect 48636 26068 48692 26078
rect 48636 25618 48692 26012
rect 48636 25566 48638 25618
rect 48690 25566 48692 25618
rect 48636 25554 48692 25566
rect 48636 24948 48692 24958
rect 48748 24948 48804 26236
rect 48860 26226 48916 26236
rect 48972 26290 49028 26302
rect 48972 26238 48974 26290
rect 49026 26238 49028 26290
rect 48860 26066 48916 26078
rect 48860 26014 48862 26066
rect 48914 26014 48916 26066
rect 48860 25506 48916 26014
rect 48972 26068 49028 26238
rect 48972 26002 49028 26012
rect 49084 26180 49140 26190
rect 48972 25620 49028 25630
rect 48972 25526 49028 25564
rect 48860 25454 48862 25506
rect 48914 25454 48916 25506
rect 48860 25442 48916 25454
rect 49084 25506 49140 26124
rect 49084 25454 49086 25506
rect 49138 25454 49140 25506
rect 48748 24892 49028 24948
rect 48636 24050 48692 24892
rect 48972 24500 49028 24892
rect 49084 24724 49140 25454
rect 49196 24946 49252 27020
rect 49420 27010 49476 27020
rect 49196 24894 49198 24946
rect 49250 24894 49252 24946
rect 49196 24882 49252 24894
rect 49420 26404 49476 26414
rect 49420 25506 49476 26348
rect 49420 25454 49422 25506
rect 49474 25454 49476 25506
rect 49084 24668 49252 24724
rect 49196 24612 49252 24668
rect 49420 24722 49476 25454
rect 49420 24670 49422 24722
rect 49474 24670 49476 24722
rect 49420 24658 49476 24670
rect 49196 24546 49252 24556
rect 49084 24500 49140 24510
rect 48972 24498 49140 24500
rect 48972 24446 49086 24498
rect 49138 24446 49140 24498
rect 48972 24444 49140 24446
rect 49084 24434 49140 24444
rect 49420 24164 49476 24174
rect 48636 23998 48638 24050
rect 48690 23998 48692 24050
rect 48636 23604 48692 23998
rect 48636 23538 48692 23548
rect 49196 24108 49420 24164
rect 49084 23042 49140 23054
rect 49084 22990 49086 23042
rect 49138 22990 49140 23042
rect 49084 22932 49140 22990
rect 48748 21700 48804 21710
rect 48748 21252 48804 21644
rect 48860 21476 48916 21486
rect 48860 21382 48916 21420
rect 48748 21186 48804 21196
rect 48972 21362 49028 21374
rect 48972 21310 48974 21362
rect 49026 21310 49028 21362
rect 48972 20802 49028 21310
rect 48972 20750 48974 20802
rect 49026 20750 49028 20802
rect 48972 20738 49028 20750
rect 48524 20638 48526 20690
rect 48578 20638 48580 20690
rect 48188 20598 48244 20636
rect 48524 20626 48580 20638
rect 47628 20524 48132 20580
rect 47628 19234 47684 20524
rect 47628 19182 47630 19234
rect 47682 19182 47684 19234
rect 47628 19170 47684 19182
rect 47964 20132 48020 20142
rect 47516 19070 47518 19122
rect 47570 19070 47572 19122
rect 47516 19058 47572 19070
rect 47516 18450 47572 18462
rect 47516 18398 47518 18450
rect 47570 18398 47572 18450
rect 47516 18340 47572 18398
rect 47516 18274 47572 18284
rect 47628 18450 47684 18462
rect 47628 18398 47630 18450
rect 47682 18398 47684 18450
rect 47292 17388 47460 17444
rect 47292 16772 47348 17388
rect 47404 17220 47460 17230
rect 47628 17220 47684 18398
rect 47740 18452 47796 18462
rect 47740 18358 47796 18396
rect 47964 17666 48020 20076
rect 49084 19908 49140 22876
rect 48412 19234 48468 19246
rect 48412 19182 48414 19234
rect 48466 19182 48468 19234
rect 48300 19122 48356 19134
rect 48300 19070 48302 19122
rect 48354 19070 48356 19122
rect 48188 18676 48244 18686
rect 47964 17614 47966 17666
rect 48018 17614 48020 17666
rect 47964 17602 48020 17614
rect 48076 18452 48132 18462
rect 48076 17554 48132 18396
rect 48188 18450 48244 18620
rect 48188 18398 48190 18450
rect 48242 18398 48244 18450
rect 48188 18386 48244 18398
rect 48300 18116 48356 19070
rect 48412 18788 48468 19182
rect 48972 19236 49028 19246
rect 48972 19142 49028 19180
rect 49084 19124 49140 19852
rect 49196 19684 49252 24108
rect 49420 24098 49476 24108
rect 49532 23268 49588 29036
rect 49644 28532 49700 28542
rect 49644 28438 49700 28476
rect 49644 27860 49700 27870
rect 49644 26962 49700 27804
rect 49756 27300 49812 30716
rect 49980 30098 50036 30110
rect 49980 30046 49982 30098
rect 50034 30046 50036 30098
rect 49980 28868 50036 30046
rect 51100 29988 51156 29998
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 51100 29426 51156 29932
rect 51100 29374 51102 29426
rect 51154 29374 51156 29426
rect 51100 29362 51156 29374
rect 50988 29316 51044 29326
rect 50876 29260 50988 29316
rect 50540 29092 50596 29102
rect 49980 28812 50484 28868
rect 49868 28642 49924 28654
rect 49868 28590 49870 28642
rect 49922 28590 49924 28642
rect 49868 28532 49924 28590
rect 49868 28466 49924 28476
rect 50092 28642 50148 28654
rect 50092 28590 50094 28642
rect 50146 28590 50148 28642
rect 49980 28420 50036 28430
rect 49980 28326 50036 28364
rect 50092 27636 50148 28590
rect 50316 28642 50372 28654
rect 50316 28590 50318 28642
rect 50370 28590 50372 28642
rect 50316 28084 50372 28590
rect 50316 28018 50372 28028
rect 50316 27860 50372 27870
rect 50316 27766 50372 27804
rect 50428 27636 50484 28812
rect 50540 28642 50596 29036
rect 50540 28590 50542 28642
rect 50594 28590 50596 28642
rect 50540 28578 50596 28590
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50540 28084 50596 28094
rect 50540 27860 50596 28028
rect 50876 28082 50932 29260
rect 50988 29250 51044 29260
rect 50876 28030 50878 28082
rect 50930 28030 50932 28082
rect 50876 28018 50932 28030
rect 50988 28532 51044 28542
rect 50988 27970 51044 28476
rect 50988 27918 50990 27970
rect 51042 27918 51044 27970
rect 50540 27858 50932 27860
rect 50540 27806 50542 27858
rect 50594 27806 50932 27858
rect 50540 27804 50932 27806
rect 50540 27794 50596 27804
rect 50764 27636 50820 27646
rect 50428 27580 50596 27636
rect 50092 27570 50148 27580
rect 49756 27234 49812 27244
rect 50428 27300 50484 27310
rect 49868 27188 49924 27198
rect 49868 27186 50148 27188
rect 49868 27134 49870 27186
rect 49922 27134 50148 27186
rect 49868 27132 50148 27134
rect 49868 27122 49924 27132
rect 49644 26910 49646 26962
rect 49698 26910 49700 26962
rect 49644 26898 49700 26910
rect 49756 27074 49812 27086
rect 49756 27022 49758 27074
rect 49810 27022 49812 27074
rect 49756 26852 49812 27022
rect 50092 27074 50148 27132
rect 50092 27022 50094 27074
rect 50146 27022 50148 27074
rect 50092 27010 50148 27022
rect 50428 27074 50484 27244
rect 50428 27022 50430 27074
rect 50482 27022 50484 27074
rect 50428 27010 50484 27022
rect 50204 26964 50260 26974
rect 50092 26852 50260 26908
rect 49756 26796 49924 26852
rect 49756 26628 49812 26638
rect 49644 26404 49700 26414
rect 49644 26310 49700 26348
rect 49308 23212 49588 23268
rect 49644 25732 49700 25742
rect 49308 21812 49364 23212
rect 49532 23044 49588 23054
rect 49532 22820 49588 22988
rect 49532 22754 49588 22764
rect 49308 21810 49588 21812
rect 49308 21758 49310 21810
rect 49362 21758 49588 21810
rect 49308 21756 49588 21758
rect 49308 21746 49364 21756
rect 49308 20804 49364 20814
rect 49308 20802 49476 20804
rect 49308 20750 49310 20802
rect 49362 20750 49476 20802
rect 49308 20748 49476 20750
rect 49308 20738 49364 20748
rect 49196 19618 49252 19628
rect 49084 19058 49140 19068
rect 49196 19236 49252 19246
rect 48412 18722 48468 18732
rect 48860 18452 48916 18462
rect 48860 18358 48916 18396
rect 48300 18050 48356 18060
rect 48076 17502 48078 17554
rect 48130 17502 48132 17554
rect 48076 17490 48132 17502
rect 48412 18004 48468 18014
rect 47404 16994 47460 17164
rect 47404 16942 47406 16994
rect 47458 16942 47460 16994
rect 47404 16930 47460 16942
rect 47516 17164 47684 17220
rect 48300 17442 48356 17454
rect 48300 17390 48302 17442
rect 48354 17390 48356 17442
rect 47292 15986 47348 16716
rect 47516 16210 47572 17164
rect 47628 16996 47684 17006
rect 47628 16902 47684 16940
rect 47852 16884 47908 16894
rect 47852 16790 47908 16828
rect 48076 16884 48132 16894
rect 48076 16790 48132 16828
rect 48300 16548 48356 17390
rect 48300 16482 48356 16492
rect 48412 17108 48468 17948
rect 48860 17668 48916 17678
rect 48860 17574 48916 17612
rect 49196 17554 49252 19180
rect 49420 18676 49476 20748
rect 49532 20802 49588 21756
rect 49644 21362 49700 25676
rect 49644 21310 49646 21362
rect 49698 21310 49700 21362
rect 49644 21298 49700 21310
rect 49532 20750 49534 20802
rect 49586 20750 49588 20802
rect 49532 20738 49588 20750
rect 49756 19348 49812 26572
rect 49868 26402 49924 26796
rect 49868 26350 49870 26402
rect 49922 26350 49924 26402
rect 49868 26180 49924 26350
rect 49868 26114 49924 26124
rect 50092 25956 50148 26852
rect 50540 26850 50596 27580
rect 50540 26798 50542 26850
rect 50594 26798 50596 26850
rect 50540 26786 50596 26798
rect 50652 27076 50708 27086
rect 50764 27076 50820 27580
rect 50652 27074 50820 27076
rect 50652 27022 50654 27074
rect 50706 27022 50820 27074
rect 50652 27020 50820 27022
rect 50876 27074 50932 27804
rect 50988 27636 51044 27918
rect 50988 27300 51044 27580
rect 51100 28418 51156 28430
rect 51100 28366 51102 28418
rect 51154 28366 51156 28418
rect 51100 27524 51156 28366
rect 51436 28084 51492 38612
rect 51996 30436 52052 30446
rect 51772 29316 51828 29326
rect 51772 29222 51828 29260
rect 51436 28018 51492 28028
rect 51100 27458 51156 27468
rect 51212 27858 51268 27870
rect 51212 27806 51214 27858
rect 51266 27806 51268 27858
rect 50988 27234 51044 27244
rect 51212 27300 51268 27806
rect 51772 27748 51828 27758
rect 51772 27654 51828 27692
rect 51212 27234 51268 27244
rect 51548 27524 51604 27534
rect 50876 27022 50878 27074
rect 50930 27022 50932 27074
rect 50652 26852 50708 27020
rect 50652 26786 50708 26796
rect 50876 26740 50932 27022
rect 51436 27076 51492 27086
rect 51436 26982 51492 27020
rect 51100 26962 51156 26974
rect 51100 26910 51102 26962
rect 51154 26910 51156 26962
rect 50988 26740 51044 26750
rect 50556 26684 50820 26694
rect 50876 26684 50988 26740
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50988 26674 51044 26684
rect 50556 26618 50820 26628
rect 49868 25900 50148 25956
rect 50204 26514 50260 26526
rect 50204 26462 50206 26514
rect 50258 26462 50260 26514
rect 49868 25060 49924 25900
rect 50092 25508 50148 25546
rect 50092 25442 50148 25452
rect 49868 25004 50148 25060
rect 49868 24612 49924 24622
rect 49868 24518 49924 24556
rect 49868 23154 49924 23166
rect 49868 23102 49870 23154
rect 49922 23102 49924 23154
rect 49868 22484 49924 23102
rect 49868 22418 49924 22428
rect 50092 23154 50148 25004
rect 50204 24164 50260 26462
rect 50316 26516 50372 26526
rect 50316 26290 50372 26460
rect 50764 26516 50820 26526
rect 50316 26238 50318 26290
rect 50370 26238 50372 26290
rect 50316 26226 50372 26238
rect 50652 26404 50708 26414
rect 50652 25620 50708 26348
rect 50764 26402 50820 26460
rect 50764 26350 50766 26402
rect 50818 26350 50820 26402
rect 50764 26338 50820 26350
rect 50988 26402 51044 26414
rect 50988 26350 50990 26402
rect 51042 26350 51044 26402
rect 50876 26292 50932 26302
rect 50876 26198 50932 26236
rect 50876 26068 50932 26078
rect 50764 25620 50820 25630
rect 50652 25564 50764 25620
rect 50540 25508 50596 25518
rect 50540 25414 50596 25452
rect 50764 25506 50820 25564
rect 50876 25618 50932 26012
rect 50876 25566 50878 25618
rect 50930 25566 50932 25618
rect 50876 25554 50932 25566
rect 50764 25454 50766 25506
rect 50818 25454 50820 25506
rect 50764 25442 50820 25454
rect 50316 25396 50372 25406
rect 50316 25302 50372 25340
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50764 24948 50820 24958
rect 50652 24892 50764 24948
rect 50652 24834 50708 24892
rect 50764 24882 50820 24892
rect 50652 24782 50654 24834
rect 50706 24782 50708 24834
rect 50652 24770 50708 24782
rect 50428 24724 50484 24734
rect 50988 24724 51044 26350
rect 51100 25508 51156 26910
rect 51100 25442 51156 25452
rect 51548 25508 51604 27468
rect 51772 27300 51828 27310
rect 51772 27206 51828 27244
rect 51996 27300 52052 30380
rect 52108 30322 52164 30334
rect 52108 30270 52110 30322
rect 52162 30270 52164 30322
rect 52108 29540 52164 30270
rect 54796 30212 54852 30222
rect 52780 29988 52836 29998
rect 52780 29894 52836 29932
rect 54124 29988 54180 29998
rect 54124 29894 54180 29932
rect 52108 29474 52164 29484
rect 54572 29540 54628 29550
rect 54572 29446 54628 29484
rect 53900 29316 53956 29326
rect 53900 29222 53956 29260
rect 54460 29202 54516 29214
rect 54460 29150 54462 29202
rect 54514 29150 54516 29202
rect 53788 29092 53844 29102
rect 53004 28644 53060 28654
rect 53004 28550 53060 28588
rect 53452 28644 53508 28654
rect 53452 28550 53508 28588
rect 53228 27860 53284 27870
rect 53228 27766 53284 27804
rect 53340 27858 53396 27870
rect 53340 27806 53342 27858
rect 53394 27806 53396 27858
rect 51996 27234 52052 27244
rect 52108 27636 52164 27646
rect 52108 27076 52164 27580
rect 51996 27020 52164 27076
rect 52668 27636 52724 27646
rect 51660 26962 51716 26974
rect 51660 26910 51662 26962
rect 51714 26910 51716 26962
rect 51660 25732 51716 26910
rect 51884 26740 51940 26750
rect 51884 26402 51940 26684
rect 51996 26514 52052 27020
rect 51996 26462 51998 26514
rect 52050 26462 52052 26514
rect 51996 26450 52052 26462
rect 51884 26350 51886 26402
rect 51938 26350 51940 26402
rect 51884 25844 51940 26350
rect 52108 26068 52164 26078
rect 52108 25974 52164 26012
rect 51884 25788 52276 25844
rect 51660 25666 51716 25676
rect 51772 25508 51828 25518
rect 51548 25506 51828 25508
rect 51548 25454 51774 25506
rect 51826 25454 51828 25506
rect 51548 25452 51828 25454
rect 51324 25282 51380 25294
rect 51324 25230 51326 25282
rect 51378 25230 51380 25282
rect 51324 25060 51380 25230
rect 51324 24994 51380 25004
rect 51548 24948 51604 25452
rect 51772 25442 51828 25452
rect 52108 25396 52164 25406
rect 51548 24882 51604 24892
rect 51996 25340 52108 25396
rect 50428 24630 50484 24668
rect 50764 24668 51044 24724
rect 51100 24722 51156 24734
rect 51100 24670 51102 24722
rect 51154 24670 51156 24722
rect 50540 24610 50596 24622
rect 50540 24558 50542 24610
rect 50594 24558 50596 24610
rect 50204 24098 50260 24108
rect 50428 24164 50484 24174
rect 50428 24070 50484 24108
rect 50092 23102 50094 23154
rect 50146 23102 50148 23154
rect 49980 21474 50036 21486
rect 49980 21422 49982 21474
rect 50034 21422 50036 21474
rect 49868 21362 49924 21374
rect 49868 21310 49870 21362
rect 49922 21310 49924 21362
rect 49868 20802 49924 21310
rect 49868 20750 49870 20802
rect 49922 20750 49924 20802
rect 49868 20738 49924 20750
rect 49980 20692 50036 21422
rect 50092 21476 50148 23102
rect 50204 23938 50260 23950
rect 50204 23886 50206 23938
rect 50258 23886 50260 23938
rect 50204 22260 50260 23886
rect 50540 23716 50596 24558
rect 50764 23940 50820 24668
rect 51100 24612 51156 24670
rect 51212 24612 51268 24622
rect 51100 24556 51212 24612
rect 51212 24546 51268 24556
rect 51660 24612 51716 24622
rect 50876 24498 50932 24510
rect 50876 24446 50878 24498
rect 50930 24446 50932 24498
rect 50876 24050 50932 24446
rect 51548 24498 51604 24510
rect 51548 24446 51550 24498
rect 51602 24446 51604 24498
rect 50876 23998 50878 24050
rect 50930 23998 50932 24050
rect 50876 23986 50932 23998
rect 50988 24276 51044 24286
rect 50988 23940 51044 24220
rect 51548 24164 51604 24446
rect 51660 24276 51716 24556
rect 51996 24610 52052 25340
rect 52108 25330 52164 25340
rect 52220 24946 52276 25788
rect 52220 24894 52222 24946
rect 52274 24894 52276 24946
rect 52220 24882 52276 24894
rect 51996 24558 51998 24610
rect 52050 24558 52052 24610
rect 51996 24546 52052 24558
rect 52556 24500 52612 24510
rect 52556 24406 52612 24444
rect 51660 24220 52164 24276
rect 51100 23940 51156 23950
rect 50988 23938 51156 23940
rect 50988 23886 51102 23938
rect 51154 23886 51156 23938
rect 50988 23884 51156 23886
rect 50764 23846 50820 23884
rect 51100 23874 51156 23884
rect 51548 23938 51604 24108
rect 51548 23886 51550 23938
rect 51602 23886 51604 23938
rect 51548 23874 51604 23886
rect 51772 23940 51828 23950
rect 51772 23846 51828 23884
rect 50428 23660 50596 23716
rect 50876 23716 50932 23726
rect 51324 23716 51380 23726
rect 50876 23714 51156 23716
rect 50876 23662 50878 23714
rect 50930 23662 51156 23714
rect 50876 23660 51156 23662
rect 50316 23268 50372 23278
rect 50316 23154 50372 23212
rect 50316 23102 50318 23154
rect 50370 23102 50372 23154
rect 50316 23090 50372 23102
rect 50204 22194 50260 22204
rect 50204 21868 50372 21924
rect 50204 21812 50260 21868
rect 50204 21746 50260 21756
rect 50316 21810 50372 21868
rect 50316 21758 50318 21810
rect 50370 21758 50372 21810
rect 50316 21746 50372 21758
rect 50428 21812 50484 23660
rect 50876 23650 50932 23660
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50876 23380 50932 23390
rect 50876 23378 51044 23380
rect 50876 23326 50878 23378
rect 50930 23326 51044 23378
rect 50876 23324 51044 23326
rect 50876 23314 50932 23324
rect 50764 23156 50820 23166
rect 50652 23154 50820 23156
rect 50652 23102 50766 23154
rect 50818 23102 50820 23154
rect 50652 23100 50820 23102
rect 50540 23042 50596 23054
rect 50540 22990 50542 23042
rect 50594 22990 50596 23042
rect 50540 22820 50596 22990
rect 50652 22932 50708 23100
rect 50764 23090 50820 23100
rect 50876 23156 50932 23166
rect 50652 22866 50708 22876
rect 50876 22932 50932 23100
rect 50988 23154 51044 23324
rect 50988 23102 50990 23154
rect 51042 23102 51044 23154
rect 50988 23090 51044 23102
rect 50876 22866 50932 22876
rect 51100 22820 51156 23660
rect 51212 23604 51268 23614
rect 51212 23044 51268 23548
rect 51324 23378 51380 23660
rect 51660 23714 51716 23726
rect 51660 23662 51662 23714
rect 51714 23662 51716 23714
rect 51324 23326 51326 23378
rect 51378 23326 51380 23378
rect 51324 23314 51380 23326
rect 51436 23604 51492 23614
rect 51324 23044 51380 23054
rect 51212 22988 51324 23044
rect 51324 22978 51380 22988
rect 51436 22932 51492 23548
rect 51548 23492 51604 23502
rect 51548 23378 51604 23436
rect 51548 23326 51550 23378
rect 51602 23326 51604 23378
rect 51548 23314 51604 23326
rect 51660 23380 51716 23662
rect 51996 23716 52052 23726
rect 51660 23314 51716 23324
rect 51772 23604 51828 23614
rect 51436 22876 51604 22932
rect 51100 22764 51492 22820
rect 50540 22754 50596 22764
rect 51324 22596 51380 22606
rect 51324 22502 51380 22540
rect 51436 22482 51492 22764
rect 51436 22430 51438 22482
rect 51490 22430 51492 22482
rect 51436 22418 51492 22430
rect 51548 22484 51604 22876
rect 51548 22418 51604 22428
rect 51660 22930 51716 22942
rect 51660 22878 51662 22930
rect 51714 22878 51716 22930
rect 50988 22372 51044 22382
rect 50876 22316 50988 22372
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50428 21756 50708 21812
rect 50540 21586 50596 21598
rect 50540 21534 50542 21586
rect 50594 21534 50596 21586
rect 50540 21476 50596 21534
rect 50092 21420 50596 21476
rect 50204 21028 50260 21038
rect 50204 20934 50260 20972
rect 50092 20692 50148 20702
rect 49980 20690 50148 20692
rect 49980 20638 50094 20690
rect 50146 20638 50148 20690
rect 49980 20636 50148 20638
rect 49868 19348 49924 19358
rect 49756 19346 49924 19348
rect 49756 19294 49870 19346
rect 49922 19294 49924 19346
rect 49756 19292 49924 19294
rect 49868 19282 49924 19292
rect 49532 19012 49588 19022
rect 49532 18918 49588 18956
rect 49756 19010 49812 19022
rect 49756 18958 49758 19010
rect 49810 18958 49812 19010
rect 49532 18676 49588 18686
rect 49420 18674 49588 18676
rect 49420 18622 49534 18674
rect 49586 18622 49588 18674
rect 49420 18620 49588 18622
rect 49308 18450 49364 18462
rect 49308 18398 49310 18450
rect 49362 18398 49364 18450
rect 49308 18116 49364 18398
rect 49420 18340 49476 18620
rect 49532 18610 49588 18620
rect 49756 18676 49812 18958
rect 49980 19012 50036 19022
rect 49980 18918 50036 18956
rect 49756 18610 49812 18620
rect 49420 18274 49476 18284
rect 49980 18450 50036 18462
rect 49980 18398 49982 18450
rect 50034 18398 50036 18450
rect 49308 18050 49364 18060
rect 49532 17668 49588 17678
rect 49532 17574 49588 17612
rect 49196 17502 49198 17554
rect 49250 17502 49252 17554
rect 49196 17490 49252 17502
rect 49868 17556 49924 17566
rect 49868 17462 49924 17500
rect 48412 16322 48468 17052
rect 49868 17108 49924 17118
rect 49868 17014 49924 17052
rect 48524 16996 48580 17006
rect 48748 16996 48804 17006
rect 48580 16940 48692 16996
rect 48524 16930 48580 16940
rect 48636 16772 48692 16940
rect 48748 16994 48916 16996
rect 48748 16942 48750 16994
rect 48802 16942 48916 16994
rect 48748 16940 48916 16942
rect 48748 16930 48804 16940
rect 48860 16772 48916 16940
rect 48636 16716 48804 16772
rect 48412 16270 48414 16322
rect 48466 16270 48468 16322
rect 48412 16258 48468 16270
rect 47516 16158 47518 16210
rect 47570 16158 47572 16210
rect 47516 16146 47572 16158
rect 47292 15934 47294 15986
rect 47346 15934 47348 15986
rect 47292 15922 47348 15934
rect 48076 16098 48132 16110
rect 48636 16100 48692 16110
rect 48076 16046 48078 16098
rect 48130 16046 48132 16098
rect 47180 15810 47236 15820
rect 47404 15876 47460 15886
rect 47404 15782 47460 15820
rect 47628 15874 47684 15886
rect 47628 15822 47630 15874
rect 47682 15822 47684 15874
rect 46396 14914 46452 14924
rect 46508 15092 46900 15148
rect 47628 15764 47684 15822
rect 48076 15764 48132 16046
rect 47628 15708 48076 15764
rect 46396 13972 46452 13982
rect 46396 13878 46452 13916
rect 45948 12238 45950 12290
rect 46002 12238 46004 12290
rect 45948 11618 46004 12238
rect 45948 11566 45950 11618
rect 46002 11566 46004 11618
rect 45948 11554 46004 11566
rect 46060 12348 46228 12404
rect 46396 12516 46452 12526
rect 46396 12402 46452 12460
rect 46396 12350 46398 12402
rect 46450 12350 46452 12402
rect 45164 11106 45220 11116
rect 45500 11170 45556 11182
rect 45500 11118 45502 11170
rect 45554 11118 45556 11170
rect 45052 10220 45332 10276
rect 45052 10052 45108 10062
rect 44940 10050 45108 10052
rect 44940 9998 45054 10050
rect 45106 9998 45108 10050
rect 44940 9996 45108 9998
rect 45052 9986 45108 9996
rect 44828 9874 44884 9884
rect 45164 9940 45220 9950
rect 45164 9846 45220 9884
rect 45276 9716 45332 10220
rect 45500 10052 45556 11118
rect 45836 11172 45892 11182
rect 45836 11078 45892 11116
rect 46060 10836 46116 12348
rect 46396 12338 46452 12350
rect 46172 12180 46228 12190
rect 46172 12086 46228 12124
rect 46284 12066 46340 12078
rect 46284 12014 46286 12066
rect 46338 12014 46340 12066
rect 46284 11396 46340 12014
rect 46060 10770 46116 10780
rect 46172 11340 46340 11396
rect 46396 11618 46452 11630
rect 46396 11566 46398 11618
rect 46450 11566 46452 11618
rect 46172 10722 46228 11340
rect 46284 11172 46340 11182
rect 46396 11172 46452 11566
rect 46284 11170 46452 11172
rect 46284 11118 46286 11170
rect 46338 11118 46452 11170
rect 46284 11116 46452 11118
rect 46284 11106 46340 11116
rect 46172 10670 46174 10722
rect 46226 10670 46228 10722
rect 46172 10658 46228 10670
rect 46060 10610 46116 10622
rect 46060 10558 46062 10610
rect 46114 10558 46116 10610
rect 45500 9986 45556 9996
rect 45612 10498 45668 10510
rect 45612 10446 45614 10498
rect 45666 10446 45668 10498
rect 44716 9090 44772 9100
rect 45164 9660 45332 9716
rect 45388 9826 45444 9838
rect 45388 9774 45390 9826
rect 45442 9774 45444 9826
rect 45388 9716 45444 9774
rect 45500 9716 45556 9726
rect 45388 9660 45500 9716
rect 44380 8194 44436 8204
rect 45052 8260 45108 8270
rect 45052 8166 45108 8204
rect 44268 7980 44436 8036
rect 44044 7868 44324 7924
rect 43932 7756 44212 7812
rect 43708 7588 43764 7598
rect 43708 6916 43764 7532
rect 43596 6860 43764 6916
rect 43596 5684 43652 6860
rect 43708 6692 43764 6702
rect 43708 5906 43764 6636
rect 44044 6580 44100 6590
rect 43708 5854 43710 5906
rect 43762 5854 43764 5906
rect 43708 5842 43764 5854
rect 43932 6578 44100 6580
rect 43932 6526 44046 6578
rect 44098 6526 44100 6578
rect 43932 6524 44100 6526
rect 43932 6468 43988 6524
rect 44044 6514 44100 6524
rect 44156 6580 44212 7756
rect 44156 6486 44212 6524
rect 43596 5628 43764 5684
rect 43708 5122 43764 5628
rect 43708 5070 43710 5122
rect 43762 5070 43764 5122
rect 43708 5058 43764 5070
rect 43596 5012 43652 5022
rect 43596 3556 43652 4956
rect 43932 4788 43988 6412
rect 44268 6468 44324 7868
rect 44380 6804 44436 7980
rect 44940 7700 44996 7710
rect 44940 7362 44996 7644
rect 44940 7310 44942 7362
rect 44994 7310 44996 7362
rect 44940 7298 44996 7310
rect 44380 6738 44436 6748
rect 44940 7028 44996 7038
rect 45164 7028 45220 9660
rect 45500 9650 45556 9660
rect 45500 9380 45556 9390
rect 45276 8372 45332 8382
rect 45332 8316 45444 8372
rect 45276 8306 45332 8316
rect 45276 8036 45332 8046
rect 45276 7942 45332 7980
rect 45388 7474 45444 8316
rect 45500 8258 45556 9324
rect 45612 9268 45668 10446
rect 45948 10052 46004 10062
rect 46060 10052 46116 10558
rect 45948 10050 46116 10052
rect 45948 9998 45950 10050
rect 46002 9998 46116 10050
rect 45948 9996 46116 9998
rect 45948 9986 46004 9996
rect 46508 9940 46564 15092
rect 47180 14868 47236 14878
rect 46844 13634 46900 13646
rect 46844 13582 46846 13634
rect 46898 13582 46900 13634
rect 46844 13524 46900 13582
rect 47068 13524 47124 13534
rect 46844 13522 47124 13524
rect 46844 13470 47070 13522
rect 47122 13470 47124 13522
rect 46844 13468 47124 13470
rect 46956 12850 47012 12862
rect 46956 12798 46958 12850
rect 47010 12798 47012 12850
rect 46956 12404 47012 12798
rect 46956 12338 47012 12348
rect 46620 12180 46676 12190
rect 46620 12086 46676 12124
rect 46956 11170 47012 11182
rect 46956 11118 46958 11170
rect 47010 11118 47012 11170
rect 46844 10834 46900 10846
rect 46844 10782 46846 10834
rect 46898 10782 46900 10834
rect 46732 10612 46788 10622
rect 46732 10388 46788 10556
rect 46732 10322 46788 10332
rect 46284 9884 46564 9940
rect 45836 9714 45892 9726
rect 45836 9662 45838 9714
rect 45890 9662 45892 9714
rect 45836 9492 45892 9662
rect 45948 9716 46004 9726
rect 46284 9716 46340 9884
rect 46004 9660 46340 9716
rect 45948 9622 46004 9660
rect 45836 9426 45892 9436
rect 46396 9602 46452 9614
rect 46396 9550 46398 9602
rect 46450 9550 46452 9602
rect 46396 9380 46452 9550
rect 46508 9380 46564 9884
rect 46732 10052 46788 10062
rect 46732 9826 46788 9996
rect 46732 9774 46734 9826
rect 46786 9774 46788 9826
rect 46732 9762 46788 9774
rect 46620 9714 46676 9726
rect 46620 9662 46622 9714
rect 46674 9662 46676 9714
rect 46620 9492 46676 9662
rect 46620 9436 46788 9492
rect 46508 9324 46676 9380
rect 46396 9314 46452 9324
rect 45612 9202 45668 9212
rect 46284 9156 46340 9166
rect 46508 9156 46564 9166
rect 46340 9100 46452 9156
rect 46284 9090 46340 9100
rect 45500 8206 45502 8258
rect 45554 8206 45556 8258
rect 45500 8194 45556 8206
rect 45612 8484 45668 8494
rect 45612 8036 45668 8428
rect 45724 8260 45780 8270
rect 45724 8166 45780 8204
rect 45388 7422 45390 7474
rect 45442 7422 45444 7474
rect 45388 7410 45444 7422
rect 45500 7980 45668 8036
rect 46284 8146 46340 8158
rect 46284 8094 46286 8146
rect 46338 8094 46340 8146
rect 44996 6972 45220 7028
rect 44380 6580 44436 6590
rect 44380 6486 44436 6524
rect 44268 6402 44324 6412
rect 44604 6468 44660 6478
rect 44828 6468 44884 6478
rect 44660 6466 44884 6468
rect 44660 6414 44830 6466
rect 44882 6414 44884 6466
rect 44660 6412 44884 6414
rect 44604 6402 44660 6412
rect 44828 6402 44884 6412
rect 43932 4722 43988 4732
rect 44044 6356 44100 6366
rect 43708 4228 43764 4238
rect 43708 4134 43764 4172
rect 43708 3556 43764 3566
rect 43596 3554 43764 3556
rect 43596 3502 43710 3554
rect 43762 3502 43764 3554
rect 43596 3500 43764 3502
rect 43708 3490 43764 3500
rect 43932 3444 43988 3454
rect 44044 3444 44100 6300
rect 44604 5682 44660 5694
rect 44604 5630 44606 5682
rect 44658 5630 44660 5682
rect 44604 4452 44660 5630
rect 44604 4386 44660 4396
rect 43932 3442 44100 3444
rect 43932 3390 43934 3442
rect 43986 3390 44100 3442
rect 43932 3388 44100 3390
rect 43932 3378 43988 3388
rect 44156 924 44436 980
rect 44156 800 44212 924
rect 43036 700 43540 756
rect 44128 0 44240 800
rect 44380 756 44436 924
rect 44940 756 44996 6972
rect 45052 6804 45108 6814
rect 45052 6690 45108 6748
rect 45052 6638 45054 6690
rect 45106 6638 45108 6690
rect 45052 6626 45108 6638
rect 45388 6690 45444 6702
rect 45388 6638 45390 6690
rect 45442 6638 45444 6690
rect 45388 6580 45444 6638
rect 45388 6514 45444 6524
rect 45388 6244 45444 6254
rect 45276 5908 45332 5918
rect 45276 5346 45332 5852
rect 45276 5294 45278 5346
rect 45330 5294 45332 5346
rect 45276 5282 45332 5294
rect 45388 5572 45444 6188
rect 45388 5346 45444 5516
rect 45388 5294 45390 5346
rect 45442 5294 45444 5346
rect 45388 5282 45444 5294
rect 45500 5124 45556 7980
rect 46060 7364 46116 7374
rect 45612 7362 46116 7364
rect 45612 7310 46062 7362
rect 46114 7310 46116 7362
rect 45612 7308 46116 7310
rect 45612 6802 45668 7308
rect 46060 7298 46116 7308
rect 45612 6750 45614 6802
rect 45666 6750 45668 6802
rect 45612 6738 45668 6750
rect 45836 7140 45892 7150
rect 45836 6690 45892 7084
rect 46284 7028 46340 8094
rect 46284 6962 46340 6972
rect 45836 6638 45838 6690
rect 45890 6638 45892 6690
rect 45836 6626 45892 6638
rect 45948 6692 46004 6702
rect 45948 6598 46004 6636
rect 46396 6692 46452 9100
rect 46396 6626 46452 6636
rect 46508 6580 46564 9100
rect 46620 8930 46676 9324
rect 46620 8878 46622 8930
rect 46674 8878 46676 8930
rect 46620 8866 46676 8878
rect 46732 7700 46788 9436
rect 46732 7634 46788 7644
rect 46508 6578 46676 6580
rect 46508 6526 46510 6578
rect 46562 6526 46676 6578
rect 46508 6524 46676 6526
rect 46508 6514 46564 6524
rect 46508 5794 46564 5806
rect 46508 5742 46510 5794
rect 46562 5742 46564 5794
rect 45612 5348 45668 5358
rect 45668 5292 45892 5348
rect 45612 5254 45668 5292
rect 45724 5124 45780 5134
rect 45500 5122 45780 5124
rect 45500 5070 45726 5122
rect 45778 5070 45780 5122
rect 45500 5068 45780 5070
rect 45724 5058 45780 5068
rect 45836 4226 45892 5292
rect 46284 5234 46340 5246
rect 46284 5182 46286 5234
rect 46338 5182 46340 5234
rect 46284 4450 46340 5182
rect 46508 4564 46564 5742
rect 46508 4498 46564 4508
rect 46284 4398 46286 4450
rect 46338 4398 46340 4450
rect 46284 4386 46340 4398
rect 45836 4174 45838 4226
rect 45890 4174 45892 4226
rect 45836 4162 45892 4174
rect 45500 3666 45556 3678
rect 45500 3614 45502 3666
rect 45554 3614 45556 3666
rect 45500 800 45556 3614
rect 46620 3388 46676 6524
rect 46844 3554 46900 10782
rect 46956 8036 47012 11118
rect 47068 9604 47124 13468
rect 47180 12516 47236 14812
rect 47404 13634 47460 13646
rect 47404 13582 47406 13634
rect 47458 13582 47460 13634
rect 47180 12402 47236 12460
rect 47180 12350 47182 12402
rect 47234 12350 47236 12402
rect 47180 12338 47236 12350
rect 47292 12740 47348 12750
rect 47180 9604 47236 9614
rect 47068 9602 47236 9604
rect 47068 9550 47182 9602
rect 47234 9550 47236 9602
rect 47068 9548 47236 9550
rect 47068 8372 47124 9548
rect 47180 9538 47236 9548
rect 47292 9492 47348 12684
rect 47404 11396 47460 13582
rect 47516 12516 47572 12526
rect 47516 12402 47572 12460
rect 47516 12350 47518 12402
rect 47570 12350 47572 12402
rect 47516 12338 47572 12350
rect 47628 11396 47684 15708
rect 48076 15670 48132 15708
rect 48188 16044 48636 16100
rect 48188 15876 48244 16044
rect 48636 16006 48692 16044
rect 48188 15202 48244 15820
rect 48188 15150 48190 15202
rect 48242 15150 48244 15202
rect 48188 15148 48244 15150
rect 47964 15092 48244 15148
rect 48300 15540 48356 15550
rect 48300 15148 48356 15484
rect 48748 15148 48804 16716
rect 48860 16706 48916 16716
rect 49084 16882 49140 16894
rect 49084 16830 49086 16882
rect 49138 16830 49140 16882
rect 49084 16100 49140 16830
rect 49532 16884 49588 16894
rect 49196 16100 49252 16110
rect 49084 16098 49252 16100
rect 49084 16046 49198 16098
rect 49250 16046 49252 16098
rect 49084 16044 49252 16046
rect 49196 15876 49252 16044
rect 49532 16098 49588 16828
rect 49868 16548 49924 16558
rect 49532 16046 49534 16098
rect 49586 16046 49588 16098
rect 49532 16034 49588 16046
rect 49644 16324 49700 16334
rect 49196 15810 49252 15820
rect 48972 15764 49028 15774
rect 48860 15540 48916 15550
rect 48860 15446 48916 15484
rect 48972 15426 49028 15708
rect 49644 15652 49700 16268
rect 49756 16100 49812 16110
rect 49756 15986 49812 16044
rect 49868 16098 49924 16492
rect 49868 16046 49870 16098
rect 49922 16046 49924 16098
rect 49868 16034 49924 16046
rect 49756 15934 49758 15986
rect 49810 15934 49812 15986
rect 49756 15922 49812 15934
rect 48972 15374 48974 15426
rect 49026 15374 49028 15426
rect 48972 15362 49028 15374
rect 49420 15596 49700 15652
rect 49420 15540 49476 15596
rect 49420 15148 49476 15484
rect 49980 15540 50036 18398
rect 50092 18452 50148 20636
rect 50204 20132 50260 20142
rect 50316 20132 50372 21420
rect 50652 21026 50708 21756
rect 50876 21252 50932 22316
rect 50988 22278 51044 22316
rect 51548 22258 51604 22270
rect 51548 22206 51550 22258
rect 51602 22206 51604 22258
rect 51548 22148 51604 22206
rect 51548 22082 51604 22092
rect 51660 22036 51716 22878
rect 51660 21970 51716 21980
rect 51772 21812 51828 23548
rect 51436 21756 51828 21812
rect 51884 23044 51940 23054
rect 51100 21700 51156 21710
rect 51100 21606 51156 21644
rect 50988 21586 51044 21598
rect 50988 21534 50990 21586
rect 51042 21534 51044 21586
rect 50988 21364 51044 21534
rect 51212 21588 51268 21598
rect 51212 21494 51268 21532
rect 51324 21476 51380 21486
rect 51324 21364 51380 21420
rect 50988 21308 51380 21364
rect 50876 21196 51156 21252
rect 50652 20974 50654 21026
rect 50706 20974 50708 21026
rect 50652 20962 50708 20974
rect 51100 20692 51156 21196
rect 51324 20804 51380 20814
rect 51324 20710 51380 20748
rect 50988 20636 51156 20692
rect 50764 20580 50820 20618
rect 50764 20514 50820 20524
rect 50876 20578 50932 20590
rect 50876 20526 50878 20578
rect 50930 20526 50932 20578
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50260 20076 50372 20132
rect 50204 20066 50260 20076
rect 50876 20020 50932 20526
rect 50876 19954 50932 19964
rect 50988 19906 51044 20636
rect 51436 20580 51492 21756
rect 51660 21586 51716 21598
rect 51660 21534 51662 21586
rect 51714 21534 51716 21586
rect 51660 20916 51716 21534
rect 51772 21588 51828 21598
rect 51772 21474 51828 21532
rect 51772 21422 51774 21474
rect 51826 21422 51828 21474
rect 51772 21410 51828 21422
rect 51660 20850 51716 20860
rect 51772 21252 51828 21262
rect 51660 20692 51716 20702
rect 51660 20598 51716 20636
rect 51772 20690 51828 21196
rect 51772 20638 51774 20690
rect 51826 20638 51828 20690
rect 51772 20626 51828 20638
rect 50988 19854 50990 19906
rect 51042 19854 51044 19906
rect 50988 19842 51044 19854
rect 51324 20524 51492 20580
rect 51548 20578 51604 20590
rect 51548 20526 51550 20578
rect 51602 20526 51604 20578
rect 50204 19684 50260 19694
rect 50204 19122 50260 19628
rect 51324 19572 51380 20524
rect 51548 20468 51604 20526
rect 51436 20412 51604 20468
rect 51436 19796 51492 20412
rect 51884 20356 51940 22988
rect 51996 21812 52052 23660
rect 52108 23044 52164 24220
rect 52220 23940 52276 23950
rect 52220 23938 52388 23940
rect 52220 23886 52222 23938
rect 52274 23886 52388 23938
rect 52220 23884 52388 23886
rect 52220 23492 52276 23884
rect 52332 23716 52388 23884
rect 52332 23650 52388 23660
rect 52220 23426 52276 23436
rect 52668 23380 52724 27580
rect 53340 27076 53396 27806
rect 53340 27010 53396 27020
rect 53676 26852 53732 26862
rect 52780 26402 52836 26414
rect 52780 26350 52782 26402
rect 52834 26350 52836 26402
rect 52780 25620 52836 26350
rect 53116 26404 53172 26414
rect 53116 26310 53172 26348
rect 52892 26068 52948 26078
rect 52948 26012 53172 26068
rect 52892 26002 52948 26012
rect 52780 25554 52836 25564
rect 53116 25620 53172 26012
rect 53116 25618 53284 25620
rect 53116 25566 53118 25618
rect 53170 25566 53284 25618
rect 53116 25564 53284 25566
rect 53116 25554 53172 25564
rect 53004 25508 53060 25518
rect 53004 25414 53060 25452
rect 52780 24612 52836 24622
rect 52780 24610 52948 24612
rect 52780 24558 52782 24610
rect 52834 24558 52948 24610
rect 52780 24556 52948 24558
rect 52780 24546 52836 24556
rect 52780 24164 52836 24174
rect 52780 24050 52836 24108
rect 52780 23998 52782 24050
rect 52834 23998 52836 24050
rect 52780 23986 52836 23998
rect 52892 23604 52948 24556
rect 52892 23538 52948 23548
rect 52668 23314 52724 23324
rect 52780 23492 52836 23502
rect 52556 23156 52612 23166
rect 52108 22596 52164 22988
rect 52332 23044 52388 23054
rect 52220 22596 52276 22606
rect 52108 22540 52220 22596
rect 52220 22482 52276 22540
rect 52220 22430 52222 22482
rect 52274 22430 52276 22482
rect 52220 22418 52276 22430
rect 52332 22148 52388 22988
rect 52332 22082 52388 22092
rect 52444 22932 52500 22942
rect 52108 22036 52164 22046
rect 52164 21980 52276 22036
rect 52108 21970 52164 21980
rect 51996 21746 52052 21756
rect 51436 19730 51492 19740
rect 51548 20300 51940 20356
rect 51996 21362 52052 21374
rect 51996 21310 51998 21362
rect 52050 21310 52052 21362
rect 51324 19516 51492 19572
rect 51324 19348 51380 19358
rect 50204 19070 50206 19122
rect 50258 19070 50260 19122
rect 50204 19058 50260 19070
rect 51100 19234 51156 19246
rect 51100 19182 51102 19234
rect 51154 19182 51156 19234
rect 50092 17444 50148 18396
rect 50316 19012 50372 19022
rect 50316 18452 50372 18956
rect 50876 19012 50932 19022
rect 51100 19012 51156 19182
rect 51324 19234 51380 19292
rect 51324 19182 51326 19234
rect 51378 19182 51380 19234
rect 51324 19170 51380 19182
rect 51436 19234 51492 19516
rect 51436 19182 51438 19234
rect 51490 19182 51492 19234
rect 50876 19010 51156 19012
rect 50876 18958 50878 19010
rect 50930 18958 51156 19010
rect 50876 18956 51156 18958
rect 51436 19012 51492 19182
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50876 18676 50932 18956
rect 51436 18946 51492 18956
rect 50764 18620 50932 18676
rect 50316 18450 50596 18452
rect 50316 18398 50318 18450
rect 50370 18398 50596 18450
rect 50316 18396 50596 18398
rect 50092 17378 50148 17388
rect 50204 17442 50260 17454
rect 50204 17390 50206 17442
rect 50258 17390 50260 17442
rect 50204 17108 50260 17390
rect 50204 17042 50260 17052
rect 50316 16996 50372 18396
rect 50540 17554 50596 18396
rect 50764 18228 50820 18620
rect 50988 18452 51044 18462
rect 50764 18172 50932 18228
rect 50540 17502 50542 17554
rect 50594 17502 50596 17554
rect 50540 17490 50596 17502
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50876 17220 50932 18172
rect 50988 17890 51044 18396
rect 51212 18450 51268 18462
rect 51212 18398 51214 18450
rect 51266 18398 51268 18450
rect 51212 18004 51268 18398
rect 51212 17938 51268 17948
rect 50988 17838 50990 17890
rect 51042 17838 51044 17890
rect 50988 17826 51044 17838
rect 50988 17556 51044 17566
rect 50988 17462 51044 17500
rect 51100 17556 51156 17566
rect 51100 17554 51268 17556
rect 51100 17502 51102 17554
rect 51154 17502 51268 17554
rect 51100 17500 51268 17502
rect 51100 17490 51156 17500
rect 51100 17332 51156 17342
rect 50876 17164 51044 17220
rect 50316 16930 50372 16940
rect 50876 16996 50932 17006
rect 49980 15474 50036 15484
rect 50204 16884 50260 16894
rect 50204 15148 50260 16828
rect 50876 16882 50932 16940
rect 50876 16830 50878 16882
rect 50930 16830 50932 16882
rect 50876 16818 50932 16830
rect 50652 16658 50708 16670
rect 50652 16606 50654 16658
rect 50706 16606 50708 16658
rect 50652 15876 50708 16606
rect 50988 16660 51044 17164
rect 51100 17106 51156 17276
rect 51100 17054 51102 17106
rect 51154 17054 51156 17106
rect 51100 16884 51156 17054
rect 51212 17106 51268 17500
rect 51212 17054 51214 17106
rect 51266 17054 51268 17106
rect 51212 17042 51268 17054
rect 51324 17220 51380 17230
rect 51324 17106 51380 17164
rect 51324 17054 51326 17106
rect 51378 17054 51380 17106
rect 51324 17042 51380 17054
rect 51100 16818 51156 16828
rect 50988 16604 51156 16660
rect 50652 15820 51044 15876
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 48300 15092 48692 15148
rect 48748 15092 48916 15148
rect 49420 15092 49588 15148
rect 47964 14530 48020 15092
rect 48636 14642 48692 15092
rect 48860 15090 48916 15092
rect 48860 15038 48862 15090
rect 48914 15038 48916 15090
rect 48860 15026 48916 15038
rect 48636 14590 48638 14642
rect 48690 14590 48692 14642
rect 48636 14578 48692 14590
rect 49196 14756 49252 14766
rect 47964 14478 47966 14530
rect 48018 14478 48020 14530
rect 47964 14466 48020 14478
rect 47740 14308 47796 14318
rect 48076 14308 48132 14318
rect 47740 14306 48020 14308
rect 47740 14254 47742 14306
rect 47794 14254 48020 14306
rect 47740 14252 48020 14254
rect 47740 14242 47796 14252
rect 47740 13634 47796 13646
rect 47740 13582 47742 13634
rect 47794 13582 47796 13634
rect 47740 13522 47796 13582
rect 47740 13470 47742 13522
rect 47794 13470 47796 13522
rect 47740 13458 47796 13470
rect 47740 12962 47796 12974
rect 47740 12910 47742 12962
rect 47794 12910 47796 12962
rect 47740 12404 47796 12910
rect 47964 12628 48020 14252
rect 48076 14306 48692 14308
rect 48076 14254 48078 14306
rect 48130 14254 48692 14306
rect 48076 14252 48692 14254
rect 48076 14242 48132 14252
rect 48188 13636 48244 13646
rect 48244 13580 48356 13636
rect 48188 13542 48244 13580
rect 48076 13524 48132 13534
rect 48076 13188 48132 13468
rect 48076 13122 48132 13132
rect 48300 12962 48356 13580
rect 48300 12910 48302 12962
rect 48354 12910 48356 12962
rect 48300 12898 48356 12910
rect 48524 12740 48580 12750
rect 48524 12646 48580 12684
rect 47964 12572 48132 12628
rect 47964 12404 48020 12414
rect 47740 12348 47964 12404
rect 47964 12310 48020 12348
rect 47852 11732 47908 11742
rect 47852 11506 47908 11676
rect 47852 11454 47854 11506
rect 47906 11454 47908 11506
rect 47852 11442 47908 11454
rect 47404 11340 47572 11396
rect 47292 9426 47348 9436
rect 47404 11170 47460 11182
rect 47404 11118 47406 11170
rect 47458 11118 47460 11170
rect 47292 9042 47348 9054
rect 47292 8990 47294 9042
rect 47346 8990 47348 9042
rect 47068 8306 47124 8316
rect 47180 8930 47236 8942
rect 47180 8878 47182 8930
rect 47234 8878 47236 8930
rect 46956 7970 47012 7980
rect 47180 7252 47236 8878
rect 47180 4676 47236 7196
rect 47292 7140 47348 8990
rect 47292 7074 47348 7084
rect 47180 4610 47236 4620
rect 47292 6692 47348 6702
rect 46844 3502 46846 3554
rect 46898 3502 46900 3554
rect 46844 3490 46900 3502
rect 47292 3444 47348 6636
rect 47404 5012 47460 11118
rect 47516 9716 47572 11340
rect 47628 10610 47684 11340
rect 47628 10558 47630 10610
rect 47682 10558 47684 10610
rect 47628 10546 47684 10558
rect 47740 10276 47796 10286
rect 47516 9650 47572 9660
rect 47628 10052 47684 10062
rect 47516 9154 47572 9166
rect 47516 9102 47518 9154
rect 47570 9102 47572 9154
rect 47516 8596 47572 9102
rect 47628 9154 47684 9996
rect 47740 9938 47796 10220
rect 47740 9886 47742 9938
rect 47794 9886 47796 9938
rect 47740 9874 47796 9886
rect 47964 10164 48020 10174
rect 47628 9102 47630 9154
rect 47682 9102 47684 9154
rect 47628 9090 47684 9102
rect 47516 8540 47684 8596
rect 47404 4946 47460 4956
rect 47516 8370 47572 8382
rect 47516 8318 47518 8370
rect 47570 8318 47572 8370
rect 47516 3556 47572 8318
rect 47628 7364 47684 8540
rect 47852 8148 47908 8158
rect 47628 7298 47684 7308
rect 47740 8146 47908 8148
rect 47740 8094 47854 8146
rect 47906 8094 47908 8146
rect 47740 8092 47908 8094
rect 47740 5348 47796 8092
rect 47852 8082 47908 8092
rect 47964 8146 48020 10108
rect 47964 8094 47966 8146
rect 48018 8094 48020 8146
rect 47964 8082 48020 8094
rect 47852 6804 47908 6814
rect 47852 6018 47908 6748
rect 47852 5966 47854 6018
rect 47906 5966 47908 6018
rect 47852 5954 47908 5966
rect 48076 5348 48132 12572
rect 48524 11396 48580 11406
rect 48524 11302 48580 11340
rect 48188 11284 48244 11294
rect 48188 11190 48244 11228
rect 48636 11284 48692 14252
rect 49196 13972 49252 14700
rect 48748 13970 49252 13972
rect 48748 13918 49198 13970
rect 49250 13918 49252 13970
rect 48748 13916 49252 13918
rect 48748 12962 48804 13916
rect 49196 13906 49252 13916
rect 49420 14306 49476 14318
rect 49420 14254 49422 14306
rect 49474 14254 49476 14306
rect 49308 13524 49364 13534
rect 49196 13522 49364 13524
rect 49196 13470 49310 13522
rect 49362 13470 49364 13522
rect 49196 13468 49364 13470
rect 48860 13076 48916 13086
rect 48860 13074 49028 13076
rect 48860 13022 48862 13074
rect 48914 13022 49028 13074
rect 48860 13020 49028 13022
rect 48860 13010 48916 13020
rect 48748 12910 48750 12962
rect 48802 12910 48804 12962
rect 48748 12898 48804 12910
rect 48860 12738 48916 12750
rect 48860 12686 48862 12738
rect 48914 12686 48916 12738
rect 48748 12292 48804 12302
rect 48748 12198 48804 12236
rect 48860 12180 48916 12686
rect 48860 12114 48916 12124
rect 48748 11284 48804 11294
rect 48636 11282 48804 11284
rect 48636 11230 48750 11282
rect 48802 11230 48804 11282
rect 48636 11228 48804 11230
rect 48636 10836 48692 11228
rect 48748 11218 48804 11228
rect 48860 11284 48916 11294
rect 48524 10780 48692 10836
rect 48188 10612 48244 10622
rect 48188 10610 48468 10612
rect 48188 10558 48190 10610
rect 48242 10558 48468 10610
rect 48188 10556 48468 10558
rect 48188 10546 48244 10556
rect 48188 9602 48244 9614
rect 48188 9550 48190 9602
rect 48242 9550 48244 9602
rect 48188 9156 48244 9550
rect 48300 9268 48356 9278
rect 48300 9174 48356 9212
rect 48188 9090 48244 9100
rect 48412 8708 48468 10556
rect 48524 10164 48580 10780
rect 48860 10724 48916 11228
rect 48524 9826 48580 10108
rect 48524 9774 48526 9826
rect 48578 9774 48580 9826
rect 48524 9762 48580 9774
rect 48636 10668 48916 10724
rect 48636 10276 48692 10668
rect 48972 10610 49028 13020
rect 49084 12180 49140 12190
rect 49084 12086 49140 12124
rect 49084 11732 49140 11742
rect 49084 11170 49140 11676
rect 49084 11118 49086 11170
rect 49138 11118 49140 11170
rect 49084 11106 49140 11118
rect 49196 10836 49252 13468
rect 49308 13458 49364 13468
rect 49420 13188 49476 14254
rect 49420 13122 49476 13132
rect 49532 12964 49588 15092
rect 50092 15092 50260 15148
rect 50764 15540 50820 15550
rect 49756 14306 49812 14318
rect 49756 14254 49758 14306
rect 49810 14254 49812 14306
rect 49420 12908 49588 12964
rect 49644 13634 49700 13646
rect 49644 13582 49646 13634
rect 49698 13582 49700 13634
rect 49644 12964 49700 13582
rect 49756 13522 49812 14254
rect 49756 13470 49758 13522
rect 49810 13470 49812 13522
rect 49756 13458 49812 13470
rect 49308 12852 49364 12862
rect 49308 12758 49364 12796
rect 49308 12292 49364 12302
rect 49420 12292 49476 12908
rect 49644 12898 49700 12908
rect 49756 13076 49812 13086
rect 49756 12962 49812 13020
rect 49756 12910 49758 12962
rect 49810 12910 49812 12962
rect 49756 12898 49812 12910
rect 49980 12962 50036 12974
rect 49980 12910 49982 12962
rect 50034 12910 50036 12962
rect 49532 12740 49588 12750
rect 49532 12646 49588 12684
rect 49644 12738 49700 12750
rect 49644 12686 49646 12738
rect 49698 12686 49700 12738
rect 49644 12402 49700 12686
rect 49644 12350 49646 12402
rect 49698 12350 49700 12402
rect 49644 12338 49700 12350
rect 49756 12292 49812 12302
rect 49420 12236 49588 12292
rect 49308 12178 49364 12236
rect 49308 12126 49310 12178
rect 49362 12126 49364 12178
rect 49308 12114 49364 12126
rect 49308 11956 49364 11966
rect 49364 11900 49476 11956
rect 49308 11890 49364 11900
rect 49196 10770 49252 10780
rect 48972 10558 48974 10610
rect 49026 10558 49028 10610
rect 48972 10546 49028 10558
rect 49196 10612 49252 10622
rect 49196 10518 49252 10556
rect 48636 9826 48692 10220
rect 48636 9774 48638 9826
rect 48690 9774 48692 9826
rect 48636 9762 48692 9774
rect 48860 10498 48916 10510
rect 48860 10446 48862 10498
rect 48914 10446 48916 10498
rect 48748 9714 48804 9726
rect 48748 9662 48750 9714
rect 48802 9662 48804 9714
rect 48748 8708 48804 9662
rect 48412 8652 48804 8708
rect 48412 8484 48468 8652
rect 48860 8596 48916 10446
rect 48972 9940 49028 9950
rect 48972 9266 49028 9884
rect 49196 9828 49252 9838
rect 49196 9734 49252 9772
rect 49420 9380 49476 11900
rect 49532 11284 49588 12236
rect 49756 12198 49812 12236
rect 49868 12180 49924 12190
rect 49980 12180 50036 12910
rect 49924 12124 50036 12180
rect 49868 12114 49924 12124
rect 49756 11954 49812 11966
rect 49756 11902 49758 11954
rect 49810 11902 49812 11954
rect 49756 11732 49812 11902
rect 50092 11956 50148 15092
rect 50316 14420 50372 14430
rect 50204 13972 50260 13982
rect 50204 13878 50260 13916
rect 50316 13076 50372 14364
rect 50764 14308 50820 15484
rect 50876 15428 50932 15438
rect 50876 15202 50932 15372
rect 50876 15150 50878 15202
rect 50930 15150 50932 15202
rect 50876 15138 50932 15150
rect 50764 14252 50932 14308
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50764 13972 50820 13982
rect 50876 13972 50932 14252
rect 50764 13970 50932 13972
rect 50764 13918 50766 13970
rect 50818 13918 50932 13970
rect 50764 13916 50932 13918
rect 50764 13906 50820 13916
rect 50876 13634 50932 13646
rect 50876 13582 50878 13634
rect 50930 13582 50932 13634
rect 50428 13076 50484 13086
rect 50372 13074 50484 13076
rect 50372 13022 50430 13074
rect 50482 13022 50484 13074
rect 50372 13020 50484 13022
rect 50316 12982 50372 13020
rect 50428 13010 50484 13020
rect 50876 12852 50932 13582
rect 50988 13412 51044 15820
rect 51100 13524 51156 16604
rect 51548 15148 51604 20300
rect 51996 20244 52052 21310
rect 52108 20916 52164 20926
rect 52108 20822 52164 20860
rect 51884 20188 52052 20244
rect 52108 20692 52164 20702
rect 51884 20020 51940 20188
rect 51772 19796 51828 19806
rect 51772 19124 51828 19740
rect 51884 19236 51940 19964
rect 51996 20018 52052 20030
rect 51996 19966 51998 20018
rect 52050 19966 52052 20018
rect 51996 19908 52052 19966
rect 51996 19842 52052 19852
rect 52108 19458 52164 20636
rect 52220 20244 52276 21980
rect 52332 21586 52388 21598
rect 52332 21534 52334 21586
rect 52386 21534 52388 21586
rect 52332 21252 52388 21534
rect 52332 21186 52388 21196
rect 52220 20188 52388 20244
rect 52108 19406 52110 19458
rect 52162 19406 52164 19458
rect 52108 19394 52164 19406
rect 52220 20020 52276 20030
rect 52220 19348 52276 19964
rect 52332 19348 52388 20188
rect 52444 19572 52500 22876
rect 52556 21588 52612 23100
rect 52780 23154 52836 23436
rect 52780 23102 52782 23154
rect 52834 23102 52836 23154
rect 52780 23090 52836 23102
rect 52892 23156 52948 23166
rect 52892 23062 52948 23100
rect 53116 23154 53172 23166
rect 53116 23102 53118 23154
rect 53170 23102 53172 23154
rect 53004 23042 53060 23054
rect 53004 22990 53006 23042
rect 53058 22990 53060 23042
rect 52668 22372 52724 22382
rect 52668 22278 52724 22316
rect 52892 21812 52948 21822
rect 53004 21812 53060 22990
rect 53116 23044 53172 23102
rect 53116 22978 53172 22988
rect 53228 22148 53284 25564
rect 53340 25508 53396 25518
rect 53340 25414 53396 25452
rect 53564 24500 53620 24510
rect 53564 24162 53620 24444
rect 53564 24110 53566 24162
rect 53618 24110 53620 24162
rect 53564 24098 53620 24110
rect 53676 23716 53732 26796
rect 53788 26178 53844 29036
rect 53900 28756 53956 28766
rect 53900 28642 53956 28700
rect 53900 28590 53902 28642
rect 53954 28590 53956 28642
rect 53900 26628 53956 28590
rect 54348 28644 54404 28654
rect 54460 28644 54516 29150
rect 54404 28588 54516 28644
rect 54236 28418 54292 28430
rect 54236 28366 54238 28418
rect 54290 28366 54292 28418
rect 53900 26562 53956 26572
rect 54012 27970 54068 27982
rect 54012 27918 54014 27970
rect 54066 27918 54068 27970
rect 53788 26126 53790 26178
rect 53842 26126 53844 26178
rect 53788 25506 53844 26126
rect 53788 25454 53790 25506
rect 53842 25454 53844 25506
rect 53788 25442 53844 25454
rect 53900 26404 53956 26414
rect 53900 25394 53956 26348
rect 54012 26290 54068 27918
rect 54236 26908 54292 28366
rect 54348 27860 54404 28588
rect 54348 27766 54404 27804
rect 54684 27076 54740 27086
rect 54796 27076 54852 30156
rect 55244 30210 55300 30222
rect 55244 30158 55246 30210
rect 55298 30158 55300 30210
rect 55020 29540 55076 29550
rect 55020 29446 55076 29484
rect 55244 29316 55300 30158
rect 55804 30210 55860 30222
rect 55804 30158 55806 30210
rect 55858 30158 55860 30210
rect 55244 29250 55300 29260
rect 55468 29988 55524 29998
rect 54908 28980 54964 28990
rect 55132 28980 55188 28990
rect 54964 28924 55076 28980
rect 54908 28914 54964 28924
rect 55020 28308 55076 28924
rect 55132 28530 55188 28924
rect 55132 28478 55134 28530
rect 55186 28478 55188 28530
rect 55132 28466 55188 28478
rect 55356 28532 55412 28542
rect 55020 28252 55300 28308
rect 55244 27970 55300 28252
rect 55244 27918 55246 27970
rect 55298 27918 55300 27970
rect 55244 27906 55300 27918
rect 55132 27860 55188 27870
rect 54684 27074 54852 27076
rect 54684 27022 54686 27074
rect 54738 27022 54852 27074
rect 54684 27020 54852 27022
rect 55020 27076 55076 27086
rect 54684 27010 54740 27020
rect 55020 26982 55076 27020
rect 54124 26852 54292 26908
rect 55132 26962 55188 27804
rect 55132 26910 55134 26962
rect 55186 26910 55188 26962
rect 55132 26898 55188 26910
rect 55356 26908 55412 28476
rect 54124 26786 54180 26796
rect 54348 26850 54404 26862
rect 54348 26798 54350 26850
rect 54402 26798 54404 26850
rect 54348 26404 54404 26798
rect 55244 26852 55412 26908
rect 54572 26628 54628 26638
rect 54460 26404 54516 26414
rect 54348 26348 54460 26404
rect 54012 26238 54014 26290
rect 54066 26238 54068 26290
rect 54012 25620 54068 26238
rect 54460 26290 54516 26348
rect 54460 26238 54462 26290
rect 54514 26238 54516 26290
rect 54460 26226 54516 26238
rect 54012 25554 54068 25564
rect 54124 26066 54180 26078
rect 54572 26068 54628 26572
rect 54124 26014 54126 26066
rect 54178 26014 54180 26066
rect 53900 25342 53902 25394
rect 53954 25342 53956 25394
rect 53900 25330 53956 25342
rect 53900 24276 53956 24286
rect 53900 24052 53956 24220
rect 53900 23986 53956 23996
rect 54124 24276 54180 26014
rect 54460 26012 54628 26068
rect 54460 25396 54516 26012
rect 54460 25302 54516 25340
rect 54236 25284 54292 25294
rect 54236 25190 54292 25228
rect 55244 25060 55300 26852
rect 55132 25004 55300 25060
rect 55020 24724 55076 24734
rect 53564 23714 53732 23716
rect 53564 23662 53678 23714
rect 53730 23662 53732 23714
rect 53564 23660 53732 23662
rect 53340 23156 53396 23166
rect 53340 23062 53396 23100
rect 53564 22932 53620 23660
rect 53676 23650 53732 23660
rect 53900 23714 53956 23726
rect 53900 23662 53902 23714
rect 53954 23662 53956 23714
rect 53676 23492 53732 23502
rect 53676 23266 53732 23436
rect 53676 23214 53678 23266
rect 53730 23214 53732 23266
rect 53676 23202 53732 23214
rect 53788 23266 53844 23278
rect 53788 23214 53790 23266
rect 53842 23214 53844 23266
rect 53564 22866 53620 22876
rect 53788 22708 53844 23214
rect 53900 23268 53956 23662
rect 53900 23202 53956 23212
rect 53788 22642 53844 22652
rect 54012 23156 54068 23166
rect 53228 22092 53396 22148
rect 53116 21812 53172 21822
rect 53004 21810 53172 21812
rect 53004 21758 53118 21810
rect 53170 21758 53172 21810
rect 53004 21756 53172 21758
rect 52892 21718 52948 21756
rect 53116 21746 53172 21756
rect 52668 21700 52724 21710
rect 52724 21644 52836 21700
rect 52668 21634 52724 21644
rect 52780 21642 52836 21644
rect 52780 21590 52782 21642
rect 52834 21590 52836 21642
rect 52780 21578 52836 21590
rect 52556 21522 52612 21532
rect 52780 21476 52836 21486
rect 52668 21474 52836 21476
rect 52668 21422 52782 21474
rect 52834 21422 52836 21474
rect 52668 21420 52836 21422
rect 52556 20916 52612 20926
rect 52556 20802 52612 20860
rect 52556 20750 52558 20802
rect 52610 20750 52612 20802
rect 52556 20738 52612 20750
rect 52556 20244 52612 20254
rect 52668 20244 52724 21420
rect 52780 21410 52836 21420
rect 53340 20804 53396 22092
rect 53676 21812 53732 21822
rect 53732 21756 53844 21812
rect 53676 21746 53732 21756
rect 53676 21362 53732 21374
rect 53676 21310 53678 21362
rect 53730 21310 53732 21362
rect 53676 21140 53732 21310
rect 53340 20738 53396 20748
rect 53452 21084 53676 21140
rect 53004 20692 53060 20702
rect 53004 20690 53172 20692
rect 53004 20638 53006 20690
rect 53058 20638 53172 20690
rect 53004 20636 53172 20638
rect 53004 20626 53060 20636
rect 52892 20580 52948 20590
rect 52892 20486 52948 20524
rect 52556 20242 52724 20244
rect 52556 20190 52558 20242
rect 52610 20190 52724 20242
rect 52556 20188 52724 20190
rect 52780 20468 52836 20478
rect 52780 20242 52836 20412
rect 52780 20190 52782 20242
rect 52834 20190 52836 20242
rect 52556 20178 52612 20188
rect 52780 20178 52836 20190
rect 52892 20130 52948 20142
rect 52892 20078 52894 20130
rect 52946 20078 52948 20130
rect 52892 19684 52948 20078
rect 53004 20132 53060 20142
rect 53004 20038 53060 20076
rect 53116 19908 53172 20636
rect 53228 20690 53284 20702
rect 53228 20638 53230 20690
rect 53282 20638 53284 20690
rect 53228 20468 53284 20638
rect 53228 20412 53396 20468
rect 53340 20244 53396 20412
rect 53340 20178 53396 20188
rect 52892 19618 52948 19628
rect 53004 19852 53172 19908
rect 53340 19906 53396 19918
rect 53340 19854 53342 19906
rect 53394 19854 53396 19906
rect 52444 19506 52500 19516
rect 52892 19348 52948 19358
rect 52332 19346 52948 19348
rect 52332 19294 52894 19346
rect 52946 19294 52948 19346
rect 52332 19292 52948 19294
rect 52220 19282 52276 19292
rect 52892 19282 52948 19292
rect 51996 19236 52052 19246
rect 51884 19180 51996 19236
rect 51996 19142 52052 19180
rect 52668 19124 52724 19134
rect 51772 19068 51940 19124
rect 51660 19010 51716 19022
rect 51660 18958 51662 19010
rect 51714 18958 51716 19010
rect 51660 18228 51716 18958
rect 51884 18450 51940 19068
rect 52668 19122 52836 19124
rect 52668 19070 52670 19122
rect 52722 19070 52836 19122
rect 52668 19068 52836 19070
rect 52668 19058 52724 19068
rect 52556 19012 52612 19022
rect 52444 19010 52612 19012
rect 52444 18958 52558 19010
rect 52610 18958 52612 19010
rect 52444 18956 52612 18958
rect 52444 18562 52500 18956
rect 52556 18946 52612 18956
rect 52444 18510 52446 18562
rect 52498 18510 52500 18562
rect 52444 18498 52500 18510
rect 51884 18398 51886 18450
rect 51938 18398 51940 18450
rect 51884 18386 51940 18398
rect 52108 18450 52164 18462
rect 52108 18398 52110 18450
rect 52162 18398 52164 18450
rect 51772 18340 51828 18350
rect 51772 18246 51828 18284
rect 51660 17556 51716 18172
rect 52108 17892 52164 18398
rect 52668 18452 52724 18462
rect 52668 18358 52724 18396
rect 52780 18116 52836 19068
rect 53004 18340 53060 19852
rect 53116 19684 53172 19694
rect 53116 19458 53172 19628
rect 53116 19406 53118 19458
rect 53170 19406 53172 19458
rect 53116 19394 53172 19406
rect 53340 19460 53396 19854
rect 53340 19394 53396 19404
rect 53340 19236 53396 19246
rect 53452 19236 53508 21084
rect 53676 21074 53732 21084
rect 53676 20916 53732 20926
rect 53788 20916 53844 21756
rect 54012 21586 54068 23100
rect 54012 21534 54014 21586
rect 54066 21534 54068 21586
rect 54012 21522 54068 21534
rect 54124 21588 54180 24220
rect 54236 24722 55076 24724
rect 54236 24670 55022 24722
rect 55074 24670 55076 24722
rect 54236 24668 55076 24670
rect 54236 23938 54292 24668
rect 55020 24658 55076 24668
rect 55132 24276 55188 25004
rect 54236 23886 54238 23938
rect 54290 23886 54292 23938
rect 54236 23874 54292 23886
rect 54460 24220 55188 24276
rect 55244 24834 55300 24846
rect 55244 24782 55246 24834
rect 55298 24782 55300 24834
rect 54348 23042 54404 23054
rect 54348 22990 54350 23042
rect 54402 22990 54404 23042
rect 54348 22932 54404 22990
rect 54348 22866 54404 22876
rect 54236 21588 54292 21598
rect 54124 21586 54292 21588
rect 54124 21534 54238 21586
rect 54290 21534 54292 21586
rect 54124 21532 54292 21534
rect 54236 21522 54292 21532
rect 53676 20914 53844 20916
rect 53676 20862 53678 20914
rect 53730 20862 53844 20914
rect 53676 20860 53844 20862
rect 53564 20244 53620 20254
rect 53564 19684 53620 20188
rect 53564 19618 53620 19628
rect 53340 19234 53508 19236
rect 53340 19182 53342 19234
rect 53394 19182 53508 19234
rect 53340 19180 53508 19182
rect 53340 19170 53396 19180
rect 53564 19124 53620 19134
rect 53564 19030 53620 19068
rect 53116 19012 53172 19022
rect 53116 18450 53172 18956
rect 53452 18674 53508 18686
rect 53452 18622 53454 18674
rect 53506 18622 53508 18674
rect 53116 18398 53118 18450
rect 53170 18398 53172 18450
rect 53116 18386 53172 18398
rect 53340 18450 53396 18462
rect 53340 18398 53342 18450
rect 53394 18398 53396 18450
rect 53004 18274 53060 18284
rect 52892 18228 52948 18238
rect 52892 18134 52948 18172
rect 52780 18050 52836 18060
rect 53340 18116 53396 18398
rect 53340 18050 53396 18060
rect 51660 17490 51716 17500
rect 51884 17836 52612 17892
rect 51884 17220 51940 17836
rect 52444 17556 52500 17566
rect 51884 17106 51940 17164
rect 51884 17054 51886 17106
rect 51938 17054 51940 17106
rect 51884 17042 51940 17054
rect 52332 17332 52388 17342
rect 52332 17106 52388 17276
rect 52332 17054 52334 17106
rect 52386 17054 52388 17106
rect 52332 17042 52388 17054
rect 51772 15874 51828 15886
rect 51772 15822 51774 15874
rect 51826 15822 51828 15874
rect 51772 15428 51828 15822
rect 51772 15362 51828 15372
rect 52220 15874 52276 15886
rect 52220 15822 52222 15874
rect 52274 15822 52276 15874
rect 51100 13458 51156 13468
rect 51436 15092 51604 15148
rect 51660 15092 51716 15102
rect 52220 15092 52276 15822
rect 50988 13346 51044 13356
rect 50876 12786 50932 12796
rect 51100 12738 51156 12750
rect 51100 12686 51102 12738
rect 51154 12686 51156 12738
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 51100 12404 51156 12686
rect 51100 12348 51380 12404
rect 50204 12290 50260 12302
rect 50204 12238 50206 12290
rect 50258 12238 50260 12290
rect 50204 12180 50260 12238
rect 50540 12292 50596 12302
rect 50764 12292 50820 12302
rect 50540 12290 50764 12292
rect 50540 12238 50542 12290
rect 50594 12238 50764 12290
rect 50540 12236 50764 12238
rect 50540 12226 50596 12236
rect 50204 12114 50260 12124
rect 50092 11900 50260 11956
rect 50092 11732 50148 11742
rect 49756 11676 50036 11732
rect 49532 11218 49588 11228
rect 49644 11508 49700 11518
rect 49308 9268 49364 9278
rect 49420 9268 49476 9324
rect 48972 9214 48974 9266
rect 49026 9214 49028 9266
rect 48972 9202 49028 9214
rect 49196 9266 49476 9268
rect 49196 9214 49310 9266
rect 49362 9214 49476 9266
rect 49196 9212 49476 9214
rect 49532 11060 49588 11070
rect 48412 8418 48468 8428
rect 48524 8540 48916 8596
rect 48188 8034 48244 8046
rect 48188 7982 48190 8034
rect 48242 7982 48244 8034
rect 48188 7588 48244 7982
rect 48300 8036 48356 8046
rect 48356 7980 48468 8036
rect 48300 7970 48356 7980
rect 48188 7522 48244 7532
rect 48188 7364 48244 7374
rect 48188 7270 48244 7308
rect 48300 6132 48356 6142
rect 48076 5292 48244 5348
rect 47740 5282 47796 5292
rect 48076 5012 48132 5022
rect 48076 4918 48132 4956
rect 47964 4788 48020 4798
rect 47964 4450 48020 4732
rect 48076 4564 48132 4574
rect 48188 4564 48244 5292
rect 48076 4562 48244 4564
rect 48076 4510 48078 4562
rect 48130 4510 48244 4562
rect 48076 4508 48244 4510
rect 48076 4498 48132 4508
rect 47964 4398 47966 4450
rect 48018 4398 48020 4450
rect 47964 4386 48020 4398
rect 47628 4340 47684 4350
rect 47628 4226 47684 4284
rect 47628 4174 47630 4226
rect 47682 4174 47684 4226
rect 47628 4162 47684 4174
rect 48188 3892 48244 4508
rect 48300 4562 48356 6076
rect 48300 4510 48302 4562
rect 48354 4510 48356 4562
rect 48300 4498 48356 4510
rect 47964 3836 48244 3892
rect 47628 3556 47684 3566
rect 47516 3554 47684 3556
rect 47516 3502 47630 3554
rect 47682 3502 47684 3554
rect 47516 3500 47684 3502
rect 47628 3490 47684 3500
rect 47404 3444 47460 3454
rect 47292 3442 47460 3444
rect 47292 3390 47406 3442
rect 47458 3390 47460 3442
rect 47292 3388 47460 3390
rect 46620 3332 46900 3388
rect 47404 3378 47460 3388
rect 47964 3388 48020 3836
rect 48412 3388 48468 7980
rect 48524 3554 48580 8540
rect 48860 8372 48916 8382
rect 48916 8316 49140 8372
rect 48860 8278 48916 8316
rect 48748 7362 48804 7374
rect 48748 7310 48750 7362
rect 48802 7310 48804 7362
rect 48636 6804 48692 6814
rect 48636 6710 48692 6748
rect 48748 6356 48804 7310
rect 48860 7250 48916 7262
rect 48860 7198 48862 7250
rect 48914 7198 48916 7250
rect 48860 6916 48916 7198
rect 48860 6850 48916 6860
rect 49084 6692 49140 8316
rect 49196 7586 49252 9212
rect 49308 9202 49364 9212
rect 49532 8372 49588 11004
rect 49644 8484 49700 11452
rect 49980 10610 50036 11676
rect 50092 11394 50148 11676
rect 50092 11342 50094 11394
rect 50146 11342 50148 11394
rect 50092 11330 50148 11342
rect 50204 10836 50260 11900
rect 50764 11506 50820 12236
rect 51100 12180 51156 12190
rect 51100 12086 51156 12124
rect 50764 11454 50766 11506
rect 50818 11454 50820 11506
rect 50764 11442 50820 11454
rect 49980 10558 49982 10610
rect 50034 10558 50036 10610
rect 49980 10546 50036 10558
rect 50092 10780 50260 10836
rect 50316 11170 50372 11182
rect 50316 11118 50318 11170
rect 50370 11118 50372 11170
rect 50316 11060 50372 11118
rect 51212 11170 51268 11182
rect 51212 11118 51214 11170
rect 51266 11118 51268 11170
rect 49756 9828 49812 9838
rect 49756 9734 49812 9772
rect 49756 9604 49812 9614
rect 49756 9266 49812 9548
rect 49756 9214 49758 9266
rect 49810 9214 49812 9266
rect 49756 8932 49812 9214
rect 49756 8866 49812 8876
rect 50092 9268 50148 10780
rect 50204 10612 50260 10622
rect 50204 10518 50260 10556
rect 50204 10388 50260 10398
rect 50204 9938 50260 10332
rect 50316 10164 50372 11004
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50652 10388 50708 10398
rect 50316 10098 50372 10108
rect 50428 10386 50708 10388
rect 50428 10334 50654 10386
rect 50706 10334 50708 10386
rect 50428 10332 50708 10334
rect 50204 9886 50206 9938
rect 50258 9886 50260 9938
rect 50204 9874 50260 9886
rect 49644 8428 49812 8484
rect 49756 8372 49812 8428
rect 49532 8316 49700 8372
rect 49420 8260 49476 8270
rect 49420 8166 49476 8204
rect 49532 8148 49588 8158
rect 49532 7698 49588 8092
rect 49532 7646 49534 7698
rect 49586 7646 49588 7698
rect 49532 7634 49588 7646
rect 49196 7534 49198 7586
rect 49250 7534 49252 7586
rect 49196 7522 49252 7534
rect 49308 7586 49364 7598
rect 49308 7534 49310 7586
rect 49362 7534 49364 7586
rect 49308 7476 49364 7534
rect 49308 7410 49364 7420
rect 49196 6692 49252 6702
rect 49084 6636 49196 6692
rect 49196 6598 49252 6636
rect 48748 6290 48804 6300
rect 48860 6580 48916 6590
rect 48860 5908 48916 6524
rect 49644 6580 49700 8316
rect 49756 8306 49812 8316
rect 49756 8146 49812 8158
rect 49756 8094 49758 8146
rect 49810 8094 49812 8146
rect 49756 8036 49812 8094
rect 49756 7970 49812 7980
rect 49644 6514 49700 6524
rect 49756 7476 49812 7486
rect 50092 7476 50148 9212
rect 50316 9604 50372 9614
rect 50316 9266 50372 9548
rect 50316 9214 50318 9266
rect 50370 9214 50372 9266
rect 50316 9202 50372 9214
rect 50204 7476 50260 7486
rect 50092 7474 50260 7476
rect 50092 7422 50206 7474
rect 50258 7422 50260 7474
rect 50092 7420 50260 7422
rect 48748 5236 48804 5246
rect 48748 5142 48804 5180
rect 48748 4340 48804 4350
rect 48748 4246 48804 4284
rect 48524 3502 48526 3554
rect 48578 3502 48580 3554
rect 48524 3490 48580 3502
rect 47964 3332 48132 3388
rect 46844 800 46900 3332
rect 48076 2996 48132 3332
rect 48076 2930 48132 2940
rect 48188 3332 48468 3388
rect 48188 800 48244 3332
rect 48860 1540 48916 5852
rect 49196 5794 49252 5806
rect 49196 5742 49198 5794
rect 49250 5742 49252 5794
rect 49196 5684 49252 5742
rect 49644 5796 49700 5806
rect 49252 5628 49476 5684
rect 49196 5618 49252 5628
rect 49308 4452 49364 4462
rect 49308 4358 49364 4396
rect 49420 2772 49476 5628
rect 49644 4450 49700 5740
rect 49756 5794 49812 7420
rect 50204 7410 50260 7420
rect 49868 7364 49924 7374
rect 49868 7270 49924 7308
rect 50092 6916 50148 6926
rect 50148 6860 50372 6916
rect 50092 6850 50148 6860
rect 49980 6580 50036 6590
rect 49980 6486 50036 6524
rect 49756 5742 49758 5794
rect 49810 5742 49812 5794
rect 49756 5730 49812 5742
rect 50316 5010 50372 6860
rect 50428 6468 50484 10332
rect 50652 10322 50708 10332
rect 50540 9828 50596 9838
rect 50540 9734 50596 9772
rect 50876 9604 50932 9614
rect 50876 9602 51044 9604
rect 50876 9550 50878 9602
rect 50930 9550 51044 9602
rect 50876 9548 51044 9550
rect 50876 9538 50932 9548
rect 50988 9492 51044 9548
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50988 9426 51044 9436
rect 50556 9370 50820 9380
rect 51212 9268 51268 11118
rect 50540 9212 51268 9268
rect 50540 8260 50596 9212
rect 51324 9154 51380 12348
rect 51324 9102 51326 9154
rect 51378 9102 51380 9154
rect 51324 9090 51380 9102
rect 51212 9044 51268 9054
rect 51100 8988 51212 9044
rect 50652 8930 50708 8942
rect 50652 8878 50654 8930
rect 50706 8878 50708 8930
rect 50652 8820 50708 8878
rect 50988 8820 51044 8830
rect 50652 8818 51044 8820
rect 50652 8766 50990 8818
rect 51042 8766 51044 8818
rect 50652 8764 51044 8766
rect 50540 8194 50596 8204
rect 50876 8370 50932 8382
rect 50876 8318 50878 8370
rect 50930 8318 50932 8370
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50652 7700 50708 7710
rect 50652 7606 50708 7644
rect 50540 6468 50596 6478
rect 50428 6412 50540 6468
rect 50540 6402 50596 6412
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50876 5236 50932 8318
rect 50988 6804 51044 8764
rect 51100 8820 51156 8988
rect 51212 8950 51268 8988
rect 51100 8754 51156 8764
rect 51324 8708 51380 8718
rect 50988 6738 51044 6748
rect 51212 8652 51324 8708
rect 50876 5180 51156 5236
rect 50316 4958 50318 5010
rect 50370 4958 50372 5010
rect 50316 4946 50372 4958
rect 50428 5122 50484 5134
rect 50428 5070 50430 5122
rect 50482 5070 50484 5122
rect 50428 4562 50484 5070
rect 50876 5012 50932 5022
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50428 4510 50430 4562
rect 50482 4510 50484 4562
rect 50428 4498 50484 4510
rect 49644 4398 49646 4450
rect 49698 4398 49700 4450
rect 49644 4386 49700 4398
rect 49644 3442 49700 3454
rect 49644 3390 49646 3442
rect 49698 3390 49700 3442
rect 49644 3388 49700 3390
rect 49420 2706 49476 2716
rect 49532 3332 49700 3388
rect 48860 1474 48916 1484
rect 49532 800 49588 3332
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 50876 800 50932 4956
rect 51100 3556 51156 5180
rect 51212 4452 51268 8652
rect 51324 8642 51380 8652
rect 51436 7698 51492 15092
rect 51716 15036 51828 15092
rect 51660 15026 51716 15036
rect 51660 12740 51716 12750
rect 51548 12738 51716 12740
rect 51548 12686 51662 12738
rect 51714 12686 51716 12738
rect 51548 12684 51716 12686
rect 51548 10948 51604 12684
rect 51660 12674 51716 12684
rect 51772 12516 51828 15036
rect 52220 15026 52276 15036
rect 52108 13860 52164 13870
rect 51660 12460 51828 12516
rect 51884 13634 51940 13646
rect 51884 13582 51886 13634
rect 51938 13582 51940 13634
rect 51660 11506 51716 12460
rect 51660 11454 51662 11506
rect 51714 11454 51716 11506
rect 51660 11396 51716 11454
rect 51772 12066 51828 12078
rect 51772 12014 51774 12066
rect 51826 12014 51828 12066
rect 51772 11508 51828 12014
rect 51772 11442 51828 11452
rect 51660 11330 51716 11340
rect 51548 10882 51604 10892
rect 51884 10724 51940 13582
rect 52108 11620 52164 13804
rect 52220 12738 52276 12750
rect 52220 12686 52222 12738
rect 52274 12686 52276 12738
rect 52220 12404 52276 12686
rect 52220 12338 52276 12348
rect 52108 11506 52164 11564
rect 52108 11454 52110 11506
rect 52162 11454 52164 11506
rect 52108 11442 52164 11454
rect 51772 10668 51940 10724
rect 51996 10836 52052 10846
rect 51548 10498 51604 10510
rect 51548 10446 51550 10498
rect 51602 10446 51604 10498
rect 51548 9156 51604 10446
rect 51660 9716 51716 9726
rect 51660 9622 51716 9660
rect 51548 9100 51716 9156
rect 51548 8930 51604 8942
rect 51548 8878 51550 8930
rect 51602 8878 51604 8930
rect 51548 8708 51604 8878
rect 51548 8642 51604 8652
rect 51436 7646 51438 7698
rect 51490 7646 51492 7698
rect 51436 7634 51492 7646
rect 51548 8372 51604 8382
rect 51548 8034 51604 8316
rect 51548 7982 51550 8034
rect 51602 7982 51604 8034
rect 51548 6916 51604 7982
rect 51548 5796 51604 6860
rect 51660 6356 51716 9100
rect 51660 6290 51716 6300
rect 51548 5730 51604 5740
rect 51772 5124 51828 10668
rect 51884 10500 51940 10510
rect 51884 10406 51940 10444
rect 51884 9828 51940 9838
rect 51884 8708 51940 9772
rect 51996 9492 52052 10780
rect 52332 10498 52388 10510
rect 52332 10446 52334 10498
rect 52386 10446 52388 10498
rect 51996 9266 52052 9436
rect 51996 9214 51998 9266
rect 52050 9214 52052 9266
rect 51996 9202 52052 9214
rect 52220 9602 52276 9614
rect 52220 9550 52222 9602
rect 52274 9550 52276 9602
rect 52220 8818 52276 9550
rect 52220 8766 52222 8818
rect 52274 8766 52276 8818
rect 52220 8754 52276 8766
rect 52332 9604 52388 10446
rect 51884 8642 51940 8652
rect 52332 8484 52388 9548
rect 52332 8418 52388 8428
rect 52444 9940 52500 17500
rect 52556 17444 52612 17836
rect 52892 17668 52948 17678
rect 52780 17444 52836 17454
rect 52556 17442 52836 17444
rect 52556 17390 52782 17442
rect 52834 17390 52836 17442
rect 52556 17388 52836 17390
rect 52556 17108 52612 17118
rect 52556 15148 52612 17052
rect 52780 16100 52836 17388
rect 52892 16882 52948 17612
rect 53452 16996 53508 18622
rect 53564 16996 53620 17006
rect 53452 16994 53620 16996
rect 53452 16942 53566 16994
rect 53618 16942 53620 16994
rect 53452 16940 53620 16942
rect 53564 16930 53620 16940
rect 52892 16830 52894 16882
rect 52946 16830 52948 16882
rect 52892 16818 52948 16830
rect 52780 16034 52836 16044
rect 52892 16548 52948 16558
rect 52892 16098 52948 16492
rect 53676 16548 53732 20860
rect 54348 20804 54404 20814
rect 54348 20710 54404 20748
rect 54124 20578 54180 20590
rect 54124 20526 54126 20578
rect 54178 20526 54180 20578
rect 54124 20244 54180 20526
rect 54124 20178 54180 20188
rect 53900 19908 53956 19918
rect 53900 16996 53956 19852
rect 54012 19124 54068 19134
rect 54012 19030 54068 19068
rect 53900 16930 53956 16940
rect 54012 17780 54068 17790
rect 53004 16212 53060 16222
rect 53564 16212 53620 16222
rect 53676 16212 53732 16492
rect 53004 16210 53284 16212
rect 53004 16158 53006 16210
rect 53058 16158 53284 16210
rect 53004 16156 53284 16158
rect 53004 16146 53060 16156
rect 52892 16046 52894 16098
rect 52946 16046 52948 16098
rect 52892 16034 52948 16046
rect 53116 15986 53172 15998
rect 53116 15934 53118 15986
rect 53170 15934 53172 15986
rect 52668 15876 52724 15886
rect 52668 15428 52724 15820
rect 52668 15362 52724 15372
rect 52892 15204 52948 15214
rect 52556 15092 52724 15148
rect 52668 14530 52724 15092
rect 52668 14478 52670 14530
rect 52722 14478 52724 14530
rect 52668 14466 52724 14478
rect 52780 14644 52836 14654
rect 52668 13748 52724 13758
rect 52668 13654 52724 13692
rect 52780 12628 52836 14588
rect 52892 14530 52948 15148
rect 52892 14478 52894 14530
rect 52946 14478 52948 14530
rect 52892 14466 52948 14478
rect 53004 15202 53060 15214
rect 53004 15150 53006 15202
rect 53058 15150 53060 15202
rect 53004 14306 53060 15150
rect 53004 14254 53006 14306
rect 53058 14254 53060 14306
rect 53004 14242 53060 14254
rect 53116 15092 53172 15934
rect 53116 13860 53172 15036
rect 53228 14530 53284 16156
rect 53564 16210 53732 16212
rect 53564 16158 53566 16210
rect 53618 16158 53732 16210
rect 53564 16156 53732 16158
rect 53564 16146 53620 16156
rect 53228 14478 53230 14530
rect 53282 14478 53284 14530
rect 53228 14466 53284 14478
rect 53788 15314 53844 15326
rect 53788 15262 53790 15314
rect 53842 15262 53844 15314
rect 53788 14308 53844 15262
rect 54012 14868 54068 17724
rect 54124 15876 54180 15886
rect 54180 15820 54404 15876
rect 54124 15782 54180 15820
rect 54124 15540 54180 15550
rect 54124 15446 54180 15484
rect 54348 15538 54404 15820
rect 54348 15486 54350 15538
rect 54402 15486 54404 15538
rect 54348 15474 54404 15486
rect 54236 15204 54292 15242
rect 54236 15138 54292 15148
rect 54460 15148 54516 24220
rect 54684 24052 54740 24062
rect 54684 23938 54740 23996
rect 54684 23886 54686 23938
rect 54738 23886 54740 23938
rect 54684 23874 54740 23886
rect 54796 23826 54852 23838
rect 54796 23774 54798 23826
rect 54850 23774 54852 23826
rect 54684 23268 54740 23278
rect 54684 23174 54740 23212
rect 54796 21364 54852 23774
rect 54684 21308 54852 21364
rect 54908 23714 54964 23726
rect 54908 23662 54910 23714
rect 54962 23662 54964 23714
rect 54908 21586 54964 23662
rect 55132 23604 55188 23614
rect 55020 23156 55076 23166
rect 55020 22596 55076 23100
rect 55020 22530 55076 22540
rect 55132 21810 55188 23548
rect 55244 23268 55300 24782
rect 55356 24724 55412 24734
rect 55356 24630 55412 24668
rect 55244 23202 55300 23212
rect 55356 23716 55412 23726
rect 55132 21758 55134 21810
rect 55186 21758 55188 21810
rect 55132 21746 55188 21758
rect 55356 23042 55412 23660
rect 55356 22990 55358 23042
rect 55410 22990 55412 23042
rect 55356 21588 55412 22990
rect 55468 22484 55524 29932
rect 55580 29316 55636 29326
rect 55580 29314 55748 29316
rect 55580 29262 55582 29314
rect 55634 29262 55748 29314
rect 55580 29260 55748 29262
rect 55580 29250 55636 29260
rect 55692 28756 55748 29260
rect 55804 29092 55860 30158
rect 55804 29026 55860 29036
rect 55916 30212 55972 30222
rect 55580 27972 55636 27982
rect 55580 27878 55636 27916
rect 55692 26908 55748 28700
rect 55916 28644 55972 30156
rect 56252 30098 56308 30110
rect 56252 30046 56254 30098
rect 56306 30046 56308 30098
rect 55916 28550 55972 28588
rect 56028 28756 56084 28766
rect 56252 28756 56308 30046
rect 56028 28754 56308 28756
rect 56028 28702 56030 28754
rect 56082 28702 56308 28754
rect 56028 28700 56308 28702
rect 55580 26850 55636 26862
rect 55692 26852 55860 26908
rect 55580 26798 55582 26850
rect 55634 26798 55636 26850
rect 55580 23828 55636 26798
rect 55692 26292 55748 26302
rect 55692 26198 55748 26236
rect 55804 25620 55860 26852
rect 55916 26404 55972 26414
rect 55916 26310 55972 26348
rect 56028 26290 56084 28700
rect 56364 28084 56420 38612
rect 61068 38612 61796 38668
rect 60956 32004 61012 32014
rect 60508 29988 60564 29998
rect 59948 29986 60564 29988
rect 59948 29934 60510 29986
rect 60562 29934 60564 29986
rect 59948 29932 60564 29934
rect 59500 29652 59556 29662
rect 59164 29650 59556 29652
rect 59164 29598 59502 29650
rect 59554 29598 59556 29650
rect 59164 29596 59556 29598
rect 56588 29426 56644 29438
rect 56588 29374 56590 29426
rect 56642 29374 56644 29426
rect 56588 29316 56644 29374
rect 56588 29250 56644 29260
rect 57036 29314 57092 29326
rect 57036 29262 57038 29314
rect 57090 29262 57092 29314
rect 56812 29204 56868 29214
rect 56476 28980 56532 28990
rect 56476 28754 56532 28924
rect 56476 28702 56478 28754
rect 56530 28702 56532 28754
rect 56476 28690 56532 28702
rect 56812 28754 56868 29148
rect 56812 28702 56814 28754
rect 56866 28702 56868 28754
rect 56364 28018 56420 28028
rect 56812 26908 56868 28702
rect 56924 28644 56980 28654
rect 56924 27860 56980 28588
rect 57036 28420 57092 29262
rect 57820 28756 57876 28766
rect 58492 28756 58548 28766
rect 57876 28700 57988 28756
rect 57820 28690 57876 28700
rect 57260 28644 57316 28654
rect 57708 28644 57764 28654
rect 57036 28354 57092 28364
rect 57148 28642 57764 28644
rect 57148 28590 57262 28642
rect 57314 28590 57710 28642
rect 57762 28590 57764 28642
rect 57148 28588 57764 28590
rect 57148 27972 57204 28588
rect 57260 28578 57316 28588
rect 57708 28578 57764 28588
rect 56924 27858 57092 27860
rect 56924 27806 56926 27858
rect 56978 27806 57092 27858
rect 56924 27804 57092 27806
rect 56924 27794 56980 27804
rect 56812 26852 56980 26908
rect 56924 26628 56980 26852
rect 56924 26562 56980 26572
rect 56924 26404 56980 26414
rect 56812 26402 56980 26404
rect 56812 26350 56926 26402
rect 56978 26350 56980 26402
rect 56812 26348 56980 26350
rect 56028 26238 56030 26290
rect 56082 26238 56084 26290
rect 55916 25620 55972 25630
rect 55804 25618 55972 25620
rect 55804 25566 55918 25618
rect 55970 25566 55972 25618
rect 55804 25564 55972 25566
rect 55916 25554 55972 25564
rect 56028 25172 56084 26238
rect 56028 25106 56084 25116
rect 56140 26292 56196 26302
rect 55804 24948 55860 24958
rect 55804 24854 55860 24892
rect 55916 24836 55972 24846
rect 55916 24742 55972 24780
rect 56028 24836 56084 24846
rect 56140 24836 56196 26236
rect 56812 25508 56868 26348
rect 56924 26338 56980 26348
rect 57036 25620 57092 27804
rect 57148 27746 57204 27916
rect 57820 28420 57876 28430
rect 57372 27860 57428 27870
rect 57708 27860 57764 27870
rect 57372 27858 57764 27860
rect 57372 27806 57374 27858
rect 57426 27806 57710 27858
rect 57762 27806 57764 27858
rect 57372 27804 57764 27806
rect 57820 27860 57876 28364
rect 57932 27972 57988 28700
rect 58492 28642 58548 28700
rect 58492 28590 58494 28642
rect 58546 28590 58548 28642
rect 58492 28578 58548 28590
rect 59052 28644 59108 28654
rect 59164 28644 59220 29596
rect 59500 29586 59556 29596
rect 59388 29426 59444 29438
rect 59388 29374 59390 29426
rect 59442 29374 59444 29426
rect 59388 28980 59444 29374
rect 59500 29204 59556 29214
rect 59500 29202 59668 29204
rect 59500 29150 59502 29202
rect 59554 29150 59668 29202
rect 59500 29148 59668 29150
rect 59500 29138 59556 29148
rect 59444 28924 59556 28980
rect 59388 28914 59444 28924
rect 59052 28642 59220 28644
rect 59052 28590 59054 28642
rect 59106 28590 59220 28642
rect 59052 28588 59220 28590
rect 59052 28578 59108 28588
rect 58044 28420 58100 28430
rect 58044 28326 58100 28364
rect 59052 28420 59108 28430
rect 58044 27972 58100 27982
rect 57932 27970 58100 27972
rect 57932 27918 58046 27970
rect 58098 27918 58100 27970
rect 57932 27916 58100 27918
rect 58044 27906 58100 27916
rect 58828 27860 58884 27870
rect 57820 27804 57988 27860
rect 57372 27794 57428 27804
rect 57148 27694 57150 27746
rect 57202 27694 57204 27746
rect 57148 27074 57204 27694
rect 57708 27412 57764 27804
rect 57932 27748 57988 27804
rect 57932 27692 58100 27748
rect 57820 27636 57876 27646
rect 57820 27542 57876 27580
rect 57708 27356 57988 27412
rect 57148 27022 57150 27074
rect 57202 27022 57204 27074
rect 57148 27010 57204 27022
rect 57708 27076 57764 27086
rect 57148 26292 57204 26302
rect 57148 26198 57204 26236
rect 57708 26290 57764 27020
rect 57708 26238 57710 26290
rect 57762 26238 57764 26290
rect 57708 26226 57764 26238
rect 57036 25564 57316 25620
rect 57260 25508 57316 25564
rect 57596 25508 57652 25518
rect 57260 25506 57652 25508
rect 57260 25454 57598 25506
rect 57650 25454 57652 25506
rect 57260 25452 57652 25454
rect 56028 24834 56196 24836
rect 56028 24782 56030 24834
rect 56082 24782 56196 24834
rect 56028 24780 56196 24782
rect 56252 25282 56308 25294
rect 56252 25230 56254 25282
rect 56306 25230 56308 25282
rect 56028 24770 56084 24780
rect 55580 23772 55748 23828
rect 55692 23716 55748 23772
rect 55692 23650 55748 23660
rect 55692 23380 55748 23390
rect 55692 23154 55748 23324
rect 55692 23102 55694 23154
rect 55746 23102 55748 23154
rect 55692 23090 55748 23102
rect 55804 23268 55860 23278
rect 55804 22708 55860 23212
rect 56252 23156 56308 25230
rect 56812 24946 56868 25452
rect 57596 25442 57652 25452
rect 57148 25394 57204 25406
rect 57148 25342 57150 25394
rect 57202 25342 57204 25394
rect 57148 25172 57204 25342
rect 57148 25060 57204 25116
rect 57148 25004 57540 25060
rect 56812 24894 56814 24946
rect 56866 24894 56868 24946
rect 56812 24882 56868 24894
rect 57036 24836 57092 24874
rect 57092 24780 57204 24836
rect 57036 24770 57092 24780
rect 56476 24722 56532 24734
rect 56476 24670 56478 24722
rect 56530 24670 56532 24722
rect 56476 23604 56532 24670
rect 56924 24724 56980 24734
rect 56924 24388 56980 24668
rect 56476 23538 56532 23548
rect 56812 24332 56980 24388
rect 57036 24610 57092 24622
rect 57036 24558 57038 24610
rect 57090 24558 57092 24610
rect 55524 22428 55636 22484
rect 55468 22418 55524 22428
rect 55468 21588 55524 21598
rect 54908 21534 54910 21586
rect 54962 21534 54964 21586
rect 54908 21364 54964 21534
rect 54684 20692 54740 21308
rect 54908 21298 54964 21308
rect 55020 21586 55524 21588
rect 55020 21534 55470 21586
rect 55522 21534 55524 21586
rect 55020 21532 55524 21534
rect 54796 20804 54852 20814
rect 54796 20710 54852 20748
rect 54684 20626 54740 20636
rect 54684 19012 54740 19022
rect 54908 19012 54964 19022
rect 54684 19010 54964 19012
rect 54684 18958 54686 19010
rect 54738 18958 54910 19010
rect 54962 18958 54964 19010
rect 54684 18956 54964 18958
rect 54684 17892 54740 18956
rect 54908 18946 54964 18956
rect 55020 18788 55076 21532
rect 55468 21522 55524 21532
rect 55132 21140 55188 21150
rect 55132 20690 55188 21084
rect 55132 20638 55134 20690
rect 55186 20638 55188 20690
rect 55132 20626 55188 20638
rect 55132 19460 55188 19470
rect 55132 19234 55188 19404
rect 55132 19182 55134 19234
rect 55186 19182 55188 19234
rect 55132 19170 55188 19182
rect 55244 19346 55300 19358
rect 55244 19294 55246 19346
rect 55298 19294 55300 19346
rect 54684 17826 54740 17836
rect 54796 18732 55076 18788
rect 54796 15314 54852 18732
rect 55244 17780 55300 19294
rect 55356 19124 55412 19134
rect 55356 19030 55412 19068
rect 55244 17714 55300 17724
rect 55468 17668 55524 17678
rect 55580 17668 55636 22428
rect 55804 21924 55860 22652
rect 55804 21698 55860 21868
rect 55804 21646 55806 21698
rect 55858 21646 55860 21698
rect 55804 21634 55860 21646
rect 56140 23100 56308 23156
rect 56812 23154 56868 24332
rect 56812 23102 56814 23154
rect 56866 23102 56868 23154
rect 56028 21140 56084 21150
rect 55916 20802 55972 20814
rect 55916 20750 55918 20802
rect 55970 20750 55972 20802
rect 55916 20692 55972 20750
rect 55916 20626 55972 20636
rect 56028 19234 56084 21084
rect 56028 19182 56030 19234
rect 56082 19182 56084 19234
rect 55692 19124 55748 19134
rect 55692 19030 55748 19068
rect 55916 19010 55972 19022
rect 55916 18958 55918 19010
rect 55970 18958 55972 19010
rect 55916 18452 55972 18958
rect 56028 19012 56084 19182
rect 56028 18946 56084 18956
rect 55916 18386 55972 18396
rect 56140 18004 56196 23100
rect 56812 23090 56868 23102
rect 56924 23156 56980 23166
rect 56924 23062 56980 23100
rect 56588 23044 56644 23054
rect 55468 17666 55580 17668
rect 55468 17614 55470 17666
rect 55522 17614 55580 17666
rect 55468 17612 55580 17614
rect 55468 17602 55524 17612
rect 55580 17574 55636 17612
rect 56028 17948 56196 18004
rect 56252 23042 56644 23044
rect 56252 22990 56590 23042
rect 56642 22990 56644 23042
rect 56252 22988 56644 22990
rect 56252 18004 56308 22988
rect 56588 22978 56644 22988
rect 57036 22708 57092 24558
rect 57148 23940 57204 24780
rect 57148 23874 57204 23884
rect 57372 24498 57428 24510
rect 57372 24446 57374 24498
rect 57426 24446 57428 24498
rect 57036 22642 57092 22652
rect 57036 22484 57092 22494
rect 57036 22390 57092 22428
rect 57148 22148 57204 22158
rect 56588 21924 56644 21934
rect 56588 21586 56644 21868
rect 57148 21812 57204 22092
rect 56588 21534 56590 21586
rect 56642 21534 56644 21586
rect 56588 21522 56644 21534
rect 56700 21810 57204 21812
rect 56700 21758 57150 21810
rect 57202 21758 57204 21810
rect 56700 21756 57204 21758
rect 56700 21140 56756 21756
rect 57148 21746 57204 21756
rect 57372 21812 57428 24446
rect 57484 23940 57540 25004
rect 57932 24834 57988 27356
rect 58044 27076 58100 27692
rect 58044 27010 58100 27020
rect 58716 26962 58772 26974
rect 58716 26910 58718 26962
rect 58770 26910 58772 26962
rect 58156 26628 58212 26638
rect 58156 26402 58212 26572
rect 58156 26350 58158 26402
rect 58210 26350 58212 26402
rect 58156 26338 58212 26350
rect 58716 26404 58772 26910
rect 58716 26338 58772 26348
rect 58044 26292 58100 26302
rect 58044 25506 58100 26236
rect 58828 25620 58884 27804
rect 59052 27188 59108 28364
rect 59164 27860 59220 28588
rect 59388 28756 59444 28766
rect 59388 28642 59444 28700
rect 59388 28590 59390 28642
rect 59442 28590 59444 28642
rect 59388 28578 59444 28590
rect 59276 27860 59332 27870
rect 59164 27858 59332 27860
rect 59164 27806 59278 27858
rect 59330 27806 59332 27858
rect 59164 27804 59332 27806
rect 58828 25564 58996 25620
rect 58044 25454 58046 25506
rect 58098 25454 58100 25506
rect 58044 25442 58100 25454
rect 58492 25506 58548 25518
rect 58492 25454 58494 25506
rect 58546 25454 58548 25506
rect 57932 24782 57934 24834
rect 57986 24782 57988 24834
rect 57708 24724 57764 24734
rect 57708 24630 57764 24668
rect 57708 24052 57764 24062
rect 57596 23940 57652 23950
rect 57484 23938 57652 23940
rect 57484 23886 57598 23938
rect 57650 23886 57652 23938
rect 57484 23884 57652 23886
rect 57596 23874 57652 23884
rect 57372 21252 57428 21756
rect 57708 21700 57764 23996
rect 57820 23268 57876 23278
rect 57820 23174 57876 23212
rect 57932 23156 57988 24782
rect 58156 25396 58212 25406
rect 58156 23938 58212 25340
rect 58492 24948 58548 25454
rect 58268 24836 58324 24846
rect 58268 24742 58324 24780
rect 58492 24722 58548 24892
rect 58492 24670 58494 24722
rect 58546 24670 58548 24722
rect 58492 24658 58548 24670
rect 58828 25394 58884 25406
rect 58828 25342 58830 25394
rect 58882 25342 58884 25394
rect 58828 24724 58884 25342
rect 58828 24658 58884 24668
rect 58604 24052 58660 24062
rect 58604 23958 58660 23996
rect 58156 23886 58158 23938
rect 58210 23886 58212 23938
rect 58156 23874 58212 23886
rect 58380 23828 58436 23838
rect 57932 23090 57988 23100
rect 58268 23380 58324 23390
rect 58268 22258 58324 23324
rect 58380 23266 58436 23772
rect 58380 23214 58382 23266
rect 58434 23214 58436 23266
rect 58380 23202 58436 23214
rect 58604 23154 58660 23166
rect 58604 23102 58606 23154
rect 58658 23102 58660 23154
rect 58604 22372 58660 23102
rect 58268 22206 58270 22258
rect 58322 22206 58324 22258
rect 58268 22194 58324 22206
rect 58380 22316 58660 22372
rect 58828 23154 58884 23166
rect 58828 23102 58830 23154
rect 58882 23102 58884 23154
rect 58380 22260 58436 22316
rect 57372 21186 57428 21196
rect 57484 21644 57764 21700
rect 56588 21084 56756 21140
rect 56364 20802 56420 20814
rect 56364 20750 56366 20802
rect 56418 20750 56420 20802
rect 56364 20020 56420 20750
rect 56476 20244 56532 20254
rect 56588 20244 56644 21084
rect 57372 20916 57428 20926
rect 57484 20916 57540 21644
rect 57372 20914 57484 20916
rect 57372 20862 57374 20914
rect 57426 20862 57484 20914
rect 57372 20860 57484 20862
rect 57372 20850 57428 20860
rect 57484 20822 57540 20860
rect 58268 20916 58324 20926
rect 58268 20822 58324 20860
rect 56476 20242 56644 20244
rect 56476 20190 56478 20242
rect 56530 20190 56644 20242
rect 56476 20188 56644 20190
rect 56812 20578 56868 20590
rect 56812 20526 56814 20578
rect 56866 20526 56868 20578
rect 56476 20178 56532 20188
rect 56700 20132 56756 20142
rect 56588 20130 56756 20132
rect 56588 20078 56702 20130
rect 56754 20078 56756 20130
rect 56588 20076 56756 20078
rect 56588 20020 56644 20076
rect 56700 20066 56756 20076
rect 56364 19964 56644 20020
rect 56588 19236 56644 19964
rect 56812 20018 56868 20526
rect 56812 19966 56814 20018
rect 56866 19966 56868 20018
rect 56812 19572 56868 19966
rect 56588 19170 56644 19180
rect 56700 19516 56868 19572
rect 57484 20580 57540 20590
rect 56700 18674 56756 19516
rect 57484 19348 57540 20524
rect 58268 19572 58324 19582
rect 58380 19572 58436 22204
rect 58604 22148 58660 22158
rect 58604 22054 58660 22092
rect 58828 21812 58884 23102
rect 58940 22820 58996 25564
rect 59052 25506 59108 27132
rect 59276 26908 59332 27804
rect 59500 27858 59556 28924
rect 59500 27806 59502 27858
rect 59554 27806 59556 27858
rect 59500 27794 59556 27806
rect 59388 27412 59444 27422
rect 59388 27186 59444 27356
rect 59612 27300 59668 29148
rect 59724 28418 59780 28430
rect 59724 28366 59726 28418
rect 59778 28366 59780 28418
rect 59724 27412 59780 28366
rect 59836 27860 59892 27870
rect 59836 27766 59892 27804
rect 59724 27356 59892 27412
rect 59612 27244 59780 27300
rect 59388 27134 59390 27186
rect 59442 27134 59444 27186
rect 59388 27122 59444 27134
rect 59612 27074 59668 27086
rect 59612 27022 59614 27074
rect 59666 27022 59668 27074
rect 59500 26964 59556 26974
rect 59276 26852 59556 26908
rect 59388 26290 59444 26852
rect 59388 26238 59390 26290
rect 59442 26238 59444 26290
rect 59388 26226 59444 26238
rect 59612 26068 59668 27022
rect 59612 26002 59668 26012
rect 59052 25454 59054 25506
rect 59106 25454 59108 25506
rect 59052 25442 59108 25454
rect 59500 25508 59556 25518
rect 59724 25508 59780 27244
rect 59556 25452 59780 25508
rect 59500 25414 59556 25452
rect 59164 25172 59220 25182
rect 59164 24610 59220 25116
rect 59500 24948 59556 24958
rect 59836 24948 59892 27356
rect 59948 27298 60004 29932
rect 60508 29922 60564 29932
rect 60732 28642 60788 28654
rect 60732 28590 60734 28642
rect 60786 28590 60788 28642
rect 60620 27860 60676 27870
rect 60620 27766 60676 27804
rect 59948 27246 59950 27298
rect 60002 27246 60004 27298
rect 59948 27234 60004 27246
rect 60508 27412 60564 27422
rect 60732 27412 60788 28590
rect 60564 27356 60788 27412
rect 60844 27858 60900 27870
rect 60844 27806 60846 27858
rect 60898 27806 60900 27858
rect 60844 27524 60900 27806
rect 60508 26740 60564 27356
rect 60844 27186 60900 27468
rect 60844 27134 60846 27186
rect 60898 27134 60900 27186
rect 60844 27122 60900 27134
rect 60956 26908 61012 31948
rect 61068 30210 61124 38612
rect 61068 30158 61070 30210
rect 61122 30158 61124 30210
rect 61068 30146 61124 30158
rect 62076 29876 62132 29886
rect 61068 27860 61124 27870
rect 61068 27766 61124 27804
rect 62076 27746 62132 29820
rect 62972 29876 63028 55244
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 68012 30548 68068 56140
rect 70588 56082 70644 56094
rect 70588 56030 70590 56082
rect 70642 56030 70644 56082
rect 70588 55468 70644 56030
rect 74172 55972 74228 59200
rect 77980 56196 78036 59200
rect 81276 56476 81540 56486
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81276 56410 81540 56420
rect 81788 56308 81844 59200
rect 81788 56242 81844 56252
rect 83020 56308 83076 56318
rect 83020 56214 83076 56252
rect 78204 56196 78260 56206
rect 77980 56194 78260 56196
rect 77980 56142 78206 56194
rect 78258 56142 78260 56194
rect 77980 56140 78260 56142
rect 76972 56082 77028 56094
rect 76972 56030 76974 56082
rect 77026 56030 77028 56082
rect 74620 55972 74676 55982
rect 74172 55970 74676 55972
rect 74172 55918 74622 55970
rect 74674 55918 74676 55970
rect 74172 55916 74676 55918
rect 74620 55906 74676 55916
rect 70476 55412 70644 55468
rect 76972 55468 77028 56030
rect 76972 55412 77252 55468
rect 69804 55300 69860 55310
rect 69804 55206 69860 55244
rect 70140 55298 70196 55310
rect 70140 55246 70142 55298
rect 70194 55246 70196 55298
rect 70140 55188 70196 55246
rect 70140 55122 70196 55132
rect 70364 55188 70420 55198
rect 70476 55188 70532 55412
rect 71036 55300 71092 55310
rect 71036 55206 71092 55244
rect 70364 55186 70532 55188
rect 70364 55134 70366 55186
rect 70418 55134 70532 55186
rect 70364 55132 70532 55134
rect 70700 55188 70756 55198
rect 70364 55122 70420 55132
rect 70700 55094 70756 55132
rect 71484 55188 71540 55198
rect 71484 55094 71540 55132
rect 77196 55074 77252 55412
rect 77980 55410 78036 56140
rect 78204 56130 78260 56140
rect 78540 56194 78596 56206
rect 78540 56142 78542 56194
rect 78594 56142 78596 56194
rect 78540 55468 78596 56142
rect 82012 56082 82068 56094
rect 82012 56030 82014 56082
rect 82066 56030 82068 56082
rect 82012 55468 82068 56030
rect 85596 55972 85652 59200
rect 89404 56308 89460 59200
rect 89628 56308 89684 56318
rect 89404 56306 89684 56308
rect 89404 56254 89630 56306
rect 89682 56254 89684 56306
rect 89404 56252 89684 56254
rect 88396 56082 88452 56094
rect 88396 56030 88398 56082
rect 88450 56030 88452 56082
rect 86044 55972 86100 55982
rect 85596 55970 86100 55972
rect 85596 55918 86046 55970
rect 86098 55918 86100 55970
rect 85596 55916 86100 55918
rect 86044 55906 86100 55916
rect 78540 55412 78708 55468
rect 77980 55358 77982 55410
rect 78034 55358 78036 55410
rect 77980 55346 78036 55358
rect 77196 55022 77198 55074
rect 77250 55022 77252 55074
rect 74620 30996 74676 31006
rect 74060 30884 74116 30894
rect 68012 30482 68068 30492
rect 69468 30772 69524 30782
rect 62972 29810 63028 29820
rect 65324 29314 65380 29326
rect 65324 29262 65326 29314
rect 65378 29262 65380 29314
rect 62636 28644 62692 28654
rect 62860 28644 62916 28654
rect 62076 27694 62078 27746
rect 62130 27694 62132 27746
rect 62076 27682 62132 27694
rect 62524 28642 62916 28644
rect 62524 28590 62638 28642
rect 62690 28590 62862 28642
rect 62914 28590 62916 28642
rect 62524 28588 62916 28590
rect 60508 26674 60564 26684
rect 60620 26852 61012 26908
rect 61180 27300 61236 27310
rect 60508 26290 60564 26302
rect 60508 26238 60510 26290
rect 60562 26238 60564 26290
rect 59556 24892 59892 24948
rect 59948 26178 60004 26190
rect 59948 26126 59950 26178
rect 60002 26126 60004 26178
rect 59500 24722 59556 24892
rect 59500 24670 59502 24722
rect 59554 24670 59556 24722
rect 59500 24658 59556 24670
rect 59164 24558 59166 24610
rect 59218 24558 59220 24610
rect 59164 24546 59220 24558
rect 59388 23716 59444 23726
rect 59276 23714 59444 23716
rect 59276 23662 59390 23714
rect 59442 23662 59444 23714
rect 59276 23660 59444 23662
rect 59052 23268 59108 23278
rect 59276 23268 59332 23660
rect 59388 23650 59444 23660
rect 59052 23266 59332 23268
rect 59052 23214 59054 23266
rect 59106 23214 59332 23266
rect 59052 23212 59332 23214
rect 59052 23202 59108 23212
rect 59164 23044 59220 23054
rect 59164 22950 59220 22988
rect 59276 22820 59332 23212
rect 59948 23268 60004 26126
rect 60508 25508 60564 26238
rect 60508 25442 60564 25452
rect 60284 24948 60340 24958
rect 59948 23202 60004 23212
rect 60060 23828 60116 23838
rect 58940 22754 58996 22764
rect 59164 22764 59332 22820
rect 59836 23156 59892 23166
rect 58828 21746 58884 21756
rect 59052 22708 59108 22718
rect 59052 21924 59108 22652
rect 59052 21586 59108 21868
rect 59052 21534 59054 21586
rect 59106 21534 59108 21586
rect 59052 21522 59108 21534
rect 59164 21140 59220 22764
rect 59836 22484 59892 23100
rect 59836 22418 59892 22428
rect 60060 22370 60116 23772
rect 60284 23156 60340 24892
rect 60620 24164 60676 26852
rect 61180 26292 61236 27244
rect 61628 27188 61684 27198
rect 61628 27094 61684 27132
rect 61964 27186 62020 27198
rect 61964 27134 61966 27186
rect 62018 27134 62020 27186
rect 61292 27074 61348 27086
rect 61292 27022 61294 27074
rect 61346 27022 61348 27074
rect 61292 26852 61348 27022
rect 61852 26964 61908 27002
rect 61852 26898 61908 26908
rect 61292 26786 61348 26796
rect 61964 26852 62020 27134
rect 62524 26908 62580 28588
rect 62636 28578 62692 28588
rect 62860 28578 62916 28588
rect 63644 28642 63700 28654
rect 63644 28590 63646 28642
rect 63698 28590 63700 28642
rect 63196 28084 63252 28094
rect 62748 27524 62804 27534
rect 62748 27186 62804 27468
rect 62748 27134 62750 27186
rect 62802 27134 62804 27186
rect 62748 27122 62804 27134
rect 63196 27186 63252 28028
rect 63644 28084 63700 28590
rect 65324 28196 65380 29262
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 68236 28868 68292 28878
rect 64988 28140 65380 28196
rect 65996 28418 66052 28430
rect 65996 28366 65998 28418
rect 66050 28366 66052 28418
rect 63644 28018 63700 28028
rect 63980 28084 64036 28094
rect 64764 28084 64820 28094
rect 63980 28082 64708 28084
rect 63980 28030 63982 28082
rect 64034 28030 64708 28082
rect 63980 28028 64708 28030
rect 63980 28018 64036 28028
rect 63756 27972 63812 27982
rect 63756 27878 63812 27916
rect 64652 27970 64708 28028
rect 64764 27990 64820 28028
rect 64652 27918 64654 27970
rect 64706 27918 64708 27970
rect 64652 27906 64708 27918
rect 63644 27858 63700 27870
rect 63644 27806 63646 27858
rect 63698 27806 63700 27858
rect 63308 27748 63364 27758
rect 63644 27748 63700 27806
rect 63308 27746 63700 27748
rect 63308 27694 63310 27746
rect 63362 27694 63700 27746
rect 63308 27692 63700 27694
rect 64540 27858 64596 27870
rect 64540 27806 64542 27858
rect 64594 27806 64596 27858
rect 64540 27748 64596 27806
rect 64988 27748 65044 28140
rect 65660 28084 65716 28094
rect 65324 27972 65380 27982
rect 65324 27878 65380 27916
rect 65100 27860 65156 27870
rect 65100 27766 65156 27804
rect 65660 27858 65716 28028
rect 65996 27972 66052 28366
rect 66444 28418 66500 28430
rect 66444 28366 66446 28418
rect 66498 28366 66500 28418
rect 66108 28196 66164 28206
rect 66444 28196 66500 28366
rect 66164 28140 66500 28196
rect 67676 28420 67732 28430
rect 66108 28082 66164 28140
rect 66108 28030 66110 28082
rect 66162 28030 66164 28082
rect 66108 28018 66164 28030
rect 65996 27906 66052 27916
rect 65660 27806 65662 27858
rect 65714 27806 65716 27858
rect 65660 27794 65716 27806
rect 65884 27860 65940 27870
rect 65884 27766 65940 27804
rect 66220 27860 66276 27870
rect 66220 27766 66276 27804
rect 67116 27858 67172 27870
rect 67116 27806 67118 27858
rect 67170 27806 67172 27858
rect 64540 27692 65044 27748
rect 63308 27636 63364 27692
rect 63308 27570 63364 27580
rect 63196 27134 63198 27186
rect 63250 27134 63252 27186
rect 63196 27076 63252 27134
rect 63644 27188 63700 27692
rect 63644 27094 63700 27132
rect 64316 27186 64372 27198
rect 64316 27134 64318 27186
rect 64370 27134 64372 27186
rect 63196 27010 63252 27020
rect 63980 27076 64036 27086
rect 64316 27076 64372 27134
rect 64652 27076 64708 27086
rect 64316 27074 64708 27076
rect 64316 27022 64654 27074
rect 64706 27022 64708 27074
rect 64316 27020 64708 27022
rect 63980 26982 64036 27020
rect 64652 27010 64708 27020
rect 64764 27076 64820 27692
rect 64764 27010 64820 27020
rect 65660 27634 65716 27646
rect 65660 27582 65662 27634
rect 65714 27582 65716 27634
rect 65660 26962 65716 27582
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 66444 27188 66500 27198
rect 66444 27094 66500 27132
rect 65660 26910 65662 26962
rect 65714 26910 65716 26962
rect 62524 26852 62916 26908
rect 65660 26898 65716 26910
rect 67116 26964 67172 27806
rect 67116 26908 67284 26964
rect 67564 26962 67620 26974
rect 67564 26910 67566 26962
rect 67618 26910 67620 26962
rect 61180 26226 61236 26236
rect 61964 26292 62020 26796
rect 62636 26740 62692 26750
rect 62412 26292 62468 26302
rect 61964 26226 62020 26236
rect 62188 26290 62468 26292
rect 62188 26238 62414 26290
rect 62466 26238 62468 26290
rect 62188 26236 62468 26238
rect 60956 26178 61012 26190
rect 60956 26126 60958 26178
rect 61010 26126 61012 26178
rect 60956 26068 61012 26126
rect 60732 25284 60788 25294
rect 60732 25190 60788 25228
rect 60284 23062 60340 23100
rect 60508 24108 60676 24164
rect 60956 24164 61012 26012
rect 61516 26178 61572 26190
rect 61516 26126 61518 26178
rect 61570 26126 61572 26178
rect 61516 26068 61572 26126
rect 61516 26002 61572 26012
rect 61180 25956 61236 25966
rect 61180 25620 61236 25900
rect 62188 25844 62244 26236
rect 62412 26226 62468 26236
rect 62188 25730 62244 25788
rect 62188 25678 62190 25730
rect 62242 25678 62244 25730
rect 62188 25666 62244 25678
rect 61180 25618 61460 25620
rect 61180 25566 61182 25618
rect 61234 25566 61460 25618
rect 61180 25564 61460 25566
rect 61180 25554 61236 25564
rect 60060 22318 60062 22370
rect 60114 22318 60116 22370
rect 60060 22306 60116 22318
rect 60396 23044 60452 23054
rect 60396 22370 60452 22988
rect 60396 22318 60398 22370
rect 60450 22318 60452 22370
rect 60396 22306 60452 22318
rect 59724 22260 59780 22270
rect 59612 22258 59780 22260
rect 59612 22206 59726 22258
rect 59778 22206 59780 22258
rect 59612 22204 59780 22206
rect 59388 22148 59444 22158
rect 58940 21084 59220 21140
rect 59276 22092 59388 22148
rect 58828 20580 58884 20590
rect 58324 19516 58436 19572
rect 58492 19516 58772 19572
rect 58268 19506 58324 19516
rect 57484 19282 57540 19292
rect 58268 19124 58324 19134
rect 58268 19030 58324 19068
rect 56700 18622 56702 18674
rect 56754 18622 56756 18674
rect 56700 18610 56756 18622
rect 58156 18900 58212 18910
rect 56924 18452 56980 18462
rect 56812 18450 56980 18452
rect 56812 18398 56926 18450
rect 56978 18398 56980 18450
rect 56812 18396 56980 18398
rect 56812 18340 56868 18396
rect 56924 18386 56980 18396
rect 54796 15262 54798 15314
rect 54850 15262 54852 15314
rect 54796 15250 54852 15262
rect 55020 16996 55076 17006
rect 55020 15148 55076 16940
rect 55692 16884 55748 16894
rect 55692 16770 55748 16828
rect 55692 16718 55694 16770
rect 55746 16718 55748 16770
rect 55692 16706 55748 16718
rect 55916 16436 55972 16446
rect 55916 16210 55972 16380
rect 56028 16324 56084 17948
rect 56252 17938 56308 17948
rect 56588 18228 56644 18238
rect 56140 17780 56196 17790
rect 56140 17686 56196 17724
rect 56588 16884 56644 18172
rect 56700 17668 56756 17678
rect 56700 17108 56756 17612
rect 56812 17556 56868 18284
rect 57372 18338 57428 18350
rect 57372 18286 57374 18338
rect 57426 18286 57428 18338
rect 56812 17490 56868 17500
rect 57260 18226 57316 18238
rect 57260 18174 57262 18226
rect 57314 18174 57316 18226
rect 57260 18116 57316 18174
rect 57372 18228 57428 18286
rect 57820 18340 57876 18350
rect 57820 18246 57876 18284
rect 57372 18162 57428 18172
rect 57260 17220 57316 18060
rect 57260 17154 57316 17164
rect 57596 17332 57652 17342
rect 56700 17014 56756 17052
rect 57596 16994 57652 17276
rect 57596 16942 57598 16994
rect 57650 16942 57652 16994
rect 57596 16930 57652 16942
rect 56588 16818 56644 16828
rect 57036 16884 57092 16894
rect 57036 16790 57092 16828
rect 56028 16258 56084 16268
rect 56588 16436 56644 16446
rect 55916 16158 55918 16210
rect 55970 16158 55972 16210
rect 55916 16146 55972 16158
rect 56588 15988 56644 16380
rect 57484 16100 57540 16110
rect 57484 16006 57540 16044
rect 56924 15988 56980 15998
rect 56588 15986 57204 15988
rect 56588 15934 56590 15986
rect 56642 15934 56926 15986
rect 56978 15934 57204 15986
rect 56588 15932 57204 15934
rect 56588 15922 56644 15932
rect 56924 15922 56980 15932
rect 56252 15874 56308 15886
rect 56252 15822 56254 15874
rect 56306 15822 56308 15874
rect 56252 15764 56308 15822
rect 56252 15698 56308 15708
rect 55132 15540 55188 15550
rect 55132 15446 55188 15484
rect 57148 15540 57204 15932
rect 57372 15540 57428 15550
rect 57148 15538 57428 15540
rect 57148 15486 57150 15538
rect 57202 15486 57374 15538
rect 57426 15486 57428 15538
rect 57148 15484 57428 15486
rect 57148 15474 57204 15484
rect 57372 15474 57428 15484
rect 57708 15426 57764 15438
rect 57708 15374 57710 15426
rect 57762 15374 57764 15426
rect 54460 15092 54852 15148
rect 55020 15092 55188 15148
rect 54012 14802 54068 14812
rect 54012 14308 54068 14318
rect 53788 14306 54068 14308
rect 53788 14254 54014 14306
rect 54066 14254 54068 14306
rect 53788 14252 54068 14254
rect 53116 13794 53172 13804
rect 53004 12964 53060 12974
rect 53788 12964 53844 12974
rect 52780 12562 52836 12572
rect 52892 12908 53004 12964
rect 52892 12180 52948 12908
rect 53004 12870 53060 12908
rect 53228 12962 53844 12964
rect 53228 12910 53790 12962
rect 53842 12910 53844 12962
rect 53228 12908 53844 12910
rect 54012 12964 54068 14252
rect 54572 14308 54628 14318
rect 54572 14214 54628 14252
rect 54460 13636 54516 13646
rect 54460 13634 54628 13636
rect 54460 13582 54462 13634
rect 54514 13582 54628 13634
rect 54460 13580 54628 13582
rect 54460 13570 54516 13580
rect 54348 12964 54404 12974
rect 54012 12908 54348 12964
rect 52668 11956 52724 11966
rect 52668 11394 52724 11900
rect 52780 11508 52836 11518
rect 52780 11414 52836 11452
rect 52668 11342 52670 11394
rect 52722 11342 52724 11394
rect 52668 11330 52724 11342
rect 52892 10948 52948 12124
rect 53004 11396 53060 11406
rect 53004 11302 53060 11340
rect 53228 11394 53284 12908
rect 53788 12898 53844 12908
rect 53452 12738 53508 12750
rect 53452 12686 53454 12738
rect 53506 12686 53508 12738
rect 53452 12628 53508 12686
rect 53452 12562 53508 12572
rect 53676 12738 53732 12750
rect 53676 12686 53678 12738
rect 53730 12686 53732 12738
rect 53564 12516 53620 12526
rect 53228 11342 53230 11394
rect 53282 11342 53284 11394
rect 53228 11330 53284 11342
rect 53452 12404 53508 12414
rect 52444 8260 52500 9884
rect 52780 10892 52948 10948
rect 52780 9826 52836 10892
rect 52892 10500 52948 10510
rect 53340 10500 53396 10510
rect 52892 10498 53396 10500
rect 52892 10446 52894 10498
rect 52946 10446 53342 10498
rect 53394 10446 53396 10498
rect 52892 10444 53396 10446
rect 52892 10434 52948 10444
rect 53340 10388 53396 10444
rect 53340 10322 53396 10332
rect 52780 9774 52782 9826
rect 52834 9774 52836 9826
rect 52780 9762 52836 9774
rect 52556 9268 52612 9278
rect 52556 9174 52612 9212
rect 52892 9154 52948 9166
rect 52892 9102 52894 9154
rect 52946 9102 52948 9154
rect 52780 9044 52836 9054
rect 52780 8950 52836 8988
rect 52556 8818 52612 8830
rect 52556 8766 52558 8818
rect 52610 8766 52612 8818
rect 52556 8484 52612 8766
rect 52556 8428 52836 8484
rect 52108 8204 52500 8260
rect 52780 8260 52836 8428
rect 51884 8146 51940 8158
rect 51884 8094 51886 8146
rect 51938 8094 51940 8146
rect 51884 7364 51940 8094
rect 51996 8034 52052 8046
rect 51996 7982 51998 8034
rect 52050 7982 52052 8034
rect 51996 7924 52052 7982
rect 51996 7858 52052 7868
rect 52108 7474 52164 8204
rect 52780 8194 52836 8204
rect 52668 8146 52724 8158
rect 52668 8094 52670 8146
rect 52722 8094 52724 8146
rect 52220 8034 52276 8046
rect 52220 7982 52222 8034
rect 52274 7982 52276 8034
rect 52220 7924 52276 7982
rect 52220 7868 52388 7924
rect 52108 7422 52110 7474
rect 52162 7422 52164 7474
rect 52108 7410 52164 7422
rect 52220 7700 52276 7710
rect 51884 7298 51940 7308
rect 52108 6804 52164 6814
rect 52108 6710 52164 6748
rect 52108 6468 52164 6478
rect 51884 6020 51940 6030
rect 51884 5926 51940 5964
rect 51772 5122 52052 5124
rect 51772 5070 51774 5122
rect 51826 5070 52052 5122
rect 51772 5068 52052 5070
rect 51772 5058 51828 5068
rect 51548 5010 51604 5022
rect 51548 4958 51550 5010
rect 51602 4958 51604 5010
rect 51548 4788 51604 4958
rect 51548 4722 51604 4732
rect 51268 4396 51380 4452
rect 51212 4386 51268 4396
rect 51324 4338 51380 4396
rect 51324 4286 51326 4338
rect 51378 4286 51380 4338
rect 51324 4274 51380 4286
rect 51884 4340 51940 4350
rect 51884 4246 51940 4284
rect 51212 3556 51268 3566
rect 51100 3554 51268 3556
rect 51100 3502 51214 3554
rect 51266 3502 51268 3554
rect 51100 3500 51268 3502
rect 51212 3490 51268 3500
rect 51548 3444 51604 3454
rect 51548 3350 51604 3388
rect 51996 2884 52052 5068
rect 52108 3554 52164 6412
rect 52108 3502 52110 3554
rect 52162 3502 52164 3554
rect 52108 3490 52164 3502
rect 51996 2818 52052 2828
rect 52220 800 52276 7644
rect 52332 7588 52388 7868
rect 52332 7532 52500 7588
rect 52332 7364 52388 7374
rect 52332 7140 52388 7308
rect 52332 5124 52388 7084
rect 52444 6468 52500 7532
rect 52556 7476 52612 7486
rect 52556 7382 52612 7420
rect 52668 6916 52724 8094
rect 52444 6402 52500 6412
rect 52556 6860 52724 6916
rect 52780 8034 52836 8046
rect 52780 7982 52782 8034
rect 52834 7982 52836 8034
rect 52556 6132 52612 6860
rect 52556 6066 52612 6076
rect 52668 6692 52724 6702
rect 52668 5908 52724 6636
rect 52780 6020 52836 7982
rect 52892 6804 52948 9102
rect 53116 9042 53172 9054
rect 53116 8990 53118 9042
rect 53170 8990 53172 9042
rect 53004 8148 53060 8158
rect 53004 8054 53060 8092
rect 53116 8036 53172 8990
rect 53228 8372 53284 8382
rect 53228 8148 53284 8316
rect 53228 8054 53284 8092
rect 53116 7970 53172 7980
rect 52892 6738 52948 6748
rect 53004 7364 53060 7374
rect 52780 5954 52836 5964
rect 53004 6018 53060 7308
rect 53452 7364 53508 12348
rect 53564 11956 53620 12460
rect 53676 12068 53732 12686
rect 53900 12740 53956 12750
rect 53900 12738 54068 12740
rect 53900 12686 53902 12738
rect 53954 12686 54068 12738
rect 53900 12684 54068 12686
rect 53900 12674 53956 12684
rect 53900 12068 53956 12078
rect 53676 12066 53956 12068
rect 53676 12014 53902 12066
rect 53954 12014 53956 12066
rect 53676 12012 53956 12014
rect 53564 11394 53620 11900
rect 53900 11956 53956 12012
rect 53900 11890 53956 11900
rect 53564 11342 53566 11394
rect 53618 11342 53620 11394
rect 53564 11330 53620 11342
rect 53788 11620 53844 11630
rect 53788 11394 53844 11564
rect 53788 11342 53790 11394
rect 53842 11342 53844 11394
rect 53788 11330 53844 11342
rect 53676 11170 53732 11182
rect 53676 11118 53678 11170
rect 53730 11118 53732 11170
rect 53676 10836 53732 11118
rect 53564 10780 53732 10836
rect 54012 10836 54068 12684
rect 54124 11284 54180 11294
rect 54124 11190 54180 11228
rect 53564 9938 53620 10780
rect 54012 10770 54068 10780
rect 54124 10836 54180 10846
rect 54236 10836 54292 12908
rect 54348 12870 54404 12908
rect 54460 12628 54516 12638
rect 54460 12402 54516 12572
rect 54460 12350 54462 12402
rect 54514 12350 54516 12402
rect 54460 12338 54516 12350
rect 54572 11394 54628 13580
rect 54684 12516 54740 12526
rect 54684 12290 54740 12460
rect 54684 12238 54686 12290
rect 54738 12238 54740 12290
rect 54684 12226 54740 12238
rect 54572 11342 54574 11394
rect 54626 11342 54628 11394
rect 54124 10834 54292 10836
rect 54124 10782 54126 10834
rect 54178 10782 54292 10834
rect 54124 10780 54292 10782
rect 54460 10836 54516 10846
rect 54124 10770 54180 10780
rect 54460 10742 54516 10780
rect 53788 10724 53844 10734
rect 53788 10630 53844 10668
rect 53564 9886 53566 9938
rect 53618 9886 53620 9938
rect 53564 9874 53620 9886
rect 53676 10612 53732 10622
rect 53564 8930 53620 8942
rect 53564 8878 53566 8930
rect 53618 8878 53620 8930
rect 53564 8258 53620 8878
rect 53564 8206 53566 8258
rect 53618 8206 53620 8258
rect 53564 8194 53620 8206
rect 53452 7298 53508 7308
rect 53564 7474 53620 7486
rect 53564 7422 53566 7474
rect 53618 7422 53620 7474
rect 53340 6804 53396 6814
rect 53564 6804 53620 7422
rect 53396 6748 53620 6804
rect 53340 6738 53396 6748
rect 53676 6690 53732 10556
rect 54572 10612 54628 11342
rect 54572 10546 54628 10556
rect 54796 10834 54852 15092
rect 55132 13748 55188 15092
rect 57708 14754 57764 15374
rect 58156 14980 58212 18844
rect 58380 18676 58436 18686
rect 58380 18450 58436 18620
rect 58380 18398 58382 18450
rect 58434 18398 58436 18450
rect 58380 18386 58436 18398
rect 58492 18340 58548 19516
rect 58604 19346 58660 19358
rect 58604 19294 58606 19346
rect 58658 19294 58660 19346
rect 58604 18564 58660 19294
rect 58716 19234 58772 19516
rect 58716 19182 58718 19234
rect 58770 19182 58772 19234
rect 58716 19170 58772 19182
rect 58604 18470 58660 18508
rect 58716 18562 58772 18574
rect 58716 18510 58718 18562
rect 58770 18510 58772 18562
rect 58380 17780 58436 17790
rect 58492 17780 58548 18284
rect 58380 17778 58548 17780
rect 58380 17726 58382 17778
rect 58434 17726 58548 17778
rect 58380 17724 58548 17726
rect 58716 17780 58772 18510
rect 58828 17892 58884 20524
rect 58940 19572 58996 21084
rect 59052 20916 59108 20926
rect 59052 20802 59108 20860
rect 59052 20750 59054 20802
rect 59106 20750 59108 20802
rect 59052 20468 59108 20750
rect 59052 20402 59108 20412
rect 59164 20578 59220 20590
rect 59164 20526 59166 20578
rect 59218 20526 59220 20578
rect 59164 20020 59220 20526
rect 59164 19954 59220 19964
rect 59052 19572 59108 19582
rect 58940 19516 59052 19572
rect 59052 19506 59108 19516
rect 59276 19460 59332 22092
rect 59388 22054 59444 22092
rect 59612 21810 59668 22204
rect 59724 22194 59780 22204
rect 59836 22260 59892 22270
rect 59836 22166 59892 22204
rect 59612 21758 59614 21810
rect 59666 21758 59668 21810
rect 59612 21746 59668 21758
rect 60060 21924 60116 21934
rect 60060 21698 60116 21868
rect 60060 21646 60062 21698
rect 60114 21646 60116 21698
rect 60060 21634 60116 21646
rect 59500 21588 59556 21598
rect 59500 21494 59556 21532
rect 59724 21586 59780 21598
rect 60284 21588 60340 21598
rect 59724 21534 59726 21586
rect 59778 21534 59780 21586
rect 59388 20804 59444 20814
rect 59388 20710 59444 20748
rect 59612 20802 59668 20814
rect 59612 20750 59614 20802
rect 59666 20750 59668 20802
rect 59388 20580 59444 20590
rect 59612 20580 59668 20750
rect 59724 20804 59780 21534
rect 60172 21586 60340 21588
rect 60172 21534 60286 21586
rect 60338 21534 60340 21586
rect 60172 21532 60340 21534
rect 60172 21140 60228 21532
rect 60284 21522 60340 21532
rect 60508 21586 60564 24108
rect 60956 24098 61012 24108
rect 60956 23828 61012 23838
rect 60956 23734 61012 23772
rect 61068 23714 61124 23726
rect 61292 23716 61348 23726
rect 61068 23662 61070 23714
rect 61122 23662 61124 23714
rect 60956 23044 61012 23054
rect 60620 23042 61012 23044
rect 60620 22990 60958 23042
rect 61010 22990 61012 23042
rect 60620 22988 61012 22990
rect 60620 22482 60676 22988
rect 60956 22978 61012 22988
rect 61068 23044 61124 23662
rect 61068 22978 61124 22988
rect 61180 23714 61348 23716
rect 61180 23662 61294 23714
rect 61346 23662 61348 23714
rect 61180 23660 61348 23662
rect 61180 22820 61236 23660
rect 61292 23650 61348 23660
rect 61404 23380 61460 25564
rect 62636 25618 62692 26684
rect 62636 25566 62638 25618
rect 62690 25566 62692 25618
rect 62636 25554 62692 25566
rect 61852 25508 61908 25518
rect 61852 25506 62244 25508
rect 61852 25454 61854 25506
rect 61906 25454 62244 25506
rect 61852 25452 62244 25454
rect 61852 25442 61908 25452
rect 61628 25394 61684 25406
rect 61628 25342 61630 25394
rect 61682 25342 61684 25394
rect 61628 25284 61684 25342
rect 61628 25218 61684 25228
rect 62188 24612 62244 25452
rect 62860 24948 62916 26852
rect 64204 26852 64260 26862
rect 64204 26758 64260 26796
rect 67004 26850 67060 26862
rect 67228 26852 67508 26908
rect 67004 26798 67006 26850
rect 67058 26798 67060 26850
rect 64428 26740 64484 26750
rect 63644 26628 63700 26638
rect 63644 26402 63700 26572
rect 63644 26350 63646 26402
rect 63698 26350 63700 26402
rect 63644 26338 63700 26350
rect 63756 26516 63812 26526
rect 63196 26292 63252 26302
rect 63196 26198 63252 26236
rect 63756 26290 63812 26460
rect 64428 26514 64484 26684
rect 64428 26462 64430 26514
rect 64482 26462 64484 26514
rect 64428 26450 64484 26462
rect 65436 26740 65492 26750
rect 65436 26514 65492 26684
rect 65436 26462 65438 26514
rect 65490 26462 65492 26514
rect 65436 26450 65492 26462
rect 67004 26516 67060 26798
rect 67004 26450 67060 26460
rect 67452 26740 67508 26852
rect 63756 26238 63758 26290
rect 63810 26238 63812 26290
rect 63756 26226 63812 26238
rect 67452 26290 67508 26684
rect 67564 26628 67620 26910
rect 67676 26962 67732 28364
rect 67676 26910 67678 26962
rect 67730 26910 67732 26962
rect 67676 26898 67732 26910
rect 67900 26964 67956 26974
rect 67900 26870 67956 26908
rect 67788 26852 67844 26862
rect 67788 26628 67844 26796
rect 67564 26562 67620 26572
rect 67676 26572 67844 26628
rect 67452 26238 67454 26290
rect 67506 26238 67508 26290
rect 67452 26226 67508 26238
rect 67676 26290 67732 26572
rect 67676 26238 67678 26290
rect 67730 26238 67732 26290
rect 67676 26226 67732 26238
rect 64988 26178 65044 26190
rect 64988 26126 64990 26178
rect 65042 26126 65044 26178
rect 64988 25508 65044 26126
rect 67788 26178 67844 26190
rect 67788 26126 67790 26178
rect 67842 26126 67844 26178
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 64764 25396 64820 25406
rect 64764 25394 64932 25396
rect 64764 25342 64766 25394
rect 64818 25342 64932 25394
rect 64764 25340 64932 25342
rect 64764 25330 64820 25340
rect 62860 24854 62916 24892
rect 64316 24948 64372 24958
rect 62412 24612 62468 24622
rect 62188 24610 62468 24612
rect 62188 24558 62414 24610
rect 62466 24558 62468 24610
rect 62188 24556 62468 24558
rect 62412 24498 62468 24556
rect 62412 24446 62414 24498
rect 62466 24446 62468 24498
rect 62412 24434 62468 24446
rect 62972 24498 63028 24510
rect 62972 24446 62974 24498
rect 63026 24446 63028 24498
rect 61404 23314 61460 23324
rect 60620 22430 60622 22482
rect 60674 22430 60676 22482
rect 60620 22418 60676 22430
rect 60844 22764 61236 22820
rect 60844 22370 60900 22764
rect 60844 22318 60846 22370
rect 60898 22318 60900 22370
rect 60844 22306 60900 22318
rect 60956 22370 61012 22382
rect 60956 22318 60958 22370
rect 61010 22318 61012 22370
rect 60956 22148 61012 22318
rect 60956 22082 61012 22092
rect 60844 21812 60900 21822
rect 60844 21718 60900 21756
rect 60508 21534 60510 21586
rect 60562 21534 60564 21586
rect 60508 21522 60564 21534
rect 60732 21586 60788 21598
rect 60732 21534 60734 21586
rect 60786 21534 60788 21586
rect 59836 21084 60228 21140
rect 59836 20914 59892 21084
rect 59836 20862 59838 20914
rect 59890 20862 59892 20914
rect 59836 20850 59892 20862
rect 59948 20916 60004 20926
rect 59948 20822 60004 20860
rect 60508 20916 60564 20926
rect 60508 20822 60564 20860
rect 59724 20738 59780 20748
rect 60620 20804 60676 20814
rect 60620 20710 60676 20748
rect 59444 20524 59668 20580
rect 59388 20514 59444 20524
rect 59724 20468 59780 20478
rect 59388 20244 59444 20254
rect 59724 20244 59780 20412
rect 59388 20242 59780 20244
rect 59388 20190 59390 20242
rect 59442 20190 59780 20242
rect 59388 20188 59780 20190
rect 59388 20178 59444 20188
rect 59724 20018 59780 20188
rect 60732 20244 60788 21534
rect 60956 21588 61012 21598
rect 60956 20804 61012 21532
rect 60956 20710 61012 20748
rect 60732 20178 60788 20188
rect 62524 20244 62580 20254
rect 59724 19966 59726 20018
rect 59778 19966 59780 20018
rect 59724 19954 59780 19966
rect 60060 20132 60116 20142
rect 59836 19906 59892 19918
rect 59836 19854 59838 19906
rect 59890 19854 59892 19906
rect 59836 19796 59892 19854
rect 59836 19730 59892 19740
rect 59276 19394 59332 19404
rect 59388 19572 59444 19582
rect 58828 17836 59332 17892
rect 58716 17724 59108 17780
rect 58380 17714 58436 17724
rect 58828 17554 58884 17566
rect 58828 17502 58830 17554
rect 58882 17502 58884 17554
rect 58716 17108 58772 17118
rect 58716 17014 58772 17052
rect 58828 16884 58884 17502
rect 58940 17556 58996 17566
rect 58940 17462 58996 17500
rect 59052 17444 59108 17724
rect 59164 17444 59220 17454
rect 59052 17442 59220 17444
rect 59052 17390 59166 17442
rect 59218 17390 59220 17442
rect 59052 17388 59220 17390
rect 58828 16818 58884 16828
rect 59164 16884 59220 17388
rect 59164 16818 59220 16828
rect 59276 16100 59332 17836
rect 59276 16034 59332 16044
rect 59388 15540 59444 19516
rect 60060 18674 60116 20076
rect 60172 20130 60228 20142
rect 60172 20078 60174 20130
rect 60226 20078 60228 20130
rect 60172 20020 60228 20078
rect 60956 20132 61012 20142
rect 60956 20038 61012 20076
rect 60172 19012 60228 19964
rect 61180 20018 61236 20030
rect 61180 19966 61182 20018
rect 61234 19966 61236 20018
rect 60172 18946 60228 18956
rect 60732 19234 60788 19246
rect 60732 19182 60734 19234
rect 60786 19182 60788 19234
rect 60732 19124 60788 19182
rect 60620 18788 60676 18798
rect 60060 18622 60062 18674
rect 60114 18622 60116 18674
rect 60060 18610 60116 18622
rect 60508 18732 60620 18788
rect 59724 18564 59780 18574
rect 59500 18452 59556 18462
rect 59500 18358 59556 18396
rect 59724 18228 59780 18508
rect 59724 18134 59780 18172
rect 59500 17556 59556 17566
rect 59500 17462 59556 17500
rect 59948 17442 60004 17454
rect 59948 17390 59950 17442
rect 60002 17390 60004 17442
rect 59948 17332 60004 17390
rect 59948 17266 60004 17276
rect 60396 17332 60452 17342
rect 60396 17106 60452 17276
rect 60396 17054 60398 17106
rect 60450 17054 60452 17106
rect 60396 17042 60452 17054
rect 60508 16660 60564 18732
rect 60620 18722 60676 18732
rect 60732 18450 60788 19068
rect 61180 19234 61236 19966
rect 61180 19182 61182 19234
rect 61234 19182 61236 19234
rect 61180 18564 61236 19182
rect 62412 19236 62468 19246
rect 62300 19124 62356 19134
rect 62300 19030 62356 19068
rect 61180 18498 61236 18508
rect 61292 19012 61348 19022
rect 60732 18398 60734 18450
rect 60786 18398 60788 18450
rect 60732 18340 60788 18398
rect 60732 18274 60788 18284
rect 61068 18452 61124 18462
rect 61292 18452 61348 18956
rect 62412 19010 62468 19180
rect 62412 18958 62414 19010
rect 62466 18958 62468 19010
rect 62412 18946 62468 18958
rect 61964 18562 62020 18574
rect 61964 18510 61966 18562
rect 62018 18510 62020 18562
rect 61628 18452 61684 18462
rect 61292 18450 61684 18452
rect 61292 18398 61630 18450
rect 61682 18398 61684 18450
rect 61292 18396 61684 18398
rect 61068 18338 61124 18396
rect 61628 18386 61684 18396
rect 61068 18286 61070 18338
rect 61122 18286 61124 18338
rect 60620 18228 60676 18238
rect 60620 17778 60676 18172
rect 61068 18116 61124 18286
rect 61068 18050 61124 18060
rect 61964 18340 62020 18510
rect 62524 18562 62580 20188
rect 62524 18510 62526 18562
rect 62578 18510 62580 18562
rect 62524 18498 62580 18510
rect 62636 18562 62692 18574
rect 62636 18510 62638 18562
rect 62690 18510 62692 18562
rect 60620 17726 60622 17778
rect 60674 17726 60676 17778
rect 60620 17714 60676 17726
rect 61964 17554 62020 18284
rect 61964 17502 61966 17554
rect 62018 17502 62020 17554
rect 61964 17490 62020 17502
rect 62076 18226 62132 18238
rect 62076 18174 62078 18226
rect 62130 18174 62132 18226
rect 61068 17442 61124 17454
rect 61068 17390 61070 17442
rect 61122 17390 61124 17442
rect 60732 16884 60788 16894
rect 60732 16790 60788 16828
rect 60956 16884 61012 16894
rect 60956 16790 61012 16828
rect 60508 16604 60788 16660
rect 60620 16212 60676 16222
rect 58156 14914 58212 14924
rect 58268 15202 58324 15214
rect 58268 15150 58270 15202
rect 58322 15150 58324 15202
rect 58268 15148 58324 15150
rect 58716 15202 58772 15214
rect 58716 15150 58718 15202
rect 58770 15150 58772 15202
rect 58716 15148 58772 15150
rect 58268 15092 58772 15148
rect 58268 14756 58324 15092
rect 57708 14702 57710 14754
rect 57762 14702 57764 14754
rect 57708 14690 57764 14702
rect 57820 14700 58324 14756
rect 57820 14642 57876 14700
rect 57820 14590 57822 14642
rect 57874 14590 57876 14642
rect 57820 14578 57876 14590
rect 58380 14642 58436 14654
rect 58380 14590 58382 14642
rect 58434 14590 58436 14642
rect 58380 14532 58436 14590
rect 58156 14530 58436 14532
rect 58156 14478 58382 14530
rect 58434 14478 58436 14530
rect 58156 14476 58436 14478
rect 57036 14306 57092 14318
rect 57036 14254 57038 14306
rect 57090 14254 57092 14306
rect 55132 13654 55188 13692
rect 56588 13746 56644 13758
rect 56588 13694 56590 13746
rect 56642 13694 56644 13746
rect 55244 13636 55300 13646
rect 55020 12852 55076 12862
rect 54908 12850 55076 12852
rect 54908 12798 55022 12850
rect 55074 12798 55076 12850
rect 54908 12796 55076 12798
rect 54908 12402 54964 12796
rect 55020 12786 55076 12796
rect 54908 12350 54910 12402
rect 54962 12350 54964 12402
rect 54908 12338 54964 12350
rect 55132 12292 55188 12302
rect 54908 12180 54964 12190
rect 54908 12086 54964 12124
rect 54796 10782 54798 10834
rect 54850 10782 54852 10834
rect 54796 10500 54852 10782
rect 54796 10434 54852 10444
rect 55132 10276 55188 12236
rect 55244 12290 55300 13580
rect 55244 12238 55246 12290
rect 55298 12238 55300 12290
rect 55244 12226 55300 12238
rect 55916 13634 55972 13646
rect 55916 13582 55918 13634
rect 55970 13582 55972 13634
rect 55916 12964 55972 13582
rect 55916 12180 55972 12908
rect 56028 12404 56084 12414
rect 56028 12310 56084 12348
rect 55916 12114 55972 12124
rect 55580 11284 55636 11294
rect 55468 10836 55524 10846
rect 55468 10742 55524 10780
rect 55580 10834 55636 11228
rect 55580 10782 55582 10834
rect 55634 10782 55636 10834
rect 55580 10770 55636 10782
rect 55916 10948 55972 10958
rect 55132 10210 55188 10220
rect 55692 10610 55748 10622
rect 55692 10558 55694 10610
rect 55746 10558 55748 10610
rect 53900 10164 53956 10174
rect 53676 6638 53678 6690
rect 53730 6638 53732 6690
rect 53676 6626 53732 6638
rect 53788 10108 53900 10164
rect 53340 6468 53396 6478
rect 53396 6412 53508 6468
rect 53340 6402 53396 6412
rect 53004 5966 53006 6018
rect 53058 5966 53060 6018
rect 52668 5814 52724 5852
rect 52780 5460 52836 5470
rect 52780 5346 52836 5404
rect 52780 5294 52782 5346
rect 52834 5294 52836 5346
rect 52780 5282 52836 5294
rect 52668 5124 52724 5134
rect 52332 5122 52724 5124
rect 52332 5070 52670 5122
rect 52722 5070 52724 5122
rect 52332 5068 52724 5070
rect 52668 5058 52724 5068
rect 52780 5012 52836 5022
rect 52780 4918 52836 4956
rect 53004 4900 53060 5966
rect 53004 4834 53060 4844
rect 53116 6018 53172 6030
rect 53116 5966 53118 6018
rect 53170 5966 53172 6018
rect 53116 3444 53172 5966
rect 53340 6020 53396 6030
rect 53340 5926 53396 5964
rect 53340 5348 53396 5358
rect 53340 5122 53396 5292
rect 53340 5070 53342 5122
rect 53394 5070 53396 5122
rect 53340 5058 53396 5070
rect 53452 5122 53508 6412
rect 53452 5070 53454 5122
rect 53506 5070 53508 5122
rect 53452 5058 53508 5070
rect 53564 5794 53620 5806
rect 53564 5742 53566 5794
rect 53618 5742 53620 5794
rect 53564 4564 53620 5742
rect 53676 5124 53732 5134
rect 53676 5030 53732 5068
rect 53788 5122 53844 10108
rect 53900 10098 53956 10108
rect 55020 10052 55076 10062
rect 54348 9156 54404 9166
rect 54348 9062 54404 9100
rect 55020 8370 55076 9996
rect 55692 9938 55748 10558
rect 55692 9886 55694 9938
rect 55746 9886 55748 9938
rect 55692 9828 55748 9886
rect 55692 9762 55748 9772
rect 55804 9940 55860 9950
rect 55244 9716 55300 9726
rect 55244 9042 55300 9660
rect 55804 9268 55860 9884
rect 55916 9380 55972 10892
rect 56588 10836 56644 13694
rect 56812 13748 56868 13758
rect 56812 13654 56868 13692
rect 56700 13636 56756 13646
rect 56700 13542 56756 13580
rect 56812 12852 56868 12862
rect 56700 10836 56756 10846
rect 56644 10834 56756 10836
rect 56644 10782 56702 10834
rect 56754 10782 56756 10834
rect 56644 10780 56756 10782
rect 56588 10742 56644 10780
rect 56700 10770 56756 10780
rect 56812 10834 56868 12796
rect 57036 12740 57092 14254
rect 57484 14306 57540 14318
rect 57484 14254 57486 14306
rect 57538 14254 57540 14306
rect 57484 13972 57540 14254
rect 57484 13916 57876 13972
rect 57036 12404 57092 12684
rect 57036 12338 57092 12348
rect 57148 13746 57204 13758
rect 57148 13694 57150 13746
rect 57202 13694 57204 13746
rect 57148 13636 57204 13694
rect 56924 12180 56980 12190
rect 56924 12086 56980 12124
rect 57036 12068 57092 12078
rect 56812 10782 56814 10834
rect 56866 10782 56868 10834
rect 56812 10770 56868 10782
rect 56924 10836 56980 10846
rect 57036 10836 57092 12012
rect 57148 11060 57204 13580
rect 57596 13748 57652 13758
rect 57596 13634 57652 13692
rect 57596 13582 57598 13634
rect 57650 13582 57652 13634
rect 57260 12740 57316 12750
rect 57596 12740 57652 13582
rect 57708 12852 57764 12862
rect 57708 12758 57764 12796
rect 57260 12738 57652 12740
rect 57260 12686 57262 12738
rect 57314 12686 57652 12738
rect 57260 12684 57652 12686
rect 57260 12404 57316 12684
rect 57820 12628 57876 13916
rect 58044 13636 58100 13646
rect 58044 13542 58100 13580
rect 57932 12850 57988 12862
rect 57932 12798 57934 12850
rect 57986 12798 57988 12850
rect 57932 12628 57988 12798
rect 57260 12338 57316 12348
rect 57484 12572 57988 12628
rect 58044 12738 58100 12750
rect 58044 12686 58046 12738
rect 58098 12686 58100 12738
rect 57484 11396 57540 12572
rect 58044 12404 58100 12686
rect 57596 12348 58100 12404
rect 57596 12290 57652 12348
rect 57596 12238 57598 12290
rect 57650 12238 57652 12290
rect 57596 12226 57652 12238
rect 57484 11330 57540 11340
rect 58044 11956 58100 11966
rect 57148 10994 57204 11004
rect 56924 10834 57092 10836
rect 56924 10782 56926 10834
rect 56978 10782 57092 10834
rect 56924 10780 57092 10782
rect 57148 10780 57428 10836
rect 56924 10724 56980 10780
rect 56924 10658 56980 10668
rect 56140 10612 56196 10622
rect 56140 10518 56196 10556
rect 56700 10052 56756 10062
rect 56700 9938 56756 9996
rect 56700 9886 56702 9938
rect 56754 9886 56756 9938
rect 56700 9874 56756 9886
rect 56812 9826 56868 9838
rect 57036 9828 57092 9838
rect 56812 9774 56814 9826
rect 56866 9774 56868 9826
rect 56028 9716 56084 9726
rect 56028 9622 56084 9660
rect 56364 9716 56420 9726
rect 56588 9716 56644 9726
rect 56364 9714 56644 9716
rect 56364 9662 56366 9714
rect 56418 9662 56590 9714
rect 56642 9662 56644 9714
rect 56364 9660 56644 9662
rect 56364 9650 56420 9660
rect 56588 9650 56644 9660
rect 56140 9604 56196 9614
rect 56140 9510 56196 9548
rect 56812 9604 56868 9774
rect 56812 9538 56868 9548
rect 56924 9826 57092 9828
rect 56924 9774 57038 9826
rect 57090 9774 57092 9826
rect 56924 9772 57092 9774
rect 55916 9324 56084 9380
rect 55468 9212 55860 9268
rect 55244 8990 55246 9042
rect 55298 8990 55300 9042
rect 55244 8484 55300 8990
rect 55356 9154 55412 9166
rect 55356 9102 55358 9154
rect 55410 9102 55412 9154
rect 55356 8932 55412 9102
rect 55356 8866 55412 8876
rect 55244 8418 55300 8428
rect 55020 8318 55022 8370
rect 55074 8318 55076 8370
rect 55020 8306 55076 8318
rect 54348 8258 54404 8270
rect 54348 8206 54350 8258
rect 54402 8206 54404 8258
rect 53900 8034 53956 8046
rect 53900 7982 53902 8034
rect 53954 7982 53956 8034
rect 53900 7588 53956 7982
rect 53900 7522 53956 7532
rect 54012 7476 54068 7486
rect 54012 7382 54068 7420
rect 54236 7364 54292 7374
rect 54124 7362 54292 7364
rect 54124 7310 54238 7362
rect 54290 7310 54292 7362
rect 54124 7308 54292 7310
rect 54124 6580 54180 7308
rect 54236 7298 54292 7308
rect 54348 6692 54404 8206
rect 54684 8148 54740 8158
rect 54460 8036 54516 8046
rect 54460 7586 54516 7980
rect 54460 7534 54462 7586
rect 54514 7534 54516 7586
rect 54460 7522 54516 7534
rect 54684 7474 54740 8092
rect 54684 7422 54686 7474
rect 54738 7422 54740 7474
rect 54684 7364 54740 7422
rect 54684 7298 54740 7308
rect 55132 7474 55188 7486
rect 55132 7422 55134 7474
rect 55186 7422 55188 7474
rect 54124 6514 54180 6524
rect 54236 6636 54348 6692
rect 53788 5070 53790 5122
rect 53842 5070 53844 5122
rect 53788 5058 53844 5070
rect 54236 5908 54292 6636
rect 54348 6626 54404 6636
rect 54236 5122 54292 5852
rect 54236 5070 54238 5122
rect 54290 5070 54292 5122
rect 54236 5058 54292 5070
rect 54684 6356 54740 6366
rect 53564 4508 53956 4564
rect 53452 4452 53508 4462
rect 53452 4450 53844 4452
rect 53452 4398 53454 4450
rect 53506 4398 53844 4450
rect 53452 4396 53844 4398
rect 53452 4386 53508 4396
rect 53116 3378 53172 3388
rect 53564 3442 53620 3454
rect 53564 3390 53566 3442
rect 53618 3390 53620 3442
rect 53564 800 53620 3390
rect 53788 3220 53844 4396
rect 53900 4450 53956 4508
rect 53900 4398 53902 4450
rect 53954 4398 53956 4450
rect 53900 4386 53956 4398
rect 54684 3388 54740 6300
rect 54908 5124 54964 5134
rect 54908 5030 54964 5068
rect 55020 5012 55076 5022
rect 55020 3666 55076 4956
rect 55132 4226 55188 7422
rect 55468 7140 55524 9212
rect 55804 9154 55860 9212
rect 55804 9102 55806 9154
rect 55858 9102 55860 9154
rect 55804 9090 55860 9102
rect 55916 9156 55972 9166
rect 55916 9062 55972 9100
rect 55580 9044 55636 9054
rect 55580 9042 55748 9044
rect 55580 8990 55582 9042
rect 55634 8990 55748 9042
rect 55580 8988 55748 8990
rect 55580 8978 55636 8988
rect 55692 8596 55748 8988
rect 55692 8530 55748 8540
rect 55580 8484 55636 8494
rect 55580 7252 55636 8428
rect 56028 8484 56084 9324
rect 56924 9154 56980 9772
rect 57036 9762 57092 9772
rect 57148 9380 57204 10780
rect 57372 10724 57428 10780
rect 58044 10834 58100 11900
rect 58044 10782 58046 10834
rect 58098 10782 58100 10834
rect 58044 10770 58100 10782
rect 58156 10834 58212 14476
rect 58380 14466 58436 14476
rect 58380 12962 58436 12974
rect 58380 12910 58382 12962
rect 58434 12910 58436 12962
rect 58380 12516 58436 12910
rect 58380 12450 58436 12460
rect 58156 10782 58158 10834
rect 58210 10782 58212 10834
rect 57596 10724 57652 10734
rect 57372 10722 57652 10724
rect 57372 10670 57598 10722
rect 57650 10670 57652 10722
rect 57372 10668 57652 10670
rect 57596 10658 57652 10668
rect 57260 10612 57316 10622
rect 57260 10518 57316 10556
rect 57820 10610 57876 10622
rect 57820 10558 57822 10610
rect 57874 10558 57876 10610
rect 57708 10388 57764 10398
rect 57708 9940 57764 10332
rect 57820 10052 57876 10558
rect 57932 10500 57988 10510
rect 57932 10406 57988 10444
rect 57932 10052 57988 10062
rect 58156 10052 58212 10782
rect 57820 9996 57932 10052
rect 57708 9884 57876 9940
rect 57708 9716 57764 9726
rect 56924 9102 56926 9154
rect 56978 9102 56980 9154
rect 56140 9044 56196 9054
rect 56140 8950 56196 8988
rect 56588 9042 56644 9054
rect 56588 8990 56590 9042
rect 56642 8990 56644 9042
rect 56588 8820 56644 8990
rect 56588 8754 56644 8764
rect 56812 8596 56868 8606
rect 56028 8418 56084 8428
rect 56700 8484 56756 8494
rect 56028 7700 56084 7710
rect 55916 7644 56028 7700
rect 55692 7476 55748 7486
rect 55692 7382 55748 7420
rect 55580 7196 55748 7252
rect 55468 7074 55524 7084
rect 55580 6356 55636 6366
rect 55580 6018 55636 6300
rect 55580 5966 55582 6018
rect 55634 5966 55636 6018
rect 55580 5954 55636 5966
rect 55692 4340 55748 7196
rect 55692 4274 55748 4284
rect 55804 6580 55860 6590
rect 55804 4338 55860 6524
rect 55804 4286 55806 4338
rect 55858 4286 55860 4338
rect 55804 4274 55860 4286
rect 55132 4174 55134 4226
rect 55186 4174 55188 4226
rect 55132 4162 55188 4174
rect 55020 3614 55022 3666
rect 55074 3614 55076 3666
rect 55020 3602 55076 3614
rect 55916 3388 55972 7644
rect 56028 7634 56084 7644
rect 56476 7700 56532 7710
rect 56140 7364 56196 7374
rect 56028 6468 56084 6478
rect 56028 4562 56084 6412
rect 56028 4510 56030 4562
rect 56082 4510 56084 4562
rect 56028 4498 56084 4510
rect 54684 3332 54964 3388
rect 55916 3332 56084 3388
rect 53788 3154 53844 3164
rect 54908 800 54964 3332
rect 56028 980 56084 3332
rect 56140 1316 56196 7308
rect 56476 5572 56532 7644
rect 56700 7698 56756 8428
rect 56812 8260 56868 8540
rect 56924 8484 56980 9102
rect 56924 8418 56980 8428
rect 57036 9324 57204 9380
rect 57260 9714 57764 9716
rect 57260 9662 57710 9714
rect 57762 9662 57764 9714
rect 57260 9660 57764 9662
rect 56812 8204 56980 8260
rect 56700 7646 56702 7698
rect 56754 7646 56756 7698
rect 56700 7634 56756 7646
rect 56588 7588 56644 7598
rect 56588 7494 56644 7532
rect 56924 7474 56980 8204
rect 56924 7422 56926 7474
rect 56978 7422 56980 7474
rect 56924 7410 56980 7422
rect 57036 7924 57092 9324
rect 57148 9156 57204 9166
rect 57148 8370 57204 9100
rect 57148 8318 57150 8370
rect 57202 8318 57204 8370
rect 57148 8306 57204 8318
rect 57260 7924 57316 9660
rect 57708 9650 57764 9660
rect 57820 9268 57876 9884
rect 57932 9826 57988 9996
rect 57932 9774 57934 9826
rect 57986 9774 57988 9826
rect 57932 9762 57988 9774
rect 58044 9996 58212 10052
rect 58268 11284 58324 11294
rect 58044 9604 58100 9996
rect 58268 9938 58324 11228
rect 58492 10836 58548 15092
rect 58716 15026 58772 15036
rect 59388 14642 59444 15484
rect 60508 15764 60564 15774
rect 60508 15538 60564 15708
rect 60508 15486 60510 15538
rect 60562 15486 60564 15538
rect 60508 15474 60564 15486
rect 59500 15202 59556 15214
rect 59500 15150 59502 15202
rect 59554 15150 59556 15202
rect 59500 15148 59556 15150
rect 60284 15202 60340 15214
rect 60284 15150 60286 15202
rect 60338 15150 60340 15202
rect 59500 15092 59780 15148
rect 59388 14590 59390 14642
rect 59442 14590 59444 14642
rect 59388 14578 59444 14590
rect 59388 13746 59444 13758
rect 59388 13694 59390 13746
rect 59442 13694 59444 13746
rect 58604 13634 58660 13646
rect 58940 13636 58996 13646
rect 59388 13636 59444 13694
rect 58604 13582 58606 13634
rect 58658 13582 58660 13634
rect 58604 13524 58660 13582
rect 58604 13458 58660 13468
rect 58828 13634 59444 13636
rect 58828 13582 58942 13634
rect 58994 13582 59444 13634
rect 58828 13580 59444 13582
rect 58716 13076 58772 13086
rect 58828 13076 58884 13580
rect 58940 13570 58996 13580
rect 58716 13074 58884 13076
rect 58716 13022 58718 13074
rect 58770 13022 58884 13074
rect 58716 13020 58884 13022
rect 59276 13412 59332 13422
rect 58716 12180 58772 13020
rect 58716 11508 58772 12124
rect 58716 11414 58772 11452
rect 58828 12740 58884 12750
rect 58268 9886 58270 9938
rect 58322 9886 58324 9938
rect 58268 9874 58324 9886
rect 58380 10780 58548 10836
rect 58828 11060 58884 12684
rect 58156 9828 58212 9838
rect 58156 9734 58212 9772
rect 58268 9604 58324 9614
rect 58044 9548 58268 9604
rect 58268 9510 58324 9548
rect 56812 7140 56868 7150
rect 56700 7028 56756 7038
rect 56476 5506 56532 5516
rect 56588 6972 56700 7028
rect 56588 5236 56644 6972
rect 56700 6962 56756 6972
rect 56812 6244 56868 7084
rect 57036 7028 57092 7868
rect 57036 6962 57092 6972
rect 57148 7868 57316 7924
rect 57372 9212 57876 9268
rect 56700 6188 56868 6244
rect 56700 5796 56756 6188
rect 56812 6020 56868 6030
rect 56812 5926 56868 5964
rect 57036 5906 57092 5918
rect 57036 5854 57038 5906
rect 57090 5854 57092 5906
rect 56700 5740 56868 5796
rect 56588 5170 56644 5180
rect 56588 4900 56644 4910
rect 56588 4450 56644 4844
rect 56588 4398 56590 4450
rect 56642 4398 56644 4450
rect 56588 4386 56644 4398
rect 56700 4452 56756 4462
rect 56812 4452 56868 5740
rect 56924 5794 56980 5806
rect 56924 5742 56926 5794
rect 56978 5742 56980 5794
rect 56924 4676 56980 5742
rect 57036 5460 57092 5854
rect 57036 5394 57092 5404
rect 57036 5236 57092 5246
rect 57036 5142 57092 5180
rect 57148 5012 57204 7868
rect 57260 7700 57316 7710
rect 57260 7606 57316 7644
rect 57372 7586 57428 9212
rect 58268 9156 58324 9166
rect 57708 9154 58324 9156
rect 57708 9102 58270 9154
rect 58322 9102 58324 9154
rect 57708 9100 58324 9102
rect 57372 7534 57374 7586
rect 57426 7534 57428 7586
rect 57372 7522 57428 7534
rect 57484 8930 57540 8942
rect 57484 8878 57486 8930
rect 57538 8878 57540 8930
rect 57484 6580 57540 8878
rect 57484 6514 57540 6524
rect 57596 8484 57652 8494
rect 57596 7474 57652 8428
rect 57708 8370 57764 9100
rect 58268 9090 58324 9100
rect 57708 8318 57710 8370
rect 57762 8318 57764 8370
rect 57708 8306 57764 8318
rect 57596 7422 57598 7474
rect 57650 7422 57652 7474
rect 57260 5908 57316 5918
rect 57596 5908 57652 7422
rect 58044 7476 58100 7486
rect 58380 7476 58436 10780
rect 58716 10724 58772 10734
rect 58044 7474 58436 7476
rect 58044 7422 58046 7474
rect 58098 7422 58436 7474
rect 58044 7420 58436 7422
rect 58044 7410 58100 7420
rect 57708 6804 57764 6814
rect 58380 6804 58436 7420
rect 57764 6748 57876 6804
rect 57708 6710 57764 6748
rect 57260 5906 57652 5908
rect 57260 5854 57262 5906
rect 57314 5854 57652 5906
rect 57260 5852 57652 5854
rect 57260 5348 57316 5852
rect 57708 5796 57764 5806
rect 57708 5702 57764 5740
rect 57260 5282 57316 5292
rect 57148 4946 57204 4956
rect 57372 4898 57428 4910
rect 57372 4846 57374 4898
rect 57426 4846 57428 4898
rect 56924 4620 57204 4676
rect 56924 4452 56980 4462
rect 56812 4450 56980 4452
rect 56812 4398 56926 4450
rect 56978 4398 56980 4450
rect 56812 4396 56980 4398
rect 56700 4358 56756 4396
rect 56924 4386 56980 4396
rect 57148 3666 57204 4620
rect 57372 4450 57428 4846
rect 57372 4398 57374 4450
rect 57426 4398 57428 4450
rect 57372 4386 57428 4398
rect 57148 3614 57150 3666
rect 57202 3614 57204 3666
rect 57148 3602 57204 3614
rect 57596 3668 57652 3678
rect 56140 1250 56196 1260
rect 56028 924 56308 980
rect 56252 800 56308 924
rect 57596 800 57652 3612
rect 57820 3554 57876 6748
rect 58380 6738 58436 6748
rect 58492 10722 58772 10724
rect 58492 10670 58718 10722
rect 58770 10670 58772 10722
rect 58492 10668 58772 10670
rect 58492 6468 58548 10668
rect 58716 10658 58772 10668
rect 58828 10722 58884 11004
rect 59276 10836 59332 13356
rect 59388 13076 59444 13580
rect 59500 13076 59556 13086
rect 59388 13020 59500 13076
rect 59500 12982 59556 13020
rect 59276 10742 59332 10780
rect 58828 10670 58830 10722
rect 58882 10670 58884 10722
rect 58828 10658 58884 10670
rect 59388 10610 59444 10622
rect 59388 10558 59390 10610
rect 59442 10558 59444 10610
rect 59052 10500 59108 10510
rect 58716 10386 58772 10398
rect 58716 10334 58718 10386
rect 58770 10334 58772 10386
rect 58716 10164 58772 10334
rect 58716 10098 58772 10108
rect 59052 9938 59108 10444
rect 59276 10388 59332 10398
rect 59276 10294 59332 10332
rect 59052 9886 59054 9938
rect 59106 9886 59108 9938
rect 59052 9874 59108 9886
rect 59388 9940 59444 10558
rect 59388 9874 59444 9884
rect 59724 9828 59780 15092
rect 60060 13634 60116 13646
rect 60060 13582 60062 13634
rect 60114 13582 60116 13634
rect 59948 13300 60004 13310
rect 59836 12964 59892 12974
rect 59836 12402 59892 12908
rect 59836 12350 59838 12402
rect 59890 12350 59892 12402
rect 59836 12068 59892 12350
rect 59836 12002 59892 12012
rect 59948 12740 60004 13244
rect 60060 13188 60116 13582
rect 60060 13122 60116 13132
rect 60060 12740 60116 12750
rect 59948 12738 60116 12740
rect 59948 12686 60062 12738
rect 60114 12686 60116 12738
rect 59948 12684 60116 12686
rect 59836 11620 59892 11630
rect 59836 10050 59892 11564
rect 59948 11172 60004 12684
rect 60060 12674 60116 12684
rect 59948 11106 60004 11116
rect 60060 11508 60116 11518
rect 60060 10610 60116 11452
rect 60060 10558 60062 10610
rect 60114 10558 60116 10610
rect 60060 10546 60116 10558
rect 59836 9998 59838 10050
rect 59890 9998 59892 10050
rect 59836 9986 59892 9998
rect 59948 9828 60004 9838
rect 59724 9772 59892 9828
rect 59388 9714 59444 9726
rect 59388 9662 59390 9714
rect 59442 9662 59444 9714
rect 59052 9604 59108 9614
rect 59052 9042 59108 9548
rect 59164 9156 59220 9166
rect 59164 9062 59220 9100
rect 59052 8990 59054 9042
rect 59106 8990 59108 9042
rect 59052 8978 59108 8990
rect 59276 8930 59332 8942
rect 59276 8878 59278 8930
rect 59330 8878 59332 8930
rect 58716 7700 58772 7710
rect 58716 7586 58772 7644
rect 58716 7534 58718 7586
rect 58770 7534 58772 7586
rect 58716 7522 58772 7534
rect 58492 6402 58548 6412
rect 58604 6578 58660 6590
rect 58604 6526 58606 6578
rect 58658 6526 58660 6578
rect 58268 5906 58324 5918
rect 58268 5854 58270 5906
rect 58322 5854 58324 5906
rect 58268 4228 58324 5854
rect 58604 5794 58660 6526
rect 58604 5742 58606 5794
rect 58658 5742 58660 5794
rect 58604 5730 58660 5742
rect 58940 5012 58996 5022
rect 58380 4228 58436 4238
rect 58268 4226 58436 4228
rect 58268 4174 58382 4226
rect 58434 4174 58436 4226
rect 58268 4172 58436 4174
rect 58380 4162 58436 4172
rect 58940 4226 58996 4956
rect 58940 4174 58942 4226
rect 58994 4174 58996 4226
rect 58940 4162 58996 4174
rect 59052 3668 59108 3678
rect 59052 3574 59108 3612
rect 57820 3502 57822 3554
rect 57874 3502 57876 3554
rect 57820 3490 57876 3502
rect 59276 1204 59332 8878
rect 59388 1652 59444 9662
rect 59836 9714 59892 9772
rect 59948 9734 60004 9772
rect 59836 9662 59838 9714
rect 59890 9662 59892 9714
rect 59724 9604 59780 9614
rect 59500 8148 59556 8158
rect 59500 8054 59556 8092
rect 59724 5010 59780 9548
rect 59836 9492 59892 9662
rect 59836 7700 59892 9436
rect 59836 7634 59892 7644
rect 60284 7588 60340 15150
rect 60620 14756 60676 16156
rect 60620 14690 60676 14700
rect 60732 14532 60788 16604
rect 61068 16324 61124 17390
rect 61964 17220 62020 17230
rect 61068 16210 61124 16268
rect 61068 16158 61070 16210
rect 61122 16158 61124 16210
rect 61068 16146 61124 16158
rect 61404 16884 61460 16894
rect 61404 16098 61460 16828
rect 61516 16772 61572 16782
rect 61516 16770 61796 16772
rect 61516 16718 61518 16770
rect 61570 16718 61796 16770
rect 61516 16716 61796 16718
rect 61516 16706 61572 16716
rect 61404 16046 61406 16098
rect 61458 16046 61460 16098
rect 61404 16034 61460 16046
rect 61516 15874 61572 15886
rect 61516 15822 61518 15874
rect 61570 15822 61572 15874
rect 61404 15764 61460 15774
rect 61516 15764 61572 15822
rect 61460 15708 61572 15764
rect 61404 15698 61460 15708
rect 61404 15316 61460 15326
rect 61628 15316 61684 15326
rect 60732 14466 60788 14476
rect 61068 15314 61460 15316
rect 61068 15262 61406 15314
rect 61458 15262 61460 15314
rect 61068 15260 61460 15262
rect 61068 15202 61124 15260
rect 61404 15250 61460 15260
rect 61516 15260 61628 15316
rect 61068 15150 61070 15202
rect 61122 15150 61124 15202
rect 60732 14308 60788 14318
rect 60732 14306 61012 14308
rect 60732 14254 60734 14306
rect 60786 14254 61012 14306
rect 60732 14252 61012 14254
rect 60732 14242 60788 14252
rect 60508 13524 60564 13534
rect 60508 12962 60564 13468
rect 60732 13300 60788 13310
rect 60620 13188 60676 13198
rect 60620 13074 60676 13132
rect 60620 13022 60622 13074
rect 60674 13022 60676 13074
rect 60620 13010 60676 13022
rect 60732 13076 60788 13244
rect 60956 13300 61012 14252
rect 61068 14306 61124 15150
rect 61404 14532 61460 14542
rect 61516 14532 61572 15260
rect 61628 15250 61684 15260
rect 61740 15148 61796 16716
rect 61964 16098 62020 17164
rect 62076 16884 62132 18174
rect 62076 16770 62132 16828
rect 62188 17666 62244 17678
rect 62188 17614 62190 17666
rect 62242 17614 62244 17666
rect 62188 17332 62244 17614
rect 62188 16882 62244 17276
rect 62412 16884 62468 16894
rect 62636 16884 62692 18510
rect 62860 18450 62916 18462
rect 62860 18398 62862 18450
rect 62914 18398 62916 18450
rect 62860 17780 62916 18398
rect 62860 17714 62916 17724
rect 62188 16830 62190 16882
rect 62242 16830 62244 16882
rect 62188 16818 62244 16830
rect 62300 16828 62412 16884
rect 62468 16828 62692 16884
rect 62748 17220 62804 17230
rect 62076 16718 62078 16770
rect 62130 16718 62132 16770
rect 62076 16706 62132 16718
rect 62076 16324 62132 16334
rect 62076 16230 62132 16268
rect 62300 16100 62356 16828
rect 62412 16790 62468 16828
rect 61964 16046 61966 16098
rect 62018 16046 62020 16098
rect 61964 16034 62020 16046
rect 62076 16044 62356 16100
rect 62076 15986 62132 16044
rect 62076 15934 62078 15986
rect 62130 15934 62132 15986
rect 62076 15922 62132 15934
rect 62636 15874 62692 15886
rect 62636 15822 62638 15874
rect 62690 15822 62692 15874
rect 62188 15428 62244 15438
rect 62188 15202 62244 15372
rect 62188 15150 62190 15202
rect 62242 15150 62244 15202
rect 61740 15092 61908 15148
rect 62188 15138 62244 15150
rect 61460 14476 61572 14532
rect 61628 14532 61684 14542
rect 61404 14438 61460 14476
rect 61628 14438 61684 14476
rect 61068 14254 61070 14306
rect 61122 14254 61124 14306
rect 61068 14084 61124 14254
rect 61068 14018 61124 14028
rect 61516 14306 61572 14318
rect 61516 14254 61518 14306
rect 61570 14254 61572 14306
rect 60956 13234 61012 13244
rect 61068 13412 61124 13422
rect 60732 13020 60900 13076
rect 60508 12910 60510 12962
rect 60562 12910 60564 12962
rect 60508 12898 60564 12910
rect 60844 12962 60900 13020
rect 60844 12910 60846 12962
rect 60898 12910 60900 12962
rect 60844 12898 60900 12910
rect 61068 12962 61124 13356
rect 61516 13412 61572 14254
rect 61516 13346 61572 13356
rect 61628 13524 61684 13534
rect 61068 12910 61070 12962
rect 61122 12910 61124 12962
rect 61068 12898 61124 12910
rect 61404 13300 61460 13310
rect 60620 12852 60676 12862
rect 60508 12516 60564 12526
rect 60508 12402 60564 12460
rect 60508 12350 60510 12402
rect 60562 12350 60564 12402
rect 60508 12338 60564 12350
rect 60620 11618 60676 12796
rect 60844 12516 60900 12526
rect 60844 12402 60900 12460
rect 60844 12350 60846 12402
rect 60898 12350 60900 12402
rect 60844 12338 60900 12350
rect 61292 12292 61348 12302
rect 61292 12198 61348 12236
rect 60620 11566 60622 11618
rect 60674 11566 60676 11618
rect 60620 11554 60676 11566
rect 61180 11954 61236 11966
rect 61180 11902 61182 11954
rect 61234 11902 61236 11954
rect 60732 11508 60788 11518
rect 60508 11284 60564 11294
rect 60508 11190 60564 11228
rect 60396 10052 60452 10062
rect 60396 9266 60452 9996
rect 60396 9214 60398 9266
rect 60450 9214 60452 9266
rect 60396 9202 60452 9214
rect 60732 9714 60788 11452
rect 60844 10836 60900 10846
rect 60900 10780 61012 10836
rect 60844 10770 60900 10780
rect 60844 10498 60900 10510
rect 60844 10446 60846 10498
rect 60898 10446 60900 10498
rect 60844 9938 60900 10446
rect 60844 9886 60846 9938
rect 60898 9886 60900 9938
rect 60844 9874 60900 9886
rect 60732 9662 60734 9714
rect 60786 9662 60788 9714
rect 60732 9156 60788 9662
rect 60844 9716 60900 9726
rect 60844 9266 60900 9660
rect 60844 9214 60846 9266
rect 60898 9214 60900 9266
rect 60844 9202 60900 9214
rect 60732 9090 60788 9100
rect 60284 7522 60340 7532
rect 60396 9042 60452 9054
rect 60396 8990 60398 9042
rect 60450 8990 60452 9042
rect 59948 6802 60004 6814
rect 59948 6750 59950 6802
rect 60002 6750 60004 6802
rect 59948 5124 60004 6750
rect 59948 5058 60004 5068
rect 60284 6020 60340 6030
rect 59724 4958 59726 5010
rect 59778 4958 59780 5010
rect 59724 3388 59780 4958
rect 59388 1586 59444 1596
rect 59500 3332 59780 3388
rect 59276 1138 59332 1148
rect 58940 924 59332 980
rect 58940 800 58996 924
rect 44380 700 44996 756
rect 45472 0 45584 800
rect 46816 0 46928 800
rect 48160 0 48272 800
rect 49504 0 49616 800
rect 50848 0 50960 800
rect 52192 0 52304 800
rect 53536 0 53648 800
rect 54880 0 54992 800
rect 56224 0 56336 800
rect 57568 0 57680 800
rect 58912 0 59024 800
rect 59276 756 59332 924
rect 59500 756 59556 3332
rect 60284 800 60340 5964
rect 60396 5012 60452 8990
rect 60620 8428 60900 8484
rect 60620 8370 60676 8428
rect 60620 8318 60622 8370
rect 60674 8318 60676 8370
rect 60620 8306 60676 8318
rect 60732 8258 60788 8270
rect 60732 8206 60734 8258
rect 60786 8206 60788 8258
rect 60508 8146 60564 8158
rect 60508 8094 60510 8146
rect 60562 8094 60564 8146
rect 60508 7140 60564 8094
rect 60508 7074 60564 7084
rect 60732 6916 60788 8206
rect 60844 7588 60900 8428
rect 60956 7700 61012 10780
rect 61068 9716 61124 9726
rect 61068 9622 61124 9660
rect 61180 9604 61236 11902
rect 61404 11394 61460 13244
rect 61628 12850 61684 13468
rect 61740 13188 61796 13198
rect 61740 13094 61796 13132
rect 61628 12798 61630 12850
rect 61682 12798 61684 12850
rect 61404 11342 61406 11394
rect 61458 11342 61460 11394
rect 61292 10388 61348 10398
rect 61404 10388 61460 11342
rect 61516 12516 61572 12526
rect 61516 11284 61572 12460
rect 61628 11508 61684 12798
rect 61740 12738 61796 12750
rect 61740 12686 61742 12738
rect 61794 12686 61796 12738
rect 61740 12292 61796 12686
rect 61740 12226 61796 12236
rect 61740 12066 61796 12078
rect 61740 12014 61742 12066
rect 61794 12014 61796 12066
rect 61740 11954 61796 12014
rect 61740 11902 61742 11954
rect 61794 11902 61796 11954
rect 61740 11890 61796 11902
rect 61628 11442 61684 11452
rect 61852 11396 61908 15092
rect 62076 14980 62132 14990
rect 62076 14530 62132 14924
rect 62524 14754 62580 14766
rect 62524 14702 62526 14754
rect 62578 14702 62580 14754
rect 62524 14642 62580 14702
rect 62524 14590 62526 14642
rect 62578 14590 62580 14642
rect 62076 14478 62078 14530
rect 62130 14478 62132 14530
rect 62076 14466 62132 14478
rect 62188 14532 62244 14542
rect 62076 14084 62132 14094
rect 61964 13972 62020 13982
rect 61964 11508 62020 13916
rect 61964 11442 62020 11452
rect 61852 11330 61908 11340
rect 62076 11396 62132 14028
rect 62188 13634 62244 14476
rect 62524 14532 62580 14590
rect 62524 14466 62580 14476
rect 62524 13860 62580 13870
rect 62188 13582 62190 13634
rect 62242 13582 62244 13634
rect 62188 13570 62244 13582
rect 62300 13804 62524 13860
rect 62300 13074 62356 13804
rect 62524 13766 62580 13804
rect 62300 13022 62302 13074
rect 62354 13022 62356 13074
rect 62300 13010 62356 13022
rect 62636 12292 62692 15822
rect 62748 14868 62804 17164
rect 62972 17108 63028 24446
rect 64316 24052 64372 24892
rect 64764 24836 64820 24846
rect 64764 24742 64820 24780
rect 64428 24722 64484 24734
rect 64428 24670 64430 24722
rect 64482 24670 64484 24722
rect 64428 24276 64484 24670
rect 64428 24210 64484 24220
rect 64428 24052 64484 24062
rect 64316 24050 64708 24052
rect 64316 23998 64430 24050
rect 64482 23998 64708 24050
rect 64316 23996 64708 23998
rect 64428 23986 64484 23996
rect 64652 23938 64708 23996
rect 64652 23886 64654 23938
rect 64706 23886 64708 23938
rect 64652 23874 64708 23886
rect 64652 23266 64708 23278
rect 64652 23214 64654 23266
rect 64706 23214 64708 23266
rect 63084 23044 63140 23054
rect 63140 22988 63476 23044
rect 63084 22950 63140 22988
rect 63308 21028 63364 21038
rect 63308 20802 63364 20972
rect 63308 20750 63310 20802
rect 63362 20750 63364 20802
rect 63308 20738 63364 20750
rect 63420 18676 63476 22988
rect 63868 23042 63924 23054
rect 63868 22990 63870 23042
rect 63922 22990 63924 23042
rect 63868 22820 63924 22990
rect 64428 22932 64484 22942
rect 64428 22930 64596 22932
rect 64428 22878 64430 22930
rect 64482 22878 64596 22930
rect 64428 22876 64596 22878
rect 64428 22866 64484 22876
rect 63420 18450 63476 18620
rect 63420 18398 63422 18450
rect 63474 18398 63476 18450
rect 63420 18386 63476 18398
rect 63532 22372 63588 22382
rect 63084 18340 63140 18350
rect 63084 18246 63140 18284
rect 63420 17666 63476 17678
rect 63420 17614 63422 17666
rect 63474 17614 63476 17666
rect 63084 17108 63140 17118
rect 62972 17106 63140 17108
rect 62972 17054 63086 17106
rect 63138 17054 63140 17106
rect 62972 17052 63140 17054
rect 62748 14802 62804 14812
rect 62860 16772 62916 16782
rect 62860 14980 62916 16716
rect 63084 16324 63140 17052
rect 63420 16884 63476 17614
rect 63420 16790 63476 16828
rect 63084 16258 63140 16268
rect 63196 15316 63252 15354
rect 63196 15250 63252 15260
rect 63084 15204 63140 15214
rect 63532 15148 63588 22316
rect 63868 22148 63924 22764
rect 63868 22082 63924 22092
rect 63644 21812 63700 21822
rect 63644 20802 63700 21756
rect 64428 21474 64484 21486
rect 64428 21422 64430 21474
rect 64482 21422 64484 21474
rect 64092 21140 64148 21150
rect 64428 21140 64484 21422
rect 64540 21252 64596 22876
rect 64652 22820 64708 23214
rect 64764 23044 64820 23054
rect 64876 23044 64932 25340
rect 64764 23042 64932 23044
rect 64764 22990 64766 23042
rect 64818 22990 64932 23042
rect 64764 22988 64932 22990
rect 64764 22978 64820 22988
rect 64764 22820 64820 22830
rect 64652 22764 64764 22820
rect 64764 22754 64820 22764
rect 64988 21588 65044 25452
rect 65548 25506 65604 25518
rect 65548 25454 65550 25506
rect 65602 25454 65604 25506
rect 65436 24948 65492 24958
rect 65548 24948 65604 25454
rect 65492 24892 65604 24948
rect 65436 24882 65492 24892
rect 67564 24722 67620 24734
rect 67564 24670 67566 24722
rect 67618 24670 67620 24722
rect 65772 24612 65828 24622
rect 65436 23938 65492 23950
rect 65436 23886 65438 23938
rect 65490 23886 65492 23938
rect 65436 23042 65492 23886
rect 65436 22990 65438 23042
rect 65490 22990 65492 23042
rect 65436 22978 65492 22990
rect 65548 23266 65604 23278
rect 65548 23214 65550 23266
rect 65602 23214 65604 23266
rect 65324 22820 65380 22830
rect 65548 22820 65604 23214
rect 65772 23266 65828 24556
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 67564 24052 67620 24670
rect 67788 24724 67844 26126
rect 67788 24658 67844 24668
rect 68012 25172 68068 25182
rect 68012 24722 68068 25116
rect 68012 24670 68014 24722
rect 68066 24670 68068 24722
rect 68012 24658 68068 24670
rect 67788 24052 67844 24062
rect 67564 23996 67788 24052
rect 67788 23958 67844 23996
rect 65772 23214 65774 23266
rect 65826 23214 65828 23266
rect 65772 23202 65828 23214
rect 68012 23828 68068 23838
rect 65380 22764 65604 22820
rect 65916 22764 66180 22774
rect 65100 22148 65156 22158
rect 65324 22148 65380 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 65100 22146 65380 22148
rect 65100 22094 65102 22146
rect 65154 22094 65380 22146
rect 65100 22092 65380 22094
rect 65100 22082 65156 22092
rect 64988 21532 65156 21588
rect 64540 21196 65044 21252
rect 64428 21084 64820 21140
rect 63644 20750 63646 20802
rect 63698 20750 63700 20802
rect 63644 20738 63700 20750
rect 63868 20804 63924 20814
rect 63868 20802 64036 20804
rect 63868 20750 63870 20802
rect 63922 20750 64036 20802
rect 63868 20748 64036 20750
rect 63868 20738 63924 20748
rect 63868 19796 63924 19806
rect 63868 19234 63924 19740
rect 63980 19460 64036 20748
rect 64092 20802 64148 21084
rect 64092 20750 64094 20802
rect 64146 20750 64148 20802
rect 64092 20468 64148 20750
rect 64428 20916 64484 20926
rect 64092 20402 64148 20412
rect 64316 20690 64372 20702
rect 64316 20638 64318 20690
rect 64370 20638 64372 20690
rect 64316 20244 64372 20638
rect 64428 20578 64484 20860
rect 64428 20526 64430 20578
rect 64482 20526 64484 20578
rect 64428 20514 64484 20526
rect 64652 20804 64708 20814
rect 64428 20244 64484 20254
rect 64316 20242 64484 20244
rect 64316 20190 64430 20242
rect 64482 20190 64484 20242
rect 64316 20188 64484 20190
rect 64428 20178 64484 20188
rect 64540 19908 64596 19918
rect 64652 19908 64708 20748
rect 64428 19906 64708 19908
rect 64428 19854 64542 19906
rect 64594 19854 64708 19906
rect 64428 19852 64708 19854
rect 64764 20802 64820 21084
rect 64764 20750 64766 20802
rect 64818 20750 64820 20802
rect 63980 19404 64372 19460
rect 64204 19236 64260 19246
rect 63868 19182 63870 19234
rect 63922 19182 63924 19234
rect 63868 19170 63924 19182
rect 63980 19180 64204 19236
rect 63980 19012 64036 19180
rect 64204 19142 64260 19180
rect 63756 18956 64036 19012
rect 63756 18338 63812 18956
rect 63756 18286 63758 18338
rect 63810 18286 63812 18338
rect 63756 18274 63812 18286
rect 64204 18564 64260 18574
rect 64204 17780 64260 18508
rect 64316 18004 64372 19404
rect 64428 18450 64484 19852
rect 64540 19842 64596 19852
rect 64764 19796 64820 20750
rect 64988 20132 65044 21196
rect 64652 19740 64820 19796
rect 64876 20076 65044 20132
rect 64652 19236 64708 19740
rect 64652 19170 64708 19180
rect 64428 18398 64430 18450
rect 64482 18398 64484 18450
rect 64428 18386 64484 18398
rect 64540 19124 64596 19134
rect 64316 17938 64372 17948
rect 64428 17892 64484 17902
rect 64540 17892 64596 19068
rect 64764 19122 64820 19134
rect 64764 19070 64766 19122
rect 64818 19070 64820 19122
rect 64764 18676 64820 19070
rect 64764 18610 64820 18620
rect 64428 17890 64596 17892
rect 64428 17838 64430 17890
rect 64482 17838 64596 17890
rect 64428 17836 64596 17838
rect 64428 17826 64484 17836
rect 64316 17780 64372 17790
rect 64204 17778 64372 17780
rect 64204 17726 64318 17778
rect 64370 17726 64372 17778
rect 64204 17724 64372 17726
rect 63868 17668 63924 17678
rect 63868 17574 63924 17612
rect 63756 17108 63812 17118
rect 63756 16994 63812 17052
rect 63756 16942 63758 16994
rect 63810 16942 63812 16994
rect 63756 16930 63812 16942
rect 64316 16210 64372 17724
rect 64540 17108 64596 17118
rect 64540 17014 64596 17052
rect 64316 16158 64318 16210
rect 64370 16158 64372 16210
rect 64316 16146 64372 16158
rect 64540 16884 64596 16894
rect 64540 16098 64596 16828
rect 64540 16046 64542 16098
rect 64594 16046 64596 16098
rect 64540 16034 64596 16046
rect 64092 15876 64148 15886
rect 63868 15874 64148 15876
rect 63868 15822 64094 15874
rect 64146 15822 64148 15874
rect 63868 15820 64148 15822
rect 63084 15092 63252 15148
rect 62860 14642 62916 14924
rect 62860 14590 62862 14642
rect 62914 14590 62916 14642
rect 62860 14578 62916 14590
rect 62860 14084 62916 14094
rect 62860 13970 62916 14028
rect 62860 13918 62862 13970
rect 62914 13918 62916 13970
rect 62860 13906 62916 13918
rect 63084 13524 63140 13534
rect 62860 13522 63140 13524
rect 62860 13470 63086 13522
rect 63138 13470 63140 13522
rect 62860 13468 63140 13470
rect 62748 13300 62804 13310
rect 62748 13074 62804 13244
rect 62748 13022 62750 13074
rect 62802 13022 62804 13074
rect 62748 13010 62804 13022
rect 62076 11330 62132 11340
rect 62300 12236 62692 12292
rect 61628 11284 61684 11294
rect 61516 11282 61684 11284
rect 61516 11230 61630 11282
rect 61682 11230 61684 11282
rect 61516 11228 61684 11230
rect 61628 11172 61684 11228
rect 61628 11106 61684 11116
rect 61964 11172 62020 11182
rect 61964 11078 62020 11116
rect 62076 11170 62132 11182
rect 62076 11118 62078 11170
rect 62130 11118 62132 11170
rect 61964 10948 62020 10958
rect 61404 10332 61796 10388
rect 61292 9826 61348 10332
rect 61292 9774 61294 9826
rect 61346 9774 61348 9826
rect 61292 9762 61348 9774
rect 61180 9538 61236 9548
rect 61628 9602 61684 9614
rect 61628 9550 61630 9602
rect 61682 9550 61684 9602
rect 61180 9268 61236 9278
rect 61180 9174 61236 9212
rect 61628 9156 61684 9550
rect 61404 9100 61684 9156
rect 61740 9380 61796 10332
rect 61964 10164 62020 10892
rect 62076 10388 62132 11118
rect 62188 11170 62244 11182
rect 62188 11118 62190 11170
rect 62242 11118 62244 11170
rect 62188 10724 62244 11118
rect 62188 10658 62244 10668
rect 62076 10322 62132 10332
rect 61964 10108 62132 10164
rect 61964 9716 62020 9726
rect 62076 9716 62132 10108
rect 61740 9154 61796 9324
rect 61740 9102 61742 9154
rect 61794 9102 61796 9154
rect 61068 8148 61124 8158
rect 61404 8148 61460 9100
rect 61740 8596 61796 9102
rect 61852 9714 62132 9716
rect 61852 9662 61966 9714
rect 62018 9662 62132 9714
rect 61852 9660 62132 9662
rect 61852 9044 61908 9660
rect 61964 9650 62020 9660
rect 61852 8978 61908 8988
rect 62076 9154 62132 9166
rect 62076 9102 62078 9154
rect 62130 9102 62132 9154
rect 62076 9044 62132 9102
rect 61740 8540 62020 8596
rect 61740 8372 61796 8382
rect 61628 8316 61740 8372
rect 61068 8146 61460 8148
rect 61068 8094 61070 8146
rect 61122 8094 61460 8146
rect 61068 8092 61460 8094
rect 61516 8146 61572 8158
rect 61516 8094 61518 8146
rect 61570 8094 61572 8146
rect 61068 8082 61124 8092
rect 60956 7644 61124 7700
rect 60844 7532 61012 7588
rect 60844 7364 60900 7402
rect 60844 7298 60900 7308
rect 60508 6860 60788 6916
rect 60844 7140 60900 7150
rect 60508 5348 60564 6860
rect 60732 6692 60788 6702
rect 60732 6598 60788 6636
rect 60620 6020 60676 6030
rect 60620 5926 60676 5964
rect 60620 5348 60676 5358
rect 60508 5346 60676 5348
rect 60508 5294 60622 5346
rect 60674 5294 60676 5346
rect 60508 5292 60676 5294
rect 60620 5282 60676 5292
rect 60732 5124 60788 5134
rect 60844 5124 60900 7084
rect 60956 6692 61012 7532
rect 61068 7364 61124 7644
rect 61068 7298 61124 7308
rect 61068 6916 61124 6926
rect 61068 6822 61124 6860
rect 60956 6636 61124 6692
rect 60732 5122 60900 5124
rect 60732 5070 60734 5122
rect 60786 5070 60900 5122
rect 60732 5068 60900 5070
rect 60732 5058 60788 5068
rect 60620 5012 60676 5022
rect 60452 5010 60676 5012
rect 60452 4958 60622 5010
rect 60674 4958 60676 5010
rect 60452 4956 60676 4958
rect 60396 4918 60452 4956
rect 60620 4946 60676 4956
rect 61068 4450 61124 6636
rect 61180 6580 61236 8092
rect 61292 7588 61348 7598
rect 61292 6914 61348 7532
rect 61516 7362 61572 8094
rect 61516 7310 61518 7362
rect 61570 7310 61572 7362
rect 61516 7298 61572 7310
rect 61292 6862 61294 6914
rect 61346 6862 61348 6914
rect 61292 6850 61348 6862
rect 61516 7140 61572 7150
rect 61180 6514 61236 6524
rect 61516 6018 61572 7084
rect 61628 6802 61684 8316
rect 61740 8306 61796 8316
rect 61852 8260 61908 8270
rect 61852 7140 61908 8204
rect 61964 7588 62020 8540
rect 61964 7522 62020 7532
rect 61852 7074 61908 7084
rect 61628 6750 61630 6802
rect 61682 6750 61684 6802
rect 61628 6738 61684 6750
rect 61852 6804 61908 6814
rect 62076 6804 62132 8988
rect 62300 8820 62356 12236
rect 62636 12068 62692 12078
rect 62524 12066 62692 12068
rect 62524 12014 62638 12066
rect 62690 12014 62692 12066
rect 62524 12012 62692 12014
rect 62412 11170 62468 11182
rect 62412 11118 62414 11170
rect 62466 11118 62468 11170
rect 62412 10836 62468 11118
rect 62412 10770 62468 10780
rect 62524 10052 62580 12012
rect 62636 12002 62692 12012
rect 62860 11284 62916 13468
rect 63084 13458 63140 13468
rect 63196 12404 63252 15092
rect 63308 15092 63364 15102
rect 63308 14642 63364 15036
rect 63420 15092 63588 15148
rect 63644 15428 63700 15438
rect 63420 14754 63476 15092
rect 63420 14702 63422 14754
rect 63474 14702 63476 14754
rect 63420 14690 63476 14702
rect 63308 14590 63310 14642
rect 63362 14590 63364 14642
rect 63308 14578 63364 14590
rect 63644 14532 63700 15372
rect 63756 15316 63812 15326
rect 63756 15222 63812 15260
rect 63868 15148 63924 15820
rect 64092 15810 64148 15820
rect 64428 15314 64484 15326
rect 64428 15262 64430 15314
rect 64482 15262 64484 15314
rect 63868 15092 64036 15148
rect 63644 14466 63700 14476
rect 63756 14644 63812 14654
rect 63756 13972 63812 14588
rect 63756 13878 63812 13916
rect 63308 13634 63364 13646
rect 63308 13582 63310 13634
rect 63362 13582 63364 13634
rect 63308 13522 63364 13582
rect 63308 13470 63310 13522
rect 63362 13470 63364 13522
rect 63308 13458 63364 13470
rect 63420 13076 63476 13086
rect 63420 12982 63476 13020
rect 63868 13076 63924 13086
rect 63868 12962 63924 13020
rect 63868 12910 63870 12962
rect 63922 12910 63924 12962
rect 63868 12898 63924 12910
rect 63196 12348 63700 12404
rect 63084 12180 63140 12190
rect 62972 12066 63028 12078
rect 62972 12014 62974 12066
rect 63026 12014 63028 12066
rect 62972 11844 63028 12014
rect 62972 11618 63028 11788
rect 62972 11566 62974 11618
rect 63026 11566 63028 11618
rect 62972 11554 63028 11566
rect 62412 9996 62580 10052
rect 62636 11228 62916 11284
rect 62412 9492 62468 9996
rect 62524 9828 62580 9838
rect 62524 9734 62580 9772
rect 62636 9714 62692 11228
rect 62972 11172 63028 11182
rect 62860 11170 63028 11172
rect 62860 11118 62974 11170
rect 63026 11118 63028 11170
rect 62860 11116 63028 11118
rect 62860 10836 62916 11116
rect 62972 11106 63028 11116
rect 62860 10770 62916 10780
rect 62972 10724 63028 10734
rect 62972 10498 63028 10668
rect 63084 10612 63140 12124
rect 63420 12066 63476 12078
rect 63420 12014 63422 12066
rect 63474 12014 63476 12066
rect 63308 11618 63364 11630
rect 63308 11566 63310 11618
rect 63362 11566 63364 11618
rect 63308 11060 63364 11566
rect 63420 11172 63476 12014
rect 63532 11618 63588 11630
rect 63532 11566 63534 11618
rect 63586 11566 63588 11618
rect 63532 11506 63588 11566
rect 63532 11454 63534 11506
rect 63586 11454 63588 11506
rect 63532 11442 63588 11454
rect 63420 11116 63588 11172
rect 63308 11004 63476 11060
rect 63420 10778 63476 11004
rect 63420 10726 63422 10778
rect 63474 10726 63476 10778
rect 63420 10714 63476 10726
rect 63084 10546 63140 10556
rect 63308 10610 63364 10622
rect 63308 10558 63310 10610
rect 63362 10558 63364 10610
rect 62972 10446 62974 10498
rect 63026 10446 63028 10498
rect 62972 10434 63028 10446
rect 62636 9662 62638 9714
rect 62690 9662 62692 9714
rect 62412 9436 62580 9492
rect 62412 9268 62468 9278
rect 62412 9174 62468 9212
rect 61852 6802 62132 6804
rect 61852 6750 61854 6802
rect 61906 6750 62132 6802
rect 61852 6748 62132 6750
rect 62188 8764 62356 8820
rect 61852 6738 61908 6748
rect 61740 6690 61796 6702
rect 61740 6638 61742 6690
rect 61794 6638 61796 6690
rect 61740 6468 61796 6638
rect 61740 6402 61796 6412
rect 62188 6468 62244 8764
rect 62300 8596 62356 8606
rect 62300 6690 62356 8540
rect 62524 7812 62580 9436
rect 62636 8596 62692 9662
rect 63084 9828 63140 9838
rect 63308 9828 63364 10558
rect 63420 10612 63476 10622
rect 63420 10386 63476 10556
rect 63420 10334 63422 10386
rect 63474 10334 63476 10386
rect 63420 10322 63476 10334
rect 63420 9828 63476 9838
rect 63308 9772 63420 9828
rect 62860 9604 62916 9614
rect 62860 9510 62916 9548
rect 63084 9266 63140 9772
rect 63420 9734 63476 9772
rect 63084 9214 63086 9266
rect 63138 9214 63140 9266
rect 63084 9202 63140 9214
rect 63532 9714 63588 11116
rect 63644 9828 63700 12348
rect 63868 12066 63924 12078
rect 63868 12014 63870 12066
rect 63922 12014 63924 12066
rect 63756 9828 63812 9838
rect 63644 9826 63812 9828
rect 63644 9774 63758 9826
rect 63810 9774 63812 9826
rect 63644 9772 63812 9774
rect 63756 9762 63812 9772
rect 63532 9662 63534 9714
rect 63586 9662 63588 9714
rect 62748 9044 62804 9054
rect 62748 8950 62804 8988
rect 63420 9044 63476 9054
rect 62636 8530 62692 8540
rect 62524 7746 62580 7756
rect 62860 8370 62916 8382
rect 62860 8318 62862 8370
rect 62914 8318 62916 8370
rect 62860 7700 62916 8318
rect 63420 8372 63476 8988
rect 63420 8306 63476 8316
rect 62860 7634 62916 7644
rect 63196 8258 63252 8270
rect 63196 8206 63198 8258
rect 63250 8206 63252 8258
rect 63196 6804 63252 8206
rect 63532 8148 63588 9662
rect 63420 8092 63588 8148
rect 63196 6738 63252 6748
rect 63308 7364 63364 7374
rect 62300 6638 62302 6690
rect 62354 6638 62356 6690
rect 62300 6626 62356 6638
rect 62188 6402 62244 6412
rect 63084 6468 63140 6478
rect 61516 5966 61518 6018
rect 61570 5966 61572 6018
rect 61516 4676 61572 5966
rect 61516 4610 61572 4620
rect 61628 5234 61684 5246
rect 61628 5182 61630 5234
rect 61682 5182 61684 5234
rect 61068 4398 61070 4450
rect 61122 4398 61124 4450
rect 61068 4386 61124 4398
rect 61404 3554 61460 3566
rect 61404 3502 61406 3554
rect 61458 3502 61460 3554
rect 61404 2548 61460 3502
rect 61404 2482 61460 2492
rect 61628 800 61684 5182
rect 61964 5124 62020 5134
rect 61740 5012 61796 5022
rect 61740 4338 61796 4956
rect 61740 4286 61742 4338
rect 61794 4286 61796 4338
rect 61740 4274 61796 4286
rect 61964 3554 62020 5068
rect 61964 3502 61966 3554
rect 62018 3502 62020 3554
rect 61964 3490 62020 3502
rect 62524 4452 62580 4462
rect 61740 3444 61796 3482
rect 62524 3444 62580 4396
rect 62636 4228 62692 4238
rect 62636 4226 62916 4228
rect 62636 4174 62638 4226
rect 62690 4174 62916 4226
rect 62636 4172 62916 4174
rect 62636 4162 62692 4172
rect 62860 3554 62916 4172
rect 62860 3502 62862 3554
rect 62914 3502 62916 3554
rect 62860 3490 62916 3502
rect 62636 3444 62692 3454
rect 62524 3442 62692 3444
rect 62524 3390 62638 3442
rect 62690 3390 62692 3442
rect 62524 3388 62692 3390
rect 61740 3378 61796 3388
rect 62636 3378 62692 3388
rect 63084 2996 63140 6412
rect 63308 4116 63364 7308
rect 63420 7140 63476 8092
rect 63420 6578 63476 7084
rect 63420 6526 63422 6578
rect 63474 6526 63476 6578
rect 63420 6514 63476 6526
rect 63532 7812 63588 7822
rect 63532 7586 63588 7756
rect 63532 7534 63534 7586
rect 63586 7534 63588 7586
rect 63308 4050 63364 4060
rect 63532 3388 63588 7534
rect 63868 5908 63924 12014
rect 63980 11618 64036 15092
rect 64092 14308 64148 14318
rect 64428 14308 64484 15262
rect 64876 15148 64932 20076
rect 64988 19906 65044 19918
rect 64988 19854 64990 19906
rect 65042 19854 65044 19906
rect 64988 19796 65044 19854
rect 64988 19730 65044 19740
rect 65100 19124 65156 21532
rect 65212 20804 65268 20814
rect 65212 20710 65268 20748
rect 65324 20132 65380 22092
rect 65324 20066 65380 20076
rect 65436 22596 65492 22606
rect 65436 19908 65492 22540
rect 67340 21586 67396 21598
rect 67340 21534 67342 21586
rect 67394 21534 67396 21586
rect 66556 21474 66612 21486
rect 66556 21422 66558 21474
rect 66610 21422 66612 21474
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 66556 20916 66612 21422
rect 67340 21476 67396 21534
rect 67788 21476 67844 21486
rect 67340 21474 67844 21476
rect 67340 21422 67790 21474
rect 67842 21422 67844 21474
rect 67340 21420 67844 21422
rect 66556 20850 66612 20860
rect 64652 15092 64932 15148
rect 64988 19068 65156 19124
rect 65212 19852 65492 19908
rect 65548 20802 65604 20814
rect 65548 20750 65550 20802
rect 65602 20750 65604 20802
rect 64092 14306 64484 14308
rect 64092 14254 64094 14306
rect 64146 14254 64484 14306
rect 64092 14252 64484 14254
rect 64540 14868 64596 14878
rect 64540 14306 64596 14812
rect 64540 14254 64542 14306
rect 64594 14254 64596 14306
rect 64092 13076 64148 14252
rect 64540 14196 64596 14254
rect 64316 14140 64596 14196
rect 64316 13524 64372 14140
rect 64540 13972 64596 13982
rect 64652 13972 64708 15092
rect 64988 14644 65044 19068
rect 65212 18900 65268 19852
rect 65436 19684 65492 19694
rect 65212 18844 65380 18900
rect 65100 18676 65156 18686
rect 65100 18562 65156 18620
rect 65100 18510 65102 18562
rect 65154 18510 65156 18562
rect 65100 18498 65156 18510
rect 65100 17668 65156 17678
rect 65100 15986 65156 17612
rect 65100 15934 65102 15986
rect 65154 15934 65156 15986
rect 65100 15922 65156 15934
rect 64540 13970 64708 13972
rect 64540 13918 64542 13970
rect 64594 13918 64708 13970
rect 64540 13916 64708 13918
rect 64764 14588 65044 14644
rect 65212 15202 65268 15214
rect 65212 15150 65214 15202
rect 65266 15150 65268 15202
rect 64764 14196 64820 14588
rect 64988 14420 65044 14430
rect 64540 13906 64596 13916
rect 64428 13748 64484 13758
rect 64428 13654 64484 13692
rect 64652 13748 64708 13758
rect 64764 13748 64820 14140
rect 64652 13746 64820 13748
rect 64652 13694 64654 13746
rect 64706 13694 64820 13746
rect 64652 13692 64820 13694
rect 64876 14418 65044 14420
rect 64876 14366 64990 14418
rect 65042 14366 65044 14418
rect 64876 14364 65044 14366
rect 64652 13682 64708 13692
rect 64316 13468 64484 13524
rect 64092 13010 64148 13020
rect 64316 11956 64372 11966
rect 63980 11566 63982 11618
rect 64034 11566 64036 11618
rect 63980 11554 64036 11566
rect 64092 11954 64372 11956
rect 64092 11902 64318 11954
rect 64370 11902 64372 11954
rect 64092 11900 64372 11902
rect 63980 11170 64036 11182
rect 63980 11118 63982 11170
rect 64034 11118 64036 11170
rect 63980 10612 64036 11118
rect 63980 10546 64036 10556
rect 64092 10050 64148 11900
rect 64316 11890 64372 11900
rect 64204 11396 64260 11406
rect 64204 11172 64260 11340
rect 64316 11172 64372 11182
rect 64204 11170 64372 11172
rect 64204 11118 64318 11170
rect 64370 11118 64372 11170
rect 64204 11116 64372 11118
rect 64316 11060 64372 11116
rect 64316 10994 64372 11004
rect 64092 9998 64094 10050
rect 64146 9998 64148 10050
rect 64092 9986 64148 9998
rect 64204 9716 64260 9726
rect 64204 9622 64260 9660
rect 64092 9602 64148 9614
rect 64092 9550 64094 9602
rect 64146 9550 64148 9602
rect 63980 8932 64036 8942
rect 63980 8838 64036 8876
rect 63980 8484 64036 8494
rect 63980 8370 64036 8428
rect 63980 8318 63982 8370
rect 64034 8318 64036 8370
rect 63980 8306 64036 8318
rect 63868 5842 63924 5852
rect 63756 5794 63812 5806
rect 63756 5742 63758 5794
rect 63810 5742 63812 5794
rect 63644 5122 63700 5134
rect 63644 5070 63646 5122
rect 63698 5070 63700 5122
rect 63644 4900 63700 5070
rect 63644 4834 63700 4844
rect 63756 4450 63812 5742
rect 64092 5796 64148 9550
rect 64316 9604 64372 9614
rect 64316 9042 64372 9548
rect 64316 8990 64318 9042
rect 64370 8990 64372 9042
rect 64316 8978 64372 8990
rect 64428 8820 64484 13468
rect 64876 13188 64932 14364
rect 64988 14354 65044 14364
rect 65212 14306 65268 15150
rect 65324 14868 65380 18844
rect 65436 17554 65492 19628
rect 65436 17502 65438 17554
rect 65490 17502 65492 17554
rect 65436 17490 65492 17502
rect 65548 18116 65604 20750
rect 67004 20802 67060 20814
rect 67004 20750 67006 20802
rect 67058 20750 67060 20802
rect 65772 20690 65828 20702
rect 65772 20638 65774 20690
rect 65826 20638 65828 20690
rect 65772 19124 65828 20638
rect 66220 20690 66276 20702
rect 66556 20692 66612 20702
rect 66220 20638 66222 20690
rect 66274 20638 66276 20690
rect 66220 19796 66276 20638
rect 66444 20690 66612 20692
rect 66444 20638 66558 20690
rect 66610 20638 66612 20690
rect 66444 20636 66612 20638
rect 66220 19730 66276 19740
rect 66332 20468 66388 20478
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 66332 19234 66388 20412
rect 66332 19182 66334 19234
rect 66386 19182 66388 19234
rect 66332 19170 66388 19182
rect 65772 19058 65828 19068
rect 66444 18564 66500 20636
rect 66556 20626 66612 20636
rect 66892 20132 66948 20142
rect 66780 19348 66836 19358
rect 66780 19254 66836 19292
rect 66892 19236 66948 20076
rect 67004 19908 67060 20750
rect 67788 20020 67844 21420
rect 68012 21028 68068 23772
rect 68236 22484 68292 28812
rect 69132 28642 69188 28654
rect 69132 28590 69134 28642
rect 69186 28590 69188 28642
rect 69132 27186 69188 28590
rect 69356 28420 69412 28430
rect 69356 28326 69412 28364
rect 69132 27134 69134 27186
rect 69186 27134 69188 27186
rect 68460 27076 68516 27086
rect 68460 26964 68516 27020
rect 68460 26962 69076 26964
rect 68460 26910 68462 26962
rect 68514 26910 69076 26962
rect 68460 26908 69076 26910
rect 68460 26898 68516 26908
rect 68796 26628 68852 26638
rect 68348 26404 68404 26414
rect 68348 26310 68404 26348
rect 68796 25508 68852 26572
rect 69020 26292 69076 26908
rect 69132 26628 69188 27134
rect 69132 26562 69188 26572
rect 69244 27074 69300 27086
rect 69244 27022 69246 27074
rect 69298 27022 69300 27074
rect 69020 26236 69188 26292
rect 68908 26180 68964 26190
rect 68908 26178 69076 26180
rect 68908 26126 68910 26178
rect 68962 26126 69076 26178
rect 68908 26124 69076 26126
rect 68908 26114 68964 26124
rect 68908 25508 68964 25518
rect 68796 25506 68964 25508
rect 68796 25454 68910 25506
rect 68962 25454 68964 25506
rect 68796 25452 68964 25454
rect 68908 25284 68964 25452
rect 68908 25218 68964 25228
rect 68684 25172 68740 25182
rect 68684 24834 68740 25116
rect 68908 24948 68964 24986
rect 68908 24882 68964 24892
rect 68684 24782 68686 24834
rect 68738 24782 68740 24834
rect 68684 24770 68740 24782
rect 68348 24724 68404 24734
rect 68348 24630 68404 24668
rect 68908 24724 68964 24734
rect 68908 23938 68964 24668
rect 69020 24052 69076 26124
rect 69020 23986 69076 23996
rect 68908 23886 68910 23938
rect 68962 23886 68964 23938
rect 68908 23874 68964 23886
rect 68796 23828 68852 23838
rect 68796 23734 68852 23772
rect 68572 23714 68628 23726
rect 68572 23662 68574 23714
rect 68626 23662 68628 23714
rect 68572 23492 68628 23662
rect 69132 23604 69188 26236
rect 69244 25172 69300 27022
rect 69468 26964 69524 30716
rect 73388 30548 73444 30558
rect 73388 28756 73444 30492
rect 73388 28754 73780 28756
rect 73388 28702 73390 28754
rect 73442 28702 73780 28754
rect 73388 28700 73780 28702
rect 73388 28690 73444 28700
rect 72716 28644 72772 28654
rect 72716 28642 72884 28644
rect 72716 28590 72718 28642
rect 72770 28590 72884 28642
rect 72716 28588 72884 28590
rect 72716 28578 72772 28588
rect 70588 28420 70644 28430
rect 71036 28420 71092 28430
rect 70364 28418 70644 28420
rect 70364 28366 70590 28418
rect 70642 28366 70644 28418
rect 70364 28364 70644 28366
rect 69692 27858 69748 27870
rect 69692 27806 69694 27858
rect 69746 27806 69748 27858
rect 69692 27412 69748 27806
rect 70364 27860 70420 28364
rect 70588 28354 70644 28364
rect 70924 28418 71092 28420
rect 70924 28366 71038 28418
rect 71090 28366 71092 28418
rect 70924 28364 71092 28366
rect 70924 27970 70980 28364
rect 71036 28354 71092 28364
rect 72716 28420 72772 28430
rect 70924 27918 70926 27970
rect 70978 27918 70980 27970
rect 70364 27766 70420 27804
rect 70700 27858 70756 27870
rect 70700 27806 70702 27858
rect 70754 27806 70756 27858
rect 70700 27636 70756 27806
rect 70700 27570 70756 27580
rect 70812 27746 70868 27758
rect 70812 27694 70814 27746
rect 70866 27694 70868 27746
rect 70140 27412 70196 27422
rect 70812 27412 70868 27694
rect 69692 27356 69972 27412
rect 69580 27188 69636 27198
rect 69916 27188 69972 27356
rect 70028 27188 70084 27198
rect 69916 27186 70084 27188
rect 69916 27134 70030 27186
rect 70082 27134 70084 27186
rect 69916 27132 70084 27134
rect 69580 27094 69636 27132
rect 70028 27122 70084 27132
rect 69804 27074 69860 27086
rect 69804 27022 69806 27074
rect 69858 27022 69860 27074
rect 69804 26964 69860 27022
rect 69468 26908 69748 26964
rect 69468 26404 69524 26414
rect 69468 25506 69524 26348
rect 69468 25454 69470 25506
rect 69522 25454 69524 25506
rect 69468 25442 69524 25454
rect 69244 25106 69300 25116
rect 69468 25284 69524 25294
rect 69356 25060 69412 25070
rect 69244 24052 69300 24062
rect 69244 23958 69300 23996
rect 69356 23828 69412 25004
rect 69468 24946 69524 25228
rect 69468 24894 69470 24946
rect 69522 24894 69524 24946
rect 69468 24882 69524 24894
rect 69580 25172 69636 25182
rect 69580 24946 69636 25116
rect 69580 24894 69582 24946
rect 69634 24894 69636 24946
rect 69580 24882 69636 24894
rect 69468 24612 69524 24622
rect 69468 24518 69524 24556
rect 69356 23734 69412 23772
rect 68572 23426 68628 23436
rect 68908 23548 69188 23604
rect 68348 22484 68404 22494
rect 68236 22482 68404 22484
rect 68236 22430 68350 22482
rect 68402 22430 68404 22482
rect 68236 22428 68404 22430
rect 68348 22418 68404 22428
rect 68012 20962 68068 20972
rect 68908 21474 68964 23548
rect 69692 21812 69748 26908
rect 70140 26908 70196 27356
rect 70252 27356 70868 27412
rect 70252 27074 70308 27356
rect 70252 27022 70254 27074
rect 70306 27022 70308 27074
rect 70252 27010 70308 27022
rect 70364 27076 70420 27086
rect 70364 26982 70420 27020
rect 70924 26908 70980 27918
rect 71372 28084 71428 28094
rect 71148 27858 71204 27870
rect 71148 27806 71150 27858
rect 71202 27806 71204 27858
rect 71148 27412 71204 27806
rect 71148 27346 71204 27356
rect 71372 27300 71428 28028
rect 71484 27860 71540 27870
rect 72716 27860 72772 28364
rect 71484 27858 71988 27860
rect 71484 27806 71486 27858
rect 71538 27806 71988 27858
rect 71484 27804 71988 27806
rect 71484 27794 71540 27804
rect 71596 27300 71652 27310
rect 71372 27244 71596 27300
rect 71596 27206 71652 27244
rect 71708 27076 71764 27086
rect 71708 26982 71764 27020
rect 71932 27074 71988 27804
rect 72492 27858 72772 27860
rect 72492 27806 72718 27858
rect 72770 27806 72772 27858
rect 72492 27804 72772 27806
rect 71932 27022 71934 27074
rect 71986 27022 71988 27074
rect 71932 27010 71988 27022
rect 72268 27746 72324 27758
rect 72268 27694 72270 27746
rect 72322 27694 72324 27746
rect 72268 27074 72324 27694
rect 72268 27022 72270 27074
rect 72322 27022 72324 27074
rect 72268 27010 72324 27022
rect 72380 27300 72436 27310
rect 69804 26898 69860 26908
rect 69916 26852 70196 26908
rect 70252 26852 70308 26862
rect 69916 25620 69972 26852
rect 70140 26404 70196 26414
rect 70252 26404 70308 26796
rect 70700 26852 70980 26908
rect 71260 26964 71316 26974
rect 72380 26908 72436 27244
rect 71260 26852 71428 26908
rect 70140 26402 70308 26404
rect 70140 26350 70142 26402
rect 70194 26350 70308 26402
rect 70140 26348 70308 26350
rect 70476 26628 70532 26638
rect 70140 26338 70196 26348
rect 70476 26292 70532 26572
rect 70588 26292 70644 26302
rect 70476 26290 70644 26292
rect 70476 26238 70590 26290
rect 70642 26238 70644 26290
rect 70476 26236 70644 26238
rect 70588 26226 70644 26236
rect 69804 25618 69972 25620
rect 69804 25566 69918 25618
rect 69970 25566 69972 25618
rect 69804 25564 69972 25566
rect 69804 24946 69860 25564
rect 69916 25554 69972 25564
rect 70476 25620 70532 25630
rect 70476 25506 70532 25564
rect 70476 25454 70478 25506
rect 70530 25454 70532 25506
rect 70476 25442 70532 25454
rect 70700 25508 70756 26852
rect 70700 25414 70756 25452
rect 70812 25506 70868 25518
rect 71148 25508 71204 25518
rect 70812 25454 70814 25506
rect 70866 25454 70868 25506
rect 69916 25396 69972 25406
rect 69916 25302 69972 25340
rect 69804 24894 69806 24946
rect 69858 24894 69860 24946
rect 69804 24882 69860 24894
rect 70028 25284 70084 25294
rect 70028 24834 70084 25228
rect 70588 25284 70644 25294
rect 70588 25190 70644 25228
rect 70364 25172 70420 25182
rect 70420 25116 70532 25172
rect 70364 25106 70420 25116
rect 70476 24948 70532 25116
rect 70588 24948 70644 24958
rect 70476 24946 70644 24948
rect 70476 24894 70590 24946
rect 70642 24894 70644 24946
rect 70476 24892 70644 24894
rect 70588 24882 70644 24892
rect 70028 24782 70030 24834
rect 70082 24782 70084 24834
rect 70028 24770 70084 24782
rect 70364 24724 70420 24734
rect 70364 24630 70420 24668
rect 70700 24612 70756 24622
rect 70812 24612 70868 25454
rect 71036 25506 71204 25508
rect 71036 25454 71150 25506
rect 71202 25454 71204 25506
rect 71036 25452 71204 25454
rect 70924 24948 70980 24958
rect 71036 24948 71092 25452
rect 71148 25442 71204 25452
rect 70924 24946 71092 24948
rect 70924 24894 70926 24946
rect 70978 24894 71092 24946
rect 70924 24892 71092 24894
rect 71260 24948 71316 24958
rect 70924 24882 70980 24892
rect 71148 24836 71204 24846
rect 71148 24742 71204 24780
rect 71260 24834 71316 24892
rect 71260 24782 71262 24834
rect 71314 24782 71316 24834
rect 71260 24770 71316 24782
rect 70700 24610 70868 24612
rect 70700 24558 70702 24610
rect 70754 24558 70868 24610
rect 70700 24556 70868 24558
rect 70700 24546 70756 24556
rect 71372 24500 71428 26852
rect 72156 26850 72212 26862
rect 72156 26798 72158 26850
rect 72210 26798 72212 26850
rect 71708 26516 71764 26526
rect 71596 26460 71708 26516
rect 71596 25620 71652 26460
rect 71708 26422 71764 26460
rect 72156 26516 72212 26798
rect 72156 26450 72212 26460
rect 72268 26852 72436 26908
rect 72268 26402 72324 26852
rect 72492 26628 72548 27804
rect 72716 27794 72772 27804
rect 72828 27186 72884 28588
rect 72940 28418 72996 28430
rect 72940 28366 72942 28418
rect 72994 28366 72996 28418
rect 72940 27748 72996 28366
rect 73724 27970 73780 28700
rect 73724 27918 73726 27970
rect 73778 27918 73780 27970
rect 73724 27906 73780 27918
rect 73948 27858 74004 27870
rect 73948 27806 73950 27858
rect 74002 27806 74004 27858
rect 73164 27748 73220 27758
rect 72940 27746 73444 27748
rect 72940 27694 73166 27746
rect 73218 27694 73444 27746
rect 72940 27692 73444 27694
rect 73164 27682 73220 27692
rect 72828 27134 72830 27186
rect 72882 27134 72884 27186
rect 72828 26852 72884 27134
rect 73276 27076 73332 27086
rect 73276 26982 73332 27020
rect 73388 26908 73444 27692
rect 73948 27636 74004 27806
rect 73948 27570 74004 27580
rect 73612 27300 73668 27310
rect 73612 27074 73668 27244
rect 73612 27022 73614 27074
rect 73666 27022 73668 27074
rect 73612 27010 73668 27022
rect 73724 26964 73780 26974
rect 73388 26852 73668 26908
rect 73724 26870 73780 26908
rect 73948 26964 74004 26974
rect 73948 26870 74004 26908
rect 72828 26786 72884 26796
rect 72492 26572 73332 26628
rect 72492 26514 72548 26572
rect 72492 26462 72494 26514
rect 72546 26462 72548 26514
rect 72492 26450 72548 26462
rect 72716 26460 73108 26516
rect 72268 26350 72270 26402
rect 72322 26350 72324 26402
rect 72268 26338 72324 26350
rect 72716 26402 72772 26460
rect 72716 26350 72718 26402
rect 72770 26350 72772 26402
rect 71596 25526 71652 25564
rect 71708 26180 71764 26190
rect 71708 24836 71764 26124
rect 72716 25732 72772 26350
rect 73052 26402 73108 26460
rect 73276 26514 73332 26572
rect 73276 26462 73278 26514
rect 73330 26462 73332 26514
rect 73276 26450 73332 26462
rect 73052 26350 73054 26402
rect 73106 26350 73108 26402
rect 73052 26338 73108 26350
rect 72828 26292 72884 26302
rect 72828 26198 72884 26236
rect 73612 26292 73668 26852
rect 74060 26852 74116 30828
rect 74284 27748 74340 27758
rect 74284 27654 74340 27692
rect 74172 27188 74228 27198
rect 74172 27074 74228 27132
rect 74172 27022 74174 27074
rect 74226 27022 74228 27074
rect 74172 27010 74228 27022
rect 74060 26786 74116 26796
rect 74284 26850 74340 26862
rect 74284 26798 74286 26850
rect 74338 26798 74340 26850
rect 74284 26628 74340 26798
rect 73724 26572 74340 26628
rect 73724 26292 73780 26572
rect 73948 26404 74004 26442
rect 74004 26348 74116 26404
rect 73948 26338 74004 26348
rect 73612 26290 73780 26292
rect 73612 26238 73614 26290
rect 73666 26238 73780 26290
rect 73612 26236 73780 26238
rect 73836 26292 73892 26302
rect 73612 26226 73668 26236
rect 73836 26198 73892 26236
rect 72492 25676 72772 25732
rect 73388 26066 73444 26078
rect 73388 26014 73390 26066
rect 73442 26014 73444 26066
rect 72044 25508 72100 25518
rect 72044 25414 72100 25452
rect 72492 25060 72548 25676
rect 72716 25506 72772 25518
rect 72716 25454 72718 25506
rect 72770 25454 72772 25506
rect 72492 24994 72548 25004
rect 72604 25394 72660 25406
rect 72604 25342 72606 25394
rect 72658 25342 72660 25394
rect 72604 24948 72660 25342
rect 72716 25396 72772 25454
rect 72772 25340 73108 25396
rect 72716 25330 72772 25340
rect 72604 24882 72660 24892
rect 71708 24742 71764 24780
rect 72716 24722 72772 24734
rect 72716 24670 72718 24722
rect 72770 24670 72772 24722
rect 72380 24612 72436 24622
rect 72716 24612 72772 24670
rect 71372 24434 71428 24444
rect 72268 24610 72772 24612
rect 72268 24558 72382 24610
rect 72434 24558 72772 24610
rect 72268 24556 72772 24558
rect 72268 23156 72324 24556
rect 72380 24546 72436 24556
rect 73052 24052 73108 25340
rect 73388 24724 73444 26014
rect 74060 25396 74116 26348
rect 74284 26292 74340 26572
rect 74508 26850 74564 26862
rect 74508 26798 74510 26850
rect 74562 26798 74564 26850
rect 74396 26292 74452 26302
rect 74284 26236 74396 26292
rect 74396 26226 74452 26236
rect 73836 25340 74116 25396
rect 74172 26178 74228 26190
rect 74172 26126 74174 26178
rect 74226 26126 74228 26178
rect 73836 24724 73892 25340
rect 74172 25060 74228 26126
rect 74172 24994 74228 25004
rect 74396 24948 74452 24958
rect 74284 24892 74396 24948
rect 73388 24658 73444 24668
rect 73612 24722 73892 24724
rect 73612 24670 73838 24722
rect 73890 24670 73892 24722
rect 73612 24668 73892 24670
rect 73052 23958 73108 23996
rect 73612 23938 73668 24668
rect 73836 24658 73892 24668
rect 74172 24836 74228 24846
rect 73612 23886 73614 23938
rect 73666 23886 73668 23938
rect 73612 23874 73668 23886
rect 74172 24052 74228 24780
rect 74284 24610 74340 24892
rect 74396 24882 74452 24892
rect 74284 24558 74286 24610
rect 74338 24558 74340 24610
rect 74284 24546 74340 24558
rect 74172 23826 74228 23996
rect 74508 23938 74564 26798
rect 74508 23886 74510 23938
rect 74562 23886 74564 23938
rect 74508 23874 74564 23886
rect 74172 23774 74174 23826
rect 74226 23774 74228 23826
rect 74172 23762 74228 23774
rect 72268 23090 72324 23100
rect 72492 23156 72548 23166
rect 72492 23062 72548 23100
rect 73052 23154 73108 23166
rect 73052 23102 73054 23154
rect 73106 23102 73108 23154
rect 73052 23044 73108 23102
rect 73052 22978 73108 22988
rect 74620 22932 74676 30940
rect 77196 29428 77252 55022
rect 77196 29362 77252 29372
rect 78652 28084 78708 55412
rect 81788 55412 82068 55468
rect 88396 55468 88452 56030
rect 88396 55412 88676 55468
rect 81564 55298 81620 55310
rect 81564 55246 81566 55298
rect 81618 55246 81620 55298
rect 81116 55188 81172 55198
rect 81116 55094 81172 55132
rect 81564 55188 81620 55246
rect 81564 55122 81620 55132
rect 81788 55186 81844 55412
rect 81788 55134 81790 55186
rect 81842 55134 81844 55186
rect 81788 55122 81844 55134
rect 88620 55074 88676 55412
rect 89404 55410 89460 56252
rect 89628 56242 89684 56252
rect 93212 56308 93268 59200
rect 93212 56242 93268 56252
rect 94444 56308 94500 56318
rect 94444 56214 94500 56252
rect 97020 56308 97076 59200
rect 97020 56242 97076 56252
rect 98252 56308 98308 56318
rect 98252 56214 98308 56252
rect 100828 56308 100884 59200
rect 101052 56308 101108 56318
rect 100828 56306 101108 56308
rect 100828 56254 101054 56306
rect 101106 56254 101108 56306
rect 100828 56252 101108 56254
rect 89964 56194 90020 56206
rect 89964 56142 89966 56194
rect 90018 56142 90020 56194
rect 89964 55468 90020 56142
rect 93436 56082 93492 56094
rect 93436 56030 93438 56082
rect 93490 56030 93492 56082
rect 93436 55468 93492 56030
rect 97580 56082 97636 56094
rect 97580 56030 97582 56082
rect 97634 56030 97636 56082
rect 96636 55692 96900 55702
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96636 55626 96900 55636
rect 89964 55412 90356 55468
rect 89404 55358 89406 55410
rect 89458 55358 89460 55410
rect 89404 55346 89460 55358
rect 88620 55022 88622 55074
rect 88674 55022 88676 55074
rect 81276 54908 81540 54918
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81276 54842 81540 54852
rect 81276 53340 81540 53350
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81276 53274 81540 53284
rect 81276 51772 81540 51782
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81276 51706 81540 51716
rect 81276 50204 81540 50214
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81276 50138 81540 50148
rect 81276 48636 81540 48646
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81276 48570 81540 48580
rect 81276 47068 81540 47078
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81276 47002 81540 47012
rect 81276 45500 81540 45510
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81276 45434 81540 45444
rect 81276 43932 81540 43942
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81276 43866 81540 43876
rect 88620 43708 88676 55022
rect 88620 43652 88900 43708
rect 81276 42364 81540 42374
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81276 42298 81540 42308
rect 81276 40796 81540 40806
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81276 40730 81540 40740
rect 81276 39228 81540 39238
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81276 39162 81540 39172
rect 81276 37660 81540 37670
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81276 37594 81540 37604
rect 81276 36092 81540 36102
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81276 36026 81540 36036
rect 81276 34524 81540 34534
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81276 34458 81540 34468
rect 81276 32956 81540 32966
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81276 32890 81540 32900
rect 81276 31388 81540 31398
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81276 31322 81540 31332
rect 81276 29820 81540 29830
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81276 29754 81540 29764
rect 83244 29428 83300 29438
rect 81276 28252 81540 28262
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81276 28186 81540 28196
rect 78204 28082 78708 28084
rect 78204 28030 78654 28082
rect 78706 28030 78708 28082
rect 78204 28028 78708 28030
rect 78204 27970 78260 28028
rect 78652 28018 78708 28028
rect 78204 27918 78206 27970
rect 78258 27918 78260 27970
rect 78204 27906 78260 27918
rect 77308 27860 77364 27870
rect 74732 27746 74788 27758
rect 74732 27694 74734 27746
rect 74786 27694 74788 27746
rect 74732 27188 74788 27694
rect 75852 27748 75908 27758
rect 75292 27412 75348 27422
rect 74732 27122 74788 27132
rect 75180 27188 75236 27198
rect 75180 27094 75236 27132
rect 74956 27074 75012 27086
rect 74956 27022 74958 27074
rect 75010 27022 75012 27074
rect 74956 26964 75012 27022
rect 74956 26898 75012 26908
rect 75292 27074 75348 27356
rect 75292 27022 75294 27074
rect 75346 27022 75348 27074
rect 75068 26852 75124 26862
rect 75124 26796 75236 26852
rect 75068 26786 75124 26796
rect 74732 26290 74788 26302
rect 74732 26238 74734 26290
rect 74786 26238 74788 26290
rect 74732 25506 74788 26238
rect 74732 25454 74734 25506
rect 74786 25454 74788 25506
rect 74732 25060 74788 25454
rect 74844 25732 74900 25742
rect 74844 25394 74900 25676
rect 74844 25342 74846 25394
rect 74898 25342 74900 25394
rect 74844 25330 74900 25342
rect 74732 25004 75012 25060
rect 74732 24948 74788 25004
rect 74732 24882 74788 24892
rect 74844 24836 74900 24846
rect 74844 24742 74900 24780
rect 74732 24724 74788 24734
rect 74732 24630 74788 24668
rect 74956 23938 75012 25004
rect 74956 23886 74958 23938
rect 75010 23886 75012 23938
rect 74956 23874 75012 23886
rect 75068 23716 75124 23726
rect 75068 23622 75124 23660
rect 74284 22876 74676 22932
rect 75180 22932 75236 26796
rect 75292 26514 75348 27022
rect 75516 27074 75572 27086
rect 75516 27022 75518 27074
rect 75570 27022 75572 27074
rect 75292 26462 75294 26514
rect 75346 26462 75348 26514
rect 75292 26450 75348 26462
rect 75404 26516 75460 26526
rect 75516 26516 75572 27022
rect 75852 26908 75908 27692
rect 77196 27636 77252 27646
rect 76188 27076 76244 27086
rect 76188 26982 76244 27020
rect 75852 26852 76132 26908
rect 75404 26514 75572 26516
rect 75404 26462 75406 26514
rect 75458 26462 75572 26514
rect 75404 26460 75572 26462
rect 75404 26450 75460 26460
rect 75740 26404 75796 26414
rect 75628 26402 75796 26404
rect 75628 26350 75742 26402
rect 75794 26350 75796 26402
rect 75628 26348 75796 26350
rect 75516 26292 75572 26302
rect 75516 26198 75572 26236
rect 75628 25284 75684 26348
rect 75740 26338 75796 26348
rect 75516 25228 75684 25284
rect 75292 24612 75348 24622
rect 75292 24518 75348 24556
rect 71260 22370 71316 22382
rect 71260 22318 71262 22370
rect 71314 22318 71316 22370
rect 69356 21756 69748 21812
rect 70476 22258 70532 22270
rect 70476 22206 70478 22258
rect 70530 22206 70532 22258
rect 68908 21422 68910 21474
rect 68962 21422 68964 21474
rect 68908 20244 68964 21422
rect 68908 20178 68964 20188
rect 69132 21700 69188 21710
rect 67900 20020 67956 20030
rect 67788 20018 67956 20020
rect 67788 19966 67902 20018
rect 67954 19966 67956 20018
rect 67788 19964 67956 19966
rect 67004 19842 67060 19852
rect 67116 19906 67172 19918
rect 67116 19854 67118 19906
rect 67170 19854 67172 19906
rect 67004 19236 67060 19246
rect 66892 19180 67004 19236
rect 67004 19142 67060 19180
rect 66556 19124 66612 19134
rect 66556 19030 66612 19068
rect 67116 19010 67172 19854
rect 67900 19908 67956 19964
rect 69132 20018 69188 21644
rect 69356 20132 69412 21756
rect 69468 21586 69524 21598
rect 69468 21534 69470 21586
rect 69522 21534 69524 21586
rect 69468 20356 69524 21534
rect 70476 21252 70532 22206
rect 71260 22148 71316 22318
rect 73836 22260 73892 22270
rect 71708 22148 71764 22158
rect 71260 22146 71764 22148
rect 71260 22094 71710 22146
rect 71762 22094 71764 22146
rect 71260 22092 71764 22094
rect 70476 21186 70532 21196
rect 71708 20804 71764 22092
rect 73836 21698 73892 22204
rect 73836 21646 73838 21698
rect 73890 21646 73892 21698
rect 73836 21634 73892 21646
rect 74172 21588 74228 21598
rect 74172 21494 74228 21532
rect 72828 21476 72884 21486
rect 72044 20804 72100 20814
rect 71708 20802 72100 20804
rect 71708 20750 72046 20802
rect 72098 20750 72100 20802
rect 71708 20748 72100 20750
rect 69468 20300 69748 20356
rect 69692 20244 69748 20300
rect 69692 20242 69860 20244
rect 69692 20190 69694 20242
rect 69746 20190 69860 20242
rect 69692 20188 69860 20190
rect 69692 20178 69748 20188
rect 69356 20076 69636 20132
rect 69132 19966 69134 20018
rect 69186 19966 69188 20018
rect 69132 19954 69188 19966
rect 68348 19908 68404 19918
rect 67900 19906 68628 19908
rect 67900 19854 68350 19906
rect 68402 19854 68628 19906
rect 67900 19852 68628 19854
rect 68348 19842 68404 19852
rect 67676 19796 67732 19806
rect 67564 19236 67620 19246
rect 67564 19142 67620 19180
rect 67116 18958 67118 19010
rect 67170 18958 67172 19010
rect 67116 18946 67172 18958
rect 66444 18498 66500 18508
rect 66780 18674 66836 18686
rect 66780 18622 66782 18674
rect 66834 18622 66836 18674
rect 66556 18452 66612 18462
rect 66556 18358 66612 18396
rect 65548 16884 65604 18060
rect 65916 18060 66180 18070
rect 65772 18004 65828 18014
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 65660 17668 65716 17678
rect 65660 17574 65716 17612
rect 65548 16818 65604 16828
rect 65772 17556 65828 17948
rect 65324 14802 65380 14812
rect 65324 14420 65380 14430
rect 65324 14326 65380 14364
rect 65548 14418 65604 14430
rect 65548 14366 65550 14418
rect 65602 14366 65604 14418
rect 65212 14254 65214 14306
rect 65266 14254 65268 14306
rect 65212 14242 65268 14254
rect 65548 13972 65604 14366
rect 65772 14420 65828 17500
rect 66220 16884 66276 16894
rect 66444 16884 66500 16894
rect 66220 16882 66500 16884
rect 66220 16830 66222 16882
rect 66274 16830 66446 16882
rect 66498 16830 66500 16882
rect 66220 16828 66500 16830
rect 66220 16818 66276 16828
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 66444 15988 66500 16828
rect 66444 15922 66500 15932
rect 66780 15148 66836 18622
rect 67340 18564 67396 18574
rect 67004 17554 67060 17566
rect 67004 17502 67006 17554
rect 67058 17502 67060 17554
rect 66668 15092 66724 15102
rect 66780 15092 66948 15148
rect 66332 14980 66388 14990
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 65884 14420 65940 14430
rect 65772 14418 65940 14420
rect 65772 14366 65886 14418
rect 65938 14366 65940 14418
rect 65772 14364 65940 14366
rect 65548 13906 65604 13916
rect 65772 14084 65828 14094
rect 65660 13860 65716 13870
rect 65660 13766 65716 13804
rect 65772 13858 65828 14028
rect 65772 13806 65774 13858
rect 65826 13806 65828 13858
rect 65772 13794 65828 13806
rect 64988 13746 65044 13758
rect 65436 13748 65492 13758
rect 64988 13694 64990 13746
rect 65042 13694 65044 13746
rect 64988 13634 65044 13694
rect 64988 13582 64990 13634
rect 65042 13582 65044 13634
rect 64988 13570 65044 13582
rect 65100 13746 65492 13748
rect 65100 13694 65438 13746
rect 65490 13694 65492 13746
rect 65100 13692 65492 13694
rect 64652 13132 64932 13188
rect 64652 12964 64708 13132
rect 64652 12908 65044 12964
rect 64540 12850 64596 12862
rect 64540 12798 64542 12850
rect 64594 12798 64596 12850
rect 64540 12404 64596 12798
rect 64876 12404 64932 12414
rect 64540 12402 64932 12404
rect 64540 12350 64878 12402
rect 64930 12350 64932 12402
rect 64540 12348 64932 12350
rect 64876 12338 64932 12348
rect 64652 12180 64708 12190
rect 64540 12178 64708 12180
rect 64540 12126 64654 12178
rect 64706 12126 64708 12178
rect 64540 12124 64708 12126
rect 64540 11954 64596 12124
rect 64652 12114 64708 12124
rect 64540 11902 64542 11954
rect 64594 11902 64596 11954
rect 64540 11890 64596 11902
rect 64876 11732 64932 11742
rect 64652 11618 64708 11630
rect 64652 11566 64654 11618
rect 64706 11566 64708 11618
rect 64540 11284 64596 11294
rect 64540 9940 64596 11228
rect 64652 10948 64708 11566
rect 64876 11506 64932 11676
rect 64988 11620 65044 12908
rect 65100 12290 65156 13692
rect 65436 13682 65492 13692
rect 65212 13524 65268 13534
rect 65884 13524 65940 14364
rect 66220 14306 66276 14318
rect 66220 14254 66222 14306
rect 66274 14254 66276 14306
rect 66220 13972 66276 14254
rect 66220 13906 66276 13916
rect 66332 13860 66388 14924
rect 66444 14420 66500 14430
rect 66444 14326 66500 14364
rect 66668 14418 66724 15036
rect 66668 14366 66670 14418
rect 66722 14366 66724 14418
rect 66668 14354 66724 14366
rect 66780 14418 66836 14430
rect 66780 14366 66782 14418
rect 66834 14366 66836 14418
rect 66668 14196 66724 14206
rect 66668 13970 66724 14140
rect 66668 13918 66670 13970
rect 66722 13918 66724 13970
rect 66668 13906 66724 13918
rect 66780 14084 66836 14366
rect 66220 13748 66276 13758
rect 66332 13748 66388 13804
rect 66220 13746 66612 13748
rect 66220 13694 66222 13746
rect 66274 13694 66612 13746
rect 66220 13692 66612 13694
rect 66220 13682 66276 13692
rect 65212 13522 65380 13524
rect 65212 13470 65214 13522
rect 65266 13470 65380 13522
rect 65212 13468 65380 13470
rect 65212 13458 65268 13468
rect 65100 12238 65102 12290
rect 65154 12238 65156 12290
rect 65100 12226 65156 12238
rect 64988 11554 65044 11564
rect 65212 12178 65268 12190
rect 65212 12126 65214 12178
rect 65266 12126 65268 12178
rect 64876 11454 64878 11506
rect 64930 11454 64932 11506
rect 64876 11442 64932 11454
rect 64652 10882 64708 10892
rect 64988 11284 65044 11294
rect 64876 10722 64932 10734
rect 64876 10670 64878 10722
rect 64930 10670 64932 10722
rect 64540 9874 64596 9884
rect 64652 10610 64708 10622
rect 64652 10558 64654 10610
rect 64706 10558 64708 10610
rect 64652 9042 64708 10558
rect 64876 10612 64932 10670
rect 64988 10722 65044 11228
rect 64988 10670 64990 10722
rect 65042 10670 65044 10722
rect 64988 10658 65044 10670
rect 65100 11172 65156 11182
rect 65212 11172 65268 12126
rect 65156 11116 65268 11172
rect 64876 10546 64932 10556
rect 64652 8990 64654 9042
rect 64706 8990 64708 9042
rect 64652 8978 64708 8990
rect 64764 9828 64820 9838
rect 64204 8764 64484 8820
rect 64540 8930 64596 8942
rect 64540 8878 64542 8930
rect 64594 8878 64596 8930
rect 64204 6916 64260 8764
rect 64540 8484 64596 8878
rect 64540 8418 64596 8428
rect 64764 8260 64820 9772
rect 64876 9602 64932 9614
rect 64876 9550 64878 9602
rect 64930 9550 64932 9602
rect 64876 9156 64932 9550
rect 64876 9090 64932 9100
rect 64988 9044 65044 9054
rect 65100 9044 65156 11116
rect 65324 9828 65380 13468
rect 65660 13468 65940 13524
rect 65436 11396 65492 11406
rect 65660 11396 65716 13468
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 66556 13076 66612 13692
rect 66668 13076 66724 13086
rect 66556 13074 66724 13076
rect 66556 13022 66670 13074
rect 66722 13022 66724 13074
rect 66556 13020 66724 13022
rect 66668 13010 66724 13020
rect 65996 12068 66052 12078
rect 65996 11974 66052 12012
rect 66780 11956 66836 14028
rect 66556 11900 66836 11956
rect 66892 11956 66948 15092
rect 67004 12852 67060 17502
rect 67340 16772 67396 18508
rect 67676 18562 67732 19740
rect 67676 18510 67678 18562
rect 67730 18510 67732 18562
rect 67676 18498 67732 18510
rect 68460 19346 68516 19358
rect 68460 19294 68462 19346
rect 68514 19294 68516 19346
rect 67340 16706 67396 16716
rect 67788 17444 67844 17454
rect 67340 15202 67396 15214
rect 67340 15150 67342 15202
rect 67394 15150 67396 15202
rect 67340 15092 67396 15150
rect 67340 15026 67396 15036
rect 67788 14756 67844 17388
rect 68460 17108 68516 19294
rect 68572 19236 68628 19852
rect 68572 19170 68628 19180
rect 69580 18676 69636 20076
rect 69020 18620 69636 18676
rect 69020 18450 69076 18620
rect 69020 18398 69022 18450
rect 69074 18398 69076 18450
rect 69020 18386 69076 18398
rect 69468 18452 69524 18462
rect 69468 18358 69524 18396
rect 69580 18450 69636 18620
rect 69580 18398 69582 18450
rect 69634 18398 69636 18450
rect 69580 18386 69636 18398
rect 69692 18450 69748 18462
rect 69692 18398 69694 18450
rect 69746 18398 69748 18450
rect 69692 17780 69748 18398
rect 69804 18340 69860 20188
rect 70364 20132 70420 20142
rect 70364 20130 70644 20132
rect 70364 20078 70366 20130
rect 70418 20078 70644 20130
rect 70364 20076 70644 20078
rect 70364 20066 70420 20076
rect 70140 20018 70196 20030
rect 70140 19966 70142 20018
rect 70194 19966 70196 20018
rect 69804 18274 69860 18284
rect 69916 19908 69972 19918
rect 69692 17714 69748 17724
rect 68908 17668 68964 17678
rect 68908 17574 68964 17612
rect 69356 17668 69412 17678
rect 68684 17556 68740 17566
rect 68684 17462 68740 17500
rect 69356 17554 69412 17612
rect 69356 17502 69358 17554
rect 69410 17502 69412 17554
rect 69356 17490 69412 17502
rect 69580 17666 69636 17678
rect 69580 17614 69582 17666
rect 69634 17614 69636 17666
rect 69580 17444 69636 17614
rect 69580 17378 69636 17388
rect 68460 17042 68516 17052
rect 68908 16996 68964 17006
rect 68908 16902 68964 16940
rect 68460 16100 68516 16110
rect 68460 16098 68852 16100
rect 68460 16046 68462 16098
rect 68514 16046 68852 16098
rect 68460 16044 68852 16046
rect 68460 16034 68516 16044
rect 68348 15988 68404 15998
rect 68348 15538 68404 15932
rect 68348 15486 68350 15538
rect 68402 15486 68404 15538
rect 68348 15474 68404 15486
rect 68012 15314 68068 15326
rect 68012 15262 68014 15314
rect 68066 15262 68068 15314
rect 68012 15204 68068 15262
rect 68460 15316 68516 15326
rect 68460 15222 68516 15260
rect 68684 15314 68740 15326
rect 68684 15262 68686 15314
rect 68738 15262 68740 15314
rect 68012 15138 68068 15148
rect 67788 14690 67844 14700
rect 68572 14306 68628 14318
rect 68572 14254 68574 14306
rect 68626 14254 68628 14306
rect 67228 13634 67284 13646
rect 67228 13582 67230 13634
rect 67282 13582 67284 13634
rect 67004 12786 67060 12796
rect 67116 13412 67172 13422
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 66332 11732 66388 11742
rect 66220 11508 66276 11518
rect 65884 11396 65940 11406
rect 65492 11340 65716 11396
rect 65772 11394 65940 11396
rect 65772 11342 65886 11394
rect 65938 11342 65940 11394
rect 65772 11340 65940 11342
rect 65436 11302 65492 11340
rect 65324 9762 65380 9772
rect 65436 10948 65492 10958
rect 65436 10610 65492 10892
rect 65436 10558 65438 10610
rect 65490 10558 65492 10610
rect 65212 9716 65268 9726
rect 65212 9156 65268 9660
rect 65212 9090 65268 9100
rect 65324 9602 65380 9614
rect 65324 9550 65326 9602
rect 65378 9550 65380 9602
rect 64988 9042 65156 9044
rect 64988 8990 64990 9042
rect 65042 8990 65156 9042
rect 64988 8988 65156 8990
rect 64764 8194 64820 8204
rect 64876 8932 64932 8942
rect 64764 7924 64820 7934
rect 64652 7868 64764 7924
rect 64428 7700 64484 7710
rect 64428 7606 64484 7644
rect 64204 6850 64260 6860
rect 64316 7588 64372 7598
rect 64316 6690 64372 7532
rect 64316 6638 64318 6690
rect 64370 6638 64372 6690
rect 64316 6626 64372 6638
rect 64652 7476 64708 7868
rect 64764 7858 64820 7868
rect 64092 5730 64148 5740
rect 64428 5906 64484 5918
rect 64428 5854 64430 5906
rect 64482 5854 64484 5906
rect 64428 5234 64484 5854
rect 64428 5182 64430 5234
rect 64482 5182 64484 5234
rect 64428 5170 64484 5182
rect 64652 5010 64708 7420
rect 64876 6804 64932 8876
rect 64988 8260 65044 8988
rect 65324 8820 65380 9550
rect 65436 9268 65492 10558
rect 65772 10052 65828 11340
rect 65884 11330 65940 11340
rect 66220 11170 66276 11452
rect 66332 11394 66388 11676
rect 66332 11342 66334 11394
rect 66386 11342 66388 11394
rect 66332 11330 66388 11342
rect 66444 11394 66500 11406
rect 66444 11342 66446 11394
rect 66498 11342 66500 11394
rect 66220 11118 66222 11170
rect 66274 11118 66276 11170
rect 66220 11106 66276 11118
rect 66444 11172 66500 11342
rect 66556 11284 66612 11900
rect 66892 11890 66948 11900
rect 67116 12068 67172 13356
rect 66668 11732 66724 11742
rect 66724 11676 67060 11732
rect 66668 11666 66724 11676
rect 67004 11618 67060 11676
rect 67004 11566 67006 11618
rect 67058 11566 67060 11618
rect 67004 11554 67060 11566
rect 66556 11218 66612 11228
rect 66892 11284 66948 11294
rect 66892 11190 66948 11228
rect 67004 11284 67060 11294
rect 67116 11284 67172 12012
rect 67004 11282 67172 11284
rect 67004 11230 67006 11282
rect 67058 11230 67172 11282
rect 67004 11228 67172 11230
rect 67004 11218 67060 11228
rect 66444 11106 66500 11116
rect 67228 10948 67284 13582
rect 67676 13636 67732 13646
rect 68124 13636 68180 13646
rect 67676 13634 67844 13636
rect 67676 13582 67678 13634
rect 67730 13582 67844 13634
rect 67676 13580 67844 13582
rect 67676 13570 67732 13580
rect 67564 12740 67620 12750
rect 67564 12738 67732 12740
rect 67564 12686 67566 12738
rect 67618 12686 67732 12738
rect 67564 12684 67732 12686
rect 67564 12674 67620 12684
rect 67564 11732 67620 11742
rect 67564 11060 67620 11676
rect 67228 10892 67396 10948
rect 66332 10836 66388 10846
rect 66108 10834 66388 10836
rect 66108 10782 66334 10834
rect 66386 10782 66388 10834
rect 66108 10780 66388 10782
rect 65884 10500 65940 10510
rect 66108 10500 66164 10780
rect 66332 10770 66388 10780
rect 67228 10724 67284 10734
rect 67228 10630 67284 10668
rect 66220 10612 66276 10622
rect 66276 10556 66388 10612
rect 66220 10546 66276 10556
rect 65884 10498 66164 10500
rect 65884 10446 65886 10498
rect 65938 10446 66164 10498
rect 65884 10444 66164 10446
rect 65884 10388 65940 10444
rect 65884 10322 65940 10332
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 65772 9996 66052 10052
rect 65436 9202 65492 9212
rect 65548 9602 65604 9614
rect 65548 9550 65550 9602
rect 65602 9550 65604 9602
rect 64988 8194 65044 8204
rect 65100 8764 65380 8820
rect 65436 9044 65492 9054
rect 65436 8930 65492 8988
rect 65436 8878 65438 8930
rect 65490 8878 65492 8930
rect 64988 7364 65044 7374
rect 65100 7364 65156 8764
rect 65324 8372 65380 8382
rect 65324 7698 65380 8316
rect 65324 7646 65326 7698
rect 65378 7646 65380 7698
rect 65324 7634 65380 7646
rect 64988 7362 65156 7364
rect 64988 7310 64990 7362
rect 65042 7310 65156 7362
rect 64988 7308 65156 7310
rect 64988 7298 65044 7308
rect 64764 6748 64932 6804
rect 64764 6244 64820 6748
rect 64764 6178 64820 6188
rect 64876 6578 64932 6590
rect 64876 6526 64878 6578
rect 64930 6526 64932 6578
rect 64652 4958 64654 5010
rect 64706 4958 64708 5010
rect 63756 4398 63758 4450
rect 63810 4398 63812 4450
rect 63756 4386 63812 4398
rect 64316 4676 64372 4686
rect 63084 2930 63140 2940
rect 63196 3332 63588 3388
rect 63196 980 63252 3332
rect 62972 924 63252 980
rect 62972 800 63028 924
rect 64316 800 64372 4620
rect 64540 4676 64596 4686
rect 64540 4562 64596 4620
rect 64540 4510 64542 4562
rect 64594 4510 64596 4562
rect 64540 4498 64596 4510
rect 64540 4340 64596 4350
rect 64652 4340 64708 4958
rect 64876 5796 64932 6526
rect 64988 6466 65044 6478
rect 64988 6414 64990 6466
rect 65042 6414 65044 6466
rect 64988 6018 65044 6414
rect 64988 5966 64990 6018
rect 65042 5966 65044 6018
rect 64988 5954 65044 5966
rect 64876 4452 64932 5740
rect 65100 5124 65156 7308
rect 65436 7476 65492 8878
rect 65548 8820 65604 9550
rect 65884 9268 65940 9278
rect 65548 8754 65604 8764
rect 65660 9266 65940 9268
rect 65660 9214 65886 9266
rect 65938 9214 65940 9266
rect 65660 9212 65940 9214
rect 65996 9268 66052 9996
rect 66108 10050 66164 10062
rect 66108 9998 66110 10050
rect 66162 9998 66164 10050
rect 66108 9938 66164 9998
rect 66108 9886 66110 9938
rect 66162 9886 66164 9938
rect 66108 9874 66164 9886
rect 66332 9380 66388 10556
rect 66556 10610 66612 10622
rect 66556 10558 66558 10610
rect 66610 10558 66612 10610
rect 66444 9602 66500 9614
rect 66444 9550 66446 9602
rect 66498 9550 66500 9602
rect 66444 9492 66500 9550
rect 66444 9426 66500 9436
rect 66220 9324 66388 9380
rect 66108 9268 66164 9278
rect 65996 9266 66164 9268
rect 65996 9214 66110 9266
rect 66162 9214 66164 9266
rect 65996 9212 66164 9214
rect 65660 7924 65716 9212
rect 65884 9202 65940 9212
rect 66108 9202 66164 9212
rect 65660 7858 65716 7868
rect 65772 9044 65828 9054
rect 65660 7700 65716 7710
rect 65772 7700 65828 8988
rect 66220 8820 66276 9324
rect 66444 9154 66500 9166
rect 66444 9102 66446 9154
rect 66498 9102 66500 9154
rect 66332 9044 66388 9054
rect 66332 8950 66388 8988
rect 66220 8764 66388 8820
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 66332 8484 66388 8764
rect 66108 8428 66388 8484
rect 66108 8370 66164 8428
rect 66108 8318 66110 8370
rect 66162 8318 66164 8370
rect 66108 8306 66164 8318
rect 65660 7698 65828 7700
rect 65660 7646 65662 7698
rect 65714 7646 65828 7698
rect 65660 7644 65828 7646
rect 66332 8258 66388 8270
rect 66332 8206 66334 8258
rect 66386 8206 66388 8258
rect 66332 7700 66388 8206
rect 66444 7924 66500 9102
rect 66556 8370 66612 10558
rect 67004 10498 67060 10510
rect 67004 10446 67006 10498
rect 67058 10446 67060 10498
rect 67004 10164 67060 10446
rect 67004 10098 67060 10108
rect 67228 10388 67284 10398
rect 66668 9716 66724 9726
rect 66668 9266 66724 9660
rect 67004 9602 67060 9614
rect 67004 9550 67006 9602
rect 67058 9550 67060 9602
rect 67004 9380 67060 9550
rect 67004 9314 67060 9324
rect 67116 9604 67172 9614
rect 66668 9214 66670 9266
rect 66722 9214 66724 9266
rect 66668 9202 66724 9214
rect 66556 8318 66558 8370
rect 66610 8318 66612 8370
rect 66556 8306 66612 8318
rect 66892 9156 66948 9166
rect 66668 8260 66724 8270
rect 66668 8166 66724 8204
rect 66892 8036 66948 9100
rect 67004 8260 67060 8270
rect 67116 8260 67172 9548
rect 67228 9044 67284 10332
rect 67340 9380 67396 10892
rect 67564 10610 67620 11004
rect 67564 10558 67566 10610
rect 67618 10558 67620 10610
rect 67564 10546 67620 10558
rect 67452 9828 67508 9838
rect 67452 9734 67508 9772
rect 67340 9324 67620 9380
rect 67340 9156 67396 9166
rect 67340 9154 67508 9156
rect 67340 9102 67342 9154
rect 67394 9102 67508 9154
rect 67340 9100 67508 9102
rect 67340 9090 67396 9100
rect 67228 8978 67284 8988
rect 67004 8258 67172 8260
rect 67004 8206 67006 8258
rect 67058 8206 67172 8258
rect 67004 8204 67172 8206
rect 67228 8820 67284 8830
rect 67228 8258 67284 8764
rect 67228 8206 67230 8258
rect 67282 8206 67284 8258
rect 67004 8194 67060 8204
rect 67228 8194 67284 8206
rect 67340 8818 67396 8830
rect 67340 8766 67342 8818
rect 67394 8766 67396 8818
rect 66892 7980 67060 8036
rect 66444 7858 66500 7868
rect 66556 7700 66612 7710
rect 66332 7698 66612 7700
rect 66332 7646 66558 7698
rect 66610 7646 66612 7698
rect 66332 7644 66612 7646
rect 65660 7634 65716 7644
rect 65436 6916 65492 7420
rect 66220 7364 66276 7374
rect 66220 7270 66276 7308
rect 66332 7252 66388 7644
rect 66556 7634 66612 7644
rect 66668 7588 66724 7598
rect 66444 7476 66500 7486
rect 66668 7476 66724 7532
rect 66444 7474 66724 7476
rect 66444 7422 66446 7474
rect 66498 7422 66724 7474
rect 66444 7420 66724 7422
rect 66444 7410 66500 7420
rect 66332 7196 66500 7252
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 65436 6850 65492 6860
rect 66332 6580 66388 6590
rect 66332 6020 66388 6524
rect 66332 5954 66388 5964
rect 65548 5794 65604 5806
rect 65548 5742 65550 5794
rect 65602 5742 65604 5794
rect 65212 5124 65268 5134
rect 65100 5068 65212 5124
rect 65212 5058 65268 5068
rect 65548 4564 65604 5742
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 65772 5122 65828 5134
rect 65772 5070 65774 5122
rect 65826 5070 65828 5122
rect 65772 5012 65828 5070
rect 65772 4946 65828 4956
rect 65548 4498 65604 4508
rect 65100 4452 65156 4462
rect 64876 4450 65156 4452
rect 64876 4398 65102 4450
rect 65154 4398 65156 4450
rect 64876 4396 65156 4398
rect 65100 4386 65156 4396
rect 64540 4338 64708 4340
rect 64540 4286 64542 4338
rect 64594 4286 64708 4338
rect 64540 4284 64708 4286
rect 64540 4274 64596 4284
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 65884 3780 65940 3790
rect 64876 3668 64932 3678
rect 64876 3574 64932 3612
rect 65660 3668 65716 3678
rect 65660 800 65716 3612
rect 65884 3554 65940 3724
rect 66444 3666 66500 7196
rect 66556 7250 66612 7262
rect 66556 7198 66558 7250
rect 66610 7198 66612 7250
rect 66556 6690 66612 7198
rect 66668 7252 66724 7420
rect 66668 7186 66724 7196
rect 66556 6638 66558 6690
rect 66610 6638 66612 6690
rect 66556 6626 66612 6638
rect 66892 6580 66948 6590
rect 66892 6486 66948 6524
rect 66780 6466 66836 6478
rect 66780 6414 66782 6466
rect 66834 6414 66836 6466
rect 66780 6132 66836 6414
rect 66780 6076 66948 6132
rect 66780 5906 66836 5918
rect 66780 5854 66782 5906
rect 66834 5854 66836 5906
rect 66780 5348 66836 5854
rect 66780 5282 66836 5292
rect 66556 5012 66612 5022
rect 66556 4338 66612 4956
rect 66556 4286 66558 4338
rect 66610 4286 66612 4338
rect 66556 4274 66612 4286
rect 66444 3614 66446 3666
rect 66498 3614 66500 3666
rect 66444 3602 66500 3614
rect 66892 3668 66948 6076
rect 66892 3602 66948 3612
rect 65884 3502 65886 3554
rect 65938 3502 65940 3554
rect 65884 3490 65940 3502
rect 67004 800 67060 7980
rect 67116 8034 67172 8046
rect 67116 7982 67118 8034
rect 67170 7982 67172 8034
rect 67116 7700 67172 7982
rect 67116 7634 67172 7644
rect 67228 7924 67284 7934
rect 67116 7476 67172 7486
rect 67116 5796 67172 7420
rect 67116 5730 67172 5740
rect 67228 6690 67284 7868
rect 67228 6638 67230 6690
rect 67282 6638 67284 6690
rect 67228 5012 67284 6638
rect 67340 5906 67396 8766
rect 67452 8596 67508 9100
rect 67452 8530 67508 8540
rect 67452 8372 67508 8382
rect 67452 8258 67508 8316
rect 67452 8206 67454 8258
rect 67506 8206 67508 8258
rect 67452 8194 67508 8206
rect 67452 8036 67508 8046
rect 67452 6356 67508 7980
rect 67564 6692 67620 9324
rect 67676 9156 67732 12684
rect 67788 11172 67844 13580
rect 68012 13634 68180 13636
rect 68012 13582 68126 13634
rect 68178 13582 68180 13634
rect 68012 13580 68180 13582
rect 67788 10388 67844 11116
rect 67900 11170 67956 11182
rect 67900 11118 67902 11170
rect 67954 11118 67956 11170
rect 67900 11060 67956 11118
rect 67900 10994 67956 11004
rect 68012 10948 68068 13580
rect 68124 13570 68180 13580
rect 68124 12066 68180 12078
rect 68124 12014 68126 12066
rect 68178 12014 68180 12066
rect 68124 11508 68180 12014
rect 68572 11732 68628 14254
rect 68684 13972 68740 15262
rect 68796 15148 68852 16044
rect 69132 15988 69188 15998
rect 69132 15894 69188 15932
rect 69692 15540 69748 15550
rect 69692 15446 69748 15484
rect 69132 15204 69188 15242
rect 69916 15148 69972 19852
rect 70140 18674 70196 19966
rect 70588 19346 70644 20076
rect 70588 19294 70590 19346
rect 70642 19294 70644 19346
rect 70588 19282 70644 19294
rect 71260 19460 71316 19470
rect 70140 18622 70142 18674
rect 70194 18622 70196 18674
rect 70140 18610 70196 18622
rect 70700 18452 70756 18462
rect 70700 18358 70756 18396
rect 71260 17780 71316 19404
rect 71932 19346 71988 19358
rect 71932 19294 71934 19346
rect 71986 19294 71988 19346
rect 71372 19236 71428 19246
rect 71372 18340 71428 19180
rect 71932 18564 71988 19294
rect 72044 19236 72100 20748
rect 72828 20802 72884 21420
rect 73948 21476 74004 21486
rect 73948 21382 74004 21420
rect 72828 20750 72830 20802
rect 72882 20750 72884 20802
rect 72828 20738 72884 20750
rect 73948 21252 74004 21262
rect 72940 20244 72996 20254
rect 72044 19170 72100 19180
rect 72828 20188 72940 20244
rect 71932 18498 71988 18508
rect 71596 18340 71652 18350
rect 71372 18338 71652 18340
rect 71372 18286 71598 18338
rect 71650 18286 71652 18338
rect 71372 18284 71652 18286
rect 71372 17780 71428 17790
rect 71260 17778 71428 17780
rect 71260 17726 71374 17778
rect 71426 17726 71428 17778
rect 71260 17724 71428 17726
rect 71372 17714 71428 17724
rect 68796 15092 69076 15148
rect 69132 15138 69188 15148
rect 69020 14644 69076 15092
rect 69020 14530 69076 14588
rect 69020 14478 69022 14530
rect 69074 14478 69076 14530
rect 69020 14466 69076 14478
rect 69804 15092 69972 15148
rect 70028 17666 70084 17678
rect 70028 17614 70030 17666
rect 70082 17614 70084 17666
rect 69692 14420 69748 14430
rect 69468 14418 69748 14420
rect 69468 14366 69694 14418
rect 69746 14366 69748 14418
rect 69468 14364 69748 14366
rect 68684 13906 68740 13916
rect 68908 14308 68964 14318
rect 68908 13970 68964 14252
rect 68908 13918 68910 13970
rect 68962 13918 68964 13970
rect 68796 13300 68852 13310
rect 68796 13074 68852 13244
rect 68796 13022 68798 13074
rect 68850 13022 68852 13074
rect 68796 13010 68852 13022
rect 68908 12404 68964 13918
rect 69468 13970 69524 14364
rect 69692 14354 69748 14364
rect 69804 14196 69860 15092
rect 70028 14756 70084 17614
rect 70476 17668 70532 17678
rect 70476 17574 70532 17612
rect 70924 17668 70980 17678
rect 70924 17574 70980 17612
rect 71596 16996 71652 18284
rect 72268 18340 72324 18350
rect 72268 18004 72324 18284
rect 72268 17778 72324 17948
rect 72268 17726 72270 17778
rect 72322 17726 72324 17778
rect 72268 17714 72324 17726
rect 71820 17668 71876 17678
rect 71820 17574 71876 17612
rect 72716 17554 72772 17566
rect 72716 17502 72718 17554
rect 72770 17502 72772 17554
rect 72492 17444 72548 17454
rect 72716 17444 72772 17502
rect 72548 17388 72772 17444
rect 72492 17378 72548 17388
rect 71596 16930 71652 16940
rect 72492 16996 72548 17006
rect 72492 16884 72548 16940
rect 72380 16882 72548 16884
rect 72380 16830 72494 16882
rect 72546 16830 72548 16882
rect 72380 16828 72548 16830
rect 72044 16660 72100 16670
rect 71260 16212 71316 16222
rect 70924 16210 71316 16212
rect 70924 16158 71262 16210
rect 71314 16158 71316 16210
rect 70924 16156 71316 16158
rect 70588 15764 70644 15774
rect 70140 15652 70196 15662
rect 70140 15538 70196 15596
rect 70140 15486 70142 15538
rect 70194 15486 70196 15538
rect 70140 15474 70196 15486
rect 70588 15202 70644 15708
rect 70812 15652 70868 15662
rect 70700 15316 70756 15326
rect 70700 15222 70756 15260
rect 70588 15150 70590 15202
rect 70642 15150 70644 15202
rect 70588 15138 70644 15150
rect 70028 14690 70084 14700
rect 69468 13918 69470 13970
rect 69522 13918 69524 13970
rect 69468 13906 69524 13918
rect 69692 14140 69860 14196
rect 69132 13746 69188 13758
rect 69132 13694 69134 13746
rect 69186 13694 69188 13746
rect 69132 13188 69188 13694
rect 69580 13748 69636 13758
rect 69580 13654 69636 13692
rect 69132 13122 69188 13132
rect 69132 12738 69188 12750
rect 69132 12686 69134 12738
rect 69186 12686 69188 12738
rect 68908 12348 69076 12404
rect 68124 11442 68180 11452
rect 68236 11676 68628 11732
rect 68908 12178 68964 12190
rect 68908 12126 68910 12178
rect 68962 12126 68964 12178
rect 67788 10322 67844 10332
rect 67900 10724 67956 10734
rect 67900 10050 67956 10668
rect 67900 9998 67902 10050
rect 67954 9998 67956 10050
rect 67900 9986 67956 9998
rect 67788 9940 67844 9950
rect 67788 9846 67844 9884
rect 67900 9156 67956 9166
rect 67676 9100 67900 9156
rect 67900 9062 67956 9100
rect 67788 8260 67844 8270
rect 68012 8260 68068 10892
rect 67788 8258 68068 8260
rect 67788 8206 67790 8258
rect 67842 8206 68068 8258
rect 67788 8204 68068 8206
rect 68236 8260 68292 11676
rect 68908 11618 68964 12126
rect 68908 11566 68910 11618
rect 68962 11566 68964 11618
rect 68348 11508 68404 11518
rect 68348 10612 68404 11452
rect 68572 11172 68628 11182
rect 68572 11170 68852 11172
rect 68572 11118 68574 11170
rect 68626 11118 68852 11170
rect 68572 11116 68852 11118
rect 68572 11106 68628 11116
rect 68348 10546 68404 10556
rect 68572 10500 68628 10510
rect 68572 10406 68628 10444
rect 68460 9604 68516 9614
rect 67788 8194 67844 8204
rect 68236 8194 68292 8204
rect 68348 9602 68516 9604
rect 68348 9550 68462 9602
rect 68514 9550 68516 9602
rect 68348 9548 68516 9550
rect 67676 8034 67732 8046
rect 67676 7982 67678 8034
rect 67730 7982 67732 8034
rect 67676 6804 67732 7982
rect 68236 8034 68292 8046
rect 68236 7982 68238 8034
rect 68290 7982 68292 8034
rect 67788 7700 67844 7710
rect 67788 7586 67844 7644
rect 67788 7534 67790 7586
rect 67842 7534 67844 7586
rect 67788 7522 67844 7534
rect 68236 7252 68292 7982
rect 67676 6738 67732 6748
rect 67788 7196 68292 7252
rect 67564 6626 67620 6636
rect 67788 6690 67844 7196
rect 67788 6638 67790 6690
rect 67842 6638 67844 6690
rect 67788 6626 67844 6638
rect 68236 6692 68292 6702
rect 67452 6300 67732 6356
rect 67340 5854 67342 5906
rect 67394 5854 67396 5906
rect 67340 5842 67396 5854
rect 67564 5908 67620 5918
rect 67564 5814 67620 5852
rect 67676 5906 67732 6300
rect 68012 6020 68068 6030
rect 68012 5926 68068 5964
rect 67676 5854 67678 5906
rect 67730 5854 67732 5906
rect 67676 5842 67732 5854
rect 67788 5124 67844 5134
rect 67228 4946 67284 4956
rect 67676 5012 67732 5022
rect 67676 4918 67732 4956
rect 67676 4452 67732 4462
rect 67788 4452 67844 5068
rect 67676 4450 67844 4452
rect 67676 4398 67678 4450
rect 67730 4398 67844 4450
rect 67676 4396 67844 4398
rect 67676 4386 67732 4396
rect 68236 3388 68292 6636
rect 68348 5908 68404 9548
rect 68460 9538 68516 9548
rect 68684 8932 68740 8942
rect 68460 8596 68516 8606
rect 68516 8540 68628 8596
rect 68460 8530 68516 8540
rect 68460 6468 68516 6478
rect 68460 6132 68516 6412
rect 68460 6066 68516 6076
rect 68460 5908 68516 5918
rect 68348 5906 68516 5908
rect 68348 5854 68462 5906
rect 68514 5854 68516 5906
rect 68348 5852 68516 5854
rect 68460 5796 68516 5852
rect 68460 5730 68516 5740
rect 68460 5348 68516 5358
rect 68460 5254 68516 5292
rect 68572 4562 68628 8540
rect 68684 6468 68740 8876
rect 68796 6580 68852 11116
rect 68908 10610 68964 11566
rect 69020 11396 69076 12348
rect 69132 12068 69188 12686
rect 69692 12628 69748 14140
rect 69804 13972 69860 13982
rect 70812 13972 70868 15596
rect 70924 15426 70980 16156
rect 71260 16146 71316 16156
rect 72044 16210 72100 16604
rect 72044 16158 72046 16210
rect 72098 16158 72100 16210
rect 72044 16146 72100 16158
rect 70924 15374 70926 15426
rect 70978 15374 70980 15426
rect 70924 15316 70980 15374
rect 71260 15540 71316 15550
rect 70924 15250 70980 15260
rect 71036 15314 71092 15326
rect 71036 15262 71038 15314
rect 71090 15262 71092 15314
rect 71036 15148 71092 15262
rect 71260 15148 71316 15484
rect 71484 15540 71540 15550
rect 71484 15446 71540 15484
rect 72380 15540 72436 16828
rect 72492 16818 72548 16828
rect 72492 16212 72548 16222
rect 72604 16212 72660 17388
rect 72492 16210 72660 16212
rect 72492 16158 72494 16210
rect 72546 16158 72660 16210
rect 72492 16156 72660 16158
rect 72492 16146 72548 16156
rect 71036 15092 71204 15148
rect 71260 15092 71540 15148
rect 69804 13746 69860 13916
rect 69804 13694 69806 13746
rect 69858 13694 69860 13746
rect 69804 12740 69860 13694
rect 70700 13970 70868 13972
rect 70700 13918 70814 13970
rect 70866 13918 70868 13970
rect 70700 13916 70868 13918
rect 70364 13636 70420 13646
rect 70364 13634 70644 13636
rect 70364 13582 70366 13634
rect 70418 13582 70644 13634
rect 70364 13580 70644 13582
rect 70364 13570 70420 13580
rect 70252 13524 70308 13534
rect 69916 12964 69972 12974
rect 69916 12962 70084 12964
rect 69916 12910 69918 12962
rect 69970 12910 70084 12962
rect 69916 12908 70084 12910
rect 69916 12898 69972 12908
rect 69804 12684 69972 12740
rect 69692 12562 69748 12572
rect 69916 12178 69972 12684
rect 69916 12126 69918 12178
rect 69970 12126 69972 12178
rect 69916 12114 69972 12126
rect 69580 12068 69636 12078
rect 69132 12066 69636 12068
rect 69132 12014 69582 12066
rect 69634 12014 69636 12066
rect 69132 12012 69636 12014
rect 69132 11618 69188 12012
rect 69580 11956 69636 12012
rect 70028 11956 70084 12908
rect 69580 11900 70084 11956
rect 69132 11566 69134 11618
rect 69186 11566 69188 11618
rect 69132 11554 69188 11566
rect 69020 11340 69300 11396
rect 69020 11172 69076 11182
rect 69020 11078 69076 11116
rect 68908 10558 68910 10610
rect 68962 10558 68964 10610
rect 68908 10546 68964 10558
rect 69020 9602 69076 9614
rect 69020 9550 69022 9602
rect 69074 9550 69076 9602
rect 69020 8484 69076 9550
rect 69132 9604 69188 9614
rect 69132 9510 69188 9548
rect 69244 9156 69300 11340
rect 70028 11284 70084 11900
rect 70140 12628 70196 12638
rect 70140 11620 70196 12572
rect 70252 12178 70308 13468
rect 70588 13076 70644 13580
rect 70588 13010 70644 13020
rect 70588 12852 70644 12862
rect 70364 12850 70644 12852
rect 70364 12798 70590 12850
rect 70642 12798 70644 12850
rect 70364 12796 70644 12798
rect 70364 12402 70420 12796
rect 70588 12786 70644 12796
rect 70364 12350 70366 12402
rect 70418 12350 70420 12402
rect 70364 12338 70420 12350
rect 70252 12126 70254 12178
rect 70306 12126 70308 12178
rect 70252 12114 70308 12126
rect 70476 12180 70532 12190
rect 70476 12086 70532 12124
rect 70140 11564 70308 11620
rect 70140 11396 70196 11406
rect 70140 11302 70196 11340
rect 70028 11218 70084 11228
rect 69356 11170 69412 11182
rect 69356 11118 69358 11170
rect 69410 11118 69412 11170
rect 69356 10948 69412 11118
rect 69804 11170 69860 11182
rect 69804 11118 69806 11170
rect 69858 11118 69860 11170
rect 69356 10882 69412 10892
rect 69468 11060 69524 11070
rect 69468 10164 69524 11004
rect 69804 10948 69860 11118
rect 70252 11060 70308 11564
rect 70476 11172 70532 11182
rect 70476 11170 70644 11172
rect 70476 11118 70478 11170
rect 70530 11118 70644 11170
rect 70476 11116 70644 11118
rect 70476 11106 70532 11116
rect 70252 10994 70308 11004
rect 69804 10882 69860 10892
rect 69580 10500 69636 10510
rect 69580 10498 70308 10500
rect 69580 10446 69582 10498
rect 69634 10446 70308 10498
rect 69580 10444 70308 10446
rect 69580 10434 69636 10444
rect 69356 10108 69524 10164
rect 70028 10164 70084 10174
rect 69356 9714 69412 10108
rect 69356 9662 69358 9714
rect 69410 9662 69412 9714
rect 69356 9380 69412 9662
rect 69468 9714 69524 9726
rect 69468 9662 69470 9714
rect 69522 9662 69524 9714
rect 69468 9604 69524 9662
rect 69468 9538 69524 9548
rect 69356 9324 69972 9380
rect 69244 9100 69412 9156
rect 69020 8418 69076 8428
rect 69244 8930 69300 8942
rect 69244 8878 69246 8930
rect 69298 8878 69300 8930
rect 68908 8148 68964 8158
rect 68908 6802 68964 8092
rect 69244 8148 69300 8878
rect 69244 8082 69300 8092
rect 68908 6750 68910 6802
rect 68962 6750 68964 6802
rect 68908 6738 68964 6750
rect 69356 6690 69412 9100
rect 69580 8932 69636 8942
rect 69580 8838 69636 8876
rect 69916 7362 69972 9324
rect 69916 7310 69918 7362
rect 69970 7310 69972 7362
rect 69916 7298 69972 7310
rect 69916 6916 69972 6926
rect 70028 6916 70084 10108
rect 70252 9938 70308 10444
rect 70252 9886 70254 9938
rect 70306 9886 70308 9938
rect 70252 9874 70308 9886
rect 70588 9940 70644 11116
rect 70588 9826 70644 9884
rect 70588 9774 70590 9826
rect 70642 9774 70644 9826
rect 70588 9762 70644 9774
rect 70140 9716 70196 9726
rect 70140 9622 70196 9660
rect 70476 9716 70532 9726
rect 70476 9622 70532 9660
rect 70588 9154 70644 9166
rect 70588 9102 70590 9154
rect 70642 9102 70644 9154
rect 70364 8148 70420 8158
rect 70364 8054 70420 8092
rect 70476 7364 70532 7374
rect 70476 7270 70532 7308
rect 70588 6916 70644 9102
rect 70028 6860 70308 6916
rect 69916 6802 69972 6860
rect 69916 6750 69918 6802
rect 69970 6750 69972 6802
rect 69916 6738 69972 6750
rect 69356 6638 69358 6690
rect 69410 6638 69412 6690
rect 68796 6524 68964 6580
rect 68684 6412 68852 6468
rect 68684 5124 68740 5134
rect 68684 5030 68740 5068
rect 68572 4510 68574 4562
rect 68626 4510 68628 4562
rect 68572 4498 68628 4510
rect 68796 4338 68852 6412
rect 68908 4788 68964 6524
rect 69132 5908 69188 5918
rect 69132 5814 69188 5852
rect 69244 5796 69300 5806
rect 69020 5124 69076 5134
rect 69020 5030 69076 5068
rect 68908 4722 68964 4732
rect 68796 4286 68798 4338
rect 68850 4286 68852 4338
rect 68796 4274 68852 4286
rect 69244 4340 69300 5740
rect 68572 3668 68628 3678
rect 68572 3574 68628 3612
rect 69244 3554 69300 4284
rect 69244 3502 69246 3554
rect 69298 3502 69300 3554
rect 69244 3490 69300 3502
rect 69356 5460 69412 6638
rect 69356 3388 69412 5404
rect 69468 5348 69524 5358
rect 69468 5234 69524 5292
rect 69468 5182 69470 5234
rect 69522 5182 69524 5234
rect 69468 5170 69524 5182
rect 69468 4788 69524 4798
rect 69468 4450 69524 4732
rect 69468 4398 69470 4450
rect 69522 4398 69524 4450
rect 69468 4386 69524 4398
rect 69692 3668 69748 3678
rect 68236 3332 68404 3388
rect 69356 3332 69524 3388
rect 68348 800 68404 3332
rect 69468 3220 69524 3332
rect 69468 3154 69524 3164
rect 69692 800 69748 3612
rect 70252 2436 70308 6860
rect 70588 6850 70644 6860
rect 70700 6356 70756 13916
rect 70812 13906 70868 13916
rect 71036 13748 71092 13758
rect 71148 13748 71204 15092
rect 71260 13972 71316 13982
rect 71260 13878 71316 13916
rect 71372 13748 71428 13758
rect 71148 13746 71428 13748
rect 71148 13694 71374 13746
rect 71426 13694 71428 13746
rect 71148 13692 71428 13694
rect 71036 13654 71092 13692
rect 71372 13636 71428 13692
rect 71372 13570 71428 13580
rect 71260 12068 71316 12078
rect 71484 12068 71540 15092
rect 71820 14642 71876 14654
rect 71820 14590 71822 14642
rect 71874 14590 71876 14642
rect 71820 13972 71876 14590
rect 72380 14644 72436 15484
rect 72492 15428 72548 15438
rect 72492 15334 72548 15372
rect 72828 14644 72884 20188
rect 72940 20178 72996 20188
rect 73164 19908 73220 19918
rect 73612 19908 73668 19918
rect 73164 19906 73668 19908
rect 73164 19854 73166 19906
rect 73218 19854 73614 19906
rect 73666 19854 73668 19906
rect 73164 19852 73668 19854
rect 72940 19122 72996 19134
rect 72940 19070 72942 19122
rect 72994 19070 72996 19122
rect 72940 19012 72996 19070
rect 73164 19012 73220 19852
rect 73612 19842 73668 19852
rect 73948 19572 74004 21196
rect 74172 20580 74228 20590
rect 74060 20524 74172 20580
rect 74060 20130 74116 20524
rect 74172 20514 74228 20524
rect 74060 20078 74062 20130
rect 74114 20078 74116 20130
rect 74060 20066 74116 20078
rect 74284 20132 74340 22876
rect 75180 22866 75236 22876
rect 75404 23042 75460 23054
rect 75404 22990 75406 23042
rect 75458 22990 75460 23042
rect 74620 22708 74676 22718
rect 74620 22482 74676 22652
rect 75404 22596 75460 22990
rect 74620 22430 74622 22482
rect 74674 22430 74676 22482
rect 74620 22418 74676 22430
rect 74956 22540 75460 22596
rect 74732 22372 74788 22382
rect 74956 22372 75012 22540
rect 75516 22484 75572 25228
rect 75628 24948 75684 24958
rect 75628 24722 75684 24892
rect 75628 24670 75630 24722
rect 75682 24670 75684 24722
rect 75628 24658 75684 24670
rect 75628 23940 75684 23950
rect 75628 23846 75684 23884
rect 76076 23940 76132 26852
rect 77196 26290 77252 27580
rect 77196 26238 77198 26290
rect 77250 26238 77252 26290
rect 77196 26226 77252 26238
rect 77308 27076 77364 27804
rect 77644 27858 77700 27870
rect 77644 27806 77646 27858
rect 77698 27806 77700 27858
rect 77644 27636 77700 27806
rect 77644 27570 77700 27580
rect 77756 27746 77812 27758
rect 77756 27694 77758 27746
rect 77810 27694 77812 27746
rect 76860 26180 76916 26190
rect 76860 26086 76916 26124
rect 77308 25506 77364 27020
rect 77756 26908 77812 27694
rect 78540 27188 78596 27198
rect 78540 27074 78596 27132
rect 78540 27022 78542 27074
rect 78594 27022 78596 27074
rect 78540 27010 78596 27022
rect 78876 27076 78932 27086
rect 79100 27076 79156 27086
rect 79660 27076 79716 27086
rect 78932 27074 79716 27076
rect 78932 27022 79102 27074
rect 79154 27022 79662 27074
rect 79714 27022 79716 27074
rect 78932 27020 79716 27022
rect 78876 27010 78932 27020
rect 79100 27010 79156 27020
rect 77308 25454 77310 25506
rect 77362 25454 77364 25506
rect 77308 25442 77364 25454
rect 77420 26852 77812 26908
rect 76524 25060 76580 25070
rect 76524 24948 76580 25004
rect 76524 24946 76804 24948
rect 76524 24894 76526 24946
rect 76578 24894 76804 24946
rect 76524 24892 76804 24894
rect 76524 24882 76580 24892
rect 74732 22370 75012 22372
rect 74732 22318 74734 22370
rect 74786 22318 75012 22370
rect 74732 22316 75012 22318
rect 75180 22428 75572 22484
rect 75628 23156 75684 23166
rect 75628 22484 75684 23100
rect 75740 23154 75796 23166
rect 75740 23102 75742 23154
rect 75794 23102 75796 23154
rect 75740 22708 75796 23102
rect 76076 23154 76132 23884
rect 76748 23938 76804 24892
rect 76860 24834 76916 24846
rect 76860 24782 76862 24834
rect 76914 24782 76916 24834
rect 76860 24724 76916 24782
rect 76860 24658 76916 24668
rect 76748 23886 76750 23938
rect 76802 23886 76804 23938
rect 76748 23874 76804 23886
rect 76524 23714 76580 23726
rect 76524 23662 76526 23714
rect 76578 23662 76580 23714
rect 76076 23102 76078 23154
rect 76130 23102 76132 23154
rect 76076 23090 76132 23102
rect 76300 23156 76356 23166
rect 76524 23156 76580 23662
rect 76300 23154 76524 23156
rect 76300 23102 76302 23154
rect 76354 23102 76524 23154
rect 76300 23100 76524 23102
rect 76188 23044 76244 23054
rect 76188 22950 76244 22988
rect 75740 22642 75796 22652
rect 75180 22370 75236 22428
rect 75180 22318 75182 22370
rect 75234 22318 75236 22370
rect 74508 22148 74564 22158
rect 74396 21586 74452 21598
rect 74396 21534 74398 21586
rect 74450 21534 74452 21586
rect 74396 20356 74452 21534
rect 74396 20290 74452 20300
rect 74284 20076 74452 20132
rect 74172 19796 74228 19806
rect 74172 19702 74228 19740
rect 73948 19516 74228 19572
rect 73724 19346 73780 19358
rect 73724 19294 73726 19346
rect 73778 19294 73780 19346
rect 73724 19124 73780 19294
rect 73276 19012 73332 19022
rect 72940 19010 73332 19012
rect 72940 18958 73278 19010
rect 73330 18958 73332 19010
rect 72940 18956 73332 18958
rect 72940 18226 72996 18956
rect 73276 18946 73332 18956
rect 72940 18174 72942 18226
rect 72994 18174 72996 18226
rect 72940 18116 72996 18174
rect 72940 18050 72996 18060
rect 73276 18450 73332 18462
rect 73276 18398 73278 18450
rect 73330 18398 73332 18450
rect 73276 18228 73332 18398
rect 73724 18452 73780 19068
rect 73724 18386 73780 18396
rect 74060 18450 74116 18462
rect 74060 18398 74062 18450
rect 74114 18398 74116 18450
rect 73052 17780 73108 17790
rect 73276 17780 73332 18172
rect 73052 17778 73332 17780
rect 73052 17726 73054 17778
rect 73106 17726 73332 17778
rect 73052 17724 73332 17726
rect 73052 17714 73108 17724
rect 73724 17444 73780 17454
rect 74060 17444 74116 18398
rect 74172 18450 74228 19516
rect 74284 19348 74340 19358
rect 74396 19348 74452 20076
rect 74508 20018 74564 22092
rect 74732 21700 74788 22316
rect 75180 22306 75236 22318
rect 74732 21634 74788 21644
rect 74956 21700 75012 21710
rect 74956 21586 75012 21644
rect 74956 21534 74958 21586
rect 75010 21534 75012 21586
rect 74956 21522 75012 21534
rect 74844 21362 74900 21374
rect 74844 21310 74846 21362
rect 74898 21310 74900 21362
rect 74732 20580 74788 20590
rect 74732 20242 74788 20524
rect 74732 20190 74734 20242
rect 74786 20190 74788 20242
rect 74732 20178 74788 20190
rect 74844 20244 74900 21310
rect 75180 20580 75236 20590
rect 75180 20486 75236 20524
rect 74844 20178 74900 20188
rect 74620 20132 74676 20142
rect 74620 20038 74676 20076
rect 74508 19966 74510 20018
rect 74562 19966 74564 20018
rect 74508 19954 74564 19966
rect 75180 20020 75236 20030
rect 75292 20020 75348 22428
rect 75628 22390 75684 22428
rect 76300 22260 76356 23100
rect 76524 23062 76580 23100
rect 76300 22194 76356 22204
rect 76412 22484 76468 22494
rect 76412 21812 76468 22428
rect 75404 21588 75460 21598
rect 75404 21474 75460 21532
rect 76412 21586 76468 21756
rect 76412 21534 76414 21586
rect 76466 21534 76468 21586
rect 76412 21522 76468 21534
rect 77196 21586 77252 21598
rect 77196 21534 77198 21586
rect 77250 21534 77252 21586
rect 75404 21422 75406 21474
rect 75458 21422 75460 21474
rect 75404 20692 75460 21422
rect 75404 20626 75460 20636
rect 75516 21252 75572 21262
rect 75404 20020 75460 20030
rect 75180 20018 75460 20020
rect 75180 19966 75182 20018
rect 75234 19966 75406 20018
rect 75458 19966 75460 20018
rect 75180 19964 75460 19966
rect 75180 19954 75236 19964
rect 74284 19346 74452 19348
rect 74284 19294 74286 19346
rect 74338 19294 74452 19346
rect 74284 19292 74452 19294
rect 74284 19282 74340 19292
rect 74396 19124 74452 19292
rect 74172 18398 74174 18450
rect 74226 18398 74228 18450
rect 74172 18386 74228 18398
rect 74284 18450 74340 18462
rect 74284 18398 74286 18450
rect 74338 18398 74340 18450
rect 74172 17444 74228 17454
rect 74060 17442 74228 17444
rect 74060 17390 74174 17442
rect 74226 17390 74228 17442
rect 74060 17388 74228 17390
rect 73164 16770 73220 16782
rect 73164 16718 73166 16770
rect 73218 16718 73220 16770
rect 73164 16210 73220 16718
rect 73612 16772 73668 16782
rect 73164 16158 73166 16210
rect 73218 16158 73220 16210
rect 73164 16146 73220 16158
rect 73276 16660 73332 16670
rect 73276 16098 73332 16604
rect 73276 16046 73278 16098
rect 73330 16046 73332 16098
rect 73276 16034 73332 16046
rect 73612 16098 73668 16716
rect 73612 16046 73614 16098
rect 73666 16046 73668 16098
rect 73612 16034 73668 16046
rect 73052 15988 73108 15998
rect 72940 15764 72996 15774
rect 72940 15148 72996 15708
rect 73052 15428 73108 15932
rect 73724 15764 73780 17388
rect 74172 17332 74228 17388
rect 74284 17444 74340 18398
rect 74284 17378 74340 17388
rect 74172 16212 74228 17276
rect 74284 16212 74340 16222
rect 74172 16210 74340 16212
rect 74172 16158 74286 16210
rect 74338 16158 74340 16210
rect 74172 16156 74340 16158
rect 74172 15988 74228 16156
rect 74284 16146 74340 16156
rect 74172 15922 74228 15932
rect 73836 15764 73892 15774
rect 73724 15708 73836 15764
rect 73836 15538 73892 15708
rect 73836 15486 73838 15538
rect 73890 15486 73892 15538
rect 73836 15474 73892 15486
rect 74284 15428 74340 15438
rect 73052 15362 73108 15372
rect 74060 15372 74284 15428
rect 73164 15202 73220 15214
rect 74060 15204 74116 15372
rect 74284 15334 74340 15372
rect 73164 15150 73166 15202
rect 73218 15150 73220 15202
rect 72940 15092 73108 15148
rect 72940 14644 72996 14654
rect 72828 14642 72996 14644
rect 72828 14590 72942 14642
rect 72994 14590 72996 14642
rect 72828 14588 72996 14590
rect 72380 14550 72436 14588
rect 72492 14532 72548 14542
rect 72492 14438 72548 14476
rect 71820 13906 71876 13916
rect 72380 13972 72436 13982
rect 72380 13970 72660 13972
rect 72380 13918 72382 13970
rect 72434 13918 72660 13970
rect 72380 13916 72660 13918
rect 72380 13906 72436 13916
rect 72492 13746 72548 13758
rect 72492 13694 72494 13746
rect 72546 13694 72548 13746
rect 72492 13636 72548 13694
rect 72492 13570 72548 13580
rect 72380 13524 72436 13534
rect 72380 13430 72436 13468
rect 72604 13076 72660 13916
rect 72940 13860 72996 14588
rect 72940 13794 72996 13804
rect 72940 13634 72996 13646
rect 72940 13582 72942 13634
rect 72994 13582 72996 13634
rect 72716 13076 72772 13086
rect 72604 13074 72772 13076
rect 72604 13022 72718 13074
rect 72770 13022 72772 13074
rect 72604 13020 72772 13022
rect 72716 12180 72772 13020
rect 72716 12114 72772 12124
rect 72828 12516 72884 12526
rect 71260 12066 71540 12068
rect 71260 12014 71262 12066
rect 71314 12014 71540 12066
rect 71260 12012 71540 12014
rect 71708 12066 71764 12078
rect 71708 12014 71710 12066
rect 71762 12014 71764 12066
rect 71260 12002 71316 12012
rect 71036 11620 71092 11630
rect 71036 11506 71092 11564
rect 71036 11454 71038 11506
rect 71090 11454 71092 11506
rect 71036 11442 71092 11454
rect 70924 11172 70980 11182
rect 71260 11172 71316 11182
rect 70812 11116 70924 11172
rect 70812 7140 70868 11116
rect 70924 11106 70980 11116
rect 71148 11170 71316 11172
rect 71148 11118 71262 11170
rect 71314 11118 71316 11170
rect 71148 11116 71316 11118
rect 71148 10612 71204 11116
rect 71260 11106 71316 11116
rect 71372 11060 71428 12012
rect 71596 11396 71652 11406
rect 71596 11302 71652 11340
rect 71484 11172 71540 11182
rect 71484 11078 71540 11116
rect 71708 11172 71764 12014
rect 72380 12066 72436 12078
rect 72380 12014 72382 12066
rect 72434 12014 72436 12066
rect 71932 11956 71988 11966
rect 71708 11106 71764 11116
rect 71820 11900 71932 11956
rect 71372 10724 71428 11004
rect 71372 10658 71428 10668
rect 71820 10612 71876 11900
rect 71932 11890 71988 11900
rect 72380 11954 72436 12014
rect 72380 11902 72382 11954
rect 72434 11902 72436 11954
rect 72156 11396 72212 11406
rect 71932 11282 71988 11294
rect 71932 11230 71934 11282
rect 71986 11230 71988 11282
rect 71932 11172 71988 11230
rect 71932 10948 71988 11116
rect 71932 10882 71988 10892
rect 72044 11170 72100 11182
rect 72044 11118 72046 11170
rect 72098 11118 72100 11170
rect 71036 10556 71204 10612
rect 71484 10556 71876 10612
rect 70924 9716 70980 9726
rect 70924 9622 70980 9660
rect 71036 8036 71092 10556
rect 71484 10500 71540 10556
rect 71148 10444 71540 10500
rect 71708 10498 71764 10556
rect 71708 10446 71710 10498
rect 71762 10446 71764 10498
rect 71148 9714 71204 10444
rect 71708 10434 71764 10446
rect 72044 9940 72100 11118
rect 71820 9884 72100 9940
rect 71148 9662 71150 9714
rect 71202 9662 71204 9714
rect 71148 9650 71204 9662
rect 71260 9714 71316 9726
rect 71260 9662 71262 9714
rect 71314 9662 71316 9714
rect 71260 9604 71316 9662
rect 71148 9492 71204 9502
rect 71148 9044 71204 9436
rect 71260 9268 71316 9548
rect 71708 9602 71764 9614
rect 71708 9550 71710 9602
rect 71762 9550 71764 9602
rect 71708 9492 71764 9550
rect 71708 9426 71764 9436
rect 71260 9202 71316 9212
rect 71708 9268 71764 9278
rect 71708 9174 71764 9212
rect 71372 9044 71428 9054
rect 71148 9042 71428 9044
rect 71148 8990 71374 9042
rect 71426 8990 71428 9042
rect 71148 8988 71428 8990
rect 71372 8978 71428 8988
rect 71708 8372 71764 8382
rect 71820 8372 71876 9884
rect 72156 9828 72212 11340
rect 72380 11284 72436 11902
rect 72828 12066 72884 12460
rect 72828 12014 72830 12066
rect 72882 12014 72884 12066
rect 72828 11396 72884 12014
rect 72940 11954 72996 13582
rect 72940 11902 72942 11954
rect 72994 11902 72996 11954
rect 72940 11890 72996 11902
rect 73052 11620 73108 15092
rect 73164 11956 73220 15150
rect 73836 15148 74116 15204
rect 74396 15148 74452 19068
rect 75292 19124 75348 19134
rect 75404 19124 75460 19964
rect 75516 19348 75572 21196
rect 77196 20916 77252 21534
rect 77420 21588 77476 26852
rect 77756 26290 77812 26302
rect 77756 26238 77758 26290
rect 77810 26238 77812 26290
rect 77756 26180 77812 26238
rect 77756 26114 77812 26124
rect 78092 25508 78148 25518
rect 78092 25506 78708 25508
rect 78092 25454 78094 25506
rect 78146 25454 78708 25506
rect 78092 25452 78708 25454
rect 78092 25442 78148 25452
rect 78428 24948 78484 24958
rect 78428 24854 78484 24892
rect 78204 24724 78260 24734
rect 78204 23604 78260 24668
rect 77868 23548 78260 23604
rect 78316 24610 78372 24622
rect 78316 24558 78318 24610
rect 78370 24558 78372 24610
rect 77532 23156 77588 23166
rect 77588 23100 77700 23156
rect 77532 23090 77588 23100
rect 77420 21522 77476 21532
rect 77532 20916 77588 20926
rect 77196 20914 77588 20916
rect 77196 20862 77534 20914
rect 77586 20862 77588 20914
rect 77196 20860 77588 20862
rect 77532 20850 77588 20860
rect 77084 20804 77140 20814
rect 77084 20710 77140 20748
rect 77420 20692 77476 20702
rect 77644 20692 77700 23100
rect 77868 22148 77924 23548
rect 78316 23268 78372 24558
rect 78316 23202 78372 23212
rect 78540 23938 78596 23950
rect 78540 23886 78542 23938
rect 78594 23886 78596 23938
rect 78428 23156 78484 23166
rect 78428 23062 78484 23100
rect 77756 20916 77812 20926
rect 77756 20802 77812 20860
rect 77756 20750 77758 20802
rect 77810 20750 77812 20802
rect 77756 20738 77812 20750
rect 77420 20690 77700 20692
rect 77420 20638 77422 20690
rect 77474 20638 77700 20690
rect 77420 20636 77700 20638
rect 77420 20626 77476 20636
rect 75628 20580 75684 20590
rect 75628 20578 75796 20580
rect 75628 20526 75630 20578
rect 75682 20526 75796 20578
rect 75628 20524 75796 20526
rect 75628 20514 75684 20524
rect 75516 19292 75684 19348
rect 75516 19124 75572 19134
rect 75404 19122 75572 19124
rect 75404 19070 75518 19122
rect 75570 19070 75572 19122
rect 75404 19068 75572 19070
rect 75292 19030 75348 19068
rect 75516 19058 75572 19068
rect 74844 19012 74900 19022
rect 74844 18918 74900 18956
rect 75068 19012 75124 19022
rect 75068 18918 75124 18956
rect 75180 19010 75236 19022
rect 75180 18958 75182 19010
rect 75234 18958 75236 19010
rect 75180 18788 75236 18958
rect 75628 18900 75684 19292
rect 74620 18732 75236 18788
rect 75404 18844 75684 18900
rect 74620 18562 74676 18732
rect 74620 18510 74622 18562
rect 74674 18510 74676 18562
rect 74620 18498 74676 18510
rect 74956 18228 75012 18238
rect 74844 18172 74956 18228
rect 74844 16324 74900 18172
rect 74956 18162 75012 18172
rect 75292 16770 75348 16782
rect 75292 16718 75294 16770
rect 75346 16718 75348 16770
rect 75292 16324 75348 16718
rect 74844 16268 75236 16324
rect 74844 16098 74900 16268
rect 74844 16046 74846 16098
rect 74898 16046 74900 16098
rect 74844 16034 74900 16046
rect 75068 16098 75124 16110
rect 75068 16046 75070 16098
rect 75122 16046 75124 16098
rect 74956 15988 75012 15998
rect 75068 15988 75124 16046
rect 75180 16100 75236 16268
rect 75292 16258 75348 16268
rect 75292 16100 75348 16110
rect 75180 16098 75348 16100
rect 75180 16046 75294 16098
rect 75346 16046 75348 16098
rect 75180 16044 75348 16046
rect 75292 16034 75348 16044
rect 75012 15932 75124 15988
rect 74956 15922 75012 15932
rect 75180 15876 75236 15914
rect 75180 15810 75236 15820
rect 75404 15540 75460 18844
rect 75740 18452 75796 20524
rect 76524 20578 76580 20590
rect 76524 20526 76526 20578
rect 76578 20526 76580 20578
rect 75964 20020 76020 20030
rect 76300 20020 76356 20030
rect 76524 20020 76580 20526
rect 77868 20468 77924 22092
rect 78540 21700 78596 23886
rect 78652 23378 78708 25452
rect 79660 25284 79716 27020
rect 81276 26684 81540 26694
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81276 26618 81540 26628
rect 79660 25218 79716 25228
rect 80444 25282 80500 25294
rect 80444 25230 80446 25282
rect 80498 25230 80500 25282
rect 79100 24948 79156 24958
rect 78652 23326 78654 23378
rect 78706 23326 78708 23378
rect 78652 23314 78708 23326
rect 78764 24722 78820 24734
rect 78764 24670 78766 24722
rect 78818 24670 78820 24722
rect 78540 21644 78708 21700
rect 78540 21476 78596 21486
rect 77980 20972 78484 21028
rect 77980 20802 78036 20972
rect 78428 20914 78484 20972
rect 78428 20862 78430 20914
rect 78482 20862 78484 20914
rect 78428 20850 78484 20862
rect 77980 20750 77982 20802
rect 78034 20750 78036 20802
rect 77980 20738 78036 20750
rect 78540 20802 78596 21420
rect 78540 20750 78542 20802
rect 78594 20750 78596 20802
rect 77868 20402 77924 20412
rect 78092 20580 78148 20590
rect 75964 20018 76524 20020
rect 75964 19966 75966 20018
rect 76018 19966 76302 20018
rect 76354 19966 76524 20018
rect 75964 19964 76524 19966
rect 75628 18338 75684 18350
rect 75628 18286 75630 18338
rect 75682 18286 75684 18338
rect 74844 15484 75460 15540
rect 75516 17108 75572 17118
rect 73724 15092 73892 15148
rect 74172 15092 74452 15148
rect 74620 15204 74676 15214
rect 74732 15202 74788 15214
rect 74732 15150 74734 15202
rect 74786 15150 74788 15202
rect 74732 15148 74788 15150
rect 74620 15092 74788 15148
rect 73500 14754 73556 14766
rect 73500 14702 73502 14754
rect 73554 14702 73556 14754
rect 73276 14308 73332 14318
rect 73276 12738 73332 14252
rect 73388 14306 73444 14318
rect 73388 14254 73390 14306
rect 73442 14254 73444 14306
rect 73388 13522 73444 14254
rect 73500 13970 73556 14702
rect 73500 13918 73502 13970
rect 73554 13918 73556 13970
rect 73500 13906 73556 13918
rect 73388 13470 73390 13522
rect 73442 13470 73444 13522
rect 73388 13458 73444 13470
rect 73724 13300 73780 15092
rect 73948 14308 74004 14318
rect 73948 14306 74116 14308
rect 73948 14254 73950 14306
rect 74002 14254 74116 14306
rect 73948 14252 74116 14254
rect 73948 14242 74004 14252
rect 73948 13634 74004 13646
rect 73948 13582 73950 13634
rect 74002 13582 74004 13634
rect 73724 13234 73780 13244
rect 73836 13522 73892 13534
rect 73836 13470 73838 13522
rect 73890 13470 73892 13522
rect 73276 12686 73278 12738
rect 73330 12686 73332 12738
rect 73276 12628 73332 12686
rect 73724 12738 73780 12750
rect 73724 12686 73726 12738
rect 73778 12686 73780 12738
rect 73276 12572 73556 12628
rect 73388 12066 73444 12078
rect 73388 12014 73390 12066
rect 73442 12014 73444 12066
rect 73164 11900 73332 11956
rect 73052 11564 73220 11620
rect 73052 11396 73108 11406
rect 72828 11340 72996 11396
rect 72380 11218 72436 11228
rect 72716 11282 72772 11294
rect 72716 11230 72718 11282
rect 72770 11230 72772 11282
rect 72044 9772 72212 9828
rect 72268 11170 72324 11182
rect 72268 11118 72270 11170
rect 72322 11118 72324 11170
rect 72044 9714 72100 9772
rect 72044 9662 72046 9714
rect 72098 9662 72100 9714
rect 71596 8370 71876 8372
rect 71596 8318 71710 8370
rect 71762 8318 71876 8370
rect 71596 8316 71876 8318
rect 71932 8484 71988 8494
rect 71036 7970 71092 7980
rect 71148 8034 71204 8046
rect 71148 7982 71150 8034
rect 71202 7982 71204 8034
rect 71148 7364 71204 7982
rect 71484 7586 71540 7598
rect 71484 7534 71486 7586
rect 71538 7534 71540 7586
rect 71148 7298 71204 7308
rect 71260 7476 71316 7486
rect 71260 7140 71316 7420
rect 70812 7084 71316 7140
rect 70700 5236 70756 6300
rect 70700 5170 70756 5180
rect 71148 6916 71204 6926
rect 71148 5012 71204 6860
rect 71260 5794 71316 7084
rect 71260 5742 71262 5794
rect 71314 5742 71316 5794
rect 71260 5730 71316 5742
rect 71148 4918 71204 4956
rect 70700 4898 70756 4910
rect 70700 4846 70702 4898
rect 70754 4846 70756 4898
rect 70476 3668 70532 3678
rect 70476 3574 70532 3612
rect 70700 2884 70756 4846
rect 70700 2818 70756 2828
rect 71036 4788 71092 4798
rect 70252 2370 70308 2380
rect 71036 800 71092 4732
rect 71484 4226 71540 7534
rect 71596 5124 71652 8316
rect 71708 8306 71764 8316
rect 71708 6692 71764 6702
rect 71708 6578 71764 6636
rect 71708 6526 71710 6578
rect 71762 6526 71764 6578
rect 71708 6514 71764 6526
rect 71820 6132 71876 6142
rect 71932 6132 71988 8428
rect 72044 7252 72100 9662
rect 72156 9604 72212 9614
rect 72156 7700 72212 9548
rect 72268 8596 72324 11118
rect 72716 11172 72772 11230
rect 72716 11106 72772 11116
rect 72828 11170 72884 11182
rect 72828 11118 72830 11170
rect 72882 11118 72884 11170
rect 72828 11060 72884 11118
rect 72492 10612 72548 10622
rect 72492 10518 72548 10556
rect 72716 10610 72772 10622
rect 72716 10558 72718 10610
rect 72770 10558 72772 10610
rect 72716 10500 72772 10558
rect 72716 10434 72772 10444
rect 72604 9714 72660 9726
rect 72604 9662 72606 9714
rect 72658 9662 72660 9714
rect 72268 8530 72324 8540
rect 72380 9602 72436 9614
rect 72380 9550 72382 9602
rect 72434 9550 72436 9602
rect 72380 8428 72436 9550
rect 72492 9492 72548 9502
rect 72492 9266 72548 9436
rect 72492 9214 72494 9266
rect 72546 9214 72548 9266
rect 72492 9202 72548 9214
rect 72604 9268 72660 9662
rect 72716 9604 72772 9614
rect 72716 9510 72772 9548
rect 72604 9202 72660 9212
rect 72716 9380 72772 9390
rect 72716 9042 72772 9324
rect 72716 8990 72718 9042
rect 72770 8990 72772 9042
rect 72716 8978 72772 8990
rect 72828 8708 72884 11004
rect 72940 10052 72996 11340
rect 73052 11302 73108 11340
rect 73164 10164 73220 11564
rect 73276 11618 73332 11900
rect 73388 11844 73444 12014
rect 73388 11778 73444 11788
rect 73276 11566 73278 11618
rect 73330 11566 73332 11618
rect 73276 11554 73332 11566
rect 73500 11620 73556 12572
rect 73724 12516 73780 12686
rect 73724 12402 73780 12460
rect 73724 12350 73726 12402
rect 73778 12350 73780 12402
rect 73724 12338 73780 12350
rect 73500 11554 73556 11564
rect 73836 11508 73892 13470
rect 73612 11452 73892 11508
rect 73948 12740 74004 13582
rect 74060 12852 74116 14252
rect 74172 13076 74228 15092
rect 74732 15026 74788 15036
rect 74284 14980 74340 14990
rect 74284 14532 74340 14924
rect 74284 14466 74340 14476
rect 74396 14754 74452 14766
rect 74396 14702 74398 14754
rect 74450 14702 74452 14754
rect 74284 14308 74340 14318
rect 74284 14214 74340 14252
rect 74396 13634 74452 14702
rect 74844 14532 74900 15484
rect 74732 14476 74900 14532
rect 74956 15316 75012 15326
rect 74732 14084 74788 14476
rect 74844 14308 74900 14318
rect 74844 14214 74900 14252
rect 74732 14028 74900 14084
rect 74396 13582 74398 13634
rect 74450 13582 74452 13634
rect 74396 13524 74452 13582
rect 74396 13458 74452 13468
rect 74732 13860 74788 13870
rect 74172 12982 74228 13020
rect 74508 12852 74564 12862
rect 74060 12796 74228 12852
rect 73164 10098 73220 10108
rect 73276 11394 73332 11406
rect 73276 11342 73278 11394
rect 73330 11342 73332 11394
rect 73276 10498 73332 11342
rect 73276 10446 73278 10498
rect 73330 10446 73332 10498
rect 73276 10052 73332 10446
rect 73612 11170 73668 11452
rect 73612 11118 73614 11170
rect 73666 11118 73668 11170
rect 73612 10500 73668 11118
rect 73724 11284 73780 11294
rect 73724 10610 73780 11228
rect 73948 11172 74004 12684
rect 73948 11170 74116 11172
rect 73948 11118 73950 11170
rect 74002 11118 74116 11170
rect 73948 11116 74116 11118
rect 73948 11106 74004 11116
rect 73724 10558 73726 10610
rect 73778 10558 73780 10610
rect 73724 10546 73780 10558
rect 73612 10434 73668 10444
rect 73276 9996 74004 10052
rect 72940 9986 72996 9996
rect 73052 9884 73444 9940
rect 72940 9828 72996 9838
rect 73052 9828 73108 9884
rect 72940 9826 73108 9828
rect 72940 9774 72942 9826
rect 72994 9774 73108 9826
rect 72940 9772 73108 9774
rect 73388 9826 73444 9884
rect 73388 9774 73390 9826
rect 73442 9774 73444 9826
rect 72940 9762 72996 9772
rect 73388 9762 73444 9774
rect 73724 9828 73780 9838
rect 73780 9772 73892 9828
rect 73724 9734 73780 9772
rect 73164 9714 73220 9726
rect 73164 9662 73166 9714
rect 73218 9662 73220 9714
rect 73164 9380 73220 9662
rect 73276 9716 73332 9726
rect 73276 9622 73332 9660
rect 73164 9324 73332 9380
rect 72828 8642 72884 8652
rect 72940 9044 72996 9054
rect 72380 8372 72884 8428
rect 72268 8260 72324 8270
rect 72492 8260 72548 8270
rect 72268 8258 72436 8260
rect 72268 8206 72270 8258
rect 72322 8206 72436 8258
rect 72268 8204 72436 8206
rect 72268 8194 72324 8204
rect 72156 7634 72212 7644
rect 72268 7588 72324 7598
rect 72268 7494 72324 7532
rect 72380 7476 72436 8204
rect 72380 7410 72436 7420
rect 72044 7186 72100 7196
rect 72492 6804 72548 8204
rect 72828 8148 72884 8372
rect 72940 8370 72996 8988
rect 73052 9042 73108 9054
rect 73052 8990 73054 9042
rect 73106 8990 73108 9042
rect 73052 8596 73108 8990
rect 73276 8932 73332 9324
rect 73388 9268 73444 9278
rect 73388 9266 73556 9268
rect 73388 9214 73390 9266
rect 73442 9214 73556 9266
rect 73388 9212 73556 9214
rect 73388 9202 73444 9212
rect 73500 9156 73556 9212
rect 73724 9156 73780 9166
rect 73836 9156 73892 9772
rect 73500 9100 73668 9156
rect 73388 9044 73444 9054
rect 73612 9044 73668 9100
rect 73724 9154 73892 9156
rect 73724 9102 73726 9154
rect 73778 9102 73892 9154
rect 73724 9100 73892 9102
rect 73948 9268 74004 9996
rect 74060 9380 74116 11116
rect 74060 9314 74116 9324
rect 74172 9714 74228 12796
rect 74508 12740 74564 12796
rect 74620 12740 74676 12750
rect 74508 12738 74676 12740
rect 74508 12686 74622 12738
rect 74674 12686 74676 12738
rect 74508 12684 74676 12686
rect 74620 12674 74676 12684
rect 74508 12180 74564 12190
rect 74508 12086 74564 12124
rect 74172 9662 74174 9714
rect 74226 9662 74228 9714
rect 73724 9090 73780 9100
rect 73388 9042 73556 9044
rect 73388 8990 73390 9042
rect 73442 8990 73556 9042
rect 73388 8988 73556 8990
rect 73388 8978 73444 8988
rect 73052 8530 73108 8540
rect 73164 8876 73332 8932
rect 72940 8318 72942 8370
rect 72994 8318 72996 8370
rect 72940 8306 72996 8318
rect 73164 8372 73220 8876
rect 73164 8306 73220 8316
rect 73500 8372 73556 8988
rect 73612 8978 73668 8988
rect 73500 8306 73556 8316
rect 73612 8708 73668 8718
rect 72828 8092 73220 8148
rect 72604 7588 72660 7598
rect 72604 7586 72772 7588
rect 72604 7534 72606 7586
rect 72658 7534 72772 7586
rect 72604 7532 72772 7534
rect 72604 7522 72660 7532
rect 72492 6738 72548 6748
rect 72604 7252 72660 7262
rect 72268 6580 72324 6590
rect 72492 6580 72548 6590
rect 72604 6580 72660 7196
rect 72324 6524 72436 6580
rect 72268 6514 72324 6524
rect 71820 6130 71988 6132
rect 71820 6078 71822 6130
rect 71874 6078 71988 6130
rect 71820 6076 71988 6078
rect 72044 6356 72100 6366
rect 71820 6066 71876 6076
rect 71596 5030 71652 5068
rect 72044 5684 72100 6300
rect 72044 5122 72100 5628
rect 72044 5070 72046 5122
rect 72098 5070 72100 5122
rect 72044 5058 72100 5070
rect 72268 6356 72324 6366
rect 72268 5906 72324 6300
rect 72380 6132 72436 6524
rect 72492 6578 72660 6580
rect 72492 6526 72494 6578
rect 72546 6526 72660 6578
rect 72492 6524 72660 6526
rect 72492 6514 72548 6524
rect 72380 6076 72548 6132
rect 72268 5854 72270 5906
rect 72322 5854 72324 5906
rect 72268 5124 72324 5854
rect 72268 5058 72324 5068
rect 72380 5908 72436 5918
rect 71484 4174 71486 4226
rect 71538 4174 71540 4226
rect 71484 4162 71540 4174
rect 72380 3554 72436 5852
rect 72492 4562 72548 6076
rect 72604 5348 72660 5358
rect 72604 5010 72660 5292
rect 72604 4958 72606 5010
rect 72658 4958 72660 5010
rect 72604 4946 72660 4958
rect 72716 5012 72772 7532
rect 73164 7586 73220 8092
rect 73612 7700 73668 8652
rect 73948 7700 74004 9212
rect 73164 7534 73166 7586
rect 73218 7534 73220 7586
rect 73164 7522 73220 7534
rect 73276 7644 73668 7700
rect 73724 7644 74004 7700
rect 74060 8930 74116 8942
rect 74060 8878 74062 8930
rect 74114 8878 74116 8930
rect 72828 7476 72884 7486
rect 72828 7140 72884 7420
rect 72828 7074 72884 7084
rect 72940 7474 72996 7486
rect 72940 7422 72942 7474
rect 72994 7422 72996 7474
rect 72828 6580 72884 6590
rect 72828 6486 72884 6524
rect 72940 6020 72996 7422
rect 73276 7364 73332 7644
rect 73612 7474 73668 7486
rect 73612 7422 73614 7474
rect 73666 7422 73668 7474
rect 72940 5954 72996 5964
rect 73052 7308 73332 7364
rect 73388 7364 73444 7374
rect 73388 7362 73556 7364
rect 73388 7310 73390 7362
rect 73442 7310 73556 7362
rect 73388 7308 73556 7310
rect 73052 5348 73108 7308
rect 73388 7298 73444 7308
rect 73052 5282 73108 5292
rect 73164 7140 73220 7150
rect 72716 4946 72772 4956
rect 72492 4510 72494 4562
rect 72546 4510 72548 4562
rect 72492 4498 72548 4510
rect 72716 4564 72772 4574
rect 72716 4562 73108 4564
rect 72716 4510 72718 4562
rect 72770 4510 73108 4562
rect 72716 4508 73108 4510
rect 72716 4498 72772 4508
rect 72828 4338 72884 4350
rect 72828 4286 72830 4338
rect 72882 4286 72884 4338
rect 72828 4228 72884 4286
rect 72828 4162 72884 4172
rect 72380 3502 72382 3554
rect 72434 3502 72436 3554
rect 72380 3490 72436 3502
rect 73052 3444 73108 4508
rect 73164 4340 73220 7084
rect 73388 6804 73444 6814
rect 73388 6580 73444 6748
rect 73164 4246 73220 4284
rect 73276 6578 73444 6580
rect 73276 6526 73390 6578
rect 73442 6526 73444 6578
rect 73276 6524 73444 6526
rect 73164 3444 73220 3454
rect 73052 3442 73220 3444
rect 73052 3390 73166 3442
rect 73218 3390 73220 3442
rect 73052 3388 73220 3390
rect 73164 3378 73220 3388
rect 72380 924 72772 980
rect 72380 800 72436 924
rect 59276 700 59556 756
rect 60256 0 60368 800
rect 61600 0 61712 800
rect 62944 0 63056 800
rect 64288 0 64400 800
rect 65632 0 65744 800
rect 66976 0 67088 800
rect 68320 0 68432 800
rect 69664 0 69776 800
rect 71008 0 71120 800
rect 72352 0 72464 800
rect 72716 756 72772 924
rect 73276 756 73332 6524
rect 73388 6514 73444 6524
rect 73388 6020 73444 6030
rect 73388 5926 73444 5964
rect 73500 5572 73556 7308
rect 73612 7252 73668 7422
rect 73612 7186 73668 7196
rect 73724 6580 73780 7644
rect 74060 7588 74116 8878
rect 74060 7522 74116 7532
rect 73948 7476 74004 7486
rect 73948 7382 74004 7420
rect 73724 6514 73780 6524
rect 74172 6580 74228 9662
rect 74172 6514 74228 6524
rect 74284 12066 74340 12078
rect 74284 12014 74286 12066
rect 74338 12014 74340 12066
rect 74172 5684 74228 5694
rect 74060 5682 74228 5684
rect 74060 5630 74174 5682
rect 74226 5630 74228 5682
rect 74060 5628 74228 5630
rect 73500 5516 73780 5572
rect 73500 5236 73556 5246
rect 73500 3554 73556 5180
rect 73724 4900 73780 5516
rect 73724 4844 74004 4900
rect 73948 4450 74004 4844
rect 73948 4398 73950 4450
rect 74002 4398 74004 4450
rect 73948 4386 74004 4398
rect 73500 3502 73502 3554
rect 73554 3502 73556 3554
rect 73500 3490 73556 3502
rect 74060 3444 74116 5628
rect 74172 5618 74228 5628
rect 74172 5236 74228 5246
rect 74172 5142 74228 5180
rect 74284 4676 74340 12014
rect 74396 11396 74452 11406
rect 74396 11302 74452 11340
rect 74620 11170 74676 11182
rect 74620 11118 74622 11170
rect 74674 11118 74676 11170
rect 74396 10724 74452 10734
rect 74620 10724 74676 11118
rect 74396 10722 74676 10724
rect 74396 10670 74398 10722
rect 74450 10670 74676 10722
rect 74396 10668 74676 10670
rect 74396 10658 74452 10668
rect 74508 9602 74564 9614
rect 74508 9550 74510 9602
rect 74562 9550 74564 9602
rect 74508 9380 74564 9550
rect 74508 8484 74564 9324
rect 74508 8418 74564 8428
rect 74620 9044 74676 9054
rect 74620 7586 74676 8988
rect 74620 7534 74622 7586
rect 74674 7534 74676 7586
rect 74620 7522 74676 7534
rect 74284 4610 74340 4620
rect 74732 3668 74788 13804
rect 74844 12740 74900 14028
rect 74956 13746 75012 15260
rect 75180 15316 75236 15326
rect 75516 15316 75572 17052
rect 75628 16772 75684 18286
rect 75740 17108 75796 18396
rect 75740 17014 75796 17052
rect 75852 19796 75908 19806
rect 75628 16716 75796 16772
rect 75628 15988 75684 15998
rect 75628 15894 75684 15932
rect 75180 15314 75572 15316
rect 75180 15262 75182 15314
rect 75234 15262 75572 15314
rect 75180 15260 75572 15262
rect 75180 15250 75236 15260
rect 75292 14644 75348 14654
rect 74956 13694 74958 13746
rect 75010 13694 75012 13746
rect 74956 13682 75012 13694
rect 75068 14588 75292 14644
rect 75068 13636 75124 14588
rect 75292 14578 75348 14588
rect 74956 12852 75012 12862
rect 75068 12852 75124 13580
rect 74956 12850 75124 12852
rect 74956 12798 74958 12850
rect 75010 12798 75124 12850
rect 74956 12796 75124 12798
rect 75180 14418 75236 14430
rect 75180 14366 75182 14418
rect 75234 14366 75236 14418
rect 74956 12786 75012 12796
rect 74844 12674 74900 12684
rect 74844 11396 74900 11406
rect 74844 11302 74900 11340
rect 74956 11394 75012 11406
rect 74956 11342 74958 11394
rect 75010 11342 75012 11394
rect 74844 9940 74900 9950
rect 74844 9826 74900 9884
rect 74844 9774 74846 9826
rect 74898 9774 74900 9826
rect 74844 9762 74900 9774
rect 74956 9828 75012 11342
rect 75180 9938 75236 14366
rect 75292 14308 75348 14318
rect 75628 14308 75684 14318
rect 75292 14306 75460 14308
rect 75292 14254 75294 14306
rect 75346 14254 75460 14306
rect 75292 14252 75460 14254
rect 75292 14242 75348 14252
rect 75404 13748 75460 14252
rect 75404 13682 75460 13692
rect 75516 13860 75572 13870
rect 75292 12740 75348 12750
rect 75292 12646 75348 12684
rect 75404 12292 75460 12302
rect 75516 12292 75572 13804
rect 75404 12290 75572 12292
rect 75404 12238 75406 12290
rect 75458 12238 75572 12290
rect 75404 12236 75572 12238
rect 75404 12226 75460 12236
rect 75180 9886 75182 9938
rect 75234 9886 75236 9938
rect 75180 9874 75236 9886
rect 75292 11620 75348 11630
rect 74956 9762 75012 9772
rect 75292 9826 75348 11564
rect 75628 11396 75684 14252
rect 75516 11340 75684 11396
rect 75516 10612 75572 11340
rect 75628 11170 75684 11182
rect 75628 11118 75630 11170
rect 75682 11118 75684 11170
rect 75628 10836 75684 11118
rect 75740 11172 75796 16716
rect 75852 16212 75908 19740
rect 75964 18452 76020 19964
rect 76300 19954 76356 19964
rect 76524 19926 76580 19964
rect 77196 20132 77252 20142
rect 76748 19908 76804 19918
rect 76748 19814 76804 19852
rect 77196 19234 77252 20076
rect 77756 20132 77812 20142
rect 77196 19182 77198 19234
rect 77250 19182 77252 19234
rect 77196 19170 77252 19182
rect 77308 20018 77364 20030
rect 77308 19966 77310 20018
rect 77362 19966 77364 20018
rect 76188 19012 76244 19022
rect 76076 18452 76132 18462
rect 75964 18450 76132 18452
rect 75964 18398 76078 18450
rect 76130 18398 76132 18450
rect 75964 18396 76132 18398
rect 76076 18386 76132 18396
rect 76188 16882 76244 18956
rect 77308 18452 77364 19966
rect 77644 20020 77700 20030
rect 77644 19906 77700 19964
rect 77644 19854 77646 19906
rect 77698 19854 77700 19906
rect 77644 19842 77700 19854
rect 76860 18396 77364 18452
rect 77756 18450 77812 20076
rect 78092 20130 78148 20524
rect 78316 20578 78372 20590
rect 78316 20526 78318 20578
rect 78370 20526 78372 20578
rect 78316 20468 78372 20526
rect 78540 20580 78596 20750
rect 78540 20514 78596 20524
rect 78316 20402 78372 20412
rect 78092 20078 78094 20130
rect 78146 20078 78148 20130
rect 78092 20066 78148 20078
rect 78652 20132 78708 21644
rect 78764 20804 78820 24670
rect 78988 23268 79044 23278
rect 78876 23154 78932 23166
rect 78876 23102 78878 23154
rect 78930 23102 78932 23154
rect 78876 22820 78932 23102
rect 78988 23154 79044 23212
rect 78988 23102 78990 23154
rect 79042 23102 79044 23154
rect 78988 23090 79044 23102
rect 78876 22754 78932 22764
rect 79100 22482 79156 24892
rect 80444 24948 80500 25230
rect 80444 24882 80500 24892
rect 80668 25284 80724 25294
rect 80892 25284 80948 25294
rect 80724 25282 80948 25284
rect 80724 25230 80894 25282
rect 80946 25230 80948 25282
rect 80724 25228 80948 25230
rect 80332 23828 80388 23838
rect 80668 23828 80724 25228
rect 80892 25218 80948 25228
rect 81276 25116 81540 25126
rect 80332 23826 80724 23828
rect 80332 23774 80334 23826
rect 80386 23774 80724 23826
rect 80332 23772 80724 23774
rect 80220 23268 80276 23278
rect 80220 23174 80276 23212
rect 79548 23042 79604 23054
rect 79548 22990 79550 23042
rect 79602 22990 79604 23042
rect 79548 22820 79604 22990
rect 80108 22932 80164 22942
rect 79548 22754 79604 22764
rect 79884 22930 80164 22932
rect 79884 22878 80110 22930
rect 80162 22878 80164 22930
rect 79884 22876 80164 22878
rect 79100 22430 79102 22482
rect 79154 22430 79156 22482
rect 79100 22418 79156 22430
rect 79324 22372 79380 22382
rect 78988 22148 79044 22158
rect 78764 20690 78820 20748
rect 78764 20638 78766 20690
rect 78818 20638 78820 20690
rect 78764 20626 78820 20638
rect 78876 22146 79044 22148
rect 78876 22094 78990 22146
rect 79042 22094 79044 22146
rect 78876 22092 79044 22094
rect 78652 20066 78708 20076
rect 78204 19796 78260 19806
rect 77756 18398 77758 18450
rect 77810 18398 77812 18450
rect 76636 18338 76692 18350
rect 76636 18286 76638 18338
rect 76690 18286 76692 18338
rect 76636 18228 76692 18286
rect 76188 16830 76190 16882
rect 76242 16830 76244 16882
rect 76188 16548 76244 16830
rect 76412 16882 76468 16894
rect 76412 16830 76414 16882
rect 76466 16830 76468 16882
rect 76300 16772 76356 16782
rect 76300 16678 76356 16716
rect 76188 16482 76244 16492
rect 76412 16324 76468 16830
rect 76636 16884 76692 18172
rect 76860 18340 76916 18396
rect 77756 18386 77812 18398
rect 77868 19794 78260 19796
rect 77868 19742 78206 19794
rect 78258 19742 78260 19794
rect 77868 19740 78260 19742
rect 76860 17666 76916 18284
rect 77420 18116 77476 18126
rect 77196 17780 77252 17790
rect 77196 17686 77252 17724
rect 76860 17614 76862 17666
rect 76914 17614 76916 17666
rect 76860 17602 76916 17614
rect 77420 17332 77476 18060
rect 77868 17444 77924 19740
rect 78204 19730 78260 19740
rect 77420 17266 77476 17276
rect 77756 17388 77924 17444
rect 76636 16818 76692 16828
rect 76860 16884 76916 16894
rect 76860 16790 76916 16828
rect 77644 16884 77700 16894
rect 77196 16772 77252 16782
rect 77196 16770 77476 16772
rect 77196 16718 77198 16770
rect 77250 16718 77476 16770
rect 77196 16716 77476 16718
rect 77196 16706 77252 16716
rect 77420 16548 77476 16716
rect 76412 16258 76468 16268
rect 77308 16324 77364 16334
rect 75852 16156 76132 16212
rect 75852 15876 75908 15886
rect 75852 15426 75908 15820
rect 75852 15374 75854 15426
rect 75906 15374 75908 15426
rect 75852 15362 75908 15374
rect 76076 15148 76132 16156
rect 77084 16100 77140 16110
rect 76636 16098 77140 16100
rect 76636 16046 77086 16098
rect 77138 16046 77140 16098
rect 76636 16044 77140 16046
rect 76412 15988 76468 15998
rect 76636 15988 76692 16044
rect 77084 16034 77140 16044
rect 76468 15932 76692 15988
rect 76412 15922 76468 15932
rect 76300 15876 76356 15886
rect 76300 15782 76356 15820
rect 76748 15876 76804 15886
rect 75964 15092 76132 15148
rect 76636 15764 76692 15774
rect 75740 11106 75796 11116
rect 75852 12292 75908 12302
rect 75852 11060 75908 12236
rect 75852 10994 75908 11004
rect 75628 10780 75908 10836
rect 75516 10556 75684 10612
rect 75292 9774 75294 9826
rect 75346 9774 75348 9826
rect 75292 9762 75348 9774
rect 75404 9826 75460 9838
rect 75404 9774 75406 9826
rect 75458 9774 75460 9826
rect 75068 9604 75124 9614
rect 75068 8370 75124 9548
rect 75404 9380 75460 9774
rect 75068 8318 75070 8370
rect 75122 8318 75124 8370
rect 75068 8306 75124 8318
rect 75292 9324 75460 9380
rect 75292 8036 75348 9324
rect 75628 9268 75684 10556
rect 75852 9940 75908 10780
rect 75964 10052 76020 15092
rect 76412 13748 76468 13758
rect 76412 13654 76468 13692
rect 76188 12850 76244 12862
rect 76188 12798 76190 12850
rect 76242 12798 76244 12850
rect 76076 11396 76132 11406
rect 76076 11302 76132 11340
rect 76188 11172 76244 12798
rect 76300 12738 76356 12750
rect 76300 12686 76302 12738
rect 76354 12686 76356 12738
rect 76300 12178 76356 12686
rect 76300 12126 76302 12178
rect 76354 12126 76356 12178
rect 76300 12114 76356 12126
rect 76412 11844 76468 11854
rect 76300 11396 76356 11406
rect 76300 11282 76356 11340
rect 76300 11230 76302 11282
rect 76354 11230 76356 11282
rect 76300 11218 76356 11230
rect 76412 11282 76468 11788
rect 76412 11230 76414 11282
rect 76466 11230 76468 11282
rect 76188 11106 76244 11116
rect 76412 10388 76468 11230
rect 76524 11396 76580 11406
rect 76524 10498 76580 11340
rect 76524 10446 76526 10498
rect 76578 10446 76580 10498
rect 76524 10434 76580 10446
rect 76636 10388 76692 15708
rect 76748 14644 76804 15820
rect 76972 15876 77028 15886
rect 76972 15782 77028 15820
rect 77196 15874 77252 15886
rect 77196 15822 77198 15874
rect 77250 15822 77252 15874
rect 77196 15204 77252 15822
rect 77196 15138 77252 15148
rect 77308 15148 77364 16268
rect 77420 15876 77476 16492
rect 77644 16770 77700 16828
rect 77644 16718 77646 16770
rect 77698 16718 77700 16770
rect 77644 16324 77700 16718
rect 77644 16098 77700 16268
rect 77644 16046 77646 16098
rect 77698 16046 77700 16098
rect 77644 16034 77700 16046
rect 77420 15810 77476 15820
rect 77308 15092 77476 15148
rect 76748 14642 77140 14644
rect 76748 14590 76750 14642
rect 76802 14590 77140 14642
rect 76748 14588 77140 14590
rect 76748 14578 76804 14588
rect 77084 14530 77140 14588
rect 77084 14478 77086 14530
rect 77138 14478 77140 14530
rect 77084 14466 77140 14478
rect 77420 13746 77476 15092
rect 77420 13694 77422 13746
rect 77474 13694 77476 13746
rect 77420 13682 77476 13694
rect 77084 13636 77140 13646
rect 77084 12292 77140 13580
rect 76972 12236 77140 12292
rect 77196 12962 77252 12974
rect 77196 12910 77198 12962
rect 77250 12910 77252 12962
rect 77196 12292 77252 12910
rect 76972 11844 77028 12236
rect 77196 12226 77252 12236
rect 77420 12292 77476 12302
rect 76972 11788 77140 11844
rect 77084 11506 77140 11788
rect 77084 11454 77086 11506
rect 77138 11454 77140 11506
rect 77084 11442 77140 11454
rect 77196 11620 77252 11630
rect 76748 11394 76804 11406
rect 76748 11342 76750 11394
rect 76802 11342 76804 11394
rect 76748 11060 76804 11342
rect 76972 11396 77028 11434
rect 76972 11330 77028 11340
rect 77196 11396 77252 11564
rect 77196 11394 77364 11396
rect 77196 11342 77198 11394
rect 77250 11342 77364 11394
rect 77196 11340 77364 11342
rect 77196 11330 77252 11340
rect 76972 11172 77028 11182
rect 77028 11116 77140 11172
rect 76972 11106 77028 11116
rect 76748 10994 76804 11004
rect 76972 10836 77028 10846
rect 77084 10836 77140 11116
rect 77196 10836 77252 10846
rect 77084 10834 77252 10836
rect 77084 10782 77198 10834
rect 77250 10782 77252 10834
rect 77084 10780 77252 10782
rect 76972 10742 77028 10780
rect 77196 10770 77252 10780
rect 77308 10834 77364 11340
rect 77420 11394 77476 12236
rect 77420 11342 77422 11394
rect 77474 11342 77476 11394
rect 77420 11330 77476 11342
rect 77308 10782 77310 10834
rect 77362 10782 77364 10834
rect 77308 10770 77364 10782
rect 77084 10612 77140 10622
rect 77084 10610 77252 10612
rect 77084 10558 77086 10610
rect 77138 10558 77252 10610
rect 77084 10556 77252 10558
rect 77084 10546 77140 10556
rect 76636 10332 77028 10388
rect 76412 10322 76468 10332
rect 75964 9996 76580 10052
rect 75852 9884 76020 9940
rect 75964 9380 76020 9884
rect 76188 9828 76244 9838
rect 75964 9314 76020 9324
rect 76076 9826 76244 9828
rect 76076 9774 76190 9826
rect 76242 9774 76244 9826
rect 76076 9772 76244 9774
rect 75852 9268 75908 9278
rect 75628 9266 75908 9268
rect 75628 9214 75854 9266
rect 75906 9214 75908 9266
rect 75628 9212 75908 9214
rect 75852 9202 75908 9212
rect 75404 9154 75460 9166
rect 75404 9102 75406 9154
rect 75458 9102 75460 9154
rect 75404 8596 75460 9102
rect 75404 8540 75908 8596
rect 75740 8372 75796 8382
rect 75404 8260 75460 8298
rect 75404 8194 75460 8204
rect 75740 8258 75796 8316
rect 75740 8206 75742 8258
rect 75794 8206 75796 8258
rect 75740 8194 75796 8206
rect 75404 8036 75460 8046
rect 75292 7980 75404 8036
rect 75404 7970 75460 7980
rect 75516 8034 75572 8046
rect 75516 7982 75518 8034
rect 75570 7982 75572 8034
rect 75516 7364 75572 7982
rect 75516 7298 75572 7308
rect 75740 6916 75796 6926
rect 75852 6916 75908 8540
rect 75740 6914 75908 6916
rect 75740 6862 75742 6914
rect 75794 6862 75908 6914
rect 75740 6860 75908 6862
rect 75964 7700 76020 7710
rect 75740 6850 75796 6860
rect 75292 6020 75348 6030
rect 74844 3668 74900 3678
rect 74732 3666 74900 3668
rect 74732 3614 74846 3666
rect 74898 3614 74900 3666
rect 74732 3612 74900 3614
rect 74844 3602 74900 3612
rect 73724 3388 74116 3444
rect 75292 3388 75348 5964
rect 75740 5124 75796 5134
rect 75516 5010 75572 5022
rect 75516 4958 75518 5010
rect 75570 4958 75572 5010
rect 75516 4564 75572 4958
rect 75516 4498 75572 4508
rect 75740 3388 75796 5068
rect 75964 4228 76020 7644
rect 76076 6916 76132 9772
rect 76188 9762 76244 9772
rect 76076 6850 76132 6860
rect 76188 9154 76244 9166
rect 76188 9102 76190 9154
rect 76242 9102 76244 9154
rect 76188 5124 76244 9102
rect 76188 5058 76244 5068
rect 76300 7252 76356 7262
rect 76300 4562 76356 7196
rect 76412 6692 76468 6702
rect 76412 6598 76468 6636
rect 76412 6468 76468 6478
rect 76412 5906 76468 6412
rect 76412 5854 76414 5906
rect 76466 5854 76468 5906
rect 76412 5842 76468 5854
rect 76524 5236 76580 9996
rect 76748 9604 76804 9614
rect 76748 9602 76916 9604
rect 76748 9550 76750 9602
rect 76802 9550 76916 9602
rect 76748 9548 76916 9550
rect 76748 9538 76804 9548
rect 76636 8932 76692 8942
rect 76636 6580 76692 8876
rect 76860 7588 76916 9548
rect 76972 8596 77028 10332
rect 77084 9602 77140 9614
rect 77084 9550 77086 9602
rect 77138 9550 77140 9602
rect 77084 8820 77140 9550
rect 77084 8754 77140 8764
rect 76972 8540 77140 8596
rect 76972 8370 77028 8382
rect 76972 8318 76974 8370
rect 77026 8318 77028 8370
rect 76972 8148 77028 8318
rect 77084 8258 77140 8540
rect 77084 8206 77086 8258
rect 77138 8206 77140 8258
rect 77084 8194 77140 8206
rect 76972 8082 77028 8092
rect 76860 7532 77140 7588
rect 76748 7364 76804 7374
rect 76748 7270 76804 7308
rect 77084 7362 77140 7532
rect 77084 7310 77086 7362
rect 77138 7310 77140 7362
rect 77084 7298 77140 7310
rect 77196 7364 77252 10556
rect 77532 10610 77588 10622
rect 77532 10558 77534 10610
rect 77586 10558 77588 10610
rect 77532 10500 77588 10558
rect 77532 10434 77588 10444
rect 77420 9602 77476 9614
rect 77420 9550 77422 9602
rect 77474 9550 77476 9602
rect 77420 9380 77476 9550
rect 77420 9314 77476 9324
rect 77532 9044 77588 9054
rect 77588 8988 77700 9044
rect 77532 8950 77588 8988
rect 77532 8372 77588 8382
rect 77532 8258 77588 8316
rect 77532 8206 77534 8258
rect 77586 8206 77588 8258
rect 77532 8194 77588 8206
rect 77420 8034 77476 8046
rect 77420 7982 77422 8034
rect 77474 7982 77476 8034
rect 77196 7298 77252 7308
rect 77308 7588 77364 7598
rect 77308 6916 77364 7532
rect 77196 6692 77252 6702
rect 76972 6580 77028 6590
rect 76636 6578 77140 6580
rect 76636 6526 76974 6578
rect 77026 6526 77140 6578
rect 76636 6524 77140 6526
rect 76972 6514 77028 6524
rect 76972 6020 77028 6030
rect 76972 5926 77028 5964
rect 77084 5348 77140 6524
rect 77084 5282 77140 5292
rect 76972 5236 77028 5246
rect 76524 5234 77028 5236
rect 76524 5182 76974 5234
rect 77026 5182 77028 5234
rect 76524 5180 77028 5182
rect 76972 5170 77028 5180
rect 77196 5122 77252 6636
rect 77196 5070 77198 5122
rect 77250 5070 77252 5122
rect 76524 5012 76580 5022
rect 76412 4900 76468 4910
rect 76412 4806 76468 4844
rect 76300 4510 76302 4562
rect 76354 4510 76356 4562
rect 76300 4498 76356 4510
rect 76412 4676 76468 4686
rect 76076 4228 76132 4238
rect 75964 4226 76132 4228
rect 75964 4174 76078 4226
rect 76130 4174 76132 4226
rect 75964 4172 76132 4174
rect 76076 4162 76132 4172
rect 73724 800 73780 3388
rect 74284 3330 74340 3342
rect 74284 3278 74286 3330
rect 74338 3278 74340 3330
rect 74284 2548 74340 3278
rect 74284 2482 74340 2492
rect 75068 3332 75348 3388
rect 75628 3332 75796 3388
rect 76076 3444 76132 3482
rect 76076 3378 76132 3388
rect 75068 800 75124 3332
rect 75628 2436 75684 3332
rect 75628 2370 75684 2380
rect 76412 800 76468 4620
rect 76524 4562 76580 4956
rect 76524 4510 76526 4562
rect 76578 4510 76580 4562
rect 76972 4564 77028 4574
rect 76524 4498 76580 4510
rect 76636 4506 76692 4518
rect 76636 4454 76638 4506
rect 76690 4454 76692 4506
rect 76972 4470 77028 4508
rect 76636 4452 76692 4454
rect 76636 4396 76804 4452
rect 76524 4340 76580 4350
rect 76748 4340 76804 4396
rect 77196 4340 77252 5070
rect 76748 4284 77028 4340
rect 76524 3554 76580 4284
rect 76524 3502 76526 3554
rect 76578 3502 76580 3554
rect 76524 3490 76580 3502
rect 76972 4116 77028 4284
rect 77196 4274 77252 4284
rect 77196 4116 77252 4126
rect 76972 4060 77196 4116
rect 76972 3556 77028 4060
rect 77196 4050 77252 4060
rect 76972 3442 77028 3500
rect 77196 3556 77252 3566
rect 77308 3556 77364 6860
rect 77420 5796 77476 7982
rect 77644 6356 77700 8988
rect 77756 6916 77812 17388
rect 78204 16770 78260 16782
rect 78204 16718 78206 16770
rect 78258 16718 78260 16770
rect 77980 16212 78036 16222
rect 77980 15876 78036 16156
rect 77980 15810 78036 15820
rect 77980 15204 78036 15242
rect 78204 15148 78260 16718
rect 78428 16324 78484 16334
rect 78428 16210 78484 16268
rect 78428 16158 78430 16210
rect 78482 16158 78484 16210
rect 78428 16146 78484 16158
rect 78540 16322 78596 16334
rect 78540 16270 78542 16322
rect 78594 16270 78596 16322
rect 78428 15540 78484 15550
rect 78540 15540 78596 16270
rect 78428 15538 78540 15540
rect 78428 15486 78430 15538
rect 78482 15486 78540 15538
rect 78428 15484 78540 15486
rect 78428 15474 78484 15484
rect 78540 15446 78596 15484
rect 77868 15092 78036 15148
rect 78092 15092 78260 15148
rect 77868 14418 77924 15092
rect 77868 14366 77870 14418
rect 77922 14366 77924 14418
rect 77868 14354 77924 14366
rect 77868 13972 77924 13982
rect 77868 12290 77924 13916
rect 78092 13076 78148 15092
rect 78652 14980 78708 14990
rect 78428 13972 78484 13982
rect 77868 12238 77870 12290
rect 77922 12238 77924 12290
rect 77868 12226 77924 12238
rect 77980 13020 78148 13076
rect 78204 13746 78260 13758
rect 78204 13694 78206 13746
rect 78258 13694 78260 13746
rect 78204 13524 78260 13694
rect 77868 11060 77924 11070
rect 77868 10834 77924 11004
rect 77868 10782 77870 10834
rect 77922 10782 77924 10834
rect 77868 10770 77924 10782
rect 77868 9602 77924 9614
rect 77868 9550 77870 9602
rect 77922 9550 77924 9602
rect 77868 9492 77924 9550
rect 77868 9156 77924 9436
rect 77868 9090 77924 9100
rect 77980 7588 78036 13020
rect 78092 12850 78148 12862
rect 78092 12798 78094 12850
rect 78146 12798 78148 12850
rect 78092 12740 78148 12798
rect 78092 12674 78148 12684
rect 78204 12178 78260 13468
rect 78428 12402 78484 13916
rect 78652 13970 78708 14924
rect 78652 13918 78654 13970
rect 78706 13918 78708 13970
rect 78652 13906 78708 13918
rect 78540 12962 78596 12974
rect 78540 12910 78542 12962
rect 78594 12910 78596 12962
rect 78540 12852 78596 12910
rect 78596 12796 78820 12852
rect 78540 12786 78596 12796
rect 78428 12350 78430 12402
rect 78482 12350 78484 12402
rect 78428 12338 78484 12350
rect 78204 12126 78206 12178
rect 78258 12126 78260 12178
rect 78204 12114 78260 12126
rect 78540 12292 78596 12302
rect 78204 11396 78260 11406
rect 78204 10836 78260 11340
rect 78204 10742 78260 10780
rect 78204 10388 78260 10398
rect 78204 9602 78260 10332
rect 78540 9938 78596 12236
rect 78764 12180 78820 12796
rect 78764 10834 78820 12124
rect 78764 10782 78766 10834
rect 78818 10782 78820 10834
rect 78764 10770 78820 10782
rect 78540 9886 78542 9938
rect 78594 9886 78596 9938
rect 78540 9874 78596 9886
rect 78204 9550 78206 9602
rect 78258 9550 78260 9602
rect 78204 8596 78260 9550
rect 78428 9042 78484 9054
rect 78428 8990 78430 9042
rect 78482 8990 78484 9042
rect 78316 8932 78372 8942
rect 78316 8838 78372 8876
rect 78204 8530 78260 8540
rect 78092 8370 78148 8382
rect 78092 8318 78094 8370
rect 78146 8318 78148 8370
rect 78092 8036 78148 8318
rect 78428 8372 78484 8990
rect 78764 9044 78820 9054
rect 78876 9044 78932 22092
rect 78988 22082 79044 22092
rect 79324 20916 79380 22316
rect 79548 21476 79604 21486
rect 79548 21382 79604 21420
rect 79324 20822 79380 20860
rect 78988 19122 79044 19134
rect 78988 19070 78990 19122
rect 79042 19070 79044 19122
rect 78988 18452 79044 19070
rect 79044 18396 79380 18452
rect 78988 18386 79044 18396
rect 79212 18004 79268 18014
rect 79212 17108 79268 17948
rect 79212 17014 79268 17052
rect 79324 17444 79380 18396
rect 79548 18450 79604 18462
rect 79548 18398 79550 18450
rect 79602 18398 79604 18450
rect 79548 18228 79604 18398
rect 79548 18162 79604 18172
rect 79772 17668 79828 17678
rect 79772 17444 79828 17612
rect 79324 17442 79828 17444
rect 79324 17390 79326 17442
rect 79378 17390 79774 17442
rect 79826 17390 79828 17442
rect 79324 17388 79828 17390
rect 78988 16772 79044 16782
rect 78988 16770 79156 16772
rect 78988 16718 78990 16770
rect 79042 16718 79156 16770
rect 78988 16716 79156 16718
rect 78988 16706 79044 16716
rect 78988 15874 79044 15886
rect 78988 15822 78990 15874
rect 79042 15822 79044 15874
rect 78988 12404 79044 15822
rect 79100 15428 79156 16716
rect 79324 16322 79380 17388
rect 79772 17378 79828 17388
rect 79324 16270 79326 16322
rect 79378 16270 79380 16322
rect 79324 16258 79380 16270
rect 79548 16994 79604 17006
rect 79548 16942 79550 16994
rect 79602 16942 79604 16994
rect 79548 16100 79604 16942
rect 79884 16324 79940 22876
rect 80108 22866 80164 22876
rect 80220 21812 80276 21822
rect 80332 21812 80388 23772
rect 80668 23716 80724 23772
rect 80668 23650 80724 23660
rect 80780 25060 80836 25070
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81276 25050 81540 25060
rect 80780 24946 80836 25004
rect 80780 24894 80782 24946
rect 80834 24894 80836 24946
rect 80668 23156 80724 23166
rect 80780 23156 80836 24894
rect 81116 24836 81172 24846
rect 81116 24742 81172 24780
rect 81900 24836 81956 24846
rect 81452 24612 81508 24622
rect 81452 24610 81732 24612
rect 81452 24558 81454 24610
rect 81506 24558 81732 24610
rect 81452 24556 81732 24558
rect 81452 24546 81508 24556
rect 81276 23548 81540 23558
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81276 23482 81540 23492
rect 81564 23380 81620 23390
rect 81676 23380 81732 24556
rect 81564 23378 81732 23380
rect 81564 23326 81566 23378
rect 81618 23326 81732 23378
rect 81564 23324 81732 23326
rect 80668 23154 80836 23156
rect 80668 23102 80670 23154
rect 80722 23102 80836 23154
rect 80668 23100 80836 23102
rect 80892 23266 80948 23278
rect 80892 23214 80894 23266
rect 80946 23214 80948 23266
rect 80668 23090 80724 23100
rect 80892 23044 80948 23214
rect 81564 23268 81620 23324
rect 81564 23202 81620 23212
rect 81788 23268 81844 23278
rect 81900 23268 81956 24780
rect 82796 24724 82852 24734
rect 82572 24668 82796 24724
rect 82572 23378 82628 24668
rect 82796 24658 82852 24668
rect 82572 23326 82574 23378
rect 82626 23326 82628 23378
rect 82572 23314 82628 23326
rect 81788 23266 82068 23268
rect 81788 23214 81790 23266
rect 81842 23214 82068 23266
rect 81788 23212 82068 23214
rect 81788 23202 81844 23212
rect 80892 22978 80948 22988
rect 81116 23154 81172 23166
rect 81116 23102 81118 23154
rect 81170 23102 81172 23154
rect 80276 21756 80388 21812
rect 80444 22146 80500 22158
rect 80444 22094 80446 22146
rect 80498 22094 80500 22146
rect 80444 21812 80500 22094
rect 80220 21718 80276 21756
rect 80444 21746 80500 21756
rect 81116 20804 81172 23102
rect 81676 23042 81732 23054
rect 81676 22990 81678 23042
rect 81730 22990 81732 23042
rect 81676 22932 81732 22990
rect 82012 22932 82068 23212
rect 81676 22866 81732 22876
rect 81788 22876 82068 22932
rect 82124 23154 82180 23166
rect 82124 23102 82126 23154
rect 82178 23102 82180 23154
rect 82124 22932 82180 23102
rect 81276 21980 81540 21990
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81276 21914 81540 21924
rect 81676 21924 81732 21934
rect 81452 21812 81508 21822
rect 81452 20914 81508 21756
rect 81452 20862 81454 20914
rect 81506 20862 81508 20914
rect 81452 20850 81508 20862
rect 81564 21586 81620 21598
rect 81564 21534 81566 21586
rect 81618 21534 81620 21586
rect 81116 20738 81172 20748
rect 81564 20804 81620 21534
rect 81564 20738 81620 20748
rect 80556 20580 80612 20590
rect 80444 18450 80500 18462
rect 80444 18398 80446 18450
rect 80498 18398 80500 18450
rect 79996 17668 80052 17678
rect 79996 17574 80052 17612
rect 80444 17668 80500 18398
rect 80444 17602 80500 17612
rect 80108 17108 80164 17118
rect 80108 17014 80164 17052
rect 79548 16034 79604 16044
rect 79772 16268 79940 16324
rect 79996 16996 80052 17006
rect 80444 16996 80500 17006
rect 79100 15362 79156 15372
rect 79436 15874 79492 15886
rect 79436 15822 79438 15874
rect 79490 15822 79492 15874
rect 79100 15202 79156 15214
rect 79100 15150 79102 15202
rect 79154 15150 79156 15202
rect 79100 14196 79156 15150
rect 79436 15148 79492 15822
rect 79772 15764 79828 16268
rect 79996 16210 80052 16940
rect 80220 16994 80500 16996
rect 80220 16942 80446 16994
rect 80498 16942 80500 16994
rect 80220 16940 80500 16942
rect 80220 16884 80276 16940
rect 80444 16930 80500 16940
rect 79996 16158 79998 16210
rect 80050 16158 80052 16210
rect 79996 16146 80052 16158
rect 80108 16828 80276 16884
rect 79772 15698 79828 15708
rect 79884 16100 79940 16110
rect 79548 15540 79604 15550
rect 79548 15446 79604 15484
rect 79884 15148 79940 16044
rect 80108 15988 80164 16828
rect 80556 16772 80612 20524
rect 81564 20580 81620 20618
rect 81564 20514 81620 20524
rect 81276 20412 81540 20422
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81276 20346 81540 20356
rect 80892 20020 80948 20030
rect 80780 17668 80836 17678
rect 80780 17574 80836 17612
rect 80892 17106 80948 19964
rect 81228 20018 81284 20030
rect 81228 19966 81230 20018
rect 81282 19966 81284 20018
rect 81228 19684 81284 19966
rect 81564 20018 81620 20030
rect 81564 19966 81566 20018
rect 81618 19966 81620 20018
rect 81228 19618 81284 19628
rect 81340 19906 81396 19918
rect 81340 19854 81342 19906
rect 81394 19854 81396 19906
rect 81340 19236 81396 19854
rect 81564 19796 81620 19966
rect 81564 19730 81620 19740
rect 81676 19684 81732 21868
rect 81788 21588 81844 22876
rect 82124 22866 82180 22876
rect 82236 23156 82292 23166
rect 82012 21812 82068 21822
rect 82012 21718 82068 21756
rect 82124 21812 82180 21822
rect 82236 21812 82292 23100
rect 82460 23154 82516 23166
rect 82460 23102 82462 23154
rect 82514 23102 82516 23154
rect 82460 22932 82516 23102
rect 82460 22866 82516 22876
rect 82684 23156 82740 23166
rect 82908 23156 82964 23166
rect 82684 23154 82964 23156
rect 82684 23102 82686 23154
rect 82738 23102 82910 23154
rect 82962 23102 82964 23154
rect 82684 23100 82964 23102
rect 82684 23044 82740 23100
rect 82908 23090 82964 23100
rect 82684 21924 82740 22988
rect 83132 23042 83188 23054
rect 83132 22990 83134 23042
rect 83186 22990 83188 23042
rect 83132 22708 83188 22990
rect 82908 22652 83188 22708
rect 82908 22370 82964 22652
rect 82908 22318 82910 22370
rect 82962 22318 82964 22370
rect 82908 22306 82964 22318
rect 82684 21858 82740 21868
rect 82124 21810 82292 21812
rect 82124 21758 82126 21810
rect 82178 21758 82292 21810
rect 82124 21756 82292 21758
rect 83244 21812 83300 29372
rect 88060 28756 88116 28766
rect 86940 26290 86996 26302
rect 86940 26238 86942 26290
rect 86994 26238 86996 26290
rect 86156 26180 86212 26190
rect 86156 26086 86212 26124
rect 86604 26180 86660 26190
rect 86604 26086 86660 26124
rect 86940 26068 86996 26238
rect 86996 26012 87332 26068
rect 86940 26002 86996 26012
rect 87276 25620 87332 26012
rect 87276 25618 87668 25620
rect 87276 25566 87278 25618
rect 87330 25566 87668 25618
rect 87276 25564 87668 25566
rect 87276 25554 87332 25564
rect 87612 25506 87668 25564
rect 87612 25454 87614 25506
rect 87666 25454 87668 25506
rect 87612 25442 87668 25454
rect 83804 24724 83860 24734
rect 83804 24630 83860 24668
rect 84364 24722 84420 24734
rect 84364 24670 84366 24722
rect 84418 24670 84420 24722
rect 84364 24612 84420 24670
rect 84924 24612 84980 24622
rect 84364 24610 84980 24612
rect 84364 24558 84926 24610
rect 84978 24558 84980 24610
rect 84364 24556 84980 24558
rect 83356 23716 83412 23726
rect 83356 23380 83412 23660
rect 84364 23716 84420 24556
rect 84924 24546 84980 24556
rect 84364 23650 84420 23660
rect 84588 23940 84644 23950
rect 84588 23716 84644 23884
rect 86828 23938 86884 23950
rect 86828 23886 86830 23938
rect 86882 23886 86884 23938
rect 86828 23828 86884 23886
rect 86604 23716 86660 23726
rect 84588 23650 84644 23660
rect 86380 23714 86660 23716
rect 86380 23662 86606 23714
rect 86658 23662 86660 23714
rect 86380 23660 86660 23662
rect 83356 23324 83524 23380
rect 83356 23154 83412 23166
rect 83356 23102 83358 23154
rect 83410 23102 83412 23154
rect 83356 23044 83412 23102
rect 83356 22978 83412 22988
rect 83468 22484 83524 23324
rect 86380 23266 86436 23660
rect 86604 23650 86660 23660
rect 86380 23214 86382 23266
rect 86434 23214 86436 23266
rect 83580 23156 83636 23166
rect 83580 23062 83636 23100
rect 83468 22370 83524 22428
rect 83468 22318 83470 22370
rect 83522 22318 83524 22370
rect 83468 22306 83524 22318
rect 84028 23042 84084 23054
rect 84028 22990 84030 23042
rect 84082 22990 84084 23042
rect 84028 22932 84084 22990
rect 84476 23044 84532 23054
rect 84476 22950 84532 22988
rect 86156 23044 86212 23054
rect 83244 21756 83412 21812
rect 82124 21746 82180 21756
rect 82236 21588 82292 21598
rect 81788 21586 82292 21588
rect 81788 21534 82238 21586
rect 82290 21534 82292 21586
rect 81788 21532 82292 21534
rect 81788 20132 81844 20142
rect 81788 20038 81844 20076
rect 82124 20018 82180 21532
rect 82236 21522 82292 21532
rect 82236 20132 82292 20142
rect 82236 20038 82292 20076
rect 82572 20130 82628 20142
rect 82572 20078 82574 20130
rect 82626 20078 82628 20130
rect 82124 19966 82126 20018
rect 82178 19966 82180 20018
rect 81676 19618 81732 19628
rect 82012 19796 82068 19806
rect 82012 19346 82068 19740
rect 82012 19294 82014 19346
rect 82066 19294 82068 19346
rect 82012 19282 82068 19294
rect 81116 19180 81396 19236
rect 81116 18450 81172 19180
rect 82124 19124 82180 19966
rect 82348 20018 82404 20030
rect 82348 19966 82350 20018
rect 82402 19966 82404 20018
rect 81788 19068 82180 19124
rect 82236 19684 82292 19694
rect 81276 18844 81540 18854
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81276 18778 81540 18788
rect 81116 18398 81118 18450
rect 81170 18398 81172 18450
rect 81116 18386 81172 18398
rect 81276 17276 81540 17286
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81276 17210 81540 17220
rect 80892 17054 80894 17106
rect 80946 17054 80948 17106
rect 80892 16996 80948 17054
rect 81228 17108 81284 17118
rect 81228 17106 81732 17108
rect 81228 17054 81230 17106
rect 81282 17054 81732 17106
rect 81228 17052 81732 17054
rect 81228 17042 81284 17052
rect 80892 16930 80948 16940
rect 81116 16996 81172 17006
rect 81116 16902 81172 16940
rect 81676 16994 81732 17052
rect 81676 16942 81678 16994
rect 81730 16942 81732 16994
rect 81676 16930 81732 16942
rect 81340 16884 81396 16894
rect 81340 16882 81620 16884
rect 81340 16830 81342 16882
rect 81394 16830 81620 16882
rect 81340 16828 81620 16830
rect 81340 16818 81396 16828
rect 80108 15922 80164 15932
rect 80220 16716 80612 16772
rect 81564 16772 81620 16828
rect 81788 16772 81844 19068
rect 82012 18228 82068 18238
rect 81900 17220 81956 17230
rect 81900 16994 81956 17164
rect 81900 16942 81902 16994
rect 81954 16942 81956 16994
rect 81900 16930 81956 16942
rect 81564 16716 81844 16772
rect 80108 15540 80164 15550
rect 80108 15314 80164 15484
rect 80108 15262 80110 15314
rect 80162 15262 80164 15314
rect 80108 15250 80164 15262
rect 79436 15092 79716 15148
rect 79100 13524 79156 14140
rect 79212 14530 79268 14542
rect 79212 14478 79214 14530
rect 79266 14478 79268 14530
rect 79212 13970 79268 14478
rect 79212 13918 79214 13970
rect 79266 13918 79268 13970
rect 79212 13906 79268 13918
rect 79324 13636 79380 13646
rect 79324 13542 79380 13580
rect 79100 13458 79156 13468
rect 79660 12628 79716 15092
rect 78988 12348 79380 12404
rect 79212 12178 79268 12190
rect 79212 12126 79214 12178
rect 79266 12126 79268 12178
rect 78988 11284 79044 11294
rect 78988 10836 79044 11228
rect 78988 10770 79044 10780
rect 79100 11172 79156 11182
rect 79100 10610 79156 11116
rect 79212 10722 79268 12126
rect 79212 10670 79214 10722
rect 79266 10670 79268 10722
rect 79212 10658 79268 10670
rect 79100 10558 79102 10610
rect 79154 10558 79156 10610
rect 79100 10546 79156 10558
rect 78764 9042 78932 9044
rect 78764 8990 78766 9042
rect 78818 8990 78932 9042
rect 78764 8988 78932 8990
rect 78764 8978 78820 8988
rect 78652 8818 78708 8830
rect 78652 8766 78654 8818
rect 78706 8766 78708 8818
rect 78540 8372 78596 8382
rect 78428 8316 78540 8372
rect 78540 8306 78596 8316
rect 78148 7980 78372 8036
rect 78092 7942 78148 7980
rect 77980 7522 78036 7532
rect 77756 6860 78148 6916
rect 78092 6804 78148 6860
rect 78204 6804 78260 6814
rect 78092 6802 78260 6804
rect 78092 6750 78206 6802
rect 78258 6750 78260 6802
rect 78092 6748 78260 6750
rect 78204 6738 78260 6748
rect 77644 6290 77700 6300
rect 77980 6466 78036 6478
rect 77980 6414 77982 6466
rect 78034 6414 78036 6466
rect 77420 5740 77924 5796
rect 77196 3554 77364 3556
rect 77196 3502 77198 3554
rect 77250 3502 77364 3554
rect 77196 3500 77364 3502
rect 77644 5348 77700 5358
rect 77644 5012 77700 5292
rect 77756 5012 77812 5022
rect 77644 5010 77812 5012
rect 77644 4958 77758 5010
rect 77810 4958 77812 5010
rect 77644 4956 77812 4958
rect 77196 3490 77252 3500
rect 76972 3390 76974 3442
rect 77026 3390 77028 3442
rect 76972 3378 77028 3390
rect 77644 3444 77700 4956
rect 77756 4946 77812 4956
rect 77644 3378 77700 3388
rect 77756 3668 77812 3678
rect 77756 800 77812 3612
rect 77868 3556 77924 5740
rect 77980 3780 78036 6414
rect 78316 6020 78372 7980
rect 78428 7586 78484 7598
rect 78428 7534 78430 7586
rect 78482 7534 78484 7586
rect 78428 6132 78484 7534
rect 78428 6066 78484 6076
rect 78316 5954 78372 5964
rect 78652 5908 78708 8766
rect 79212 8372 79268 8382
rect 78988 7588 79044 7598
rect 78988 7474 79044 7532
rect 78988 7422 78990 7474
rect 79042 7422 79044 7474
rect 78988 7410 79044 7422
rect 78652 5842 78708 5852
rect 79212 5234 79268 8316
rect 79324 6468 79380 12348
rect 79436 12292 79492 12302
rect 79436 12198 79492 12236
rect 79660 12292 79716 12572
rect 79660 12226 79716 12236
rect 79772 15092 79940 15148
rect 79548 12178 79604 12190
rect 79548 12126 79550 12178
rect 79602 12126 79604 12178
rect 79548 11844 79604 12126
rect 79548 11778 79604 11788
rect 79772 11172 79828 15092
rect 80220 13188 80276 16716
rect 81340 16436 81396 16446
rect 80556 16100 80612 16110
rect 80444 16098 80612 16100
rect 80444 16046 80558 16098
rect 80610 16046 80612 16098
rect 80444 16044 80612 16046
rect 80332 15986 80388 15998
rect 80332 15934 80334 15986
rect 80386 15934 80388 15986
rect 80332 14644 80388 15934
rect 80444 14756 80500 16044
rect 80556 16034 80612 16044
rect 80780 16100 80836 16110
rect 80780 16006 80836 16044
rect 81340 16098 81396 16380
rect 81340 16046 81342 16098
rect 81394 16046 81396 16098
rect 81340 16034 81396 16046
rect 80556 15874 80612 15886
rect 80556 15822 80558 15874
rect 80610 15822 80612 15874
rect 80556 15540 80612 15822
rect 81676 15876 81732 15886
rect 81676 15874 81844 15876
rect 81676 15822 81678 15874
rect 81730 15822 81844 15874
rect 81676 15820 81844 15822
rect 81676 15810 81732 15820
rect 81276 15708 81540 15718
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81276 15642 81540 15652
rect 81676 15652 81732 15662
rect 80556 15484 80948 15540
rect 80892 15426 80948 15484
rect 80892 15374 80894 15426
rect 80946 15374 80948 15426
rect 80892 15362 80948 15374
rect 80444 14690 80500 14700
rect 80556 14868 80612 14878
rect 80332 14578 80388 14588
rect 80556 14532 80612 14812
rect 81452 14756 81508 14766
rect 81452 14662 81508 14700
rect 80780 14532 80836 14542
rect 80556 14530 80836 14532
rect 80556 14478 80782 14530
rect 80834 14478 80836 14530
rect 80556 14476 80836 14478
rect 80780 14466 80836 14476
rect 81228 14532 81284 14542
rect 80332 14420 80388 14430
rect 80332 13970 80388 14364
rect 81116 14418 81172 14430
rect 81116 14366 81118 14418
rect 81170 14366 81172 14418
rect 81116 14308 81172 14366
rect 81116 14242 81172 14252
rect 81228 14306 81284 14476
rect 81564 14420 81620 14430
rect 81564 14326 81620 14364
rect 81228 14254 81230 14306
rect 81282 14254 81284 14306
rect 81228 14242 81284 14254
rect 81276 14140 81540 14150
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81276 14074 81540 14084
rect 80332 13918 80334 13970
rect 80386 13918 80388 13970
rect 80332 13748 80388 13918
rect 81116 13748 81172 13758
rect 80332 13682 80388 13692
rect 81004 13746 81172 13748
rect 81004 13694 81118 13746
rect 81170 13694 81172 13746
rect 81004 13692 81172 13694
rect 80780 13636 80836 13646
rect 81004 13636 81060 13692
rect 81116 13682 81172 13692
rect 80780 13634 81060 13636
rect 80780 13582 80782 13634
rect 80834 13582 81060 13634
rect 80780 13580 81060 13582
rect 80220 13132 80388 13188
rect 79884 13076 79940 13086
rect 79884 12962 79940 13020
rect 79884 12910 79886 12962
rect 79938 12910 79940 12962
rect 79884 12898 79940 12910
rect 80220 12962 80276 12974
rect 80220 12910 80222 12962
rect 80274 12910 80276 12962
rect 80220 12740 80276 12910
rect 80220 12674 80276 12684
rect 80108 12180 80164 12190
rect 80108 12086 80164 12124
rect 79828 11116 80052 11172
rect 79772 11106 79828 11116
rect 79660 10724 79716 10734
rect 79660 10610 79716 10668
rect 79660 10558 79662 10610
rect 79714 10558 79716 10610
rect 79660 10546 79716 10558
rect 79436 10498 79492 10510
rect 79436 10446 79438 10498
rect 79490 10446 79492 10498
rect 79436 9940 79492 10446
rect 79436 9874 79492 9884
rect 79996 9716 80052 11116
rect 79772 9380 79828 9390
rect 79436 8484 79492 8494
rect 79436 7362 79492 8428
rect 79772 7588 79828 9324
rect 79996 9156 80052 9660
rect 80108 10610 80164 10622
rect 80108 10558 80110 10610
rect 80162 10558 80164 10610
rect 80108 9380 80164 10558
rect 80332 9828 80388 13132
rect 80780 12180 80836 13580
rect 81116 13524 81172 13534
rect 81116 12180 81172 13468
rect 81564 13076 81620 13086
rect 81564 12962 81620 13020
rect 81564 12910 81566 12962
rect 81618 12910 81620 12962
rect 81564 12898 81620 12910
rect 81276 12572 81540 12582
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81276 12506 81540 12516
rect 81452 12180 81508 12190
rect 81116 12178 81508 12180
rect 81116 12126 81454 12178
rect 81506 12126 81508 12178
rect 81116 12124 81508 12126
rect 80780 12114 80836 12124
rect 81452 12114 81508 12124
rect 81564 12068 81620 12078
rect 81564 11284 81620 12012
rect 81676 11620 81732 15596
rect 81788 14644 81844 15820
rect 82012 15148 82068 18172
rect 82124 17668 82180 17678
rect 82124 17106 82180 17612
rect 82124 17054 82126 17106
rect 82178 17054 82180 17106
rect 82124 17042 82180 17054
rect 82236 16994 82292 19628
rect 82348 18452 82404 19966
rect 82572 20020 82628 20078
rect 82572 19954 82628 19964
rect 82348 18386 82404 18396
rect 83132 17444 83188 17454
rect 82236 16942 82238 16994
rect 82290 16942 82292 16994
rect 82236 16930 82292 16942
rect 82684 17442 83188 17444
rect 82684 17390 83134 17442
rect 83186 17390 83188 17442
rect 82684 17388 83188 17390
rect 82684 16996 82740 17388
rect 83132 17378 83188 17388
rect 83244 17220 83300 17230
rect 83244 17106 83300 17164
rect 83244 17054 83246 17106
rect 83298 17054 83300 17106
rect 83244 17042 83300 17054
rect 82684 16902 82740 16940
rect 82796 16884 82852 16894
rect 82572 16658 82628 16670
rect 82572 16606 82574 16658
rect 82626 16606 82628 16658
rect 82124 16436 82180 16446
rect 82124 16210 82180 16380
rect 82124 16158 82126 16210
rect 82178 16158 82180 16210
rect 82124 16146 82180 16158
rect 82572 15652 82628 16606
rect 82572 15586 82628 15596
rect 82684 15874 82740 15886
rect 82684 15822 82686 15874
rect 82738 15822 82740 15874
rect 82684 15148 82740 15822
rect 82012 15092 82292 15148
rect 81788 14578 81844 14588
rect 81900 14308 81956 14318
rect 81900 13524 81956 14252
rect 81900 13458 81956 13468
rect 81676 11564 82180 11620
rect 81564 11218 81620 11228
rect 81900 11394 81956 11406
rect 81900 11342 81902 11394
rect 81954 11342 81956 11394
rect 80444 11172 80500 11182
rect 80444 10948 80500 11116
rect 81276 11004 81540 11014
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81276 10938 81540 10948
rect 80444 10834 80500 10892
rect 80444 10782 80446 10834
rect 80498 10782 80500 10834
rect 80444 10770 80500 10782
rect 81452 10836 81508 10846
rect 81228 10612 81284 10622
rect 81116 10556 81228 10612
rect 81004 10164 81060 10174
rect 80668 9940 80724 9950
rect 80668 9846 80724 9884
rect 80332 9762 80388 9772
rect 80108 9314 80164 9324
rect 80444 9266 80500 9278
rect 80444 9214 80446 9266
rect 80498 9214 80500 9266
rect 80108 9156 80164 9166
rect 79996 9154 80164 9156
rect 79996 9102 80110 9154
rect 80162 9102 80164 9154
rect 79996 9100 80164 9102
rect 80108 9090 80164 9100
rect 80332 9044 80388 9054
rect 80220 9042 80388 9044
rect 80220 8990 80334 9042
rect 80386 8990 80388 9042
rect 80220 8988 80388 8990
rect 80220 8596 80276 8988
rect 80332 8978 80388 8988
rect 79772 7522 79828 7532
rect 80108 8540 80276 8596
rect 79436 7310 79438 7362
rect 79490 7310 79492 7362
rect 79436 7140 79492 7310
rect 79436 7074 79492 7084
rect 80108 7028 80164 8540
rect 80220 8372 80276 8382
rect 80444 8372 80500 9214
rect 80220 8370 80500 8372
rect 80220 8318 80222 8370
rect 80274 8318 80500 8370
rect 80220 8316 80500 8318
rect 80780 9042 80836 9054
rect 80780 8990 80782 9042
rect 80834 8990 80836 9042
rect 80220 8306 80276 8316
rect 80668 7364 80724 7374
rect 80108 6972 80276 7028
rect 80108 6804 80164 6814
rect 79996 6802 80164 6804
rect 79996 6750 80110 6802
rect 80162 6750 80164 6802
rect 79996 6748 80164 6750
rect 79548 6692 79604 6702
rect 79996 6692 80052 6748
rect 80108 6738 80164 6748
rect 79548 6690 80052 6692
rect 79548 6638 79550 6690
rect 79602 6638 80052 6690
rect 79548 6636 80052 6638
rect 79548 6626 79604 6636
rect 80108 6580 80164 6590
rect 79324 6412 79716 6468
rect 79436 6132 79492 6142
rect 79436 6038 79492 6076
rect 79212 5182 79214 5234
rect 79266 5182 79268 5234
rect 79212 5170 79268 5182
rect 79660 5122 79716 6412
rect 79660 5070 79662 5122
rect 79714 5070 79716 5122
rect 79100 4676 79156 4686
rect 79100 4450 79156 4620
rect 79100 4398 79102 4450
rect 79154 4398 79156 4450
rect 79100 4386 79156 4398
rect 77980 3714 78036 3724
rect 79100 4116 79156 4126
rect 78988 3668 79044 3678
rect 78988 3574 79044 3612
rect 77980 3556 78036 3566
rect 77868 3554 78036 3556
rect 77868 3502 77982 3554
rect 78034 3502 78036 3554
rect 77868 3500 78036 3502
rect 77980 3490 78036 3500
rect 79100 800 79156 4060
rect 79660 3388 79716 5070
rect 79772 6466 79828 6478
rect 79772 6414 79774 6466
rect 79826 6414 79828 6466
rect 79772 4228 79828 6414
rect 79772 4162 79828 4172
rect 80108 4226 80164 6524
rect 80220 5012 80276 6972
rect 80332 6018 80388 6030
rect 80332 5966 80334 6018
rect 80386 5966 80388 6018
rect 80332 5234 80388 5966
rect 80668 5684 80724 7308
rect 80668 5618 80724 5628
rect 80332 5182 80334 5234
rect 80386 5182 80388 5234
rect 80332 5170 80388 5182
rect 80220 4946 80276 4956
rect 80108 4174 80110 4226
rect 80162 4174 80164 4226
rect 80108 4162 80164 4174
rect 80444 4900 80500 4910
rect 79660 3332 79828 3388
rect 79772 2884 79828 3332
rect 79772 2818 79828 2828
rect 80444 800 80500 4844
rect 80780 3554 80836 8990
rect 81004 8260 81060 10108
rect 81116 9268 81172 10556
rect 81228 10546 81284 10556
rect 81452 10164 81508 10780
rect 81900 10500 81956 11342
rect 81452 9826 81508 10108
rect 81452 9774 81454 9826
rect 81506 9774 81508 9826
rect 81452 9762 81508 9774
rect 81676 10498 81956 10500
rect 81676 10446 81902 10498
rect 81954 10446 81956 10498
rect 81676 10444 81956 10446
rect 81276 9436 81540 9446
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81276 9370 81540 9380
rect 81228 9268 81284 9278
rect 81116 9266 81284 9268
rect 81116 9214 81230 9266
rect 81282 9214 81284 9266
rect 81116 9212 81284 9214
rect 81228 9202 81284 9212
rect 81452 8932 81508 8942
rect 81452 8838 81508 8876
rect 81004 8166 81060 8204
rect 81452 8258 81508 8270
rect 81452 8206 81454 8258
rect 81506 8206 81508 8258
rect 81116 8148 81172 8158
rect 80780 3502 80782 3554
rect 80834 3502 80836 3554
rect 80780 3490 80836 3502
rect 81004 7028 81060 7038
rect 81004 3442 81060 6972
rect 81116 6804 81172 8092
rect 81452 8148 81508 8206
rect 81452 8082 81508 8092
rect 81276 7868 81540 7878
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81276 7802 81540 7812
rect 81564 7476 81620 7486
rect 81676 7476 81732 10444
rect 81900 10434 81956 10444
rect 81900 10164 81956 10174
rect 81900 9938 81956 10108
rect 81900 9886 81902 9938
rect 81954 9886 81956 9938
rect 81900 9874 81956 9886
rect 81900 9044 81956 9054
rect 81564 7474 81732 7476
rect 81564 7422 81566 7474
rect 81618 7422 81732 7474
rect 81564 7420 81732 7422
rect 81788 9042 81956 9044
rect 81788 8990 81902 9042
rect 81954 8990 81956 9042
rect 81788 8988 81956 8990
rect 81564 7410 81620 7420
rect 81788 7364 81844 8988
rect 81900 8978 81956 8988
rect 81900 8260 81956 8270
rect 82124 8260 82180 11564
rect 82236 10612 82292 15092
rect 82236 10546 82292 10556
rect 82460 15092 82740 15148
rect 82796 15092 82852 16828
rect 83356 16772 83412 21756
rect 84028 20020 84084 22876
rect 84140 22484 84196 22494
rect 84140 22390 84196 22428
rect 85260 22484 85316 22494
rect 85316 22428 85540 22484
rect 85260 22390 85316 22428
rect 85484 22370 85540 22428
rect 85484 22318 85486 22370
rect 85538 22318 85540 22370
rect 85484 22306 85540 22318
rect 84028 19954 84084 19964
rect 84700 22260 84756 22270
rect 83692 18676 83748 18686
rect 83468 18452 83524 18462
rect 83468 17780 83524 18396
rect 83468 17714 83524 17724
rect 83580 16884 83636 16894
rect 83580 16790 83636 16828
rect 83468 16772 83524 16782
rect 83356 16716 83468 16772
rect 83468 16706 83524 16716
rect 83132 15876 83188 15886
rect 83132 15782 83188 15820
rect 83580 15876 83636 15886
rect 83580 15782 83636 15820
rect 83468 15428 83524 15438
rect 82460 10164 82516 15092
rect 82572 14644 82628 14654
rect 82628 14588 82740 14644
rect 82572 14578 82628 14588
rect 82684 14530 82740 14588
rect 82684 14478 82686 14530
rect 82738 14478 82740 14530
rect 82684 14466 82740 14478
rect 82572 14420 82628 14430
rect 82572 13746 82628 14364
rect 82796 13748 82852 15036
rect 83020 15202 83076 15214
rect 83020 15150 83022 15202
rect 83074 15150 83076 15202
rect 83020 14420 83076 15150
rect 83468 15148 83524 15372
rect 83468 15092 83636 15148
rect 83132 14644 83188 14654
rect 83132 14550 83188 14588
rect 83020 14354 83076 14364
rect 83580 14196 83636 15092
rect 83580 14130 83636 14140
rect 83580 13972 83636 13982
rect 82572 13694 82574 13746
rect 82626 13694 82628 13746
rect 82572 13682 82628 13694
rect 82684 13692 82852 13748
rect 82908 13746 82964 13758
rect 82908 13694 82910 13746
rect 82962 13694 82964 13746
rect 82460 10098 82516 10108
rect 82348 10052 82404 10062
rect 82348 9826 82404 9996
rect 82348 9774 82350 9826
rect 82402 9774 82404 9826
rect 82348 9762 82404 9774
rect 82460 9828 82516 9838
rect 81900 8258 82180 8260
rect 81900 8206 81902 8258
rect 81954 8206 82180 8258
rect 81900 8204 82180 8206
rect 82236 8372 82292 8382
rect 82236 8258 82292 8316
rect 82236 8206 82238 8258
rect 82290 8206 82292 8258
rect 81900 8194 81956 8204
rect 82124 8036 82180 8046
rect 81116 6738 81172 6748
rect 81676 7308 81844 7364
rect 82012 8034 82180 8036
rect 82012 7982 82126 8034
rect 82178 7982 82180 8034
rect 82012 7980 82180 7982
rect 81116 6580 81172 6590
rect 81116 6486 81172 6524
rect 81276 6300 81540 6310
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81276 6234 81540 6244
rect 81676 5794 81732 7308
rect 81788 6468 81844 6478
rect 81788 6374 81844 6412
rect 81676 5742 81678 5794
rect 81730 5742 81732 5794
rect 81676 5730 81732 5742
rect 81276 4732 81540 4742
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81276 4666 81540 4676
rect 81116 4452 81172 4462
rect 81116 3554 81172 4396
rect 81116 3502 81118 3554
rect 81170 3502 81172 3554
rect 81116 3490 81172 3502
rect 81788 3668 81844 3678
rect 81004 3390 81006 3442
rect 81058 3390 81060 3442
rect 81004 3378 81060 3390
rect 81276 3164 81540 3174
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81276 3098 81540 3108
rect 80556 2884 80612 2894
rect 80556 980 80612 2828
rect 80556 914 80612 924
rect 81788 800 81844 3612
rect 82012 3554 82068 7980
rect 82124 7970 82180 7980
rect 82124 7476 82180 7486
rect 82124 5906 82180 7420
rect 82236 6690 82292 8206
rect 82348 6804 82404 6814
rect 82348 6710 82404 6748
rect 82236 6638 82238 6690
rect 82290 6638 82292 6690
rect 82236 6626 82292 6638
rect 82460 6690 82516 9772
rect 82572 9604 82628 9614
rect 82572 9510 82628 9548
rect 82684 9042 82740 13692
rect 82796 13524 82852 13534
rect 82796 12852 82852 13468
rect 82908 13188 82964 13694
rect 83468 13412 83524 13422
rect 82908 13132 83300 13188
rect 82796 12758 82852 12796
rect 83132 12962 83188 12974
rect 83132 12910 83134 12962
rect 83186 12910 83188 12962
rect 83020 12178 83076 12190
rect 83020 12126 83022 12178
rect 83074 12126 83076 12178
rect 82908 10612 82964 10622
rect 82908 10518 82964 10556
rect 82908 9716 82964 9726
rect 82908 9622 82964 9660
rect 82684 8990 82686 9042
rect 82738 8990 82740 9042
rect 82684 7924 82740 8990
rect 82908 9156 82964 9166
rect 82908 8258 82964 9100
rect 83020 8820 83076 12126
rect 83132 11956 83188 12910
rect 83244 12740 83300 13132
rect 83244 12290 83300 12684
rect 83468 12738 83524 13356
rect 83468 12686 83470 12738
rect 83522 12686 83524 12738
rect 83468 12674 83524 12686
rect 83244 12238 83246 12290
rect 83298 12238 83300 12290
rect 83244 12180 83300 12238
rect 83244 12114 83300 12124
rect 83132 11890 83188 11900
rect 83468 11844 83524 11854
rect 83244 10388 83300 10398
rect 83244 9826 83300 10332
rect 83244 9774 83246 9826
rect 83298 9774 83300 9826
rect 83244 9762 83300 9774
rect 83356 9602 83412 9614
rect 83356 9550 83358 9602
rect 83410 9550 83412 9602
rect 83356 9154 83412 9550
rect 83356 9102 83358 9154
rect 83410 9102 83412 9154
rect 83356 9090 83412 9102
rect 83132 8820 83188 8830
rect 83020 8764 83132 8820
rect 83132 8754 83188 8764
rect 83468 8372 83524 11788
rect 83580 11396 83636 13916
rect 83580 10948 83636 11340
rect 83580 10882 83636 10892
rect 83580 9828 83636 9838
rect 83580 9734 83636 9772
rect 82908 8206 82910 8258
rect 82962 8206 82964 8258
rect 82908 8194 82964 8206
rect 83244 8316 83524 8372
rect 83244 8146 83300 8316
rect 83244 8094 83246 8146
rect 83298 8094 83300 8146
rect 83244 8082 83300 8094
rect 82684 7586 82740 7868
rect 82684 7534 82686 7586
rect 82738 7534 82740 7586
rect 82684 7476 82740 7534
rect 82460 6638 82462 6690
rect 82514 6638 82516 6690
rect 82460 6626 82516 6638
rect 82572 7140 82628 7150
rect 82124 5854 82126 5906
rect 82178 5854 82180 5906
rect 82124 5842 82180 5854
rect 82460 5012 82516 5022
rect 82572 5012 82628 7084
rect 82460 5010 82628 5012
rect 82460 4958 82462 5010
rect 82514 4958 82628 5010
rect 82460 4956 82628 4958
rect 82348 4900 82404 4910
rect 82348 4450 82404 4844
rect 82348 4398 82350 4450
rect 82402 4398 82404 4450
rect 82348 4386 82404 4398
rect 82460 4116 82516 4956
rect 82684 4340 82740 7420
rect 83468 6916 83524 8316
rect 83468 6850 83524 6860
rect 83580 9044 83636 9054
rect 82796 5796 82852 5806
rect 82796 5702 82852 5740
rect 82908 5124 82964 5134
rect 82908 5030 82964 5068
rect 83244 5124 83300 5134
rect 83244 5030 83300 5068
rect 83580 5122 83636 8988
rect 83580 5070 83582 5122
rect 83634 5070 83636 5122
rect 83580 5058 83636 5070
rect 83356 4898 83412 4910
rect 83356 4846 83358 4898
rect 83410 4846 83412 4898
rect 83132 4676 83188 4686
rect 82908 4340 82964 4350
rect 82684 4338 82964 4340
rect 82684 4286 82910 4338
rect 82962 4286 82964 4338
rect 82684 4284 82964 4286
rect 82908 4274 82964 4284
rect 82460 4050 82516 4060
rect 83020 3668 83076 3678
rect 83020 3574 83076 3612
rect 82012 3502 82014 3554
rect 82066 3502 82068 3554
rect 82012 3490 82068 3502
rect 83132 800 83188 4620
rect 83356 4564 83412 4846
rect 83692 4900 83748 18620
rect 83916 18452 83972 18462
rect 83916 17108 83972 18396
rect 83916 17014 83972 17052
rect 84028 18340 84084 18350
rect 84476 18340 84532 18350
rect 84028 18338 84476 18340
rect 84028 18286 84030 18338
rect 84082 18286 84476 18338
rect 84028 18284 84476 18286
rect 84028 16884 84084 18284
rect 84476 18246 84532 18284
rect 84252 17780 84308 17790
rect 84252 17686 84308 17724
rect 84364 17444 84420 17454
rect 84364 17350 84420 17388
rect 84028 16818 84084 16828
rect 84140 16322 84196 16334
rect 84140 16270 84142 16322
rect 84194 16270 84196 16322
rect 84140 16210 84196 16270
rect 84140 16158 84142 16210
rect 84194 16158 84196 16210
rect 83916 15202 83972 15214
rect 83916 15150 83918 15202
rect 83970 15150 83972 15202
rect 83916 15148 83972 15150
rect 83804 15092 83972 15148
rect 83804 13076 83860 15092
rect 84028 14306 84084 14318
rect 84028 14254 84030 14306
rect 84082 14254 84084 14306
rect 84028 13860 84084 14254
rect 84028 13794 84084 13804
rect 83916 13746 83972 13758
rect 83916 13694 83918 13746
rect 83970 13694 83972 13746
rect 83916 13524 83972 13694
rect 83916 13458 83972 13468
rect 83804 12404 83860 13020
rect 83916 12404 83972 12414
rect 83804 12348 83916 12404
rect 83916 12338 83972 12348
rect 83804 11956 83860 11966
rect 83804 10610 83860 11900
rect 84140 11620 84196 16158
rect 84588 15874 84644 15886
rect 84588 15822 84590 15874
rect 84642 15822 84644 15874
rect 84252 14084 84308 14094
rect 84588 14084 84644 15822
rect 84700 15876 84756 22204
rect 86156 22148 86212 22988
rect 86380 22708 86436 23214
rect 86716 23154 86772 23166
rect 86716 23102 86718 23154
rect 86770 23102 86772 23154
rect 86380 22642 86436 22652
rect 86492 23042 86548 23054
rect 86492 22990 86494 23042
rect 86546 22990 86548 23042
rect 86268 22372 86324 22382
rect 86492 22372 86548 22990
rect 86716 22932 86772 23102
rect 86716 22866 86772 22876
rect 86268 22370 86548 22372
rect 86268 22318 86270 22370
rect 86322 22318 86548 22370
rect 86268 22316 86548 22318
rect 86268 22306 86324 22316
rect 86156 22092 86324 22148
rect 86156 21698 86212 21710
rect 86156 21646 86158 21698
rect 86210 21646 86212 21698
rect 85260 20578 85316 20590
rect 85260 20526 85262 20578
rect 85314 20526 85316 20578
rect 85260 19348 85316 20526
rect 86044 20132 86100 20142
rect 86156 20132 86212 21646
rect 86268 21588 86324 22092
rect 86492 21812 86548 21822
rect 86828 21812 86884 23772
rect 86492 21810 86884 21812
rect 86492 21758 86494 21810
rect 86546 21758 86830 21810
rect 86882 21758 86884 21810
rect 86492 21756 86884 21758
rect 86492 21746 86548 21756
rect 86268 21532 86548 21588
rect 86268 20804 86324 20814
rect 86268 20242 86324 20748
rect 86268 20190 86270 20242
rect 86322 20190 86324 20242
rect 86268 20178 86324 20190
rect 86044 20130 86212 20132
rect 86044 20078 86046 20130
rect 86098 20078 86212 20130
rect 86044 20076 86212 20078
rect 85260 19282 85316 19292
rect 85372 19906 85428 19918
rect 85372 19854 85374 19906
rect 85426 19854 85428 19906
rect 85036 19012 85092 19022
rect 85036 19010 85316 19012
rect 85036 18958 85038 19010
rect 85090 18958 85316 19010
rect 85036 18956 85316 18958
rect 85036 18946 85092 18956
rect 84812 18564 84868 18574
rect 84812 15988 84868 18508
rect 85036 18340 85092 18350
rect 84924 18338 85092 18340
rect 84924 18286 85038 18338
rect 85090 18286 85092 18338
rect 84924 18284 85092 18286
rect 84924 16322 84980 18284
rect 85036 18274 85092 18284
rect 85148 17444 85204 17454
rect 85148 17350 85204 17388
rect 84924 16270 84926 16322
rect 84978 16270 84980 16322
rect 84924 16258 84980 16270
rect 84812 15932 84980 15988
rect 84700 15820 84868 15876
rect 84812 14756 84868 15820
rect 84700 14644 84756 14654
rect 84700 14530 84756 14588
rect 84700 14478 84702 14530
rect 84754 14478 84756 14530
rect 84700 14466 84756 14478
rect 84588 14028 84756 14084
rect 84252 13748 84308 14028
rect 84700 13972 84756 14028
rect 84700 13906 84756 13916
rect 84588 13860 84644 13870
rect 84252 13682 84308 13692
rect 84476 13858 84644 13860
rect 84476 13806 84590 13858
rect 84642 13806 84644 13858
rect 84476 13804 84644 13806
rect 84252 12964 84308 12974
rect 84252 12850 84308 12908
rect 84252 12798 84254 12850
rect 84306 12798 84308 12850
rect 84252 12786 84308 12798
rect 84476 12852 84532 13804
rect 84588 13794 84644 13804
rect 84588 13636 84644 13646
rect 84812 13636 84868 14700
rect 84644 13580 84868 13636
rect 84588 13570 84644 13580
rect 84364 12292 84420 12302
rect 84476 12292 84532 12796
rect 84364 12290 84532 12292
rect 84364 12238 84366 12290
rect 84418 12238 84532 12290
rect 84364 12236 84532 12238
rect 84812 12964 84868 12974
rect 84924 12964 84980 15932
rect 85148 15876 85204 15886
rect 85148 15782 85204 15820
rect 84868 12908 84980 12964
rect 85148 15652 85204 15662
rect 84364 12226 84420 12236
rect 84140 11554 84196 11564
rect 84252 12180 84308 12190
rect 84140 11396 84196 11406
rect 84140 11302 84196 11340
rect 84028 11282 84084 11294
rect 84028 11230 84030 11282
rect 84082 11230 84084 11282
rect 83916 10836 83972 10846
rect 83916 10742 83972 10780
rect 83804 10558 83806 10610
rect 83858 10558 83860 10610
rect 83804 8484 83860 10558
rect 83916 10612 83972 10622
rect 83916 10386 83972 10556
rect 83916 10334 83918 10386
rect 83970 10334 83972 10386
rect 83916 10322 83972 10334
rect 83804 8418 83860 8428
rect 83916 9716 83972 9726
rect 83916 7140 83972 9660
rect 84028 8708 84084 11230
rect 84028 8652 84196 8708
rect 83916 7074 83972 7084
rect 84028 8372 84084 8382
rect 84028 8258 84084 8316
rect 84028 8206 84030 8258
rect 84082 8206 84084 8258
rect 84028 6804 84084 8206
rect 84140 8036 84196 8652
rect 84252 8258 84308 12124
rect 84700 12178 84756 12190
rect 84700 12126 84702 12178
rect 84754 12126 84756 12178
rect 84700 12068 84756 12126
rect 84700 12002 84756 12012
rect 84588 11844 84644 11854
rect 84476 11620 84532 11630
rect 84476 11508 84532 11564
rect 84364 11452 84532 11508
rect 84364 11396 84420 11452
rect 84364 11330 84420 11340
rect 84476 11284 84532 11294
rect 84476 11190 84532 11228
rect 84476 10724 84532 10734
rect 84364 10722 84532 10724
rect 84364 10670 84478 10722
rect 84530 10670 84532 10722
rect 84364 10668 84532 10670
rect 84364 10500 84420 10668
rect 84476 10658 84532 10668
rect 84588 10722 84644 11788
rect 84812 11394 84868 12908
rect 84924 12404 84980 12414
rect 85148 12404 85204 15596
rect 85260 15204 85316 18956
rect 85372 18340 85428 19854
rect 85708 19906 85764 19918
rect 85708 19854 85710 19906
rect 85762 19854 85764 19906
rect 85708 19458 85764 19854
rect 85708 19406 85710 19458
rect 85762 19406 85764 19458
rect 85484 19012 85540 19022
rect 85484 18918 85540 18956
rect 85372 18274 85428 18284
rect 85484 18338 85540 18350
rect 85484 18286 85486 18338
rect 85538 18286 85540 18338
rect 85372 17668 85428 17678
rect 85372 17574 85428 17612
rect 85484 16884 85540 18286
rect 85708 18228 85764 19406
rect 85820 19010 85876 19022
rect 85820 18958 85822 19010
rect 85874 18958 85876 19010
rect 85820 18676 85876 18958
rect 85820 18610 85876 18620
rect 85820 18452 85876 18462
rect 85820 18358 85876 18396
rect 85708 18172 85988 18228
rect 85596 17668 85652 17678
rect 85596 17666 85764 17668
rect 85596 17614 85598 17666
rect 85650 17614 85764 17666
rect 85596 17612 85764 17614
rect 85596 17602 85652 17612
rect 85484 16818 85540 16828
rect 85708 16660 85764 17612
rect 85820 17442 85876 17454
rect 85820 17390 85822 17442
rect 85874 17390 85876 17442
rect 85820 16884 85876 17390
rect 85932 17220 85988 18172
rect 86044 17780 86100 20076
rect 86380 20018 86436 20030
rect 86380 19966 86382 20018
rect 86434 19966 86436 20018
rect 86380 19458 86436 19966
rect 86380 19406 86382 19458
rect 86434 19406 86436 19458
rect 86380 19394 86436 19406
rect 86268 19348 86324 19358
rect 86268 19254 86324 19292
rect 86156 19012 86212 19022
rect 86156 18674 86212 18956
rect 86156 18622 86158 18674
rect 86210 18622 86212 18674
rect 86156 18610 86212 18622
rect 86380 18452 86436 18462
rect 86380 18358 86436 18396
rect 86044 17666 86100 17724
rect 86044 17614 86046 17666
rect 86098 17614 86100 17666
rect 86044 17602 86100 17614
rect 86268 18338 86324 18350
rect 86268 18286 86270 18338
rect 86322 18286 86324 18338
rect 86268 17668 86324 18286
rect 86268 17602 86324 17612
rect 85932 17154 85988 17164
rect 86380 17444 86436 17454
rect 86492 17444 86548 21532
rect 86828 20244 86884 21756
rect 86940 23154 86996 23166
rect 86940 23102 86942 23154
rect 86994 23102 86996 23154
rect 86940 21812 86996 23102
rect 87388 23042 87444 23054
rect 87388 22990 87390 23042
rect 87442 22990 87444 23042
rect 87388 22932 87444 22990
rect 87388 22866 87444 22876
rect 86940 21746 86996 21756
rect 87164 21700 87220 21710
rect 87164 21606 87220 21644
rect 87836 21588 87892 21598
rect 87724 21586 87892 21588
rect 87724 21534 87838 21586
rect 87890 21534 87892 21586
rect 87724 21532 87892 21534
rect 87612 20804 87668 20814
rect 87612 20710 87668 20748
rect 86940 20244 86996 20254
rect 86828 20242 86996 20244
rect 86828 20190 86942 20242
rect 86994 20190 86996 20242
rect 86828 20188 86996 20190
rect 86940 20178 86996 20188
rect 87276 20130 87332 20142
rect 87276 20078 87278 20130
rect 87330 20078 87332 20130
rect 86604 20020 86660 20030
rect 86604 20018 86772 20020
rect 86604 19966 86606 20018
rect 86658 19966 86772 20018
rect 86604 19964 86772 19966
rect 86604 19954 86660 19964
rect 86604 19460 86660 19470
rect 86604 19012 86660 19404
rect 86716 19346 86772 19964
rect 87276 19460 87332 20078
rect 87276 19394 87332 19404
rect 86716 19294 86718 19346
rect 86770 19294 86772 19346
rect 86716 19282 86772 19294
rect 86828 19348 86884 19358
rect 86828 19234 86884 19292
rect 87276 19236 87332 19246
rect 86828 19182 86830 19234
rect 86882 19182 86884 19234
rect 86828 19170 86884 19182
rect 86940 19234 87668 19236
rect 86940 19182 87278 19234
rect 87330 19182 87668 19234
rect 86940 19180 87668 19182
rect 86604 18918 86660 18956
rect 86828 18452 86884 18462
rect 86940 18452 86996 19180
rect 87276 19170 87332 19180
rect 87612 19124 87668 19180
rect 87724 19124 87780 21532
rect 87836 21522 87892 21532
rect 88060 19236 88116 28700
rect 88172 25508 88228 25518
rect 88172 25414 88228 25452
rect 88620 22146 88676 22158
rect 88620 22094 88622 22146
rect 88674 22094 88676 22146
rect 88620 22036 88676 22094
rect 88284 21980 88676 22036
rect 88284 21586 88340 21980
rect 88396 21812 88452 21822
rect 88396 21718 88452 21756
rect 88508 21700 88564 21710
rect 88508 21606 88564 21644
rect 88284 21534 88286 21586
rect 88338 21534 88340 21586
rect 88060 19180 88228 19236
rect 87612 19122 87780 19124
rect 87612 19070 87614 19122
rect 87666 19070 87780 19122
rect 87612 19068 87780 19070
rect 87612 19058 87668 19068
rect 87836 19012 87892 19022
rect 86828 18450 86996 18452
rect 86828 18398 86830 18450
rect 86882 18398 86996 18450
rect 86828 18396 86996 18398
rect 86828 18386 86884 18396
rect 86940 17778 86996 18396
rect 87724 19010 87892 19012
rect 87724 18958 87838 19010
rect 87890 18958 87892 19010
rect 87724 18956 87892 18958
rect 86940 17726 86942 17778
rect 86994 17726 86996 17778
rect 86940 17714 86996 17726
rect 87164 18338 87220 18350
rect 87164 18286 87166 18338
rect 87218 18286 87220 18338
rect 87164 17668 87220 18286
rect 87724 18004 87780 18956
rect 87836 18946 87892 18956
rect 87948 19010 88004 19022
rect 87948 18958 87950 19010
rect 88002 18958 88004 19010
rect 87948 18564 88004 18958
rect 88060 19012 88116 19022
rect 88060 18918 88116 18956
rect 88172 18788 88228 19180
rect 87724 17938 87780 17948
rect 87836 18508 88004 18564
rect 88060 18732 88228 18788
rect 88284 18788 88340 21534
rect 88732 21588 88788 21598
rect 88732 20916 88788 21532
rect 88396 20914 88788 20916
rect 88396 20862 88734 20914
rect 88786 20862 88788 20914
rect 88396 20860 88788 20862
rect 88396 20802 88452 20860
rect 88732 20850 88788 20860
rect 88396 20750 88398 20802
rect 88450 20750 88452 20802
rect 88396 20738 88452 20750
rect 88620 19012 88676 19022
rect 87276 17668 87332 17678
rect 87164 17666 87332 17668
rect 87164 17614 87278 17666
rect 87330 17614 87332 17666
rect 87164 17612 87332 17614
rect 87276 17556 87332 17612
rect 87836 17666 87892 18508
rect 87948 18338 88004 18350
rect 87948 18286 87950 18338
rect 88002 18286 88004 18338
rect 87948 18004 88004 18286
rect 87948 17938 88004 17948
rect 87836 17614 87838 17666
rect 87890 17614 87892 17666
rect 87836 17602 87892 17614
rect 87948 17668 88004 17678
rect 87948 17574 88004 17612
rect 87276 17490 87332 17500
rect 86380 17442 86548 17444
rect 86380 17390 86382 17442
rect 86434 17390 86548 17442
rect 86380 17388 86548 17390
rect 87388 17444 87444 17454
rect 86268 16884 86324 16894
rect 85820 16882 86324 16884
rect 85820 16830 86270 16882
rect 86322 16830 86324 16882
rect 85820 16828 86324 16830
rect 86268 16818 86324 16828
rect 86380 16660 86436 17388
rect 87388 17108 87444 17388
rect 85708 16604 86436 16660
rect 87052 17106 87444 17108
rect 87052 17054 87390 17106
rect 87442 17054 87444 17106
rect 87052 17052 87444 17054
rect 87052 16882 87108 17052
rect 87052 16830 87054 16882
rect 87106 16830 87108 16882
rect 85260 15138 85316 15148
rect 85596 15874 85652 15886
rect 85596 15822 85598 15874
rect 85650 15822 85652 15874
rect 85260 14644 85316 14654
rect 85260 14308 85316 14588
rect 85260 14242 85316 14252
rect 84924 12402 85204 12404
rect 84924 12350 84926 12402
rect 84978 12350 85204 12402
rect 84924 12348 85204 12350
rect 85260 13972 85316 13982
rect 84924 12338 84980 12348
rect 85148 12068 85204 12078
rect 85148 11788 85204 12012
rect 84812 11342 84814 11394
rect 84866 11342 84868 11394
rect 84812 11330 84868 11342
rect 84924 11732 85204 11788
rect 84588 10670 84590 10722
rect 84642 10670 84644 10722
rect 84588 10658 84644 10670
rect 84924 11172 84980 11732
rect 84924 10724 84980 11116
rect 85036 11396 85092 11406
rect 85036 10834 85092 11340
rect 85036 10782 85038 10834
rect 85090 10782 85092 10834
rect 85036 10770 85092 10782
rect 84924 10658 84980 10668
rect 84364 10434 84420 10444
rect 84924 10500 84980 10510
rect 84924 10498 85204 10500
rect 84924 10446 84926 10498
rect 84978 10446 85204 10498
rect 84924 10444 85204 10446
rect 84924 10434 84980 10444
rect 84476 10388 84532 10398
rect 84476 10294 84532 10332
rect 84588 9940 84644 9950
rect 84588 9826 84644 9884
rect 84588 9774 84590 9826
rect 84642 9774 84644 9826
rect 84588 9762 84644 9774
rect 85036 9714 85092 9726
rect 85036 9662 85038 9714
rect 85090 9662 85092 9714
rect 84476 9602 84532 9614
rect 84476 9550 84478 9602
rect 84530 9550 84532 9602
rect 84476 9492 84532 9550
rect 84476 9426 84532 9436
rect 84700 9602 84756 9614
rect 84700 9550 84702 9602
rect 84754 9550 84756 9602
rect 84588 9156 84644 9166
rect 84252 8206 84254 8258
rect 84306 8206 84308 8258
rect 84252 8194 84308 8206
rect 84476 8372 84532 8382
rect 84364 8036 84420 8046
rect 84140 8034 84420 8036
rect 84140 7982 84366 8034
rect 84418 7982 84420 8034
rect 84140 7980 84420 7982
rect 84364 7970 84420 7980
rect 84476 8034 84532 8316
rect 84476 7982 84478 8034
rect 84530 7982 84532 8034
rect 84476 7252 84532 7982
rect 84476 7186 84532 7196
rect 84588 7028 84644 9100
rect 84700 8596 84756 9550
rect 84700 8530 84756 8540
rect 84812 9604 84868 9614
rect 84812 8372 84868 9548
rect 85036 9380 85092 9662
rect 85036 9314 85092 9324
rect 84700 8316 85092 8372
rect 84700 8258 84756 8316
rect 84700 8206 84702 8258
rect 84754 8206 84756 8258
rect 84700 8194 84756 8206
rect 85036 8258 85092 8316
rect 85148 8370 85204 10444
rect 85148 8318 85150 8370
rect 85202 8318 85204 8370
rect 85148 8306 85204 8318
rect 85260 8372 85316 13916
rect 85484 11732 85540 11742
rect 85484 10610 85540 11676
rect 85484 10558 85486 10610
rect 85538 10558 85540 10610
rect 85484 10546 85540 10558
rect 85372 10500 85428 10510
rect 85372 8932 85428 10444
rect 85484 10052 85540 10062
rect 85484 9938 85540 9996
rect 85484 9886 85486 9938
rect 85538 9886 85540 9938
rect 85484 9874 85540 9886
rect 85484 8932 85540 8942
rect 85372 8930 85540 8932
rect 85372 8878 85486 8930
rect 85538 8878 85540 8930
rect 85372 8876 85540 8878
rect 85484 8866 85540 8876
rect 85260 8306 85316 8316
rect 85484 8484 85540 8494
rect 85036 8206 85038 8258
rect 85090 8206 85092 8258
rect 85036 8148 85092 8206
rect 85484 8258 85540 8428
rect 85484 8206 85486 8258
rect 85538 8206 85540 8258
rect 85484 8194 85540 8206
rect 85036 8082 85092 8092
rect 85148 8036 85204 8046
rect 84588 6972 84868 7028
rect 84476 6916 84532 6926
rect 83916 6748 84084 6804
rect 84364 6804 84420 6814
rect 83916 6580 83972 6748
rect 84140 6690 84196 6702
rect 84140 6638 84142 6690
rect 84194 6638 84196 6690
rect 84140 6580 84196 6638
rect 83916 6524 84084 6580
rect 83692 4834 83748 4844
rect 83356 4508 83748 4564
rect 83692 4450 83748 4508
rect 83692 4398 83694 4450
rect 83746 4398 83748 4450
rect 83692 4386 83748 4398
rect 84028 3332 84084 6524
rect 84140 6514 84196 6524
rect 84364 6578 84420 6748
rect 84364 6526 84366 6578
rect 84418 6526 84420 6578
rect 84364 6514 84420 6526
rect 84476 6580 84532 6860
rect 84476 6514 84532 6524
rect 84700 6802 84756 6814
rect 84700 6750 84702 6802
rect 84754 6750 84756 6802
rect 84700 6468 84756 6750
rect 84700 6402 84756 6412
rect 84140 6356 84196 6366
rect 84140 5122 84196 6300
rect 84812 6244 84868 6972
rect 85036 6356 85092 6366
rect 84140 5070 84142 5122
rect 84194 5070 84196 5122
rect 84140 5058 84196 5070
rect 84364 6188 84868 6244
rect 84924 6244 84980 6254
rect 84364 5010 84420 6188
rect 84924 5794 84980 6188
rect 84924 5742 84926 5794
rect 84978 5742 84980 5794
rect 84924 5730 84980 5742
rect 84364 4958 84366 5010
rect 84418 4958 84420 5010
rect 84364 4946 84420 4958
rect 85036 4676 85092 6300
rect 85148 5572 85204 7980
rect 85260 8034 85316 8046
rect 85260 7982 85262 8034
rect 85314 7982 85316 8034
rect 85260 7700 85316 7982
rect 85260 7634 85316 7644
rect 85484 6804 85540 6814
rect 85260 6692 85316 6702
rect 85260 5908 85316 6636
rect 85260 5906 85428 5908
rect 85260 5854 85262 5906
rect 85314 5854 85428 5906
rect 85260 5852 85428 5854
rect 85260 5842 85316 5852
rect 85148 5516 85316 5572
rect 85260 5122 85316 5516
rect 85372 5234 85428 5852
rect 85372 5182 85374 5234
rect 85426 5182 85428 5234
rect 85372 5170 85428 5182
rect 85260 5070 85262 5122
rect 85314 5070 85316 5122
rect 85260 5058 85316 5070
rect 85484 5124 85540 6748
rect 85596 6356 85652 15822
rect 85932 15876 85988 15886
rect 85932 15652 85988 15820
rect 86268 15764 86324 16604
rect 86940 16100 86996 16110
rect 86268 15698 86324 15708
rect 86380 16098 86996 16100
rect 86380 16046 86942 16098
rect 86994 16046 86996 16098
rect 86380 16044 86996 16046
rect 85932 15596 86212 15652
rect 86156 15316 86212 15596
rect 86268 15316 86324 15326
rect 86156 15260 86268 15316
rect 86268 15250 86324 15260
rect 86044 15202 86100 15214
rect 86044 15150 86046 15202
rect 86098 15150 86100 15202
rect 85820 14306 85876 14318
rect 85820 14254 85822 14306
rect 85874 14254 85876 14306
rect 85708 13748 85764 13758
rect 85708 13654 85764 13692
rect 85820 13188 85876 14254
rect 85932 13972 85988 13982
rect 85932 13878 85988 13916
rect 86044 13188 86100 15150
rect 86380 15092 86436 16044
rect 86940 16034 86996 16044
rect 86492 15874 86548 15886
rect 87052 15876 87108 16830
rect 86492 15822 86494 15874
rect 86546 15822 86548 15874
rect 86492 15148 86548 15822
rect 86828 15820 87108 15876
rect 87164 16210 87220 16222
rect 87164 16158 87166 16210
rect 87218 16158 87220 16210
rect 86828 15314 86884 15820
rect 86828 15262 86830 15314
rect 86882 15262 86884 15314
rect 86828 15250 86884 15262
rect 86492 15092 86772 15148
rect 86380 15026 86436 15036
rect 85820 13122 85876 13132
rect 85932 13132 86100 13188
rect 86156 14308 86212 14318
rect 85708 12404 85764 12414
rect 85708 12310 85764 12348
rect 85820 12292 85876 12302
rect 85820 12198 85876 12236
rect 85708 11954 85764 11966
rect 85708 11902 85710 11954
rect 85762 11902 85764 11954
rect 85708 10610 85764 11902
rect 85820 10836 85876 10846
rect 85932 10836 85988 13132
rect 86044 12962 86100 12974
rect 86044 12910 86046 12962
rect 86098 12910 86100 12962
rect 86044 11620 86100 12910
rect 86156 12292 86212 14252
rect 86268 14306 86324 14318
rect 86268 14254 86270 14306
rect 86322 14254 86324 14306
rect 86268 14196 86324 14254
rect 86268 14130 86324 14140
rect 86604 14084 86660 14094
rect 86492 13634 86548 13646
rect 86492 13582 86494 13634
rect 86546 13582 86548 13634
rect 86492 12964 86548 13582
rect 86492 12404 86548 12908
rect 86492 12338 86548 12348
rect 86156 12178 86212 12236
rect 86156 12126 86158 12178
rect 86210 12126 86212 12178
rect 86156 12114 86212 12126
rect 86044 11554 86100 11564
rect 86268 11396 86324 11406
rect 86268 11302 86324 11340
rect 85820 10834 85988 10836
rect 85820 10782 85822 10834
rect 85874 10782 85988 10834
rect 85820 10780 85988 10782
rect 86380 11284 86436 11294
rect 86380 10834 86436 11228
rect 86380 10782 86382 10834
rect 86434 10782 86436 10834
rect 85820 10770 85876 10780
rect 86380 10770 86436 10782
rect 85708 10558 85710 10610
rect 85762 10558 85764 10610
rect 85708 10546 85764 10558
rect 85820 10612 85876 10622
rect 85820 9210 85876 10556
rect 86044 10610 86100 10622
rect 86044 10558 86046 10610
rect 86098 10558 86100 10610
rect 86044 10276 86100 10558
rect 86044 10210 86100 10220
rect 86604 9940 86660 14028
rect 86380 9884 86660 9940
rect 86156 9826 86212 9838
rect 86156 9774 86158 9826
rect 86210 9774 86212 9826
rect 85932 9716 85988 9726
rect 85932 9622 85988 9660
rect 85820 9158 85822 9210
rect 85874 9158 85876 9210
rect 86156 9266 86212 9774
rect 86156 9214 86158 9266
rect 86210 9214 86212 9266
rect 86156 9202 86212 9214
rect 85820 9146 85876 9158
rect 85932 9154 85988 9166
rect 85932 9102 85934 9154
rect 85986 9102 85988 9154
rect 85932 9044 85988 9102
rect 86268 9044 86324 9054
rect 85820 8988 86212 9044
rect 85708 8146 85764 8158
rect 85708 8094 85710 8146
rect 85762 8094 85764 8146
rect 85708 6916 85764 8094
rect 85820 7364 85876 8988
rect 86156 8820 86212 8988
rect 86268 8950 86324 8988
rect 86380 8820 86436 9884
rect 86604 9716 86660 9726
rect 86604 9622 86660 9660
rect 86492 9604 86548 9614
rect 86492 9510 86548 9548
rect 86716 9492 86772 15092
rect 86828 14868 86884 14878
rect 86828 14530 86884 14812
rect 86828 14478 86830 14530
rect 86882 14478 86884 14530
rect 86828 14466 86884 14478
rect 86940 14644 86996 14654
rect 86940 13970 86996 14588
rect 87164 14308 87220 16158
rect 87276 15538 87332 17052
rect 87388 17042 87444 17052
rect 87388 16772 87444 16782
rect 87388 16322 87444 16716
rect 87388 16270 87390 16322
rect 87442 16270 87444 16322
rect 87388 16258 87444 16270
rect 87276 15486 87278 15538
rect 87330 15486 87332 15538
rect 87276 15474 87332 15486
rect 87948 16100 88004 16110
rect 87948 15538 88004 16044
rect 87948 15486 87950 15538
rect 88002 15486 88004 15538
rect 87948 15474 88004 15486
rect 87276 15316 87332 15326
rect 87276 15148 87332 15260
rect 88060 15316 88116 18732
rect 88284 18722 88340 18732
rect 88508 19010 88676 19012
rect 88508 18958 88622 19010
rect 88674 18958 88676 19010
rect 88508 18956 88676 18958
rect 88172 18452 88228 18462
rect 88172 17778 88228 18396
rect 88508 18004 88564 18956
rect 88620 18946 88676 18956
rect 88508 17938 88564 17948
rect 88172 17726 88174 17778
rect 88226 17726 88228 17778
rect 88172 17714 88228 17726
rect 88284 17780 88340 17790
rect 88284 17666 88340 17724
rect 88284 17614 88286 17666
rect 88338 17614 88340 17666
rect 88284 17602 88340 17614
rect 88620 17668 88676 17678
rect 88620 17556 88676 17612
rect 88732 17556 88788 17566
rect 88620 17554 88788 17556
rect 88620 17502 88734 17554
rect 88786 17502 88788 17554
rect 88620 17500 88788 17502
rect 88396 16772 88452 16782
rect 88396 16770 88564 16772
rect 88396 16718 88398 16770
rect 88450 16718 88564 16770
rect 88396 16716 88564 16718
rect 88396 16706 88452 16716
rect 88508 15876 88564 16716
rect 88620 16324 88676 17500
rect 88732 17490 88788 17500
rect 88844 16772 88900 43652
rect 89628 30436 89684 30446
rect 89180 29428 89236 29438
rect 88956 25508 89012 25518
rect 88956 25414 89012 25452
rect 89068 18116 89124 18126
rect 89068 17106 89124 18060
rect 89068 17054 89070 17106
rect 89122 17054 89124 17106
rect 89068 16996 89124 17054
rect 89068 16930 89124 16940
rect 88844 16716 89124 16772
rect 88732 16324 88788 16334
rect 88620 16268 88732 16324
rect 88732 16258 88788 16268
rect 88956 16210 89012 16222
rect 88956 16158 88958 16210
rect 89010 16158 89012 16210
rect 88844 16098 88900 16110
rect 88844 16046 88846 16098
rect 88898 16046 88900 16098
rect 88508 15820 88788 15876
rect 88172 15316 88228 15326
rect 88060 15314 88228 15316
rect 88060 15262 88174 15314
rect 88226 15262 88228 15314
rect 88060 15260 88228 15262
rect 87276 15092 87444 15148
rect 87164 14242 87220 14252
rect 87388 14756 87444 15092
rect 87388 13972 87444 14700
rect 86940 13918 86942 13970
rect 86994 13918 86996 13970
rect 86940 13906 86996 13918
rect 87052 13970 87444 13972
rect 87052 13918 87390 13970
rect 87442 13918 87444 13970
rect 87052 13916 87444 13918
rect 87052 12180 87108 13916
rect 87388 13906 87444 13916
rect 87500 13636 87556 13646
rect 87500 12852 87556 13580
rect 87948 13636 88004 13646
rect 87724 12852 87780 12862
rect 87500 12850 87780 12852
rect 87500 12798 87726 12850
rect 87778 12798 87780 12850
rect 87500 12796 87780 12798
rect 86828 12124 87108 12180
rect 86828 11732 86884 12124
rect 87276 12068 87332 12078
rect 87276 11974 87332 12012
rect 86828 9826 86884 11676
rect 86940 11956 86996 11966
rect 86940 11282 86996 11900
rect 86940 11230 86942 11282
rect 86994 11230 86996 11282
rect 86940 11218 86996 11230
rect 87724 11282 87780 12796
rect 87948 12738 88004 13580
rect 87948 12686 87950 12738
rect 88002 12686 88004 12738
rect 87948 12674 88004 12686
rect 88060 13634 88116 15260
rect 88172 15250 88228 15260
rect 88732 15314 88788 15820
rect 88732 15262 88734 15314
rect 88786 15262 88788 15314
rect 88732 15148 88788 15262
rect 88396 15092 88788 15148
rect 88844 15540 88900 16046
rect 88396 14644 88452 15092
rect 88396 14588 88676 14644
rect 88172 14530 88228 14542
rect 88172 14478 88174 14530
rect 88226 14478 88228 14530
rect 88172 14308 88228 14478
rect 88172 14242 88228 14252
rect 88060 13582 88062 13634
rect 88114 13582 88116 13634
rect 88060 12628 88116 13582
rect 88396 13188 88452 13198
rect 88284 13076 88340 13086
rect 88284 12962 88340 13020
rect 88284 12910 88286 12962
rect 88338 12910 88340 12962
rect 88284 12898 88340 12910
rect 88284 12740 88340 12750
rect 88060 12562 88116 12572
rect 88172 12684 88284 12740
rect 88060 12404 88116 12414
rect 88060 12310 88116 12348
rect 87724 11230 87726 11282
rect 87778 11230 87780 11282
rect 87724 11218 87780 11230
rect 86940 11060 86996 11070
rect 86940 10610 86996 11004
rect 86940 10558 86942 10610
rect 86994 10558 86996 10610
rect 86940 10546 86996 10558
rect 87388 10948 87444 10958
rect 87276 10500 87332 10510
rect 87276 10406 87332 10444
rect 86828 9774 86830 9826
rect 86882 9774 86884 9826
rect 86828 9762 86884 9774
rect 86716 9436 86884 9492
rect 86492 9156 86548 9166
rect 86492 9062 86548 9100
rect 86156 8764 86436 8820
rect 86604 9042 86660 9054
rect 86604 8990 86606 9042
rect 86658 8990 86660 9042
rect 86156 8484 86212 8494
rect 85932 8260 85988 8270
rect 85932 7698 85988 8204
rect 86156 8258 86212 8428
rect 86268 8372 86324 8410
rect 86604 8372 86660 8990
rect 86828 8484 86884 9436
rect 86828 8418 86884 8428
rect 86940 9380 86996 9390
rect 86268 8306 86324 8316
rect 86380 8316 86660 8372
rect 86940 8372 86996 9324
rect 87276 9156 87332 9166
rect 86156 8206 86158 8258
rect 86210 8206 86212 8258
rect 86156 8194 86212 8206
rect 86268 8146 86324 8158
rect 86268 8094 86270 8146
rect 86322 8094 86324 8146
rect 86044 8036 86100 8046
rect 86268 8036 86324 8094
rect 86100 7980 86324 8036
rect 86044 7970 86100 7980
rect 86380 7924 86436 8316
rect 86940 8306 86996 8316
rect 87052 9154 87332 9156
rect 87052 9102 87278 9154
rect 87330 9102 87332 9154
rect 87052 9100 87332 9102
rect 86492 8148 86548 8158
rect 86492 8054 86548 8092
rect 86716 8148 86772 8158
rect 86716 8146 86996 8148
rect 86716 8094 86718 8146
rect 86770 8094 86996 8146
rect 86716 8092 86996 8094
rect 86716 8082 86772 8092
rect 85932 7646 85934 7698
rect 85986 7646 85988 7698
rect 85932 7634 85988 7646
rect 86268 7868 86436 7924
rect 86604 8036 86660 8046
rect 85820 7298 85876 7308
rect 86156 7364 86212 7402
rect 86156 7298 86212 7308
rect 85708 6850 85764 6860
rect 86156 7140 86212 7150
rect 85932 6580 85988 6590
rect 85932 6486 85988 6524
rect 85596 6290 85652 6300
rect 86156 6244 86212 7084
rect 85932 6188 86212 6244
rect 85820 5908 85876 5918
rect 85820 5814 85876 5852
rect 85932 5684 85988 6188
rect 86268 6020 86324 7868
rect 86492 7812 86548 7822
rect 86492 7140 86548 7756
rect 86492 7074 86548 7084
rect 86604 6804 86660 7980
rect 86828 7924 86884 7934
rect 86716 7476 86772 7486
rect 86716 7382 86772 7420
rect 86828 7364 86884 7868
rect 86156 5964 86324 6020
rect 86380 6748 86660 6804
rect 86716 7252 86772 7262
rect 85820 5628 85988 5684
rect 86044 5906 86100 5918
rect 86044 5854 86046 5906
rect 86098 5854 86100 5906
rect 85596 5124 85652 5134
rect 85484 5122 85652 5124
rect 85484 5070 85598 5122
rect 85650 5070 85652 5122
rect 85484 5068 85652 5070
rect 85036 4610 85092 4620
rect 85484 4676 85540 5068
rect 85596 5058 85652 5068
rect 85484 4610 85540 4620
rect 85596 4898 85652 4910
rect 85596 4846 85598 4898
rect 85650 4846 85652 4898
rect 85596 4564 85652 4846
rect 85596 4498 85652 4508
rect 84028 3266 84084 3276
rect 84476 4452 84532 4462
rect 84476 800 84532 4396
rect 85484 4340 85540 4350
rect 85484 3556 85540 4284
rect 85484 3462 85540 3500
rect 85596 4228 85652 4238
rect 85596 3442 85652 4172
rect 85820 4226 85876 5628
rect 86044 4788 86100 5854
rect 85820 4174 85822 4226
rect 85874 4174 85876 4226
rect 85820 4162 85876 4174
rect 85932 4732 86100 4788
rect 85932 4004 85988 4732
rect 85820 3948 85988 4004
rect 86044 4564 86100 4574
rect 85820 3554 85876 3948
rect 85820 3502 85822 3554
rect 85874 3502 85876 3554
rect 85820 3490 85876 3502
rect 86044 3554 86100 4508
rect 86156 4340 86212 5964
rect 86268 5796 86324 5806
rect 86268 5702 86324 5740
rect 86156 4274 86212 4284
rect 86268 5572 86324 5582
rect 86268 4338 86324 5516
rect 86380 5124 86436 6748
rect 86604 6578 86660 6590
rect 86604 6526 86606 6578
rect 86658 6526 86660 6578
rect 86604 6356 86660 6526
rect 86604 6290 86660 6300
rect 86716 6132 86772 7196
rect 86604 6076 86772 6132
rect 86492 5908 86548 5918
rect 86492 5814 86548 5852
rect 86380 5058 86436 5068
rect 86492 4564 86548 4574
rect 86492 4470 86548 4508
rect 86604 4452 86660 6076
rect 86716 5906 86772 5918
rect 86716 5854 86718 5906
rect 86770 5854 86772 5906
rect 86716 5796 86772 5854
rect 86716 5730 86772 5740
rect 86716 5124 86772 5134
rect 86828 5124 86884 7308
rect 86940 6468 86996 8092
rect 87052 7700 87108 9100
rect 87276 9090 87332 9100
rect 87388 9154 87444 10892
rect 87836 10612 87892 10622
rect 87836 9826 87892 10556
rect 87836 9774 87838 9826
rect 87890 9774 87892 9826
rect 87836 9762 87892 9774
rect 87948 9714 88004 9726
rect 87948 9662 87950 9714
rect 88002 9662 88004 9714
rect 87612 9268 87668 9278
rect 87948 9268 88004 9662
rect 87668 9212 87780 9268
rect 87612 9202 87668 9212
rect 87388 9102 87390 9154
rect 87442 9102 87444 9154
rect 87388 9090 87444 9102
rect 87276 8818 87332 8830
rect 87276 8766 87278 8818
rect 87330 8766 87332 8818
rect 87164 8036 87220 8046
rect 87164 7942 87220 7980
rect 87052 7644 87220 7700
rect 87052 7474 87108 7486
rect 87052 7422 87054 7474
rect 87106 7422 87108 7474
rect 87052 7252 87108 7422
rect 87052 7186 87108 7196
rect 86940 6402 86996 6412
rect 87164 6244 87220 7644
rect 87276 7476 87332 8766
rect 87388 8372 87444 8382
rect 87388 8034 87444 8316
rect 87388 7982 87390 8034
rect 87442 7982 87444 8034
rect 87388 7924 87444 7982
rect 87388 7858 87444 7868
rect 87500 8146 87556 8158
rect 87500 8094 87502 8146
rect 87554 8094 87556 8146
rect 87388 7700 87444 7710
rect 87500 7700 87556 8094
rect 87388 7698 87668 7700
rect 87388 7646 87390 7698
rect 87442 7646 87668 7698
rect 87388 7644 87668 7646
rect 87388 7634 87444 7644
rect 87276 7420 87556 7476
rect 87164 6178 87220 6188
rect 87276 6692 87332 6702
rect 87164 6018 87220 6030
rect 87164 5966 87166 6018
rect 87218 5966 87220 6018
rect 86716 5122 86884 5124
rect 86716 5070 86718 5122
rect 86770 5070 86884 5122
rect 86716 5068 86884 5070
rect 86940 5906 86996 5918
rect 86940 5854 86942 5906
rect 86994 5854 86996 5906
rect 86716 5058 86772 5068
rect 86940 5012 86996 5854
rect 86940 4946 86996 4956
rect 87052 5796 87108 5806
rect 87052 5348 87108 5740
rect 87164 5684 87220 5966
rect 87276 6018 87332 6636
rect 87276 5966 87278 6018
rect 87330 5966 87332 6018
rect 87276 5954 87332 5966
rect 87164 5618 87220 5628
rect 86604 4386 86660 4396
rect 86268 4286 86270 4338
rect 86322 4286 86324 4338
rect 86268 4274 86324 4286
rect 86940 4340 86996 4350
rect 87052 4340 87108 5292
rect 87388 5012 87444 5022
rect 87276 5010 87444 5012
rect 87276 4958 87390 5010
rect 87442 4958 87444 5010
rect 87276 4956 87444 4958
rect 86940 4338 87108 4340
rect 86940 4286 86942 4338
rect 86994 4286 87108 4338
rect 86940 4284 87108 4286
rect 87164 4900 87220 4910
rect 87164 4338 87220 4844
rect 87276 4562 87332 4956
rect 87388 4946 87444 4956
rect 87276 4510 87278 4562
rect 87330 4510 87332 4562
rect 87276 4498 87332 4510
rect 87164 4286 87166 4338
rect 87218 4286 87220 4338
rect 86940 4274 86996 4284
rect 87164 4274 87220 4286
rect 87500 4338 87556 7420
rect 87612 6804 87668 7644
rect 87724 7252 87780 9212
rect 87724 7186 87780 7196
rect 87836 9212 88004 9268
rect 87724 6804 87780 6814
rect 87612 6748 87724 6804
rect 87724 6738 87780 6748
rect 87836 6692 87892 9212
rect 87948 9042 88004 9054
rect 87948 8990 87950 9042
rect 88002 8990 88004 9042
rect 87948 7474 88004 8990
rect 88172 8372 88228 12684
rect 88284 12674 88340 12684
rect 88284 10836 88340 10846
rect 88396 10836 88452 13132
rect 88508 12292 88564 12302
rect 88508 12198 88564 12236
rect 88508 11396 88564 11406
rect 88508 11302 88564 11340
rect 88284 10834 88452 10836
rect 88284 10782 88286 10834
rect 88338 10782 88452 10834
rect 88284 10780 88452 10782
rect 88284 10770 88340 10780
rect 87948 7422 87950 7474
rect 88002 7422 88004 7474
rect 87948 7364 88004 7422
rect 87948 7298 88004 7308
rect 88060 8316 88228 8372
rect 88508 10276 88564 10286
rect 88060 7140 88116 8316
rect 87836 6626 87892 6636
rect 87948 7084 88116 7140
rect 88284 8258 88340 8270
rect 88284 8206 88286 8258
rect 88338 8206 88340 8258
rect 87724 6580 87780 6590
rect 87724 4564 87780 6524
rect 87836 5908 87892 5918
rect 87836 5814 87892 5852
rect 87836 4564 87892 4574
rect 87724 4562 87892 4564
rect 87724 4510 87838 4562
rect 87890 4510 87892 4562
rect 87724 4508 87892 4510
rect 87836 4498 87892 4508
rect 87500 4286 87502 4338
rect 87554 4286 87556 4338
rect 87500 4274 87556 4286
rect 86044 3502 86046 3554
rect 86098 3502 86100 3554
rect 86044 3490 86100 3502
rect 87164 4116 87220 4126
rect 85596 3390 85598 3442
rect 85650 3390 85652 3442
rect 85596 3378 85652 3390
rect 85932 3444 85988 3454
rect 85932 980 85988 3388
rect 87052 3444 87108 3454
rect 87052 3330 87108 3388
rect 87052 3278 87054 3330
rect 87106 3278 87108 3330
rect 87052 3266 87108 3278
rect 85820 924 85988 980
rect 85820 800 85876 924
rect 87164 800 87220 4060
rect 87948 2660 88004 7084
rect 88172 6804 88228 6814
rect 88060 6468 88116 6478
rect 88060 6130 88116 6412
rect 88060 6078 88062 6130
rect 88114 6078 88116 6130
rect 88060 6066 88116 6078
rect 88172 6018 88228 6748
rect 88172 5966 88174 6018
rect 88226 5966 88228 6018
rect 88172 5954 88228 5966
rect 88284 5796 88340 8206
rect 88396 8148 88452 8158
rect 88396 8054 88452 8092
rect 88508 5908 88564 10220
rect 88620 8260 88676 14588
rect 88844 14530 88900 15484
rect 88844 14478 88846 14530
rect 88898 14478 88900 14530
rect 88844 14466 88900 14478
rect 88844 14308 88900 14318
rect 88844 13634 88900 14252
rect 88844 13582 88846 13634
rect 88898 13582 88900 13634
rect 88844 13570 88900 13582
rect 88956 13188 89012 16158
rect 89068 14754 89124 16716
rect 89068 14702 89070 14754
rect 89122 14702 89124 14754
rect 89068 14690 89124 14702
rect 88844 13132 89012 13188
rect 89068 13746 89124 13758
rect 89068 13694 89070 13746
rect 89122 13694 89124 13746
rect 88732 12964 88788 12974
rect 88732 12870 88788 12908
rect 88844 12740 88900 13132
rect 88956 12964 89012 12974
rect 88956 12870 89012 12908
rect 88844 12684 89012 12740
rect 88844 11172 88900 11182
rect 88732 10612 88788 10622
rect 88732 10518 88788 10556
rect 88732 9604 88788 9614
rect 88732 9154 88788 9548
rect 88732 9102 88734 9154
rect 88786 9102 88788 9154
rect 88732 9090 88788 9102
rect 88620 8194 88676 8204
rect 88844 8258 88900 11116
rect 88956 9714 89012 12684
rect 89068 11506 89124 13694
rect 89180 13522 89236 29372
rect 89516 25282 89572 25294
rect 89516 25230 89518 25282
rect 89570 25230 89572 25282
rect 89516 22260 89572 25230
rect 89516 22194 89572 22204
rect 89628 21028 89684 30380
rect 90300 25620 90356 55412
rect 93212 55412 93492 55468
rect 92988 55298 93044 55310
rect 92988 55246 92990 55298
rect 93042 55246 93044 55298
rect 92540 55188 92596 55198
rect 92540 55094 92596 55132
rect 92988 55188 93044 55246
rect 92988 55122 93044 55132
rect 93212 55186 93268 55412
rect 93212 55134 93214 55186
rect 93266 55134 93268 55186
rect 93212 55122 93268 55134
rect 94556 55076 94612 55086
rect 89852 25618 90356 25620
rect 89852 25566 90302 25618
rect 90354 25566 90356 25618
rect 89852 25564 90356 25566
rect 89740 25508 89796 25518
rect 89740 25414 89796 25452
rect 89852 25394 89908 25564
rect 90300 25554 90356 25564
rect 91084 30324 91140 30334
rect 89852 25342 89854 25394
rect 89906 25342 89908 25394
rect 89852 25330 89908 25342
rect 89740 23154 89796 23166
rect 89740 23102 89742 23154
rect 89794 23102 89796 23154
rect 89740 21588 89796 23102
rect 90300 23156 90356 23166
rect 90300 23154 90692 23156
rect 90300 23102 90302 23154
rect 90354 23102 90692 23154
rect 90300 23100 90692 23102
rect 90300 23090 90356 23100
rect 90524 22708 90580 22718
rect 90524 22370 90580 22652
rect 90636 22484 90692 23100
rect 90748 22484 90804 22494
rect 90636 22482 90804 22484
rect 90636 22430 90750 22482
rect 90802 22430 90804 22482
rect 90636 22428 90804 22430
rect 90748 22418 90804 22428
rect 90524 22318 90526 22370
rect 90578 22318 90580 22370
rect 90524 22306 90580 22318
rect 90300 22260 90356 22270
rect 90300 22166 90356 22204
rect 90972 22260 91028 22270
rect 90972 22166 91028 22204
rect 91084 21812 91140 30268
rect 92316 24612 92372 24622
rect 92092 23380 92148 23390
rect 92148 23324 92260 23380
rect 92092 23314 92148 23324
rect 91756 22708 91812 22718
rect 91644 22652 91756 22708
rect 91196 22484 91252 22494
rect 91196 22370 91252 22428
rect 91196 22318 91198 22370
rect 91250 22318 91252 22370
rect 91196 22306 91252 22318
rect 91644 22260 91700 22652
rect 91756 22642 91812 22652
rect 91980 22484 92036 22494
rect 91980 22390 92036 22428
rect 91644 22204 91812 22260
rect 90972 21756 91140 21812
rect 90524 21588 90580 21598
rect 89740 21522 89796 21532
rect 90300 21532 90524 21588
rect 89628 20972 89908 21028
rect 89628 18340 89684 18350
rect 89628 17780 89684 18284
rect 89628 17686 89684 17724
rect 89292 17442 89348 17454
rect 89292 17390 89294 17442
rect 89346 17390 89348 17442
rect 89292 17332 89348 17390
rect 89292 17266 89348 17276
rect 89628 17108 89684 17118
rect 89404 17106 89684 17108
rect 89404 17054 89630 17106
rect 89682 17054 89684 17106
rect 89404 17052 89684 17054
rect 89292 16996 89348 17006
rect 89292 16882 89348 16940
rect 89292 16830 89294 16882
rect 89346 16830 89348 16882
rect 89292 16818 89348 16830
rect 89292 15428 89348 15438
rect 89292 15204 89348 15372
rect 89404 15426 89460 17052
rect 89628 17042 89684 17052
rect 89740 16884 89796 16894
rect 89740 16790 89796 16828
rect 89404 15374 89406 15426
rect 89458 15374 89460 15426
rect 89404 15362 89460 15374
rect 89292 15138 89348 15148
rect 89180 13470 89182 13522
rect 89234 13470 89236 13522
rect 89180 13458 89236 13470
rect 89852 13860 89908 20972
rect 90300 20018 90356 21532
rect 90524 21494 90580 21532
rect 90300 19966 90302 20018
rect 90354 19966 90356 20018
rect 90300 19954 90356 19966
rect 90860 20018 90916 20030
rect 90860 19966 90862 20018
rect 90914 19966 90916 20018
rect 90860 19346 90916 19966
rect 90860 19294 90862 19346
rect 90914 19294 90916 19346
rect 90860 19282 90916 19294
rect 90636 19234 90692 19246
rect 90636 19182 90638 19234
rect 90690 19182 90692 19234
rect 90300 18452 90356 18462
rect 90300 18358 90356 18396
rect 90636 17892 90692 19182
rect 90636 17826 90692 17836
rect 90748 17780 90804 17790
rect 90076 17442 90132 17454
rect 90076 17390 90078 17442
rect 90130 17390 90132 17442
rect 89964 16882 90020 16894
rect 89964 16830 89966 16882
rect 90018 16830 90020 16882
rect 89964 16212 90020 16830
rect 89964 16146 90020 16156
rect 90076 15148 90132 17390
rect 90748 17108 90804 17724
rect 90860 17442 90916 17454
rect 90860 17390 90862 17442
rect 90914 17390 90916 17442
rect 90860 17332 90916 17390
rect 90860 17266 90916 17276
rect 90860 17108 90916 17118
rect 90748 17106 90916 17108
rect 90748 17054 90862 17106
rect 90914 17054 90916 17106
rect 90748 17052 90916 17054
rect 90860 17042 90916 17052
rect 90412 16770 90468 16782
rect 90412 16718 90414 16770
rect 90466 16718 90468 16770
rect 90412 16100 90468 16718
rect 90748 16212 90804 16222
rect 90748 16118 90804 16156
rect 90636 16100 90692 16110
rect 90412 16044 90636 16100
rect 90636 16006 90692 16044
rect 90860 15874 90916 15886
rect 90860 15822 90862 15874
rect 90914 15822 90916 15874
rect 90748 15428 90804 15438
rect 89404 13412 89460 13422
rect 89292 12740 89348 12750
rect 89292 12646 89348 12684
rect 89404 12290 89460 13356
rect 89404 12238 89406 12290
rect 89458 12238 89460 12290
rect 89404 12226 89460 12238
rect 89516 12852 89572 12862
rect 89068 11454 89070 11506
rect 89122 11454 89124 11506
rect 89068 11442 89124 11454
rect 89180 12178 89236 12190
rect 89180 12126 89182 12178
rect 89234 12126 89236 12178
rect 89180 12068 89236 12126
rect 89180 11394 89236 12012
rect 89180 11342 89182 11394
rect 89234 11342 89236 11394
rect 89180 10612 89236 11342
rect 89404 12068 89460 12078
rect 89404 11508 89460 12012
rect 89404 11282 89460 11452
rect 89404 11230 89406 11282
rect 89458 11230 89460 11282
rect 89404 11218 89460 11230
rect 89516 10948 89572 12796
rect 89628 12740 89684 12750
rect 89628 11732 89684 12684
rect 89628 11666 89684 11676
rect 89740 12740 89796 12750
rect 89852 12740 89908 13804
rect 89740 12738 89908 12740
rect 89740 12686 89742 12738
rect 89794 12686 89908 12738
rect 89740 12684 89908 12686
rect 89964 15092 90132 15148
rect 90188 15204 90244 15214
rect 89628 10948 89684 10958
rect 89516 10892 89628 10948
rect 89628 10882 89684 10892
rect 89180 10546 89236 10556
rect 89516 10610 89572 10622
rect 89516 10558 89518 10610
rect 89570 10558 89572 10610
rect 88956 9662 88958 9714
rect 89010 9662 89012 9714
rect 88956 9650 89012 9662
rect 89068 9716 89124 9726
rect 88844 8206 88846 8258
rect 88898 8206 88900 8258
rect 88844 8194 88900 8206
rect 88956 8260 89012 8270
rect 89068 8260 89124 9660
rect 88956 8258 89124 8260
rect 88956 8206 88958 8258
rect 89010 8206 89124 8258
rect 88956 8204 89124 8206
rect 89180 9492 89236 9502
rect 88956 8194 89012 8204
rect 89180 8146 89236 9436
rect 89292 8708 89348 8718
rect 89292 8258 89348 8652
rect 89292 8206 89294 8258
rect 89346 8206 89348 8258
rect 89292 8194 89348 8206
rect 89180 8094 89182 8146
rect 89234 8094 89236 8146
rect 89180 8082 89236 8094
rect 88620 8034 88676 8046
rect 88620 7982 88622 8034
rect 88674 7982 88676 8034
rect 88620 7588 88676 7982
rect 88732 7588 88788 7598
rect 88620 7586 88788 7588
rect 88620 7534 88734 7586
rect 88786 7534 88788 7586
rect 88620 7532 88788 7534
rect 88732 7522 88788 7532
rect 89516 7364 89572 10558
rect 89516 7298 89572 7308
rect 89628 10052 89684 10062
rect 89628 9826 89684 9996
rect 89628 9774 89630 9826
rect 89682 9774 89684 9826
rect 89628 7140 89684 9774
rect 89180 7084 89684 7140
rect 89068 6468 89124 6478
rect 89068 6374 89124 6412
rect 88956 6356 89012 6366
rect 88956 6244 89012 6300
rect 88956 6188 89124 6244
rect 88508 5852 88676 5908
rect 88284 5730 88340 5740
rect 87948 2594 88004 2604
rect 88508 5684 88564 5694
rect 88508 800 88564 5628
rect 88620 5124 88676 5852
rect 88620 5058 88676 5068
rect 89068 5906 89124 6188
rect 89068 5854 89070 5906
rect 89122 5854 89124 5906
rect 89068 2996 89124 5854
rect 89068 2930 89124 2940
rect 89180 1652 89236 7084
rect 89404 6802 89460 6814
rect 89404 6750 89406 6802
rect 89458 6750 89460 6802
rect 89292 6244 89348 6254
rect 89292 3442 89348 6188
rect 89404 5572 89460 6750
rect 89516 6692 89572 6702
rect 89572 6636 89684 6692
rect 89516 6626 89572 6636
rect 89404 5506 89460 5516
rect 89516 5236 89572 5246
rect 89628 5236 89684 6636
rect 89740 5794 89796 12684
rect 89852 11394 89908 11406
rect 89852 11342 89854 11394
rect 89906 11342 89908 11394
rect 89852 9492 89908 11342
rect 89852 9426 89908 9436
rect 89964 8260 90020 15092
rect 90188 14980 90244 15148
rect 90188 14924 90692 14980
rect 90076 14530 90132 14542
rect 90076 14478 90078 14530
rect 90130 14478 90132 14530
rect 90076 13188 90132 14478
rect 90524 13636 90580 13646
rect 90524 13542 90580 13580
rect 90076 13122 90132 13132
rect 90076 12964 90132 12974
rect 90076 12850 90132 12908
rect 90524 12964 90580 12974
rect 90524 12870 90580 12908
rect 90076 12798 90078 12850
rect 90130 12798 90132 12850
rect 90076 12786 90132 12798
rect 90524 12738 90580 12750
rect 90524 12686 90526 12738
rect 90578 12686 90580 12738
rect 90300 12404 90356 12414
rect 90300 12310 90356 12348
rect 90412 12290 90468 12302
rect 90412 12238 90414 12290
rect 90466 12238 90468 12290
rect 90076 11732 90132 11742
rect 90076 10610 90132 11676
rect 90412 11620 90468 12238
rect 90300 11564 90468 11620
rect 90076 10558 90078 10610
rect 90130 10558 90132 10610
rect 90076 10546 90132 10558
rect 90188 11172 90244 11182
rect 90300 11172 90356 11564
rect 90188 11170 90356 11172
rect 90188 11118 90190 11170
rect 90242 11118 90356 11170
rect 90188 11116 90356 11118
rect 90188 10500 90244 11116
rect 90244 10444 90356 10500
rect 90188 10434 90244 10444
rect 90300 9716 90356 10444
rect 90412 9716 90468 9726
rect 90300 9714 90468 9716
rect 90300 9662 90414 9714
rect 90466 9662 90468 9714
rect 90300 9660 90468 9662
rect 90412 9650 90468 9660
rect 90524 8484 90580 12686
rect 90636 12178 90692 14924
rect 90748 14532 90804 15372
rect 90860 15204 90916 15822
rect 90860 15138 90916 15148
rect 90748 14476 90916 14532
rect 90748 14306 90804 14318
rect 90748 14254 90750 14306
rect 90802 14254 90804 14306
rect 90748 14196 90804 14254
rect 90748 14130 90804 14140
rect 90748 13748 90804 13758
rect 90860 13748 90916 14476
rect 90748 13746 90916 13748
rect 90748 13694 90750 13746
rect 90802 13694 90916 13746
rect 90748 13692 90916 13694
rect 90748 13682 90804 13692
rect 90860 13524 90916 13534
rect 90636 12126 90638 12178
rect 90690 12126 90692 12178
rect 90636 12114 90692 12126
rect 90748 13468 90860 13524
rect 90636 11172 90692 11182
rect 90636 11078 90692 11116
rect 90412 8428 90580 8484
rect 90636 9156 90692 9166
rect 89964 8258 90132 8260
rect 89964 8206 89966 8258
rect 90018 8206 90132 8258
rect 89964 8204 90132 8206
rect 89964 8194 90020 8204
rect 89852 7924 89908 7934
rect 89852 5906 89908 7868
rect 90076 7588 90132 8204
rect 90188 8036 90244 8046
rect 90188 7942 90244 7980
rect 90076 7522 90132 7532
rect 89852 5854 89854 5906
rect 89906 5854 89908 5906
rect 89852 5842 89908 5854
rect 89964 7476 90020 7486
rect 89740 5742 89742 5794
rect 89794 5742 89796 5794
rect 89740 5730 89796 5742
rect 89516 5234 89628 5236
rect 89516 5182 89518 5234
rect 89570 5182 89628 5234
rect 89516 5180 89628 5182
rect 89516 5170 89572 5180
rect 89628 5142 89684 5180
rect 89964 5234 90020 7420
rect 89964 5182 89966 5234
rect 90018 5182 90020 5234
rect 89964 5170 90020 5182
rect 89964 4452 90020 4462
rect 89964 4358 90020 4396
rect 89628 4228 89684 4238
rect 89628 3554 89684 4172
rect 89628 3502 89630 3554
rect 89682 3502 89684 3554
rect 89628 3490 89684 3502
rect 90188 3666 90244 3678
rect 90188 3614 90190 3666
rect 90242 3614 90244 3666
rect 89292 3390 89294 3442
rect 89346 3390 89348 3442
rect 89292 3378 89348 3390
rect 90188 3388 90244 3614
rect 89180 1586 89236 1596
rect 89852 3332 90244 3388
rect 90412 3388 90468 8428
rect 90524 8260 90580 8270
rect 90524 7028 90580 8204
rect 90636 8148 90692 9100
rect 90748 8708 90804 13468
rect 90860 13458 90916 13468
rect 90860 12852 90916 12862
rect 90860 11732 90916 12796
rect 90972 12402 91028 21756
rect 91084 21586 91140 21598
rect 91084 21534 91086 21586
rect 91138 21534 91140 21586
rect 91084 21476 91140 21534
rect 91196 21476 91252 21486
rect 91084 21420 91196 21476
rect 91196 21410 91252 21420
rect 91084 21140 91140 21150
rect 91084 20804 91140 21084
rect 91308 20916 91364 20926
rect 91308 20822 91364 20860
rect 91756 20804 91812 22204
rect 91868 22146 91924 22158
rect 91868 22094 91870 22146
rect 91922 22094 91924 22146
rect 91868 21700 91924 22094
rect 92092 22146 92148 22158
rect 92092 22094 92094 22146
rect 92146 22094 92148 22146
rect 92092 22036 92148 22094
rect 92092 21970 92148 21980
rect 91868 21634 91924 21644
rect 91980 21476 92036 21486
rect 91980 20914 92036 21420
rect 91980 20862 91982 20914
rect 92034 20862 92036 20914
rect 91980 20850 92036 20862
rect 91868 20804 91924 20814
rect 91084 20748 91252 20804
rect 91756 20802 91924 20804
rect 91756 20750 91870 20802
rect 91922 20750 91924 20802
rect 91756 20748 91924 20750
rect 91084 19796 91140 19806
rect 91084 19124 91140 19740
rect 91084 19030 91140 19068
rect 91196 18900 91252 20748
rect 91868 20738 91924 20748
rect 92092 20804 92148 20842
rect 92092 20738 92148 20748
rect 91868 20244 91924 20254
rect 91756 19908 91812 19918
rect 91308 19124 91364 19134
rect 91308 19122 91700 19124
rect 91308 19070 91310 19122
rect 91362 19070 91700 19122
rect 91308 19068 91700 19070
rect 91308 19058 91364 19068
rect 91532 18900 91588 18910
rect 91196 18844 91364 18900
rect 91084 18450 91140 18462
rect 91084 18398 91086 18450
rect 91138 18398 91140 18450
rect 91084 17444 91140 18398
rect 91196 17444 91252 17454
rect 91084 17388 91196 17444
rect 91196 17350 91252 17388
rect 91084 16884 91140 16894
rect 91140 16828 91252 16884
rect 91084 16818 91140 16828
rect 91084 16436 91140 16446
rect 91084 15986 91140 16380
rect 91084 15934 91086 15986
rect 91138 15934 91140 15986
rect 91084 15922 91140 15934
rect 91196 14644 91252 16828
rect 91196 14578 91252 14588
rect 91196 14420 91252 14430
rect 91084 14306 91140 14318
rect 91084 14254 91086 14306
rect 91138 14254 91140 14306
rect 91084 13412 91140 14254
rect 91196 13524 91252 14364
rect 91196 13458 91252 13468
rect 91084 13346 91140 13356
rect 91308 13300 91364 18844
rect 91532 18674 91588 18844
rect 91532 18622 91534 18674
rect 91586 18622 91588 18674
rect 91532 18610 91588 18622
rect 91644 18674 91700 19068
rect 91644 18622 91646 18674
rect 91698 18622 91700 18674
rect 91644 18610 91700 18622
rect 91756 19012 91812 19852
rect 91756 18674 91812 18956
rect 91756 18622 91758 18674
rect 91810 18622 91812 18674
rect 91756 18610 91812 18622
rect 91644 16772 91700 16782
rect 91196 13244 91364 13300
rect 91420 16770 91700 16772
rect 91420 16718 91646 16770
rect 91698 16718 91700 16770
rect 91420 16716 91700 16718
rect 91084 12852 91140 12862
rect 91196 12852 91252 13244
rect 91084 12850 91252 12852
rect 91084 12798 91086 12850
rect 91138 12798 91252 12850
rect 91084 12796 91252 12798
rect 91308 12964 91364 12974
rect 91084 12786 91140 12796
rect 90972 12350 90974 12402
rect 91026 12350 91028 12402
rect 90972 12338 91028 12350
rect 91308 12178 91364 12908
rect 91308 12126 91310 12178
rect 91362 12126 91364 12178
rect 91308 12114 91364 12126
rect 90860 11666 90916 11676
rect 90972 11282 91028 11294
rect 90972 11230 90974 11282
rect 91026 11230 91028 11282
rect 90860 11170 90916 11182
rect 90860 11118 90862 11170
rect 90914 11118 90916 11170
rect 90860 9828 90916 11118
rect 90972 10948 91028 11230
rect 90972 10882 91028 10892
rect 91308 10722 91364 10734
rect 91308 10670 91310 10722
rect 91362 10670 91364 10722
rect 91308 10500 91364 10670
rect 91308 10434 91364 10444
rect 91196 9828 91252 9838
rect 91420 9828 91476 16716
rect 91644 16706 91700 16716
rect 91532 15204 91588 15242
rect 91868 15148 91924 20188
rect 91980 19124 92036 19134
rect 91980 19010 92036 19068
rect 91980 18958 91982 19010
rect 92034 18958 92036 19010
rect 91980 17892 92036 18958
rect 92204 18676 92260 23324
rect 92316 21924 92372 24556
rect 92652 23716 92708 23726
rect 92652 23622 92708 23660
rect 93212 23714 93268 23726
rect 93212 23662 93214 23714
rect 93266 23662 93268 23714
rect 92876 23154 92932 23166
rect 92876 23102 92878 23154
rect 92930 23102 92932 23154
rect 92652 23042 92708 23054
rect 92652 22990 92654 23042
rect 92706 22990 92708 23042
rect 92316 21858 92372 21868
rect 92540 22370 92596 22382
rect 92540 22318 92542 22370
rect 92594 22318 92596 22370
rect 92540 21476 92596 22318
rect 92540 21410 92596 21420
rect 92652 22036 92708 22990
rect 92876 22708 92932 23102
rect 93100 23044 93156 23054
rect 93100 22950 93156 22988
rect 92876 22642 92932 22652
rect 92988 22596 93044 22606
rect 93044 22540 93156 22596
rect 92988 22530 93044 22540
rect 92988 22148 93044 22158
rect 92428 21028 92484 21038
rect 92484 20972 92596 21028
rect 92428 20962 92484 20972
rect 92428 20804 92484 20814
rect 92428 20710 92484 20748
rect 92540 20468 92596 20972
rect 92540 20402 92596 20412
rect 92428 19012 92484 19022
rect 92428 18918 92484 18956
rect 92540 18900 92596 18910
rect 92204 18620 92372 18676
rect 92204 18450 92260 18462
rect 92204 18398 92206 18450
rect 92258 18398 92260 18450
rect 92204 18340 92260 18398
rect 92204 18274 92260 18284
rect 91980 17826 92036 17836
rect 92316 17780 92372 18620
rect 92540 18450 92596 18844
rect 92540 18398 92542 18450
rect 92594 18398 92596 18450
rect 92540 18340 92596 18398
rect 92540 18274 92596 18284
rect 92092 17724 92372 17780
rect 91980 16996 92036 17006
rect 91980 16436 92036 16940
rect 91980 16210 92036 16380
rect 91980 16158 91982 16210
rect 92034 16158 92036 16210
rect 91980 16146 92036 16158
rect 92092 16212 92148 17724
rect 92204 17556 92260 17566
rect 92260 17500 92372 17556
rect 92204 17462 92260 17500
rect 92316 17108 92372 17500
rect 92540 17108 92596 17118
rect 92316 17106 92596 17108
rect 92316 17054 92318 17106
rect 92370 17054 92542 17106
rect 92594 17054 92596 17106
rect 92316 17052 92596 17054
rect 92316 17042 92372 17052
rect 92540 17042 92596 17052
rect 91532 15138 91588 15148
rect 91644 15092 91924 15148
rect 92092 15538 92148 16156
rect 92092 15486 92094 15538
rect 92146 15486 92148 15538
rect 91532 14644 91588 14654
rect 91532 12740 91588 14588
rect 91532 12674 91588 12684
rect 91532 12180 91588 12190
rect 91644 12180 91700 15092
rect 92092 14642 92148 15486
rect 92428 15874 92484 15886
rect 92428 15822 92430 15874
rect 92482 15822 92484 15874
rect 92428 15148 92484 15822
rect 92652 15148 92708 21980
rect 92876 22146 93044 22148
rect 92876 22094 92990 22146
rect 93042 22094 93044 22146
rect 92876 22092 93044 22094
rect 92764 21700 92820 21710
rect 92764 20578 92820 21644
rect 92876 21140 92932 22092
rect 92988 22082 93044 22092
rect 92876 21074 92932 21084
rect 92988 21028 93044 21038
rect 92876 20804 92932 20814
rect 92876 20710 92932 20748
rect 92764 20526 92766 20578
rect 92818 20526 92820 20578
rect 92764 20514 92820 20526
rect 92988 20578 93044 20972
rect 92988 20526 92990 20578
rect 93042 20526 93044 20578
rect 92876 20468 92932 20478
rect 92764 17442 92820 17454
rect 92764 17390 92766 17442
rect 92818 17390 92820 17442
rect 92764 16884 92820 17390
rect 92764 16818 92820 16828
rect 92876 16210 92932 20412
rect 92988 20244 93044 20526
rect 92988 20178 93044 20188
rect 93100 18676 93156 22540
rect 93212 21588 93268 23662
rect 93324 23716 93380 23726
rect 93324 23268 93380 23660
rect 93324 23174 93380 23212
rect 93548 23156 93604 23166
rect 93548 23154 93940 23156
rect 93548 23102 93550 23154
rect 93602 23102 93940 23154
rect 93548 23100 93940 23102
rect 93548 23090 93604 23100
rect 93884 21810 93940 23100
rect 93884 21758 93886 21810
rect 93938 21758 93940 21810
rect 93884 21746 93940 21758
rect 93772 21700 93828 21710
rect 93772 21606 93828 21644
rect 93212 21364 93268 21532
rect 93996 21586 94052 21598
rect 93996 21534 93998 21586
rect 94050 21534 94052 21586
rect 93436 21474 93492 21486
rect 93436 21422 93438 21474
rect 93490 21422 93492 21474
rect 93212 21308 93380 21364
rect 93324 20580 93380 21308
rect 93436 21028 93492 21422
rect 93436 20962 93492 20972
rect 93548 21476 93604 21486
rect 93436 20804 93492 20814
rect 93548 20804 93604 21420
rect 93996 21140 94052 21534
rect 94444 21586 94500 21598
rect 94444 21534 94446 21586
rect 94498 21534 94500 21586
rect 94444 21476 94500 21534
rect 94444 21410 94500 21420
rect 93996 21074 94052 21084
rect 93436 20802 93604 20804
rect 93436 20750 93438 20802
rect 93490 20750 93604 20802
rect 93436 20748 93604 20750
rect 93436 20738 93492 20748
rect 93324 20514 93380 20524
rect 93772 20580 93828 20590
rect 93660 20244 93716 20254
rect 93772 20244 93828 20524
rect 93660 20242 93828 20244
rect 93660 20190 93662 20242
rect 93714 20190 93828 20242
rect 93660 20188 93828 20190
rect 93660 20178 93716 20188
rect 93212 19908 93268 19918
rect 93212 19814 93268 19852
rect 94332 19458 94388 19470
rect 94332 19406 94334 19458
rect 94386 19406 94388 19458
rect 94332 19348 94388 19406
rect 94220 19346 94388 19348
rect 94220 19294 94334 19346
rect 94386 19294 94388 19346
rect 94220 19292 94388 19294
rect 93548 19010 93604 19022
rect 93548 18958 93550 19010
rect 93602 18958 93604 19010
rect 93100 18620 93268 18676
rect 93100 18450 93156 18462
rect 93100 18398 93102 18450
rect 93154 18398 93156 18450
rect 92988 17556 93044 17566
rect 93100 17556 93156 18398
rect 93044 17500 93156 17556
rect 93212 17778 93268 18620
rect 93548 18564 93604 18958
rect 93548 18470 93604 18508
rect 94220 18004 94276 19292
rect 94332 19282 94388 19292
rect 94444 18340 94500 18350
rect 94444 18246 94500 18284
rect 93212 17726 93214 17778
rect 93266 17726 93268 17778
rect 92988 17490 93044 17500
rect 92988 16996 93044 17006
rect 93044 16940 93156 16996
rect 92988 16930 93044 16940
rect 93100 16882 93156 16940
rect 93100 16830 93102 16882
rect 93154 16830 93156 16882
rect 93100 16818 93156 16830
rect 92876 16158 92878 16210
rect 92930 16158 92932 16210
rect 92876 16100 92932 16158
rect 92876 16034 92932 16044
rect 92092 14590 92094 14642
rect 92146 14590 92148 14642
rect 92092 14578 92148 14590
rect 92316 15092 92484 15148
rect 92540 15092 92708 15148
rect 92316 14756 92372 15092
rect 91756 14196 91812 14206
rect 91812 14140 91924 14196
rect 91756 14130 91812 14140
rect 91756 13188 91812 13198
rect 91756 12964 91812 13132
rect 91868 12964 91924 14140
rect 92316 13300 92372 14700
rect 92428 14306 92484 14318
rect 92428 14254 92430 14306
rect 92482 14254 92484 14306
rect 92428 14084 92484 14254
rect 92428 14018 92484 14028
rect 92316 13244 92484 13300
rect 91980 13188 92036 13198
rect 92036 13132 92372 13188
rect 91980 13122 92036 13132
rect 92316 13074 92372 13132
rect 92316 13022 92318 13074
rect 92370 13022 92372 13074
rect 92316 13010 92372 13022
rect 91868 12908 92148 12964
rect 91756 12898 91812 12908
rect 91980 12740 92036 12750
rect 91532 12178 91700 12180
rect 91532 12126 91534 12178
rect 91586 12126 91700 12178
rect 91532 12124 91700 12126
rect 91756 12738 92036 12740
rect 91756 12686 91982 12738
rect 92034 12686 92036 12738
rect 91756 12684 92036 12686
rect 91532 12114 91588 12124
rect 91644 11172 91700 11182
rect 90860 9772 91140 9828
rect 90860 9492 90916 9502
rect 90860 8930 90916 9436
rect 90860 8878 90862 8930
rect 90914 8878 90916 8930
rect 90860 8866 90916 8878
rect 90748 8652 91028 8708
rect 90748 8484 90804 8494
rect 90748 8370 90804 8428
rect 90748 8318 90750 8370
rect 90802 8318 90804 8370
rect 90748 8306 90804 8318
rect 90972 8370 91028 8652
rect 90972 8318 90974 8370
rect 91026 8318 91028 8370
rect 90972 8306 91028 8318
rect 90636 8092 90804 8148
rect 90524 6962 90580 6972
rect 90636 6578 90692 6590
rect 90636 6526 90638 6578
rect 90690 6526 90692 6578
rect 90524 6244 90580 6254
rect 90524 5906 90580 6188
rect 90524 5854 90526 5906
rect 90578 5854 90580 5906
rect 90524 5842 90580 5854
rect 90636 4562 90692 6526
rect 90636 4510 90638 4562
rect 90690 4510 90692 4562
rect 90636 4498 90692 4510
rect 90412 3332 90580 3388
rect 89852 800 89908 3332
rect 90524 2324 90580 3332
rect 90748 2996 90804 8092
rect 90860 7364 90916 7374
rect 90860 7270 90916 7308
rect 90860 6468 90916 6478
rect 90860 5010 90916 6412
rect 90860 4958 90862 5010
rect 90914 4958 90916 5010
rect 90860 4946 90916 4958
rect 91084 3668 91140 9772
rect 91196 9826 91476 9828
rect 91196 9774 91198 9826
rect 91250 9774 91476 9826
rect 91196 9772 91476 9774
rect 91532 10836 91588 10846
rect 91196 9156 91252 9772
rect 91532 9716 91588 10780
rect 91196 9090 91252 9100
rect 91308 9660 91588 9716
rect 91196 8930 91252 8942
rect 91196 8878 91198 8930
rect 91250 8878 91252 8930
rect 91196 8820 91252 8878
rect 91196 8754 91252 8764
rect 91196 7362 91252 7374
rect 91196 7310 91198 7362
rect 91250 7310 91252 7362
rect 91196 6578 91252 7310
rect 91308 6690 91364 9660
rect 91532 9492 91588 9502
rect 91420 8372 91476 8382
rect 91420 8278 91476 8316
rect 91420 7476 91476 7486
rect 91532 7476 91588 9436
rect 91420 7474 91588 7476
rect 91420 7422 91422 7474
rect 91474 7422 91588 7474
rect 91420 7420 91588 7422
rect 91644 7474 91700 11116
rect 91644 7422 91646 7474
rect 91698 7422 91700 7474
rect 91420 7410 91476 7420
rect 91644 7410 91700 7422
rect 91756 7252 91812 12684
rect 91980 12674 92036 12684
rect 91868 12516 91924 12526
rect 91868 12066 91924 12460
rect 91868 12014 91870 12066
rect 91922 12014 91924 12066
rect 91868 12002 91924 12014
rect 91980 11508 92036 11518
rect 91980 11396 92036 11452
rect 91868 11394 92036 11396
rect 91868 11342 91982 11394
rect 92034 11342 92036 11394
rect 91868 11340 92036 11342
rect 91868 9826 91924 11340
rect 91980 11330 92036 11340
rect 92092 10948 92148 12908
rect 92428 12852 92484 13244
rect 92540 12962 92596 15092
rect 92876 15090 92932 15102
rect 92876 15038 92878 15090
rect 92930 15038 92932 15090
rect 92876 14530 92932 15038
rect 92876 14478 92878 14530
rect 92930 14478 92932 14530
rect 92876 14308 92932 14478
rect 92876 14242 92932 14252
rect 92988 15092 93044 15102
rect 92988 13972 93044 15036
rect 93100 14532 93156 14542
rect 93100 14438 93156 14476
rect 93100 13972 93156 13982
rect 92988 13970 93156 13972
rect 92988 13918 93102 13970
rect 93154 13918 93156 13970
rect 92988 13916 93156 13918
rect 93100 13906 93156 13916
rect 92652 13634 92708 13646
rect 92652 13582 92654 13634
rect 92706 13582 92708 13634
rect 92652 13522 92708 13582
rect 92652 13470 92654 13522
rect 92706 13470 92708 13522
rect 92652 13458 92708 13470
rect 93100 13636 93156 13646
rect 92540 12910 92542 12962
rect 92594 12910 92596 12962
rect 92540 12898 92596 12910
rect 92316 12796 92484 12852
rect 93100 12850 93156 13580
rect 93100 12798 93102 12850
rect 93154 12798 93156 12850
rect 91868 9774 91870 9826
rect 91922 9774 91924 9826
rect 91868 9762 91924 9774
rect 91980 10892 92148 10948
rect 92204 12740 92260 12750
rect 91980 8372 92036 10892
rect 92204 10836 92260 12684
rect 92316 11620 92372 12796
rect 92764 12740 92820 12750
rect 92316 11554 92372 11564
rect 92428 12738 92820 12740
rect 92428 12686 92766 12738
rect 92818 12686 92820 12738
rect 92428 12684 92820 12686
rect 92316 11396 92372 11406
rect 92428 11396 92484 12684
rect 92764 12674 92820 12684
rect 92876 12740 92932 12750
rect 92876 11732 92932 12684
rect 92988 12738 93044 12750
rect 92988 12686 92990 12738
rect 93042 12686 93044 12738
rect 92988 12516 93044 12686
rect 92988 12450 93044 12460
rect 92316 11394 92484 11396
rect 92316 11342 92318 11394
rect 92370 11342 92484 11394
rect 92316 11340 92484 11342
rect 92540 11676 92932 11732
rect 92988 11844 93044 11854
rect 92316 11330 92372 11340
rect 92540 11284 92596 11676
rect 92988 11620 93044 11788
rect 92652 11564 93044 11620
rect 92652 11394 92708 11564
rect 93100 11508 93156 12798
rect 92988 11452 93156 11508
rect 92988 11396 93044 11452
rect 92652 11342 92654 11394
rect 92706 11342 92708 11394
rect 92652 11330 92708 11342
rect 92876 11340 93044 11396
rect 92428 11228 92596 11284
rect 92428 11170 92484 11228
rect 92764 11172 92820 11182
rect 92428 11118 92430 11170
rect 92482 11118 92484 11170
rect 92428 11106 92484 11118
rect 92540 11170 92820 11172
rect 92540 11118 92766 11170
rect 92818 11118 92820 11170
rect 92540 11116 92820 11118
rect 92204 10770 92260 10780
rect 92092 10724 92148 10734
rect 92092 8820 92148 10668
rect 92204 10612 92260 10622
rect 92204 10518 92260 10556
rect 92428 10610 92484 10622
rect 92428 10558 92430 10610
rect 92482 10558 92484 10610
rect 92428 10052 92484 10558
rect 92204 9996 92484 10052
rect 92204 9826 92260 9996
rect 92204 9774 92206 9826
rect 92258 9774 92260 9826
rect 92204 9762 92260 9774
rect 92540 9826 92596 11116
rect 92764 11106 92820 11116
rect 92652 10724 92708 10734
rect 92652 10630 92708 10668
rect 92764 10612 92820 10622
rect 92876 10612 92932 11340
rect 93100 11284 93156 11294
rect 92988 11172 93044 11182
rect 92988 11078 93044 11116
rect 93100 10724 93156 11228
rect 92764 10610 92932 10612
rect 92764 10558 92766 10610
rect 92818 10558 92932 10610
rect 92764 10556 92932 10558
rect 92988 10668 93156 10724
rect 92540 9774 92542 9826
rect 92594 9774 92596 9826
rect 92540 9762 92596 9774
rect 92652 9828 92708 9838
rect 92652 9734 92708 9772
rect 92316 9602 92372 9614
rect 92316 9550 92318 9602
rect 92370 9550 92372 9602
rect 92316 9156 92372 9550
rect 92316 9090 92372 9100
rect 92652 9604 92708 9614
rect 92092 8754 92148 8764
rect 91980 8316 92372 8372
rect 91308 6638 91310 6690
rect 91362 6638 91364 6690
rect 91308 6626 91364 6638
rect 91644 7196 91812 7252
rect 91980 8146 92036 8158
rect 91980 8094 91982 8146
rect 92034 8094 92036 8146
rect 91196 6526 91198 6578
rect 91250 6526 91252 6578
rect 91196 4564 91252 6526
rect 91196 4498 91252 4508
rect 91084 3602 91140 3612
rect 91196 4004 91252 4014
rect 90860 2996 90916 3006
rect 90748 2940 90860 2996
rect 90860 2930 90916 2940
rect 90524 2258 90580 2268
rect 91196 800 91252 3948
rect 91644 868 91700 7196
rect 91980 6802 92036 8094
rect 92092 7588 92148 7598
rect 92092 7494 92148 7532
rect 91980 6750 91982 6802
rect 92034 6750 92036 6802
rect 91980 6738 92036 6750
rect 92204 7476 92260 7486
rect 92204 6804 92260 7420
rect 91868 6020 91924 6030
rect 91868 5684 91924 5964
rect 91868 5618 91924 5628
rect 91980 5236 92036 5246
rect 91980 5010 92036 5180
rect 91980 4958 91982 5010
rect 92034 4958 92036 5010
rect 91980 4946 92036 4958
rect 92092 5012 92148 5022
rect 92204 5012 92260 6748
rect 92092 5010 92260 5012
rect 92092 4958 92094 5010
rect 92146 4958 92260 5010
rect 92092 4956 92260 4958
rect 92316 5012 92372 8316
rect 92652 6020 92708 9548
rect 92764 8708 92820 10556
rect 92988 9716 93044 10668
rect 93100 10500 93156 10510
rect 93100 10406 93156 10444
rect 92988 9714 93156 9716
rect 92988 9662 92990 9714
rect 93042 9662 93156 9714
rect 92988 9660 93156 9662
rect 92988 9650 93044 9660
rect 92764 8642 92820 8652
rect 92876 9602 92932 9614
rect 92876 9550 92878 9602
rect 92930 9550 92932 9602
rect 92876 8820 92932 9550
rect 92876 8484 92932 8764
rect 92876 8418 92932 8428
rect 92988 8372 93044 8382
rect 92764 7586 92820 7598
rect 92764 7534 92766 7586
rect 92818 7534 92820 7586
rect 92764 6692 92820 7534
rect 92988 7362 93044 8316
rect 92988 7310 92990 7362
rect 93042 7310 93044 7362
rect 92988 7298 93044 7310
rect 93100 8036 93156 9660
rect 93100 6916 93156 7980
rect 93212 7924 93268 17726
rect 93996 17948 94276 18004
rect 93996 17780 94052 17948
rect 93996 17724 94108 17780
rect 94052 17668 94108 17724
rect 94052 17612 94276 17668
rect 93772 17556 93828 17566
rect 93660 17444 93716 17454
rect 93436 17442 93716 17444
rect 93436 17390 93662 17442
rect 93714 17390 93716 17442
rect 93436 17388 93716 17390
rect 93324 16100 93380 16110
rect 93324 15314 93380 16044
rect 93324 15262 93326 15314
rect 93378 15262 93380 15314
rect 93324 15250 93380 15262
rect 93436 15148 93492 17388
rect 93660 17378 93716 17388
rect 93660 17108 93716 17118
rect 93772 17108 93828 17500
rect 93884 17108 93940 17118
rect 93660 17106 93940 17108
rect 93660 17054 93662 17106
rect 93714 17054 93886 17106
rect 93938 17054 93940 17106
rect 93660 17052 93940 17054
rect 93660 17042 93716 17052
rect 93884 17042 93940 17052
rect 93996 16212 94052 16222
rect 93996 16118 94052 16156
rect 93548 16100 93604 16110
rect 93604 16044 93940 16100
rect 93548 16006 93604 16044
rect 93324 15092 93492 15148
rect 93324 9380 93380 15092
rect 93884 13970 93940 16044
rect 93996 15428 94052 15438
rect 93996 15204 94052 15372
rect 93996 15138 94052 15148
rect 93884 13918 93886 13970
rect 93938 13918 93940 13970
rect 93884 13906 93940 13918
rect 94108 15092 94164 15102
rect 93548 13860 93604 13870
rect 93548 13766 93604 13804
rect 93436 13522 93492 13534
rect 93436 13470 93438 13522
rect 93490 13470 93492 13522
rect 93436 9604 93492 13470
rect 93996 12964 94052 12974
rect 93996 12870 94052 12908
rect 93548 12740 93604 12750
rect 93996 12740 94052 12750
rect 93548 12738 93940 12740
rect 93548 12686 93550 12738
rect 93602 12686 93940 12738
rect 93548 12684 93940 12686
rect 93548 12674 93604 12684
rect 93548 11844 93604 11854
rect 93548 11618 93604 11788
rect 93548 11566 93550 11618
rect 93602 11566 93604 11618
rect 93548 11554 93604 11566
rect 93772 11844 93828 11854
rect 93660 11284 93716 11294
rect 93660 11190 93716 11228
rect 93548 11170 93604 11182
rect 93548 11118 93550 11170
rect 93602 11118 93604 11170
rect 93548 9828 93604 11118
rect 93660 10836 93716 10846
rect 93772 10836 93828 11788
rect 93660 10834 93828 10836
rect 93660 10782 93662 10834
rect 93714 10782 93828 10834
rect 93660 10780 93828 10782
rect 93660 10770 93716 10780
rect 93884 10276 93940 12684
rect 93996 12290 94052 12684
rect 93996 12238 93998 12290
rect 94050 12238 94052 12290
rect 93996 12226 94052 12238
rect 94108 11620 94164 15036
rect 94220 11732 94276 17612
rect 94332 17666 94388 17678
rect 94332 17614 94334 17666
rect 94386 17614 94388 17666
rect 94332 17444 94388 17614
rect 94332 17378 94388 17388
rect 94444 17220 94500 17230
rect 94444 16994 94500 17164
rect 94444 16942 94446 16994
rect 94498 16942 94500 16994
rect 94444 16930 94500 16942
rect 94556 16548 94612 55020
rect 96908 55076 96964 55086
rect 96908 54982 96964 55020
rect 97580 55076 97636 56030
rect 100828 55410 100884 56252
rect 101052 56242 101108 56252
rect 104636 56308 104692 59200
rect 104636 56242 104692 56252
rect 105868 56308 105924 56318
rect 105868 56214 105924 56252
rect 108444 56308 108500 59200
rect 112252 56644 112308 59200
rect 112252 56588 112420 56644
rect 111996 56476 112260 56486
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 111996 56410 112260 56420
rect 108444 56242 108500 56252
rect 109676 56308 109732 56318
rect 109676 56214 109732 56252
rect 101388 56194 101444 56206
rect 101388 56142 101390 56194
rect 101442 56142 101444 56194
rect 101388 55468 101444 56142
rect 110012 56196 110068 56206
rect 104860 56082 104916 56094
rect 104860 56030 104862 56082
rect 104914 56030 104916 56082
rect 104860 55468 104916 56030
rect 108668 56082 108724 56094
rect 108668 56030 108670 56082
rect 108722 56030 108724 56082
rect 108668 55468 108724 56030
rect 101388 55412 101892 55468
rect 100828 55358 100830 55410
rect 100882 55358 100884 55410
rect 100828 55346 100884 55358
rect 97580 55010 97636 55020
rect 96636 54124 96900 54134
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96636 54058 96900 54068
rect 96636 52556 96900 52566
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96636 52490 96900 52500
rect 96636 50988 96900 50998
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96636 50922 96900 50932
rect 96636 49420 96900 49430
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96636 49354 96900 49364
rect 96636 47852 96900 47862
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96636 47786 96900 47796
rect 96636 46284 96900 46294
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96636 46218 96900 46228
rect 96636 44716 96900 44726
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96636 44650 96900 44660
rect 96636 43148 96900 43158
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96636 43082 96900 43092
rect 96636 41580 96900 41590
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96636 41514 96900 41524
rect 96636 40012 96900 40022
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96636 39946 96900 39956
rect 96636 38444 96900 38454
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96636 38378 96900 38388
rect 96636 36876 96900 36886
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96636 36810 96900 36820
rect 96636 35308 96900 35318
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96636 35242 96900 35252
rect 96636 33740 96900 33750
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96636 33674 96900 33684
rect 96636 32172 96900 32182
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96636 32106 96900 32116
rect 96636 30604 96900 30614
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96636 30538 96900 30548
rect 96636 29036 96900 29046
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96636 28970 96900 28980
rect 96636 27468 96900 27478
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96636 27402 96900 27412
rect 96636 25900 96900 25910
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96636 25834 96900 25844
rect 101836 25620 101892 55412
rect 104636 55412 104916 55468
rect 108332 55412 108724 55468
rect 103964 55188 104020 55198
rect 104300 55188 104356 55198
rect 104020 55186 104356 55188
rect 104020 55134 104302 55186
rect 104354 55134 104356 55186
rect 104020 55132 104356 55134
rect 103964 55094 104020 55132
rect 104300 55122 104356 55132
rect 104636 55186 104692 55412
rect 104636 55134 104638 55186
rect 104690 55134 104692 55186
rect 104636 55122 104692 55134
rect 108332 55074 108388 55412
rect 108332 55022 108334 55074
rect 108386 55022 108388 55074
rect 107100 32788 107156 32798
rect 105756 27748 105812 27758
rect 105756 27188 105812 27692
rect 105532 27186 105812 27188
rect 105532 27134 105758 27186
rect 105810 27134 105812 27186
rect 105532 27132 105812 27134
rect 105532 26402 105588 27132
rect 105756 27122 105812 27132
rect 107100 26516 107156 32732
rect 108332 29428 108388 55022
rect 108332 29362 108388 29372
rect 105532 26350 105534 26402
rect 105586 26350 105588 26402
rect 105532 26338 105588 26350
rect 106540 26514 107156 26516
rect 106540 26462 107102 26514
rect 107154 26462 107156 26514
rect 106540 26460 107156 26462
rect 106540 26402 106596 26460
rect 107100 26450 107156 26460
rect 108668 28644 108724 28654
rect 106540 26350 106542 26402
rect 106594 26350 106596 26402
rect 106540 26338 106596 26350
rect 104972 26290 105028 26302
rect 104972 26238 104974 26290
rect 105026 26238 105028 26290
rect 104524 26180 104580 26190
rect 104524 26086 104580 26124
rect 104860 26178 104916 26190
rect 104860 26126 104862 26178
rect 104914 26126 104916 26178
rect 101388 25618 101892 25620
rect 101388 25566 101838 25618
rect 101890 25566 101892 25618
rect 101388 25564 101892 25566
rect 100492 25508 100548 25518
rect 100492 25414 100548 25452
rect 100940 25508 100996 25518
rect 100940 25414 100996 25452
rect 101388 25394 101444 25564
rect 101836 25554 101892 25564
rect 104076 25732 104132 25742
rect 101388 25342 101390 25394
rect 101442 25342 101444 25394
rect 101388 25330 101444 25342
rect 100828 25282 100884 25294
rect 100828 25230 100830 25282
rect 100882 25230 100884 25282
rect 96636 24332 96900 24342
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96636 24266 96900 24276
rect 97468 23268 97524 23278
rect 95340 23044 95396 23054
rect 95340 22370 95396 22988
rect 97132 22932 97188 22942
rect 96636 22764 96900 22774
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96636 22698 96900 22708
rect 95340 22318 95342 22370
rect 95394 22318 95396 22370
rect 95340 22306 95396 22318
rect 96124 22370 96180 22382
rect 96124 22318 96126 22370
rect 96178 22318 96180 22370
rect 96124 22148 96180 22318
rect 96460 22148 96516 22158
rect 96124 22146 96516 22148
rect 96124 22094 96462 22146
rect 96514 22094 96516 22146
rect 96124 22092 96516 22094
rect 95228 21924 95284 21934
rect 95004 21252 95060 21262
rect 94892 19906 94948 19918
rect 94892 19854 94894 19906
rect 94946 19854 94948 19906
rect 94892 19458 94948 19854
rect 94892 19406 94894 19458
rect 94946 19406 94948 19458
rect 94892 19394 94948 19406
rect 94780 19012 94836 19022
rect 94444 16492 94612 16548
rect 94668 19010 94836 19012
rect 94668 18958 94782 19010
rect 94834 18958 94836 19010
rect 94668 18956 94836 18958
rect 94668 18564 94724 18956
rect 94780 18946 94836 18956
rect 94332 16212 94388 16222
rect 94332 15538 94388 16156
rect 94332 15486 94334 15538
rect 94386 15486 94388 15538
rect 94332 15474 94388 15486
rect 94444 14754 94500 16492
rect 94444 14702 94446 14754
rect 94498 14702 94500 14754
rect 94444 14690 94500 14702
rect 94556 15874 94612 15886
rect 94556 15822 94558 15874
rect 94610 15822 94612 15874
rect 94556 13860 94612 15822
rect 94668 14308 94724 18508
rect 94780 18338 94836 18350
rect 94780 18286 94782 18338
rect 94834 18286 94836 18338
rect 94780 18228 94836 18286
rect 94780 18162 94836 18172
rect 94892 18340 94948 18350
rect 94892 17666 94948 18284
rect 94892 17614 94894 17666
rect 94946 17614 94948 17666
rect 94892 17602 94948 17614
rect 95004 17106 95060 21196
rect 95228 20130 95284 21868
rect 95788 20916 95844 20926
rect 95564 20802 95620 20814
rect 95564 20750 95566 20802
rect 95618 20750 95620 20802
rect 95564 20580 95620 20750
rect 95564 20514 95620 20524
rect 95788 20244 95844 20860
rect 96348 20802 96404 20814
rect 96348 20750 96350 20802
rect 96402 20750 96404 20802
rect 96348 20356 96404 20750
rect 96460 20580 96516 22092
rect 96636 21196 96900 21206
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96636 21130 96900 21140
rect 96460 20514 96516 20524
rect 96684 20916 96740 20926
rect 96348 20300 96628 20356
rect 95228 20078 95230 20130
rect 95282 20078 95284 20130
rect 95228 20020 95284 20078
rect 95228 19348 95284 19964
rect 95676 20188 95788 20244
rect 95676 19796 95732 20188
rect 95788 20178 95844 20188
rect 96572 20242 96628 20300
rect 96572 20190 96574 20242
rect 96626 20190 96628 20242
rect 96572 20178 96628 20190
rect 96124 20130 96180 20142
rect 96124 20078 96126 20130
rect 96178 20078 96180 20130
rect 95788 20020 95844 20030
rect 96124 20020 96180 20078
rect 96460 20020 96516 20030
rect 96684 20020 96740 20860
rect 95788 19926 95844 19964
rect 95900 20018 96740 20020
rect 95900 19966 96462 20018
rect 96514 19966 96740 20018
rect 95900 19964 96740 19966
rect 96796 20244 96852 20254
rect 96796 20130 96852 20188
rect 96796 20078 96798 20130
rect 96850 20078 96852 20130
rect 95676 19740 95844 19796
rect 95228 19254 95284 19292
rect 95788 19346 95844 19740
rect 95788 19294 95790 19346
rect 95842 19294 95844 19346
rect 95788 19282 95844 19294
rect 95788 18564 95844 18574
rect 95900 18564 95956 19964
rect 96460 19954 96516 19964
rect 96796 19796 96852 20078
rect 97020 20020 97076 20030
rect 97020 19926 97076 19964
rect 97132 19796 97188 22876
rect 97468 21700 97524 23212
rect 100828 22932 100884 25230
rect 100828 22866 100884 22876
rect 99820 22370 99876 22382
rect 99820 22318 99822 22370
rect 99874 22318 99876 22370
rect 97468 21606 97524 21644
rect 98028 21810 98084 21822
rect 98028 21758 98030 21810
rect 98082 21758 98084 21810
rect 97692 21586 97748 21598
rect 97692 21534 97694 21586
rect 97746 21534 97748 21586
rect 97692 20916 97748 21534
rect 97692 20850 97748 20860
rect 97916 20468 97972 20478
rect 97580 20412 97916 20468
rect 97580 20242 97636 20412
rect 97580 20190 97582 20242
rect 97634 20190 97636 20242
rect 97580 20178 97636 20190
rect 96796 19730 96852 19740
rect 97020 19740 97188 19796
rect 97356 20018 97412 20030
rect 97356 19966 97358 20018
rect 97410 19966 97412 20018
rect 96636 19628 96900 19638
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96636 19562 96900 19572
rect 96012 19348 96068 19358
rect 96012 19234 96068 19292
rect 96012 19182 96014 19234
rect 96066 19182 96068 19234
rect 96012 18788 96068 19182
rect 96348 19012 96404 19022
rect 96684 19012 96740 19022
rect 96348 19010 96684 19012
rect 96348 18958 96350 19010
rect 96402 18958 96684 19010
rect 96348 18956 96684 18958
rect 96348 18946 96404 18956
rect 96684 18918 96740 18956
rect 96796 19010 96852 19022
rect 96796 18958 96798 19010
rect 96850 18958 96852 19010
rect 96012 18722 96068 18732
rect 96796 18676 96852 18958
rect 96348 18620 96852 18676
rect 96908 19010 96964 19022
rect 96908 18958 96910 19010
rect 96962 18958 96964 19010
rect 95788 18562 96068 18564
rect 95788 18510 95790 18562
rect 95842 18510 96068 18562
rect 95788 18508 96068 18510
rect 95788 18498 95844 18508
rect 95340 18452 95396 18462
rect 95340 18358 95396 18396
rect 95900 18340 95956 18350
rect 95900 18246 95956 18284
rect 95004 17054 95006 17106
rect 95058 17054 95060 17106
rect 95004 16772 95060 17054
rect 95004 16706 95060 16716
rect 95340 17332 95396 17342
rect 95340 16322 95396 17276
rect 96012 16884 96068 18508
rect 96348 18562 96404 18620
rect 96348 18510 96350 18562
rect 96402 18510 96404 18562
rect 96348 18498 96404 18510
rect 96124 18452 96180 18462
rect 96124 17780 96180 18396
rect 96684 18450 96740 18462
rect 96684 18398 96686 18450
rect 96738 18398 96740 18450
rect 96684 18228 96740 18398
rect 96908 18452 96964 18958
rect 96908 18386 96964 18396
rect 96684 18162 96740 18172
rect 96636 18060 96900 18070
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96636 17994 96900 18004
rect 97020 17892 97076 19740
rect 97244 19234 97300 19246
rect 97244 19182 97246 19234
rect 97298 19182 97300 19234
rect 97244 18900 97300 19182
rect 97244 18834 97300 18844
rect 97356 19012 97412 19966
rect 97468 20020 97524 20030
rect 97468 19926 97524 19964
rect 96124 17714 96180 17724
rect 96908 17836 97076 17892
rect 97244 18452 97300 18462
rect 96236 17108 96292 17118
rect 96236 17106 96628 17108
rect 96236 17054 96238 17106
rect 96290 17054 96628 17106
rect 96236 17052 96628 17054
rect 96236 17042 96292 17052
rect 96572 16996 96628 17052
rect 96908 16996 96964 17836
rect 96572 16940 96964 16996
rect 97244 17778 97300 18396
rect 97244 17726 97246 17778
rect 97298 17726 97300 17778
rect 97244 16996 97300 17726
rect 97356 17106 97412 18956
rect 97692 17778 97748 20412
rect 97916 20402 97972 20412
rect 97804 20130 97860 20142
rect 97804 20078 97806 20130
rect 97858 20078 97860 20130
rect 97804 19122 97860 20078
rect 98028 20132 98084 21758
rect 98140 21700 98196 21710
rect 98140 21606 98196 21644
rect 98028 20066 98084 20076
rect 98252 21586 98308 21598
rect 98252 21534 98254 21586
rect 98306 21534 98308 21586
rect 98140 19348 98196 19358
rect 98252 19348 98308 21534
rect 98700 20578 98756 20590
rect 98700 20526 98702 20578
rect 98754 20526 98756 20578
rect 98700 20468 98756 20526
rect 99148 20580 99204 20590
rect 99148 20486 99204 20524
rect 98700 20402 98756 20412
rect 98140 19346 98308 19348
rect 98140 19294 98142 19346
rect 98194 19294 98308 19346
rect 98140 19292 98308 19294
rect 98364 19906 98420 19918
rect 98364 19854 98366 19906
rect 98418 19854 98420 19906
rect 98140 19282 98196 19292
rect 97804 19070 97806 19122
rect 97858 19070 97860 19122
rect 97804 18900 97860 19070
rect 97804 18834 97860 18844
rect 98028 19010 98084 19022
rect 98028 18958 98030 19010
rect 98082 18958 98084 19010
rect 98028 18788 98084 18958
rect 98252 19012 98308 19022
rect 98252 18918 98308 18956
rect 98364 18788 98420 19854
rect 99260 19124 99316 19134
rect 98812 19012 98868 19022
rect 99260 19012 99316 19068
rect 98812 18918 98868 18956
rect 99148 19010 99316 19012
rect 99148 18958 99262 19010
rect 99314 18958 99316 19010
rect 99148 18956 99316 18958
rect 98028 18732 98420 18788
rect 97692 17726 97694 17778
rect 97746 17726 97748 17778
rect 97692 17714 97748 17726
rect 98140 17778 98196 18732
rect 98924 18452 98980 18462
rect 98924 18338 98980 18396
rect 98924 18286 98926 18338
rect 98978 18286 98980 18338
rect 98924 18274 98980 18286
rect 98140 17726 98142 17778
rect 98194 17726 98196 17778
rect 98140 17714 98196 17726
rect 97356 17054 97358 17106
rect 97410 17054 97412 17106
rect 97356 17042 97412 17054
rect 97804 17442 97860 17454
rect 97804 17390 97806 17442
rect 97858 17390 97860 17442
rect 96012 16828 96180 16884
rect 96124 16772 96180 16828
rect 96348 16882 96404 16894
rect 96348 16830 96350 16882
rect 96402 16830 96404 16882
rect 96348 16772 96404 16830
rect 96684 16882 96740 16940
rect 97244 16930 97300 16940
rect 96684 16830 96686 16882
rect 96738 16830 96740 16882
rect 96684 16818 96740 16830
rect 97020 16882 97076 16894
rect 97020 16830 97022 16882
rect 97074 16830 97076 16882
rect 96124 16716 96404 16772
rect 96572 16770 96628 16782
rect 96572 16718 96574 16770
rect 96626 16718 96628 16770
rect 96572 16660 96628 16718
rect 97020 16772 97076 16830
rect 97580 16882 97636 16894
rect 97580 16830 97582 16882
rect 97634 16830 97636 16882
rect 97020 16706 97076 16716
rect 97468 16772 97524 16782
rect 97468 16678 97524 16716
rect 95340 16270 95342 16322
rect 95394 16270 95396 16322
rect 95340 16210 95396 16270
rect 95340 16158 95342 16210
rect 95394 16158 95396 16210
rect 95340 16146 95396 16158
rect 96460 16604 96628 16660
rect 95788 16098 95844 16110
rect 95788 16046 95790 16098
rect 95842 16046 95844 16098
rect 94668 14242 94724 14252
rect 94780 15986 94836 15998
rect 94780 15934 94782 15986
rect 94834 15934 94836 15986
rect 94220 11666 94276 11676
rect 94444 13804 94612 13860
rect 93996 11564 94164 11620
rect 94332 11620 94388 11630
rect 93996 10500 94052 11564
rect 94108 11396 94164 11406
rect 94332 11396 94388 11564
rect 94108 11394 94388 11396
rect 94108 11342 94110 11394
rect 94162 11342 94388 11394
rect 94108 11340 94388 11342
rect 94108 11060 94164 11340
rect 94108 10994 94164 11004
rect 94220 11172 94276 11182
rect 94220 10500 94276 11116
rect 94444 10724 94500 13804
rect 94668 13524 94724 13534
rect 94668 13430 94724 13468
rect 94556 12962 94612 12974
rect 94556 12910 94558 12962
rect 94610 12910 94612 12962
rect 94556 12404 94612 12910
rect 94780 12404 94836 15934
rect 94892 15876 94948 15886
rect 94892 15782 94948 15820
rect 94892 15204 94948 15214
rect 94892 14530 94948 15148
rect 95116 15204 95172 15242
rect 95116 15138 95172 15148
rect 95228 14644 95284 14654
rect 95228 14642 95732 14644
rect 95228 14590 95230 14642
rect 95282 14590 95732 14642
rect 95228 14588 95732 14590
rect 95228 14578 95284 14588
rect 94892 14478 94894 14530
rect 94946 14478 94948 14530
rect 94892 14466 94948 14478
rect 95452 14308 95508 14318
rect 95004 13860 95060 13870
rect 94780 12348 94948 12404
rect 94556 12338 94612 12348
rect 94780 12180 94836 12190
rect 94780 12086 94836 12124
rect 94892 11956 94948 12348
rect 94780 11900 94948 11956
rect 94556 11620 94612 11630
rect 94556 11394 94612 11564
rect 94556 11342 94558 11394
rect 94610 11342 94612 11394
rect 94556 11330 94612 11342
rect 94668 11508 94724 11518
rect 94668 10948 94724 11452
rect 94668 10882 94724 10892
rect 94444 10658 94500 10668
rect 94556 10836 94612 10846
rect 94052 10444 94164 10500
rect 93996 10434 94052 10444
rect 93884 10210 93940 10220
rect 93772 9828 93828 9838
rect 93548 9826 93940 9828
rect 93548 9774 93774 9826
rect 93826 9774 93940 9826
rect 93548 9772 93940 9774
rect 93772 9762 93828 9772
rect 93436 9538 93492 9548
rect 93772 9602 93828 9614
rect 93772 9550 93774 9602
rect 93826 9550 93828 9602
rect 93324 9324 93492 9380
rect 93324 9156 93380 9166
rect 93324 9062 93380 9100
rect 93212 7858 93268 7868
rect 93324 8370 93380 8382
rect 93324 8318 93326 8370
rect 93378 8318 93380 8370
rect 93212 6916 93268 6926
rect 93100 6860 93212 6916
rect 93212 6850 93268 6860
rect 92764 6626 92820 6636
rect 92652 5954 92708 5964
rect 93100 6244 93156 6254
rect 92428 5236 92484 5246
rect 92428 5142 92484 5180
rect 92316 4956 92820 5012
rect 92092 4946 92148 4956
rect 91756 4900 91812 4910
rect 91756 4806 91812 4844
rect 92764 4450 92820 4956
rect 92764 4398 92766 4450
rect 92818 4398 92820 4450
rect 92540 4340 92596 4350
rect 92316 3780 92372 3790
rect 92316 3554 92372 3724
rect 92316 3502 92318 3554
rect 92370 3502 92372 3554
rect 92316 3490 92372 3502
rect 91644 802 91700 812
rect 92540 800 92596 4284
rect 92764 4116 92820 4398
rect 92764 4050 92820 4060
rect 93100 3666 93156 6188
rect 93324 6132 93380 8318
rect 93436 6468 93492 9324
rect 93436 6402 93492 6412
rect 93660 8260 93716 8270
rect 93660 8146 93716 8204
rect 93660 8094 93662 8146
rect 93714 8094 93716 8146
rect 93324 6066 93380 6076
rect 93548 4228 93604 4238
rect 93548 4134 93604 4172
rect 93212 3780 93268 3790
rect 93660 3780 93716 8094
rect 93772 6356 93828 9550
rect 93884 8258 93940 9772
rect 93884 8206 93886 8258
rect 93938 8206 93940 8258
rect 93884 6692 93940 8206
rect 93996 9826 94052 9838
rect 93996 9774 93998 9826
rect 94050 9774 94052 9826
rect 93996 8260 94052 9774
rect 94108 9604 94164 10444
rect 94220 10406 94276 10444
rect 94332 10612 94388 10622
rect 94108 9538 94164 9548
rect 94220 9938 94276 9950
rect 94220 9886 94222 9938
rect 94274 9886 94276 9938
rect 94108 9044 94164 9054
rect 94108 8950 94164 8988
rect 94108 8484 94164 8494
rect 94220 8484 94276 9886
rect 94332 9492 94388 10556
rect 94556 10610 94612 10780
rect 94556 10558 94558 10610
rect 94610 10558 94612 10610
rect 94556 10546 94612 10558
rect 94556 10052 94612 10062
rect 94332 9426 94388 9436
rect 94444 9996 94556 10052
rect 94444 9266 94500 9996
rect 94556 9986 94612 9996
rect 94444 9214 94446 9266
rect 94498 9214 94500 9266
rect 94444 9202 94500 9214
rect 94556 9604 94612 9614
rect 94556 9044 94612 9548
rect 94108 8482 94276 8484
rect 94108 8430 94110 8482
rect 94162 8430 94276 8482
rect 94108 8428 94276 8430
rect 94444 8988 94612 9044
rect 94108 8372 94164 8428
rect 94108 8306 94164 8316
rect 94332 8260 94388 8270
rect 93996 8194 94052 8204
rect 94220 8258 94388 8260
rect 94220 8206 94334 8258
rect 94386 8206 94388 8258
rect 94220 8204 94388 8206
rect 94220 7700 94276 8204
rect 94332 8194 94388 8204
rect 93996 7644 94276 7700
rect 93996 7588 94052 7644
rect 93996 7474 94052 7532
rect 93996 7422 93998 7474
rect 94050 7422 94052 7474
rect 93996 7410 94052 7422
rect 93884 6626 93940 6636
rect 94220 7252 94276 7262
rect 94220 6580 94276 7196
rect 94108 6578 94276 6580
rect 94108 6526 94222 6578
rect 94274 6526 94276 6578
rect 94108 6524 94276 6526
rect 93772 6300 94052 6356
rect 93884 5794 93940 5806
rect 93884 5742 93886 5794
rect 93938 5742 93940 5794
rect 93884 4452 93940 5742
rect 93996 5010 94052 6300
rect 93996 4958 93998 5010
rect 94050 4958 94052 5010
rect 93996 4946 94052 4958
rect 93884 4386 93940 4396
rect 93212 3778 93716 3780
rect 93212 3726 93214 3778
rect 93266 3726 93716 3778
rect 93212 3724 93716 3726
rect 93884 4116 93940 4126
rect 93212 3714 93268 3724
rect 93100 3614 93102 3666
rect 93154 3614 93156 3666
rect 93100 3602 93156 3614
rect 93884 800 93940 4060
rect 94108 4004 94164 6524
rect 94220 6514 94276 6524
rect 94332 7250 94388 7262
rect 94332 7198 94334 7250
rect 94386 7198 94388 7250
rect 94220 6132 94276 6142
rect 94220 6038 94276 6076
rect 94220 5908 94276 5918
rect 94220 5122 94276 5852
rect 94220 5070 94222 5122
rect 94274 5070 94276 5122
rect 94220 5058 94276 5070
rect 94108 3938 94164 3948
rect 94108 3666 94164 3678
rect 94108 3614 94110 3666
rect 94162 3614 94164 3666
rect 94108 3556 94164 3614
rect 94108 1540 94164 3500
rect 94332 3442 94388 7198
rect 94332 3390 94334 3442
rect 94386 3390 94388 3442
rect 94332 3378 94388 3390
rect 94108 1474 94164 1484
rect 94444 1316 94500 8988
rect 94556 8820 94612 8830
rect 94780 8820 94836 11900
rect 95004 11788 95060 13804
rect 95228 13636 95284 13646
rect 95284 13580 95396 13636
rect 95228 13542 95284 13580
rect 95228 12068 95284 12078
rect 95228 11974 95284 12012
rect 95004 11732 95172 11788
rect 95116 10052 95172 11732
rect 95340 11732 95396 13580
rect 95340 11666 95396 11676
rect 95228 11508 95284 11518
rect 95228 11414 95284 11452
rect 95340 10836 95396 10846
rect 95116 9986 95172 9996
rect 95228 10780 95340 10836
rect 95228 9828 95284 10780
rect 95340 10770 95396 10780
rect 95228 9762 95284 9772
rect 95340 10610 95396 10622
rect 95340 10558 95342 10610
rect 95394 10558 95396 10610
rect 95228 9604 95284 9614
rect 94612 8764 94836 8820
rect 94892 9156 94948 9166
rect 94892 8930 94948 9100
rect 94892 8878 94894 8930
rect 94946 8878 94948 8930
rect 94556 7812 94612 8764
rect 94556 7746 94612 7756
rect 94668 8148 94724 8158
rect 94668 7698 94724 8092
rect 94780 8036 94836 8046
rect 94780 7942 94836 7980
rect 94892 7812 94948 8878
rect 95228 8932 95284 9548
rect 95228 8258 95284 8876
rect 95228 8206 95230 8258
rect 95282 8206 95284 8258
rect 95228 8194 95284 8206
rect 94668 7646 94670 7698
rect 94722 7646 94724 7698
rect 94668 7634 94724 7646
rect 94780 7756 94948 7812
rect 94556 7588 94612 7598
rect 94556 7474 94612 7532
rect 94556 7422 94558 7474
rect 94610 7422 94612 7474
rect 94556 6356 94612 7422
rect 94556 6290 94612 6300
rect 94668 6692 94724 6702
rect 94668 5794 94724 6636
rect 94668 5742 94670 5794
rect 94722 5742 94724 5794
rect 94668 5730 94724 5742
rect 94556 4452 94612 4462
rect 94556 4358 94612 4396
rect 94780 1428 94836 7756
rect 94892 7586 94948 7598
rect 94892 7534 94894 7586
rect 94946 7534 94948 7586
rect 94892 7364 94948 7534
rect 95004 7476 95060 7486
rect 95004 7382 95060 7420
rect 94892 7298 94948 7308
rect 95228 6578 95284 6590
rect 95228 6526 95230 6578
rect 95282 6526 95284 6578
rect 94892 6468 94948 6478
rect 95228 6468 95284 6526
rect 94892 6374 94948 6412
rect 95004 6412 95228 6468
rect 95004 5908 95060 6412
rect 95228 6402 95284 6412
rect 95228 6132 95284 6142
rect 95228 6038 95284 6076
rect 95116 6020 95172 6030
rect 95116 5926 95172 5964
rect 95004 5460 95060 5852
rect 95004 5404 95172 5460
rect 95004 5124 95060 5134
rect 95004 3554 95060 5068
rect 95004 3502 95006 3554
rect 95058 3502 95060 3554
rect 95004 3490 95060 3502
rect 95116 3556 95172 5404
rect 95228 5012 95284 5022
rect 95340 5012 95396 10558
rect 95452 7588 95508 14252
rect 95564 12292 95620 12302
rect 95564 11394 95620 12236
rect 95564 11342 95566 11394
rect 95618 11342 95620 11394
rect 95564 11330 95620 11342
rect 95676 10834 95732 14588
rect 95788 12180 95844 16046
rect 96460 16098 96516 16604
rect 97244 16548 97300 16558
rect 96636 16492 96900 16502
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96636 16426 96900 16436
rect 96460 16046 96462 16098
rect 96514 16046 96516 16098
rect 96460 16034 96516 16046
rect 96012 15652 96068 15662
rect 96012 15314 96068 15596
rect 96012 15262 96014 15314
rect 96066 15262 96068 15314
rect 96012 15250 96068 15262
rect 95788 12114 95844 12124
rect 95900 15204 95956 15242
rect 95900 13634 95956 15148
rect 96636 14924 96900 14934
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96636 14858 96900 14868
rect 97132 14644 97188 14654
rect 97020 14588 97132 14644
rect 96908 14308 96964 14318
rect 96460 14306 96964 14308
rect 96460 14254 96910 14306
rect 96962 14254 96964 14306
rect 96460 14252 96964 14254
rect 96124 13972 96180 13982
rect 96012 13748 96068 13758
rect 96012 13654 96068 13692
rect 95900 13582 95902 13634
rect 95954 13582 95956 13634
rect 95900 12962 95956 13582
rect 95900 12910 95902 12962
rect 95954 12910 95956 12962
rect 95900 12066 95956 12910
rect 96124 12178 96180 13916
rect 96348 13412 96404 13422
rect 96124 12126 96126 12178
rect 96178 12126 96180 12178
rect 96124 12114 96180 12126
rect 96236 12962 96292 12974
rect 96236 12910 96238 12962
rect 96290 12910 96292 12962
rect 95900 12014 95902 12066
rect 95954 12014 95956 12066
rect 95900 12002 95956 12014
rect 96124 11956 96180 11966
rect 96236 11956 96292 12910
rect 96348 12964 96404 13356
rect 96348 12870 96404 12908
rect 96180 11900 96292 11956
rect 96124 11890 96180 11900
rect 96460 11732 96516 14252
rect 96908 14242 96964 14252
rect 96636 13356 96900 13366
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96636 13290 96900 13300
rect 96236 11676 96516 11732
rect 96636 11788 96900 11798
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96636 11722 96900 11732
rect 95676 10782 95678 10834
rect 95730 10782 95732 10834
rect 95676 10770 95732 10782
rect 95788 11508 95844 11518
rect 95788 10722 95844 11452
rect 95788 10670 95790 10722
rect 95842 10670 95844 10722
rect 95564 10052 95620 10062
rect 95564 8258 95620 9996
rect 95788 9714 95844 10670
rect 95788 9662 95790 9714
rect 95842 9662 95844 9714
rect 95788 9156 95844 9662
rect 96124 10610 96180 10622
rect 96124 10558 96126 10610
rect 96178 10558 96180 10610
rect 96012 9492 96068 9502
rect 95900 9156 95956 9166
rect 95788 9100 95900 9156
rect 95900 9090 95956 9100
rect 95788 8930 95844 8942
rect 95788 8878 95790 8930
rect 95842 8878 95844 8930
rect 95676 8484 95732 8494
rect 95788 8484 95844 8878
rect 95900 8820 95956 8830
rect 95900 8726 95956 8764
rect 95732 8428 95844 8484
rect 95676 8418 95732 8428
rect 95564 8206 95566 8258
rect 95618 8206 95620 8258
rect 95564 8194 95620 8206
rect 95676 8260 95732 8270
rect 95676 8146 95732 8204
rect 95676 8094 95678 8146
rect 95730 8094 95732 8146
rect 95676 8082 95732 8094
rect 95788 8146 95844 8158
rect 95788 8094 95790 8146
rect 95842 8094 95844 8146
rect 95788 8036 95844 8094
rect 95788 7970 95844 7980
rect 95452 7522 95508 7532
rect 95788 7700 95844 7710
rect 95788 7586 95844 7644
rect 95900 7700 95956 7710
rect 96012 7700 96068 9436
rect 96124 8372 96180 10558
rect 96236 10052 96292 11676
rect 96908 11396 96964 11406
rect 97020 11396 97076 14588
rect 97132 14578 97188 14588
rect 96908 11394 97076 11396
rect 96908 11342 96910 11394
rect 96962 11342 97076 11394
rect 96908 11340 97076 11342
rect 96348 11172 96404 11182
rect 96572 11172 96628 11182
rect 96348 11078 96404 11116
rect 96460 11170 96628 11172
rect 96460 11118 96574 11170
rect 96626 11118 96628 11170
rect 96460 11116 96628 11118
rect 96460 10052 96516 11116
rect 96572 11106 96628 11116
rect 96796 11170 96852 11182
rect 96796 11118 96798 11170
rect 96850 11118 96852 11170
rect 96796 10836 96852 11118
rect 96796 10770 96852 10780
rect 96908 10500 96964 11340
rect 97244 11284 97300 16492
rect 97580 16212 97636 16830
rect 97580 16146 97636 16156
rect 97580 15314 97636 15326
rect 97580 15262 97582 15314
rect 97634 15262 97636 15314
rect 97580 15148 97636 15262
rect 97580 15092 97748 15148
rect 97468 14308 97524 14318
rect 97468 14214 97524 14252
rect 97692 13748 97748 15092
rect 97804 14532 97860 17390
rect 98252 17442 98308 17454
rect 98252 17390 98254 17442
rect 98306 17390 98308 17442
rect 98252 17332 98308 17390
rect 98700 17444 98756 17454
rect 98700 17350 98756 17388
rect 98252 17266 98308 17276
rect 97916 17220 97972 17230
rect 97916 16882 97972 17164
rect 98252 16996 98308 17006
rect 98252 16902 98308 16940
rect 97916 16830 97918 16882
rect 97970 16830 97972 16882
rect 97916 15988 97972 16830
rect 98812 16772 98868 16782
rect 98588 16770 98868 16772
rect 98588 16718 98814 16770
rect 98866 16718 98868 16770
rect 98588 16716 98868 16718
rect 97916 15922 97972 15932
rect 98364 16658 98420 16670
rect 98364 16606 98366 16658
rect 98418 16606 98420 16658
rect 97804 14466 97860 14476
rect 97916 15314 97972 15326
rect 97916 15262 97918 15314
rect 97970 15262 97972 15314
rect 97916 14420 97972 15262
rect 98252 14756 98308 14766
rect 98252 14642 98308 14700
rect 98252 14590 98254 14642
rect 98306 14590 98308 14642
rect 98252 14578 98308 14590
rect 97916 14364 98308 14420
rect 97804 14306 97860 14318
rect 97804 14254 97806 14306
rect 97858 14254 97860 14306
rect 97804 13972 97860 14254
rect 97804 13916 98196 13972
rect 97468 13692 97748 13748
rect 97804 13748 97860 13758
rect 97356 13188 97412 13198
rect 97356 13094 97412 13132
rect 97468 12068 97524 13692
rect 97804 12964 97860 13692
rect 97804 12178 97860 12908
rect 97804 12126 97806 12178
rect 97858 12126 97860 12178
rect 97804 12114 97860 12126
rect 98028 13634 98084 13646
rect 98028 13582 98030 13634
rect 98082 13582 98084 13634
rect 97468 12012 97636 12068
rect 97132 11282 97300 11284
rect 97132 11230 97246 11282
rect 97298 11230 97300 11282
rect 97132 11228 97300 11230
rect 96908 10434 96964 10444
rect 97020 11172 97076 11182
rect 96636 10220 96900 10230
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96636 10154 96900 10164
rect 96236 9996 96404 10052
rect 96124 8306 96180 8316
rect 96236 9828 96292 9838
rect 96236 8370 96292 9772
rect 96348 9380 96404 9996
rect 96460 9986 96516 9996
rect 97020 10052 97076 11116
rect 97020 9986 97076 9996
rect 96684 9826 96740 9838
rect 96684 9774 96686 9826
rect 96738 9774 96740 9826
rect 96684 9492 96740 9774
rect 96684 9426 96740 9436
rect 96348 9324 96516 9380
rect 96236 8318 96238 8370
rect 96290 8318 96292 8370
rect 96236 8306 96292 8318
rect 96348 9156 96404 9166
rect 95900 7698 96068 7700
rect 95900 7646 95902 7698
rect 95954 7646 96068 7698
rect 95900 7644 96068 7646
rect 95900 7634 95956 7644
rect 95788 7534 95790 7586
rect 95842 7534 95844 7586
rect 95788 7522 95844 7534
rect 96348 7586 96404 9100
rect 96460 8148 96516 9324
rect 96572 9042 96628 9054
rect 96572 8990 96574 9042
rect 96626 8990 96628 9042
rect 96572 8820 96628 8990
rect 96572 8754 96628 8764
rect 96636 8652 96900 8662
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96636 8586 96900 8596
rect 96460 8092 96628 8148
rect 96348 7534 96350 7586
rect 96402 7534 96404 7586
rect 96348 7522 96404 7534
rect 96236 7474 96292 7486
rect 96236 7422 96238 7474
rect 96290 7422 96292 7474
rect 96012 6804 96068 6814
rect 96236 6804 96292 7422
rect 96572 7252 96628 8092
rect 96572 7186 96628 7196
rect 97020 7812 97076 7822
rect 96636 7084 96900 7094
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96636 7018 96900 7028
rect 96012 6802 96292 6804
rect 96012 6750 96014 6802
rect 96066 6750 96292 6802
rect 96012 6748 96292 6750
rect 95452 6690 95508 6702
rect 95452 6638 95454 6690
rect 95506 6638 95508 6690
rect 95452 5908 95508 6638
rect 95564 5908 95620 5918
rect 95452 5852 95564 5908
rect 95564 5124 95620 5852
rect 95564 5030 95620 5068
rect 95228 5010 95396 5012
rect 95228 4958 95230 5010
rect 95282 4958 95396 5010
rect 95228 4956 95396 4958
rect 96012 5012 96068 6748
rect 96236 6356 96292 6366
rect 96236 6020 96292 6300
rect 95228 4946 95284 4956
rect 96012 4946 96068 4956
rect 96124 6018 96292 6020
rect 96124 5966 96238 6018
rect 96290 5966 96292 6018
rect 96124 5964 96292 5966
rect 95340 4788 95396 4798
rect 95228 3556 95284 3566
rect 95116 3554 95284 3556
rect 95116 3502 95230 3554
rect 95282 3502 95284 3554
rect 95116 3500 95284 3502
rect 95228 3490 95284 3500
rect 95340 3388 95396 4732
rect 96124 4788 96180 5964
rect 96236 5954 96292 5964
rect 96636 5516 96900 5526
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96636 5450 96900 5460
rect 96124 4722 96180 4732
rect 96236 5010 96292 5022
rect 96236 4958 96238 5010
rect 96290 4958 96292 5010
rect 96236 4900 96292 4958
rect 96236 4340 96292 4844
rect 96236 4274 96292 4284
rect 96012 4116 96068 4126
rect 96012 4022 96068 4060
rect 96636 3948 96900 3958
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96636 3882 96900 3892
rect 97020 3892 97076 7756
rect 97020 3826 97076 3836
rect 96908 3668 96964 3678
rect 94780 1362 94836 1372
rect 95228 3332 95396 3388
rect 96572 3444 96628 3454
rect 94444 1250 94500 1260
rect 95228 800 95284 3332
rect 96572 800 96628 3388
rect 96908 3442 96964 3612
rect 96908 3390 96910 3442
rect 96962 3390 96964 3442
rect 96908 3378 96964 3390
rect 97132 2548 97188 11228
rect 97244 11218 97300 11228
rect 97356 11170 97412 11182
rect 97356 11118 97358 11170
rect 97410 11118 97412 11170
rect 97244 10500 97300 10510
rect 97244 9716 97300 10444
rect 97244 9650 97300 9660
rect 97356 9604 97412 11118
rect 97356 9538 97412 9548
rect 97468 10610 97524 10622
rect 97468 10558 97470 10610
rect 97522 10558 97524 10610
rect 97468 8484 97524 10558
rect 97580 9938 97636 12012
rect 97804 11844 97860 11854
rect 97804 11172 97860 11788
rect 97916 11732 97972 11742
rect 97916 11508 97972 11676
rect 97916 11442 97972 11452
rect 97580 9886 97582 9938
rect 97634 9886 97636 9938
rect 97580 9874 97636 9886
rect 97692 11170 97860 11172
rect 97692 11118 97806 11170
rect 97858 11118 97860 11170
rect 97692 11116 97860 11118
rect 97580 9716 97636 9726
rect 97580 9268 97636 9660
rect 97692 9380 97748 11116
rect 97804 11106 97860 11116
rect 97692 9314 97748 9324
rect 97804 10388 97860 10398
rect 97580 9202 97636 9212
rect 97468 8418 97524 8428
rect 97244 6468 97300 6478
rect 97244 5460 97300 6412
rect 97804 5572 97860 10332
rect 97916 9604 97972 9614
rect 97916 9042 97972 9548
rect 97916 8990 97918 9042
rect 97970 8990 97972 9042
rect 97916 8978 97972 8990
rect 97916 8372 97972 8382
rect 97916 7812 97972 8316
rect 97916 7746 97972 7756
rect 98028 7586 98084 13582
rect 98140 12292 98196 13916
rect 98252 13748 98308 14364
rect 98252 13682 98308 13692
rect 98364 12964 98420 16606
rect 98588 16548 98644 16716
rect 98812 16706 98868 16716
rect 99148 16548 99204 18956
rect 99260 18946 99316 18956
rect 99708 18788 99764 18798
rect 99708 18450 99764 18732
rect 99708 18398 99710 18450
rect 99762 18398 99764 18450
rect 99484 18340 99540 18350
rect 98588 16482 98644 16492
rect 98700 16492 99204 16548
rect 99260 17442 99316 17454
rect 99260 17390 99262 17442
rect 99314 17390 99316 17442
rect 98140 12226 98196 12236
rect 98252 12908 98420 12964
rect 98700 14642 98756 16492
rect 98812 16212 98868 16222
rect 98868 16156 99092 16212
rect 98812 16118 98868 16156
rect 98812 15092 98868 15102
rect 98812 14998 98868 15036
rect 98700 14590 98702 14642
rect 98754 14590 98756 14642
rect 98140 12066 98196 12078
rect 98140 12014 98142 12066
rect 98194 12014 98196 12066
rect 98140 9154 98196 12014
rect 98252 11396 98308 12908
rect 98364 12738 98420 12750
rect 98364 12686 98366 12738
rect 98418 12686 98420 12738
rect 98364 11732 98420 12686
rect 98364 11666 98420 11676
rect 98476 11620 98532 11630
rect 98532 11564 98644 11620
rect 98476 11554 98532 11564
rect 98252 11340 98420 11396
rect 98252 11170 98308 11182
rect 98252 11118 98254 11170
rect 98306 11118 98308 11170
rect 98252 11060 98308 11118
rect 98252 10276 98308 11004
rect 98252 10210 98308 10220
rect 98140 9102 98142 9154
rect 98194 9102 98196 9154
rect 98140 9090 98196 9102
rect 98252 9268 98308 9278
rect 98028 7534 98030 7586
rect 98082 7534 98084 7586
rect 98028 7522 98084 7534
rect 98140 8932 98196 8942
rect 97916 7474 97972 7486
rect 97916 7422 97918 7474
rect 97970 7422 97972 7474
rect 97916 6132 97972 7422
rect 98140 6690 98196 8876
rect 98140 6638 98142 6690
rect 98194 6638 98196 6690
rect 98140 6626 98196 6638
rect 97916 6066 97972 6076
rect 97804 5506 97860 5516
rect 97244 5394 97300 5404
rect 98252 5124 98308 9212
rect 98364 8372 98420 11340
rect 98588 11172 98644 11564
rect 98700 11396 98756 14590
rect 99036 14642 99092 16156
rect 99036 14590 99038 14642
rect 99090 14590 99092 14642
rect 99036 14578 99092 14590
rect 98924 14532 98980 14542
rect 98812 13524 98868 13534
rect 98812 13430 98868 13468
rect 98812 13300 98868 13310
rect 98812 12738 98868 13244
rect 98812 12686 98814 12738
rect 98866 12686 98868 12738
rect 98812 12180 98868 12686
rect 98812 12114 98868 12124
rect 98812 11956 98868 11966
rect 98812 11862 98868 11900
rect 98700 11340 98868 11396
rect 98700 11172 98756 11182
rect 98588 11170 98756 11172
rect 98588 11118 98702 11170
rect 98754 11118 98756 11170
rect 98588 11116 98756 11118
rect 98700 11106 98756 11116
rect 98812 9380 98868 11340
rect 98924 10612 98980 14476
rect 99260 14532 99316 17390
rect 99484 16212 99540 18284
rect 99708 18340 99764 18398
rect 99708 18274 99764 18284
rect 99820 18452 99876 22318
rect 103516 22258 103572 22270
rect 103516 22206 103518 22258
rect 103570 22206 103572 22258
rect 103068 21474 103124 21486
rect 103068 21422 103070 21474
rect 103122 21422 103124 21474
rect 101276 20580 101332 20590
rect 100828 20132 100884 20142
rect 100828 20018 100884 20076
rect 100828 19966 100830 20018
rect 100882 19966 100884 20018
rect 100828 19954 100884 19966
rect 101276 20132 101332 20524
rect 103068 20244 103124 21422
rect 103516 20802 103572 22206
rect 103964 21476 104020 21486
rect 103964 21382 104020 21420
rect 103516 20750 103518 20802
rect 103570 20750 103572 20802
rect 103292 20580 103348 20590
rect 103516 20580 103572 20750
rect 103348 20524 103572 20580
rect 103292 20486 103348 20524
rect 103068 20178 103124 20188
rect 101836 20132 101892 20142
rect 101276 20130 101892 20132
rect 101276 20078 101838 20130
rect 101890 20078 101892 20130
rect 101276 20076 101892 20078
rect 101276 20018 101332 20076
rect 101836 20066 101892 20076
rect 101276 19966 101278 20018
rect 101330 19966 101332 20018
rect 101276 19954 101332 19966
rect 99932 19124 99988 19134
rect 99932 19030 99988 19068
rect 104076 19124 104132 25676
rect 104412 21588 104468 21598
rect 104188 21586 104468 21588
rect 104188 21534 104414 21586
rect 104466 21534 104468 21586
rect 104188 21532 104468 21534
rect 104188 20244 104244 21532
rect 104412 21522 104468 21532
rect 104300 20804 104356 20814
rect 104300 20802 104804 20804
rect 104300 20750 104302 20802
rect 104354 20750 104804 20802
rect 104300 20748 104804 20750
rect 104300 20738 104356 20748
rect 104188 20178 104244 20188
rect 104748 20242 104804 20748
rect 104748 20190 104750 20242
rect 104802 20190 104804 20242
rect 104748 20178 104804 20190
rect 104860 20244 104916 26126
rect 104972 26180 105028 26238
rect 105980 26290 106036 26302
rect 105980 26238 105982 26290
rect 106034 26238 106036 26290
rect 104972 26114 105028 26124
rect 105532 26180 105588 26190
rect 105532 25618 105588 26124
rect 105980 26180 106036 26238
rect 105980 26114 106036 26124
rect 107548 26178 107604 26190
rect 107548 26126 107550 26178
rect 107602 26126 107604 26178
rect 106428 26068 106484 26078
rect 106428 26066 106708 26068
rect 106428 26014 106430 26066
rect 106482 26014 106708 26066
rect 106428 26012 106708 26014
rect 106428 26002 106484 26012
rect 105532 25566 105534 25618
rect 105586 25566 105588 25618
rect 105532 25554 105588 25566
rect 106092 25508 106148 25518
rect 106092 25414 106148 25452
rect 106540 25508 106596 25518
rect 106540 25414 106596 25452
rect 105420 21476 105476 21486
rect 104860 20188 105364 20244
rect 104076 19058 104132 19068
rect 104636 20020 104692 20030
rect 104860 20020 104916 20188
rect 104636 20018 104916 20020
rect 104636 19966 104638 20018
rect 104690 19966 104916 20018
rect 104636 19964 104916 19966
rect 104972 20018 105028 20030
rect 104972 19966 104974 20018
rect 105026 19966 105028 20018
rect 100268 19010 100324 19022
rect 100268 18958 100270 19010
rect 100322 18958 100324 19010
rect 99820 17666 99876 18396
rect 99820 17614 99822 17666
rect 99874 17614 99876 17666
rect 99820 17602 99876 17614
rect 100044 18450 100100 18462
rect 100044 18398 100046 18450
rect 100098 18398 100100 18450
rect 100044 18340 100100 18398
rect 99596 17108 99652 17118
rect 99820 17108 99876 17118
rect 99596 17106 99820 17108
rect 99596 17054 99598 17106
rect 99650 17054 99820 17106
rect 99596 17052 99820 17054
rect 99596 17042 99652 17052
rect 99820 17014 99876 17052
rect 100044 17108 100100 18284
rect 100044 17042 100100 17052
rect 100156 16994 100212 17006
rect 100156 16942 100158 16994
rect 100210 16942 100212 16994
rect 100044 16772 100100 16782
rect 100156 16772 100212 16942
rect 100100 16716 100212 16772
rect 100044 16706 100100 16716
rect 100268 16660 100324 18958
rect 100828 19012 100884 19022
rect 100380 18562 100436 18574
rect 100380 18510 100382 18562
rect 100434 18510 100436 18562
rect 100380 18452 100436 18510
rect 100380 18386 100436 18396
rect 100828 18338 100884 18956
rect 101388 18452 101444 18462
rect 100828 18286 100830 18338
rect 100882 18286 100884 18338
rect 100828 17108 100884 18286
rect 100716 17052 100884 17108
rect 100940 18450 101444 18452
rect 100940 18398 101390 18450
rect 101442 18398 101444 18450
rect 100940 18396 101444 18398
rect 100940 17106 100996 18396
rect 101388 18386 101444 18396
rect 101724 18450 101780 18462
rect 101724 18398 101726 18450
rect 101778 18398 101780 18450
rect 101724 18340 101780 18398
rect 101948 18452 102004 18462
rect 101724 18274 101780 18284
rect 101836 18338 101892 18350
rect 101836 18286 101838 18338
rect 101890 18286 101892 18338
rect 101724 17554 101780 17566
rect 101724 17502 101726 17554
rect 101778 17502 101780 17554
rect 101724 17444 101780 17502
rect 101612 17388 101724 17444
rect 100940 17054 100942 17106
rect 100994 17054 100996 17106
rect 99260 14466 99316 14476
rect 99372 16156 99540 16212
rect 100156 16604 100324 16660
rect 100380 16884 100436 16894
rect 99148 14308 99204 14318
rect 99148 14306 99316 14308
rect 99148 14254 99150 14306
rect 99202 14254 99316 14306
rect 99148 14252 99316 14254
rect 99148 14242 99204 14252
rect 99148 11620 99204 11630
rect 99148 11506 99204 11564
rect 99148 11454 99150 11506
rect 99202 11454 99204 11506
rect 99148 11442 99204 11454
rect 99260 10836 99316 14252
rect 99372 13748 99428 16156
rect 99820 15874 99876 15886
rect 99820 15822 99822 15874
rect 99874 15822 99876 15874
rect 99372 13682 99428 13692
rect 99596 14532 99652 14542
rect 99820 14532 99876 15822
rect 100044 15314 100100 15326
rect 100044 15262 100046 15314
rect 100098 15262 100100 15314
rect 100044 14644 100100 15262
rect 100156 14756 100212 16604
rect 100268 16212 100324 16222
rect 100380 16212 100436 16828
rect 100268 16210 100436 16212
rect 100268 16158 100270 16210
rect 100322 16158 100436 16210
rect 100268 16156 100436 16158
rect 100492 16772 100548 16782
rect 100268 16146 100324 16156
rect 100380 15652 100436 15662
rect 100156 14690 100212 14700
rect 100268 15538 100324 15550
rect 100268 15486 100270 15538
rect 100322 15486 100324 15538
rect 100044 14578 100100 14588
rect 99596 14530 99876 14532
rect 99596 14478 99598 14530
rect 99650 14478 99876 14530
rect 99596 14476 99876 14478
rect 99932 14532 99988 14542
rect 99596 13300 99652 14476
rect 99596 13234 99652 13244
rect 99708 12964 99764 12974
rect 99708 12066 99764 12908
rect 99708 12014 99710 12066
rect 99762 12014 99764 12066
rect 99708 12002 99764 12014
rect 99820 11172 99876 11182
rect 99820 11078 99876 11116
rect 99820 10836 99876 10846
rect 99260 10780 99428 10836
rect 99036 10612 99092 10622
rect 99260 10612 99316 10622
rect 98924 10556 99036 10612
rect 99036 10546 99092 10556
rect 99148 10610 99316 10612
rect 99148 10558 99262 10610
rect 99314 10558 99316 10610
rect 99148 10556 99316 10558
rect 99148 10052 99204 10556
rect 99260 10546 99316 10556
rect 99148 9826 99204 9996
rect 99148 9774 99150 9826
rect 99202 9774 99204 9826
rect 99036 9716 99092 9726
rect 99036 9622 99092 9660
rect 99148 9380 99204 9774
rect 98812 9324 99092 9380
rect 99036 9044 99092 9324
rect 99148 9314 99204 9324
rect 98364 8306 98420 8316
rect 98476 8820 98532 8830
rect 98364 8148 98420 8158
rect 98364 8054 98420 8092
rect 98252 5058 98308 5068
rect 97244 4788 97300 4798
rect 97244 3554 97300 4732
rect 98364 4340 98420 4350
rect 98476 4340 98532 8764
rect 98700 8708 98756 8718
rect 98588 8652 98700 8708
rect 98588 5796 98644 8652
rect 98700 8642 98756 8652
rect 99036 8260 99092 8988
rect 99148 8260 99204 8270
rect 99036 8204 99148 8260
rect 98924 6692 98980 6702
rect 99036 6692 99092 8204
rect 99148 8166 99204 8204
rect 98924 6690 99092 6692
rect 98924 6638 98926 6690
rect 98978 6638 99092 6690
rect 98924 6636 99092 6638
rect 98924 6626 98980 6636
rect 98700 6020 98756 6030
rect 99036 6020 99092 6030
rect 98700 6018 99092 6020
rect 98700 5966 98702 6018
rect 98754 5966 99038 6018
rect 99090 5966 99092 6018
rect 98700 5964 99092 5966
rect 98700 5954 98756 5964
rect 99036 5954 99092 5964
rect 98588 5740 99092 5796
rect 98700 5348 98756 5358
rect 98700 5254 98756 5292
rect 99036 5346 99092 5740
rect 99036 5294 99038 5346
rect 99090 5294 99092 5346
rect 99036 5282 99092 5294
rect 98924 5124 98980 5134
rect 98924 5030 98980 5068
rect 99036 5012 99092 5022
rect 99036 4918 99092 4956
rect 98364 4338 98532 4340
rect 98364 4286 98366 4338
rect 98418 4286 98532 4338
rect 98364 4284 98532 4286
rect 99036 4452 99092 4462
rect 98364 4274 98420 4284
rect 97244 3502 97246 3554
rect 97298 3502 97300 3554
rect 97244 3490 97300 3502
rect 97916 3666 97972 3678
rect 97916 3614 97918 3666
rect 97970 3614 97972 3666
rect 97132 2482 97188 2492
rect 97916 800 97972 3614
rect 99036 3444 99092 4396
rect 99036 3378 99092 3388
rect 99372 3220 99428 10780
rect 99820 10724 99876 10780
rect 99708 10722 99876 10724
rect 99708 10670 99822 10722
rect 99874 10670 99876 10722
rect 99708 10668 99876 10670
rect 99708 9938 99764 10668
rect 99820 10658 99876 10668
rect 99708 9886 99710 9938
rect 99762 9886 99764 9938
rect 99708 9874 99764 9886
rect 99820 10500 99876 10510
rect 99708 9380 99764 9390
rect 99708 9042 99764 9324
rect 99708 8990 99710 9042
rect 99762 8990 99764 9042
rect 99596 8034 99652 8046
rect 99596 7982 99598 8034
rect 99650 7982 99652 8034
rect 99596 3556 99652 7982
rect 99708 7474 99764 8990
rect 99708 7422 99710 7474
rect 99762 7422 99764 7474
rect 99708 7410 99764 7422
rect 99708 6916 99764 6926
rect 99708 6690 99764 6860
rect 99708 6638 99710 6690
rect 99762 6638 99764 6690
rect 99708 6626 99764 6638
rect 99820 6578 99876 10444
rect 99820 6526 99822 6578
rect 99874 6526 99876 6578
rect 99820 6514 99876 6526
rect 99932 5012 99988 14476
rect 100268 14530 100324 15486
rect 100380 15426 100436 15596
rect 100380 15374 100382 15426
rect 100434 15374 100436 15426
rect 100380 15362 100436 15374
rect 100492 15540 100548 16716
rect 100716 16660 100772 17052
rect 100940 17042 100996 17054
rect 101388 17220 101444 17230
rect 100828 16884 100884 16894
rect 100828 16790 100884 16828
rect 101052 16882 101108 16894
rect 101052 16830 101054 16882
rect 101106 16830 101108 16882
rect 101052 16772 101108 16830
rect 101052 16706 101108 16716
rect 101388 16882 101444 17164
rect 101388 16830 101390 16882
rect 101442 16830 101444 16882
rect 100716 16604 100996 16660
rect 100828 15874 100884 15886
rect 100828 15822 100830 15874
rect 100882 15822 100884 15874
rect 100828 15652 100884 15822
rect 100828 15586 100884 15596
rect 100268 14478 100270 14530
rect 100322 14478 100324 14530
rect 100268 14466 100324 14478
rect 100044 14084 100100 14094
rect 100044 11956 100100 14028
rect 100268 13748 100324 13758
rect 100268 13654 100324 13692
rect 100156 13188 100212 13198
rect 100156 13186 100436 13188
rect 100156 13134 100158 13186
rect 100210 13134 100436 13186
rect 100156 13132 100436 13134
rect 100156 13122 100212 13132
rect 100156 12964 100212 12974
rect 100156 12850 100212 12908
rect 100156 12798 100158 12850
rect 100210 12798 100212 12850
rect 100156 12786 100212 12798
rect 100268 12852 100324 12862
rect 100268 12758 100324 12796
rect 100044 11890 100100 11900
rect 100156 12068 100212 12078
rect 100044 8258 100100 8270
rect 100044 8206 100046 8258
rect 100098 8206 100100 8258
rect 100044 7812 100100 8206
rect 100156 8036 100212 12012
rect 100268 11394 100324 11406
rect 100268 11342 100270 11394
rect 100322 11342 100324 11394
rect 100268 10612 100324 11342
rect 100380 11394 100436 13132
rect 100492 12964 100548 15484
rect 100604 15314 100660 15326
rect 100604 15262 100606 15314
rect 100658 15262 100660 15314
rect 100604 15148 100660 15262
rect 100604 15092 100772 15148
rect 100716 13074 100772 15092
rect 100716 13022 100718 13074
rect 100770 13022 100772 13074
rect 100716 13010 100772 13022
rect 100604 12964 100660 12974
rect 100492 12962 100660 12964
rect 100492 12910 100606 12962
rect 100658 12910 100660 12962
rect 100492 12908 100660 12910
rect 100604 12898 100660 12908
rect 100828 12964 100884 12974
rect 100828 12870 100884 12908
rect 100940 11620 100996 16604
rect 101052 15988 101108 15998
rect 101052 15314 101108 15932
rect 101052 15262 101054 15314
rect 101106 15262 101108 15314
rect 101052 12850 101108 15262
rect 101388 14644 101444 16830
rect 101500 16770 101556 16782
rect 101500 16718 101502 16770
rect 101554 16718 101556 16770
rect 101500 16324 101556 16718
rect 101500 16258 101556 16268
rect 101500 16100 101556 16110
rect 101612 16100 101668 17388
rect 101724 17378 101780 17388
rect 101724 17108 101780 17118
rect 101724 16994 101780 17052
rect 101724 16942 101726 16994
rect 101778 16942 101780 16994
rect 101724 16930 101780 16942
rect 101500 16098 101668 16100
rect 101500 16046 101502 16098
rect 101554 16046 101668 16098
rect 101500 16044 101668 16046
rect 101836 16100 101892 18286
rect 101948 17220 102004 18396
rect 102508 18452 102564 18462
rect 102508 18358 102564 18396
rect 104636 18452 104692 19964
rect 104972 19348 105028 19966
rect 105196 20020 105252 20030
rect 105196 19926 105252 19964
rect 105308 19348 105364 20188
rect 105420 20018 105476 21420
rect 106652 20804 106708 26012
rect 106764 25620 106820 25630
rect 106764 25618 107492 25620
rect 106764 25566 106766 25618
rect 106818 25566 107492 25618
rect 106764 25564 107492 25566
rect 106764 25554 106820 25564
rect 106988 25396 107044 25406
rect 106988 25302 107044 25340
rect 107324 25396 107380 25406
rect 107324 24946 107380 25340
rect 107324 24894 107326 24946
rect 107378 24894 107380 24946
rect 107324 24882 107380 24894
rect 106652 20748 107044 20804
rect 106652 20578 106708 20590
rect 106652 20526 106654 20578
rect 106706 20526 106708 20578
rect 105420 19966 105422 20018
rect 105474 19966 105476 20018
rect 105420 19954 105476 19966
rect 105756 20244 105812 20254
rect 105420 19348 105476 19358
rect 105308 19346 105476 19348
rect 105308 19294 105422 19346
rect 105474 19294 105476 19346
rect 105308 19292 105476 19294
rect 104972 19282 105028 19292
rect 105420 19282 105476 19292
rect 104972 19124 105028 19134
rect 104972 19030 105028 19068
rect 104636 18386 104692 18396
rect 105756 18340 105812 20188
rect 106316 20188 106596 20244
rect 105868 20132 105924 20142
rect 105868 20038 105924 20076
rect 106092 20132 106148 20142
rect 106316 20132 106372 20188
rect 106092 20130 106372 20132
rect 106092 20078 106094 20130
rect 106146 20078 106372 20130
rect 106092 20076 106372 20078
rect 106092 20066 106148 20076
rect 105980 20020 106036 20030
rect 106428 20020 106484 20030
rect 105980 19926 106036 19964
rect 106316 19964 106428 20020
rect 105868 19348 105924 19358
rect 105868 19122 105924 19292
rect 105868 19070 105870 19122
rect 105922 19070 105924 19122
rect 105868 19058 105924 19070
rect 106092 19236 106148 19246
rect 106316 19236 106372 19964
rect 106428 19926 106484 19964
rect 106540 19908 106596 20188
rect 106652 20132 106708 20526
rect 106652 20066 106708 20076
rect 106764 20130 106820 20142
rect 106764 20078 106766 20130
rect 106818 20078 106820 20130
rect 106764 19908 106820 20078
rect 106540 19852 106820 19908
rect 106428 19348 106484 19358
rect 106484 19292 106596 19348
rect 106428 19282 106484 19292
rect 106092 19234 106372 19236
rect 106092 19182 106094 19234
rect 106146 19182 106372 19234
rect 106092 19180 106372 19182
rect 106092 19124 106148 19180
rect 106092 19058 106148 19068
rect 106428 18562 106484 18574
rect 106428 18510 106430 18562
rect 106482 18510 106484 18562
rect 106092 18450 106148 18462
rect 106092 18398 106094 18450
rect 106146 18398 106148 18450
rect 106092 18340 106148 18398
rect 105756 18338 106148 18340
rect 105756 18286 105758 18338
rect 105810 18286 106148 18338
rect 105756 18284 106148 18286
rect 106204 18452 106260 18462
rect 101948 17154 102004 17164
rect 102508 17668 102564 17678
rect 102508 17108 102564 17612
rect 102508 17014 102564 17052
rect 104860 17444 104916 17454
rect 104860 16996 104916 17388
rect 105420 17108 105476 17118
rect 105420 17014 105476 17052
rect 104972 16996 105028 17006
rect 104860 16994 105028 16996
rect 104860 16942 104974 16994
rect 105026 16942 105028 16994
rect 104860 16940 105028 16942
rect 101948 16884 102004 16894
rect 103964 16884 104020 16894
rect 104860 16884 104916 16940
rect 104972 16930 105028 16940
rect 105308 16996 105364 17006
rect 105308 16902 105364 16940
rect 101948 16882 102228 16884
rect 101948 16830 101950 16882
rect 102002 16830 102228 16882
rect 101948 16828 102228 16830
rect 101948 16818 102004 16828
rect 101948 16100 102004 16110
rect 101836 16098 102004 16100
rect 101836 16046 101950 16098
rect 102002 16046 102004 16098
rect 101836 16044 102004 16046
rect 101500 16034 101556 16044
rect 101948 16034 102004 16044
rect 101724 15540 101780 15550
rect 102060 15540 102116 15550
rect 101780 15538 102116 15540
rect 101780 15486 102062 15538
rect 102114 15486 102116 15538
rect 101780 15484 102116 15486
rect 101724 15446 101780 15484
rect 102060 15474 102116 15484
rect 102172 15538 102228 16828
rect 104020 16828 104132 16884
rect 103964 16818 104020 16828
rect 102956 16772 103012 16782
rect 102844 16770 103012 16772
rect 102844 16718 102958 16770
rect 103010 16718 103012 16770
rect 102844 16716 103012 16718
rect 102172 15486 102174 15538
rect 102226 15486 102228 15538
rect 102172 15474 102228 15486
rect 102508 15988 102564 15998
rect 102508 15538 102564 15932
rect 102508 15486 102510 15538
rect 102562 15486 102564 15538
rect 102508 15474 102564 15486
rect 101612 15428 101668 15438
rect 101612 15334 101668 15372
rect 101500 15314 101556 15326
rect 101500 15262 101502 15314
rect 101554 15262 101556 15314
rect 101500 14756 101556 15262
rect 102284 15316 102340 15326
rect 102284 15222 102340 15260
rect 101500 14690 101556 14700
rect 101388 14578 101444 14588
rect 102844 14420 102900 16716
rect 102956 16706 103012 16716
rect 103852 16770 103908 16782
rect 103852 16718 103854 16770
rect 103906 16718 103908 16770
rect 102956 16212 103012 16222
rect 102956 14868 103012 16156
rect 103516 15314 103572 15326
rect 103516 15262 103518 15314
rect 103570 15262 103572 15314
rect 102956 14802 103012 14812
rect 103068 15204 103124 15214
rect 103516 15204 103572 15262
rect 103068 15202 103572 15204
rect 103068 15150 103070 15202
rect 103122 15150 103572 15202
rect 103068 15148 103572 15150
rect 103068 14532 103124 15148
rect 103516 15092 103572 15148
rect 103516 15026 103572 15036
rect 103628 14644 103684 14654
rect 103180 14532 103236 14542
rect 103068 14530 103236 14532
rect 103068 14478 103182 14530
rect 103234 14478 103236 14530
rect 103068 14476 103236 14478
rect 102844 14364 103124 14420
rect 102732 14308 102788 14318
rect 102732 14306 102900 14308
rect 102732 14254 102734 14306
rect 102786 14254 102900 14306
rect 102732 14252 102900 14254
rect 102732 14242 102788 14252
rect 101388 13860 101444 13870
rect 101052 12798 101054 12850
rect 101106 12798 101108 12850
rect 101052 12786 101108 12798
rect 101276 12852 101332 12862
rect 100940 11554 100996 11564
rect 101276 12180 101332 12796
rect 100604 11508 100660 11518
rect 100604 11414 100660 11452
rect 100380 11342 100382 11394
rect 100434 11342 100436 11394
rect 100380 11330 100436 11342
rect 101276 11394 101332 12124
rect 101276 11342 101278 11394
rect 101330 11342 101332 11394
rect 101276 11330 101332 11342
rect 100716 11284 100772 11294
rect 100492 11282 100772 11284
rect 100492 11230 100718 11282
rect 100770 11230 100772 11282
rect 100492 11228 100772 11230
rect 100380 10612 100436 10622
rect 100268 10610 100436 10612
rect 100268 10558 100382 10610
rect 100434 10558 100436 10610
rect 100268 10556 100436 10558
rect 100380 10388 100436 10556
rect 100380 10322 100436 10332
rect 100380 9268 100436 9278
rect 100380 9154 100436 9212
rect 100380 9102 100382 9154
rect 100434 9102 100436 9154
rect 100380 9090 100436 9102
rect 100268 8372 100324 8382
rect 100268 8258 100324 8316
rect 100268 8206 100270 8258
rect 100322 8206 100324 8258
rect 100268 8194 100324 8206
rect 100156 7970 100212 7980
rect 100380 8148 100436 8158
rect 100044 7756 100212 7812
rect 100156 7588 100212 7756
rect 100044 6466 100100 6478
rect 100044 6414 100046 6466
rect 100098 6414 100100 6466
rect 100044 5236 100100 6414
rect 100044 5170 100100 5180
rect 100044 5012 100100 5022
rect 99932 5010 100100 5012
rect 99932 4958 100046 5010
rect 100098 4958 100100 5010
rect 99932 4956 100100 4958
rect 99708 3556 99764 3566
rect 99596 3554 99764 3556
rect 99596 3502 99710 3554
rect 99762 3502 99764 3554
rect 99596 3500 99764 3502
rect 99708 3490 99764 3500
rect 99372 3154 99428 3164
rect 99260 924 99652 980
rect 99260 800 99316 924
rect 72716 700 73332 756
rect 73696 0 73808 800
rect 75040 0 75152 800
rect 76384 0 76496 800
rect 77728 0 77840 800
rect 79072 0 79184 800
rect 80416 0 80528 800
rect 81760 0 81872 800
rect 83104 0 83216 800
rect 84448 0 84560 800
rect 85792 0 85904 800
rect 87136 0 87248 800
rect 88480 0 88592 800
rect 89824 0 89936 800
rect 91168 0 91280 800
rect 92512 0 92624 800
rect 93856 0 93968 800
rect 95200 0 95312 800
rect 96544 0 96656 800
rect 97888 0 98000 800
rect 99232 0 99344 800
rect 99596 756 99652 924
rect 100044 756 100100 4956
rect 100156 4676 100212 7532
rect 100268 7700 100324 7710
rect 100268 6804 100324 7644
rect 100380 7586 100436 8092
rect 100380 7534 100382 7586
rect 100434 7534 100436 7586
rect 100380 7522 100436 7534
rect 100268 6710 100324 6748
rect 100492 6468 100548 11228
rect 100716 11218 100772 11228
rect 100940 11172 100996 11182
rect 100828 11170 100996 11172
rect 100828 11118 100942 11170
rect 100994 11118 100996 11170
rect 100828 11116 100996 11118
rect 100828 10836 100884 11116
rect 100940 11106 100996 11116
rect 101164 11170 101220 11182
rect 101164 11118 101166 11170
rect 101218 11118 101220 11170
rect 100604 10780 100884 10836
rect 101164 10836 101220 11118
rect 100604 10610 100660 10780
rect 101164 10770 101220 10780
rect 100604 10558 100606 10610
rect 100658 10558 100660 10610
rect 100604 10546 100660 10558
rect 100940 10610 100996 10622
rect 100940 10558 100942 10610
rect 100994 10558 100996 10610
rect 100716 10498 100772 10510
rect 100716 10446 100718 10498
rect 100770 10446 100772 10498
rect 100716 9940 100772 10446
rect 100716 9874 100772 9884
rect 100828 8820 100884 8830
rect 100828 8726 100884 8764
rect 100604 8370 100660 8382
rect 100604 8318 100606 8370
rect 100658 8318 100660 8370
rect 100604 8036 100660 8318
rect 100604 7970 100660 7980
rect 100716 8372 100772 8382
rect 100716 7362 100772 8316
rect 100716 7310 100718 7362
rect 100770 7310 100772 7362
rect 100716 7298 100772 7310
rect 100940 6580 100996 10558
rect 101164 10610 101220 10622
rect 101164 10558 101166 10610
rect 101218 10558 101220 10610
rect 101164 10164 101220 10558
rect 101164 10098 101220 10108
rect 101276 10612 101332 10622
rect 101052 9042 101108 9054
rect 101052 8990 101054 9042
rect 101106 8990 101108 9042
rect 101052 7588 101108 8990
rect 101276 9042 101332 10556
rect 101276 8990 101278 9042
rect 101330 8990 101332 9042
rect 101276 8978 101332 8990
rect 101388 8370 101444 13804
rect 102732 13748 102788 13758
rect 102732 13654 102788 13692
rect 102060 13634 102116 13646
rect 102060 13582 102062 13634
rect 102114 13582 102116 13634
rect 102060 12964 102116 13582
rect 102620 13522 102676 13534
rect 102620 13470 102622 13522
rect 102674 13470 102676 13522
rect 102508 13300 102564 13310
rect 102620 13300 102676 13470
rect 102564 13244 102676 13300
rect 102508 13234 102564 13244
rect 102396 12964 102452 12974
rect 102060 12962 102452 12964
rect 102060 12910 102398 12962
rect 102450 12910 102452 12962
rect 102060 12908 102452 12910
rect 101836 12066 101892 12078
rect 101836 12014 101838 12066
rect 101890 12014 101892 12066
rect 101836 11508 101892 12014
rect 101836 11442 101892 11452
rect 101612 11170 101668 11182
rect 101612 11118 101614 11170
rect 101666 11118 101668 11170
rect 101388 8318 101390 8370
rect 101442 8318 101444 8370
rect 101388 7700 101444 8318
rect 101388 7634 101444 7644
rect 101500 10722 101556 10734
rect 101500 10670 101502 10722
rect 101554 10670 101556 10722
rect 101500 9604 101556 10670
rect 101612 10612 101668 11118
rect 101948 11170 102004 11182
rect 101948 11118 101950 11170
rect 102002 11118 102004 11170
rect 101836 10612 101892 10622
rect 101612 10546 101668 10556
rect 101724 10610 101892 10612
rect 101724 10558 101838 10610
rect 101890 10558 101892 10610
rect 101724 10556 101892 10558
rect 101052 7522 101108 7532
rect 101500 7476 101556 9548
rect 101500 7410 101556 7420
rect 101612 8930 101668 8942
rect 101612 8878 101614 8930
rect 101666 8878 101668 8930
rect 101612 8036 101668 8878
rect 101724 8708 101780 10556
rect 101836 10546 101892 10556
rect 101836 9940 101892 9950
rect 101836 9846 101892 9884
rect 101724 8652 101892 8708
rect 101724 8260 101780 8270
rect 101724 8166 101780 8204
rect 100940 6514 100996 6524
rect 100492 6402 100548 6412
rect 100380 5796 100436 5806
rect 100380 5794 100660 5796
rect 100380 5742 100382 5794
rect 100434 5742 100660 5794
rect 100380 5740 100660 5742
rect 100380 5730 100436 5740
rect 100156 4610 100212 4620
rect 100492 5572 100548 5582
rect 100492 4452 100548 5516
rect 100604 4564 100660 5740
rect 100716 5794 100772 5806
rect 100716 5742 100718 5794
rect 100770 5742 100772 5794
rect 100716 4788 100772 5742
rect 101612 5572 101668 7980
rect 101612 5506 101668 5516
rect 101724 6018 101780 6030
rect 101724 5966 101726 6018
rect 101778 5966 101780 6018
rect 101724 5348 101780 5966
rect 101724 5282 101780 5292
rect 101836 4788 101892 8652
rect 101948 8372 102004 11118
rect 102284 11170 102340 11182
rect 102284 11118 102286 11170
rect 102338 11118 102340 11170
rect 101948 8306 102004 8316
rect 102172 10722 102228 10734
rect 102172 10670 102174 10722
rect 102226 10670 102228 10722
rect 102060 7586 102116 7598
rect 102060 7534 102062 7586
rect 102114 7534 102116 7586
rect 102060 6804 102116 7534
rect 102060 6738 102116 6748
rect 102172 5012 102228 10670
rect 102284 9154 102340 11118
rect 102396 10612 102452 12908
rect 102508 12404 102564 12414
rect 102508 11788 102564 12348
rect 102620 12292 102676 13244
rect 102844 12964 102900 14252
rect 103068 12964 103124 14364
rect 103180 13522 103236 14476
rect 103180 13470 103182 13522
rect 103234 13470 103236 13522
rect 103180 13412 103236 13470
rect 103180 13346 103236 13356
rect 103292 14532 103348 14542
rect 103292 13188 103348 14476
rect 103628 13858 103684 14588
rect 103740 14530 103796 14542
rect 103740 14478 103742 14530
rect 103794 14478 103796 14530
rect 103740 13970 103796 14478
rect 103740 13918 103742 13970
rect 103794 13918 103796 13970
rect 103740 13906 103796 13918
rect 103628 13806 103630 13858
rect 103682 13806 103684 13858
rect 103628 13794 103684 13806
rect 103292 13122 103348 13132
rect 103516 13412 103572 13422
rect 103516 13074 103572 13356
rect 103516 13022 103518 13074
rect 103570 13022 103572 13074
rect 103516 13010 103572 13022
rect 103068 12908 103460 12964
rect 102844 12404 102900 12908
rect 102844 12348 103012 12404
rect 102620 12178 102676 12236
rect 102620 12126 102622 12178
rect 102674 12126 102676 12178
rect 102620 12114 102676 12126
rect 102956 12178 103012 12348
rect 102956 12126 102958 12178
rect 103010 12126 103012 12178
rect 102956 12114 103012 12126
rect 103068 12068 103124 12078
rect 103068 12066 103348 12068
rect 103068 12014 103070 12066
rect 103122 12014 103348 12066
rect 103068 12012 103348 12014
rect 103068 12002 103124 12012
rect 102956 11844 103012 11854
rect 103292 11844 103348 12012
rect 102732 11788 102788 11798
rect 102508 11732 102676 11788
rect 102620 11338 102676 11732
rect 102508 11282 102564 11294
rect 102508 11230 102510 11282
rect 102562 11230 102564 11282
rect 102620 11286 102622 11338
rect 102674 11286 102676 11338
rect 102620 11274 102676 11286
rect 102508 11172 102564 11230
rect 102508 11106 102564 11116
rect 102396 10546 102452 10556
rect 102620 10610 102676 10622
rect 102620 10558 102622 10610
rect 102674 10558 102676 10610
rect 102620 10500 102676 10558
rect 102620 10434 102676 10444
rect 102620 9828 102676 9838
rect 102732 9828 102788 11732
rect 102844 11788 102956 11844
rect 103180 11788 103348 11844
rect 102844 11284 102900 11788
rect 102956 11778 103012 11788
rect 103068 11732 103236 11788
rect 102956 11506 103012 11518
rect 102956 11454 102958 11506
rect 103010 11454 103012 11506
rect 102956 11396 103012 11454
rect 102956 11330 103012 11340
rect 102844 11218 102900 11228
rect 102844 10948 102900 10958
rect 102844 10834 102900 10892
rect 102844 10782 102846 10834
rect 102898 10782 102900 10834
rect 102844 10770 102900 10782
rect 102844 10500 102900 10510
rect 102844 10164 102900 10444
rect 102844 10098 102900 10108
rect 103068 10164 103124 11732
rect 103404 11284 103460 12908
rect 103628 12628 103684 12638
rect 103684 12572 103796 12628
rect 103628 12562 103684 12572
rect 103628 12404 103684 12414
rect 103628 11844 103684 12348
rect 103628 11778 103684 11788
rect 103292 10948 103348 10958
rect 103068 10098 103124 10108
rect 103180 10892 103292 10948
rect 102620 9826 102788 9828
rect 102620 9774 102622 9826
rect 102674 9774 102788 9826
rect 102620 9772 102788 9774
rect 102844 9940 102900 9950
rect 102620 9762 102676 9772
rect 102284 9102 102286 9154
rect 102338 9102 102340 9154
rect 102284 9090 102340 9102
rect 102844 9156 102900 9884
rect 103068 9828 103124 9838
rect 103068 9380 103124 9772
rect 103068 9314 103124 9324
rect 102844 9062 102900 9100
rect 102508 9042 102564 9054
rect 102508 8990 102510 9042
rect 102562 8990 102564 9042
rect 102396 8932 102452 8942
rect 102396 8838 102452 8876
rect 102508 8708 102564 8990
rect 102508 8642 102564 8652
rect 102844 8820 102900 8830
rect 102508 8146 102564 8158
rect 102508 8094 102510 8146
rect 102562 8094 102564 8146
rect 102508 7812 102564 8094
rect 102396 7756 102564 7812
rect 102396 7252 102452 7756
rect 102508 7476 102564 7486
rect 102508 7382 102564 7420
rect 102396 7196 102676 7252
rect 102508 7028 102564 7038
rect 102396 6692 102452 6702
rect 102396 6598 102452 6636
rect 102508 6018 102564 6972
rect 102620 6130 102676 7196
rect 102620 6078 102622 6130
rect 102674 6078 102676 6130
rect 102620 6066 102676 6078
rect 102732 6804 102788 6814
rect 102508 5966 102510 6018
rect 102562 5966 102564 6018
rect 102508 5954 102564 5966
rect 102508 5348 102564 5358
rect 102732 5348 102788 6748
rect 102844 6580 102900 8764
rect 102956 8260 103012 8270
rect 102956 7476 103012 8204
rect 102956 6692 103012 7420
rect 103068 7700 103124 7710
rect 103068 7474 103124 7644
rect 103068 7422 103070 7474
rect 103122 7422 103124 7474
rect 103068 7410 103124 7422
rect 103068 6692 103124 6702
rect 102956 6690 103124 6692
rect 102956 6638 103070 6690
rect 103122 6638 103124 6690
rect 102956 6636 103124 6638
rect 103068 6626 103124 6636
rect 102844 6524 103012 6580
rect 102844 6244 102900 6254
rect 102844 6018 102900 6188
rect 102844 5966 102846 6018
rect 102898 5966 102900 6018
rect 102844 5954 102900 5966
rect 102956 5906 103012 6524
rect 102956 5854 102958 5906
rect 103010 5854 103012 5906
rect 102956 5842 103012 5854
rect 102508 5346 102788 5348
rect 102508 5294 102510 5346
rect 102562 5294 102788 5346
rect 102508 5292 102788 5294
rect 102844 5572 102900 5582
rect 102508 5282 102564 5292
rect 102844 5234 102900 5516
rect 102844 5182 102846 5234
rect 102898 5182 102900 5234
rect 102844 5170 102900 5182
rect 103180 5122 103236 10892
rect 103292 10882 103348 10892
rect 103404 10500 103460 11228
rect 103628 10612 103684 10622
rect 103628 10518 103684 10556
rect 103516 10500 103572 10510
rect 103404 10444 103516 10500
rect 103292 10052 103348 10062
rect 103292 9714 103348 9996
rect 103292 9662 103294 9714
rect 103346 9662 103348 9714
rect 103292 9650 103348 9662
rect 103516 9044 103572 10444
rect 103740 9826 103796 12572
rect 103852 11172 103908 16718
rect 104076 16548 104132 16828
rect 104188 16772 104244 16782
rect 104188 16770 104692 16772
rect 104188 16718 104190 16770
rect 104242 16718 104692 16770
rect 104188 16716 104692 16718
rect 104188 16706 104244 16716
rect 104076 16492 104468 16548
rect 104188 16324 104244 16334
rect 103964 16100 104020 16110
rect 103964 15148 104020 16044
rect 104188 15314 104244 16268
rect 104412 16210 104468 16492
rect 104636 16322 104692 16716
rect 104636 16270 104638 16322
rect 104690 16270 104692 16322
rect 104636 16258 104692 16270
rect 104412 16158 104414 16210
rect 104466 16158 104468 16210
rect 104412 16146 104468 16158
rect 104860 16210 104916 16828
rect 105644 16884 105700 16894
rect 105644 16790 105700 16828
rect 105756 16660 105812 18284
rect 106204 17668 106260 18396
rect 106204 17574 106260 17612
rect 106428 17668 106484 18510
rect 106428 17602 106484 17612
rect 106540 17666 106596 19292
rect 106764 17780 106820 19852
rect 106988 18452 107044 20748
rect 107212 20020 107268 20030
rect 107212 19926 107268 19964
rect 106988 18358 107044 18396
rect 106764 17714 106820 17724
rect 106540 17614 106542 17666
rect 106594 17614 106596 17666
rect 106316 17442 106372 17454
rect 106316 17390 106318 17442
rect 106370 17390 106372 17442
rect 106316 16882 106372 17390
rect 106316 16830 106318 16882
rect 106370 16830 106372 16882
rect 106316 16818 106372 16830
rect 105756 16594 105812 16604
rect 104860 16158 104862 16210
rect 104914 16158 104916 16210
rect 104860 16146 104916 16158
rect 105308 16322 105364 16334
rect 105308 16270 105310 16322
rect 105362 16270 105364 16322
rect 105308 16210 105364 16270
rect 105308 16158 105310 16210
rect 105362 16158 105364 16210
rect 104188 15262 104190 15314
rect 104242 15262 104244 15314
rect 104188 15250 104244 15262
rect 104300 15428 104356 15438
rect 104300 15148 104356 15372
rect 103964 15092 104132 15148
rect 103964 14868 104020 14878
rect 103964 14420 104020 14812
rect 103964 13858 104020 14364
rect 103964 13806 103966 13858
rect 104018 13806 104020 13858
rect 103964 13794 104020 13806
rect 103964 13524 104020 13534
rect 104076 13524 104132 15092
rect 104188 15092 104356 15148
rect 104748 15316 104804 15326
rect 104748 15148 104804 15260
rect 104748 15092 105252 15148
rect 104188 13858 104244 15092
rect 104188 13806 104190 13858
rect 104242 13806 104244 13858
rect 104188 13794 104244 13806
rect 104636 13860 104692 13870
rect 104636 13766 104692 13804
rect 105196 13858 105252 15092
rect 105196 13806 105198 13858
rect 105250 13806 105252 13858
rect 105196 13794 105252 13806
rect 104524 13746 104580 13758
rect 104524 13694 104526 13746
rect 104578 13694 104580 13746
rect 104524 13636 104580 13694
rect 104020 13468 104132 13524
rect 104188 13580 104524 13636
rect 103964 13458 104020 13468
rect 104076 12290 104132 12302
rect 104076 12238 104078 12290
rect 104130 12238 104132 12290
rect 103964 12180 104020 12190
rect 103964 12086 104020 12124
rect 103852 11106 103908 11116
rect 103964 11844 104020 11854
rect 103740 9774 103742 9826
rect 103794 9774 103796 9826
rect 103740 9762 103796 9774
rect 103852 10836 103908 10846
rect 103852 10276 103908 10780
rect 103628 9044 103684 9054
rect 103516 9042 103684 9044
rect 103516 8990 103630 9042
rect 103682 8990 103684 9042
rect 103516 8988 103684 8990
rect 103628 8978 103684 8988
rect 103740 6692 103796 6702
rect 103852 6692 103908 10220
rect 103964 9714 104020 11788
rect 104076 11396 104132 12238
rect 104076 11330 104132 11340
rect 104188 10052 104244 13580
rect 104524 13570 104580 13580
rect 104860 13746 104916 13758
rect 104860 13694 104862 13746
rect 104914 13694 104916 13746
rect 104860 12852 104916 13694
rect 105084 13634 105140 13646
rect 105084 13582 105086 13634
rect 105138 13582 105140 13634
rect 105084 13524 105140 13582
rect 105308 13524 105364 16158
rect 105644 16212 105700 16222
rect 105644 15204 105700 16156
rect 105756 15876 105812 15886
rect 105756 15782 105812 15820
rect 106316 15876 106372 15886
rect 106316 15782 106372 15820
rect 106540 15764 106596 17614
rect 106764 17556 106820 17566
rect 106764 17462 106820 17500
rect 105644 15138 105700 15148
rect 106428 15540 106484 15550
rect 105532 14756 105588 14766
rect 105532 13858 105588 14700
rect 106092 14756 106148 14766
rect 106092 14642 106148 14700
rect 106092 14590 106094 14642
rect 106146 14590 106148 14642
rect 106092 14578 106148 14590
rect 106428 14530 106484 15484
rect 106428 14478 106430 14530
rect 106482 14478 106484 14530
rect 106428 14466 106484 14478
rect 106540 14532 106596 15708
rect 106876 17332 106932 17342
rect 106652 15316 106708 15326
rect 106652 15222 106708 15260
rect 106652 14532 106708 14542
rect 106540 14530 106708 14532
rect 106540 14478 106654 14530
rect 106706 14478 106708 14530
rect 106540 14476 106708 14478
rect 106652 14466 106708 14476
rect 106652 14308 106708 14318
rect 106652 14214 106708 14252
rect 105532 13806 105534 13858
rect 105586 13806 105588 13858
rect 105532 13794 105588 13806
rect 106092 13858 106148 13870
rect 106092 13806 106094 13858
rect 106146 13806 106148 13858
rect 106092 13748 106148 13806
rect 106652 13860 106708 13870
rect 106652 13766 106708 13804
rect 105756 13692 106148 13748
rect 106204 13746 106260 13758
rect 106204 13694 106206 13746
rect 106258 13694 106260 13746
rect 105644 13524 105700 13534
rect 105084 13468 105252 13524
rect 105308 13468 105588 13524
rect 104860 12796 105140 12852
rect 104860 12628 104916 12638
rect 104860 12402 104916 12572
rect 104860 12350 104862 12402
rect 104914 12350 104916 12402
rect 104860 12338 104916 12350
rect 104300 12180 104356 12190
rect 104636 12180 104692 12190
rect 104300 12178 104468 12180
rect 104300 12126 104302 12178
rect 104354 12126 104468 12178
rect 104300 12124 104468 12126
rect 104300 12114 104356 12124
rect 104188 9986 104244 9996
rect 104300 11172 104356 11182
rect 104300 9828 104356 11116
rect 104412 10836 104468 12124
rect 104636 12178 104804 12180
rect 104636 12126 104638 12178
rect 104690 12126 104804 12178
rect 104636 12124 104804 12126
rect 104636 12114 104692 12124
rect 104412 10780 104692 10836
rect 103964 9662 103966 9714
rect 104018 9662 104020 9714
rect 103964 8372 104020 9662
rect 103964 8306 104020 8316
rect 104188 9772 104356 9828
rect 104524 10612 104580 10622
rect 104524 10388 104580 10556
rect 104524 9826 104580 10332
rect 104524 9774 104526 9826
rect 104578 9774 104580 9826
rect 103964 7700 104020 7710
rect 104188 7700 104244 9772
rect 104524 9762 104580 9774
rect 104636 9826 104692 10780
rect 104636 9774 104638 9826
rect 104690 9774 104692 9826
rect 104636 9762 104692 9774
rect 104748 9156 104804 12124
rect 105084 11508 105140 12796
rect 105196 11620 105252 13468
rect 105308 13188 105364 13198
rect 105308 12178 105364 13132
rect 105308 12126 105310 12178
rect 105362 12126 105364 12178
rect 105308 11956 105364 12126
rect 105308 11890 105364 11900
rect 105196 11554 105252 11564
rect 105084 11442 105140 11452
rect 105420 11508 105476 11518
rect 105084 11284 105140 11294
rect 104860 11282 105140 11284
rect 104860 11230 105086 11282
rect 105138 11230 105140 11282
rect 104860 11228 105140 11230
rect 104860 9938 104916 11228
rect 105084 11218 105140 11228
rect 104860 9886 104862 9938
rect 104914 9886 104916 9938
rect 104860 9874 104916 9886
rect 104972 9716 105028 9726
rect 104412 9100 104804 9156
rect 104860 9714 105028 9716
rect 104860 9662 104974 9714
rect 105026 9662 105028 9714
rect 104860 9660 105028 9662
rect 104020 7644 104244 7700
rect 104300 8036 104356 8046
rect 103964 7474 104020 7644
rect 103964 7422 103966 7474
rect 104018 7422 104020 7474
rect 103964 7410 104020 7422
rect 104300 7474 104356 7980
rect 104300 7422 104302 7474
rect 104354 7422 104356 7474
rect 104300 7410 104356 7422
rect 103740 6690 103908 6692
rect 103740 6638 103742 6690
rect 103794 6638 103908 6690
rect 103740 6636 103908 6638
rect 103740 6626 103796 6636
rect 103404 6580 103460 6590
rect 103404 6486 103460 6524
rect 103180 5070 103182 5122
rect 103234 5070 103236 5122
rect 103180 5058 103236 5070
rect 103516 6468 103572 6478
rect 103516 5122 103572 6412
rect 103516 5070 103518 5122
rect 103570 5070 103572 5122
rect 103516 5058 103572 5070
rect 103628 6466 103684 6478
rect 103628 6414 103630 6466
rect 103682 6414 103684 6466
rect 102172 4946 102228 4956
rect 103628 4900 103684 6414
rect 103740 5796 103796 5806
rect 103740 5702 103796 5740
rect 103852 5122 103908 6636
rect 103852 5070 103854 5122
rect 103906 5070 103908 5122
rect 103852 5058 103908 5070
rect 103964 7250 104020 7262
rect 103964 7198 103966 7250
rect 104018 7198 104020 7250
rect 103740 5012 103796 5022
rect 103740 4918 103796 4956
rect 103628 4834 103684 4844
rect 101948 4788 102004 4798
rect 101836 4732 101948 4788
rect 100716 4722 100772 4732
rect 101948 4722 102004 4732
rect 103740 4788 103796 4798
rect 100604 4508 100996 4564
rect 100492 4396 100772 4452
rect 100604 3444 100660 3454
rect 100604 800 100660 3388
rect 100716 3442 100772 4396
rect 100940 3554 100996 4508
rect 101276 4452 101332 4462
rect 101612 4452 101668 4462
rect 101276 4450 101668 4452
rect 101276 4398 101278 4450
rect 101330 4398 101614 4450
rect 101666 4398 101668 4450
rect 101276 4396 101668 4398
rect 101276 4386 101332 4396
rect 101612 4386 101668 4396
rect 102956 4228 103012 4238
rect 102956 4134 103012 4172
rect 103740 4226 103796 4732
rect 103740 4174 103742 4226
rect 103794 4174 103796 4226
rect 103740 4162 103796 4174
rect 103292 4004 103348 4014
rect 100940 3502 100942 3554
rect 100994 3502 100996 3554
rect 100940 3490 100996 3502
rect 101948 3666 102004 3678
rect 101948 3614 101950 3666
rect 102002 3614 102004 3666
rect 100716 3390 100718 3442
rect 100770 3390 100772 3442
rect 100716 3378 100772 3390
rect 101948 800 102004 3614
rect 103292 800 103348 3948
rect 103964 3780 104020 7198
rect 104188 6580 104244 6590
rect 104188 4788 104244 6524
rect 104300 5796 104356 5806
rect 104412 5796 104468 9100
rect 104300 5794 104468 5796
rect 104300 5742 104302 5794
rect 104354 5742 104468 5794
rect 104300 5740 104468 5742
rect 104524 8930 104580 8942
rect 104524 8878 104526 8930
rect 104578 8878 104580 8930
rect 104300 5730 104356 5740
rect 104188 4722 104244 4732
rect 104524 5124 104580 8878
rect 104636 8596 104692 8606
rect 104636 8370 104692 8540
rect 104636 8318 104638 8370
rect 104690 8318 104692 8370
rect 104636 8306 104692 8318
rect 104860 8260 104916 9660
rect 104972 9650 105028 9660
rect 105308 9604 105364 9614
rect 105308 9510 105364 9548
rect 105420 9154 105476 11452
rect 105532 11060 105588 13468
rect 105644 13430 105700 13468
rect 105644 12290 105700 12302
rect 105644 12238 105646 12290
rect 105698 12238 105700 12290
rect 105644 12180 105700 12238
rect 105644 12114 105700 12124
rect 105756 11844 105812 13692
rect 106204 13636 106260 13694
rect 106204 13570 106260 13580
rect 106092 13522 106148 13534
rect 106092 13470 106094 13522
rect 106146 13470 106148 13522
rect 105980 12404 106036 12414
rect 105980 12310 106036 12348
rect 105532 10994 105588 11004
rect 105644 11788 105812 11844
rect 105420 9102 105422 9154
rect 105474 9102 105476 9154
rect 105420 9090 105476 9102
rect 105532 9266 105588 9278
rect 105532 9214 105534 9266
rect 105586 9214 105588 9266
rect 105196 9042 105252 9054
rect 105196 8990 105198 9042
rect 105250 8990 105252 9042
rect 105196 8820 105252 8990
rect 105196 8754 105252 8764
rect 104860 8194 104916 8204
rect 105196 8372 105252 8382
rect 105196 8258 105252 8316
rect 105196 8206 105198 8258
rect 105250 8206 105252 8258
rect 105196 8194 105252 8206
rect 104860 8034 104916 8046
rect 104860 7982 104862 8034
rect 104914 7982 104916 8034
rect 104748 7362 104804 7374
rect 104748 7310 104750 7362
rect 104802 7310 104804 7362
rect 104748 5572 104804 7310
rect 104860 7028 104916 7982
rect 105084 8034 105140 8046
rect 105084 7982 105086 8034
rect 105138 7982 105140 8034
rect 105084 7588 105140 7982
rect 105532 7700 105588 9214
rect 105644 8596 105700 11788
rect 105868 11396 105924 11406
rect 105868 11394 106036 11396
rect 105868 11342 105870 11394
rect 105922 11342 106036 11394
rect 105868 11340 106036 11342
rect 105868 11330 105924 11340
rect 105980 10498 106036 11340
rect 106092 10724 106148 13470
rect 106540 12964 106596 12974
rect 106428 12740 106484 12750
rect 106316 12290 106372 12302
rect 106316 12238 106318 12290
rect 106370 12238 106372 12290
rect 106316 11620 106372 12238
rect 106092 10658 106148 10668
rect 106204 11284 106260 11294
rect 106204 10612 106260 11228
rect 106316 10836 106372 11564
rect 106428 11732 106484 12684
rect 106428 11394 106484 11676
rect 106428 11342 106430 11394
rect 106482 11342 106484 11394
rect 106428 11330 106484 11342
rect 106316 10770 106372 10780
rect 106204 10546 106260 10556
rect 105980 10446 105982 10498
rect 106034 10446 106036 10498
rect 105868 9828 105924 9838
rect 105868 9734 105924 9772
rect 105756 9156 105812 9166
rect 105756 9062 105812 9100
rect 105980 9044 106036 10446
rect 105980 8820 106036 8988
rect 105644 8530 105700 8540
rect 105756 8764 106036 8820
rect 106092 10164 106148 10174
rect 105084 7522 105140 7532
rect 105420 7644 105588 7700
rect 104860 6962 104916 6972
rect 104860 6804 104916 6814
rect 104860 6710 104916 6748
rect 105420 6692 105476 7644
rect 105532 7476 105588 7486
rect 105756 7476 105812 8764
rect 106092 8708 106148 10108
rect 106540 9940 106596 12908
rect 106540 9874 106596 9884
rect 106652 12290 106708 12302
rect 106652 12238 106654 12290
rect 106706 12238 106708 12290
rect 106652 10724 106708 12238
rect 106876 10948 106932 17276
rect 106988 15876 107044 15886
rect 107044 15820 107156 15876
rect 106988 15782 107044 15820
rect 106988 15428 107044 15438
rect 106988 14530 107044 15372
rect 107100 15204 107156 15820
rect 107436 15540 107492 25564
rect 107548 25508 107604 26126
rect 108668 25620 108724 28588
rect 108220 25618 108724 25620
rect 108220 25566 108670 25618
rect 108722 25566 108724 25618
rect 108220 25564 108724 25566
rect 107660 25508 107716 25546
rect 107548 25452 107660 25508
rect 107660 25442 107716 25452
rect 108220 25394 108276 25564
rect 108668 25554 108724 25564
rect 108220 25342 108222 25394
rect 108274 25342 108276 25394
rect 108220 25330 108276 25342
rect 110012 25396 110068 56140
rect 112364 55972 112420 56588
rect 116060 56308 116116 59200
rect 116060 56242 116116 56252
rect 117292 56308 117348 56318
rect 117292 56214 117348 56252
rect 119868 56308 119924 59200
rect 119868 56242 119924 56252
rect 121100 56308 121156 56318
rect 121100 56214 121156 56252
rect 112476 56196 112532 56206
rect 112476 56102 112532 56140
rect 115052 56196 115108 56206
rect 112700 56082 112756 56094
rect 112700 56030 112702 56082
rect 112754 56030 112756 56082
rect 112700 55972 112756 56030
rect 112364 55916 112756 55972
rect 112364 55468 112420 55916
rect 112252 55412 112420 55468
rect 112252 55410 112308 55412
rect 112252 55358 112254 55410
rect 112306 55358 112308 55410
rect 112252 55346 112308 55358
rect 111996 54908 112260 54918
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 111996 54842 112260 54852
rect 111996 53340 112260 53350
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 111996 53274 112260 53284
rect 111996 51772 112260 51782
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 111996 51706 112260 51716
rect 111996 50204 112260 50214
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 111996 50138 112260 50148
rect 111996 48636 112260 48646
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 111996 48570 112260 48580
rect 111996 47068 112260 47078
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 111996 47002 112260 47012
rect 111996 45500 112260 45510
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 111996 45434 112260 45444
rect 111996 43932 112260 43942
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 111996 43866 112260 43876
rect 111996 42364 112260 42374
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 111996 42298 112260 42308
rect 111996 40796 112260 40806
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 111996 40730 112260 40740
rect 111996 39228 112260 39238
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 111996 39162 112260 39172
rect 111996 37660 112260 37670
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 111996 37594 112260 37604
rect 111996 36092 112260 36102
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 111996 36026 112260 36036
rect 111996 34524 112260 34534
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 111996 34458 112260 34468
rect 111996 32956 112260 32966
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 111996 32890 112260 32900
rect 111996 31388 112260 31398
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 111996 31322 112260 31332
rect 111996 29820 112260 29830
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 111996 29754 112260 29764
rect 115052 28644 115108 56140
rect 116284 56082 116340 56094
rect 116284 56030 116286 56082
rect 116338 56030 116340 56082
rect 116284 55468 116340 56030
rect 120092 56082 120148 56094
rect 120092 56030 120094 56082
rect 120146 56030 120148 56082
rect 120092 55468 120148 56030
rect 116060 55412 116340 55468
rect 119756 55412 120148 55468
rect 123676 55972 123732 59200
rect 127484 56308 127540 59200
rect 127484 56242 127540 56252
rect 128716 56308 128772 56318
rect 128716 56214 128772 56252
rect 131292 56308 131348 59200
rect 131292 56242 131348 56252
rect 132524 56308 132580 56318
rect 132524 56214 132580 56252
rect 135100 56308 135156 59200
rect 135324 56308 135380 56318
rect 135100 56306 135380 56308
rect 135100 56254 135326 56306
rect 135378 56254 135380 56306
rect 135100 56252 135380 56254
rect 123900 56196 123956 56206
rect 123900 56102 123956 56140
rect 124124 56082 124180 56094
rect 124124 56030 124126 56082
rect 124178 56030 124180 56082
rect 124124 55972 124180 56030
rect 127708 56082 127764 56094
rect 127708 56030 127710 56082
rect 127762 56030 127764 56082
rect 123676 55916 124180 55972
rect 125132 55972 125188 55982
rect 115724 55300 115780 55310
rect 115948 55300 116004 55310
rect 115780 55298 116004 55300
rect 115780 55246 115950 55298
rect 116002 55246 116004 55298
rect 115780 55244 116004 55246
rect 115724 55206 115780 55244
rect 115948 55234 116004 55244
rect 116060 54738 116116 55412
rect 116060 54686 116062 54738
rect 116114 54686 116116 54738
rect 116060 54674 116116 54686
rect 116508 55186 116564 55198
rect 116508 55134 116510 55186
rect 116562 55134 116564 55186
rect 115836 54514 115892 54526
rect 115836 54462 115838 54514
rect 115890 54462 115892 54514
rect 115836 54404 115892 54462
rect 116508 54404 116564 55134
rect 119756 55074 119812 55412
rect 123676 55410 123732 55916
rect 123676 55358 123678 55410
rect 123730 55358 123732 55410
rect 123676 55346 123732 55358
rect 119756 55022 119758 55074
rect 119810 55022 119812 55074
rect 116620 54404 116676 54414
rect 116508 54348 116620 54404
rect 115836 54338 115892 54348
rect 116620 54310 116676 54348
rect 115052 28578 115108 28588
rect 111996 28252 112260 28262
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 111996 28186 112260 28196
rect 111996 26684 112260 26694
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 111996 26618 112260 26628
rect 110012 25330 110068 25340
rect 107884 25282 107940 25294
rect 107884 25230 107886 25282
rect 107938 25230 107940 25282
rect 107772 20132 107828 20142
rect 107772 20038 107828 20076
rect 107884 20020 107940 25230
rect 111996 25116 112260 25126
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 111996 25050 112260 25060
rect 111996 23548 112260 23558
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 111996 23482 112260 23492
rect 108892 22932 108948 22942
rect 108668 21586 108724 21598
rect 108668 21534 108670 21586
rect 108722 21534 108724 21586
rect 108332 21476 108388 21486
rect 108668 21476 108724 21534
rect 108332 21474 108724 21476
rect 108332 21422 108334 21474
rect 108386 21422 108724 21474
rect 108332 21420 108724 21422
rect 108220 20802 108276 20814
rect 108220 20750 108222 20802
rect 108274 20750 108276 20802
rect 107996 20580 108052 20590
rect 108220 20580 108276 20750
rect 108052 20524 108276 20580
rect 107996 20486 108052 20524
rect 108220 20020 108276 20030
rect 108332 20020 108388 21420
rect 108556 20132 108612 20142
rect 108556 20038 108612 20076
rect 107884 19964 108164 20020
rect 107884 19796 107940 19806
rect 107884 19702 107940 19740
rect 107884 19124 107940 19134
rect 107884 19030 107940 19068
rect 107548 17780 107604 17790
rect 107548 17666 107604 17724
rect 107548 17614 107550 17666
rect 107602 17614 107604 17666
rect 107548 16884 107604 17614
rect 107996 17668 108052 17678
rect 107660 17556 107716 17566
rect 107660 17462 107716 17500
rect 107996 17554 108052 17612
rect 107996 17502 107998 17554
rect 108050 17502 108052 17554
rect 107996 17490 108052 17502
rect 107772 17442 107828 17454
rect 107772 17390 107774 17442
rect 107826 17390 107828 17442
rect 107548 16828 107716 16884
rect 107660 16100 107716 16828
rect 107772 16772 107828 17390
rect 107772 16706 107828 16716
rect 107884 16100 107940 16110
rect 107660 16098 107940 16100
rect 107660 16046 107886 16098
rect 107938 16046 107940 16098
rect 107660 16044 107940 16046
rect 108108 16100 108164 19964
rect 108276 19964 108388 20020
rect 108780 20018 108836 20030
rect 108780 19966 108782 20018
rect 108834 19966 108836 20018
rect 108220 19926 108276 19964
rect 108780 19908 108836 19966
rect 108668 19852 108780 19908
rect 108668 19346 108724 19852
rect 108780 19842 108836 19852
rect 108668 19294 108670 19346
rect 108722 19294 108724 19346
rect 108668 19282 108724 19294
rect 108668 18452 108724 18462
rect 108892 18452 108948 22876
rect 111996 21980 112260 21990
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 111996 21914 112260 21924
rect 109004 21700 109060 21710
rect 109004 21698 109172 21700
rect 109004 21646 109006 21698
rect 109058 21646 109172 21698
rect 109004 21644 109172 21646
rect 109004 21634 109060 21644
rect 109004 20802 109060 20814
rect 109004 20750 109006 20802
rect 109058 20750 109060 20802
rect 109004 20242 109060 20750
rect 109004 20190 109006 20242
rect 109058 20190 109060 20242
rect 109004 20178 109060 20190
rect 109116 20018 109172 21644
rect 110796 21588 110852 21598
rect 109452 20132 109956 20188
rect 109452 20130 109508 20132
rect 109452 20078 109454 20130
rect 109506 20078 109508 20130
rect 109452 20066 109508 20078
rect 109900 20130 109956 20132
rect 109900 20078 109902 20130
rect 109954 20078 109956 20130
rect 109900 20066 109956 20078
rect 110236 20130 110292 20142
rect 110236 20078 110238 20130
rect 110290 20078 110292 20130
rect 109116 19966 109118 20018
rect 109170 19966 109172 20018
rect 109116 18564 109172 19966
rect 109788 20020 109844 20030
rect 109788 19684 109844 19964
rect 110012 20020 110068 20030
rect 110012 19926 110068 19964
rect 109452 19236 109508 19246
rect 109788 19236 109844 19628
rect 110236 19908 110292 20078
rect 110236 19236 110292 19852
rect 110796 19796 110852 21532
rect 111692 20802 111748 20814
rect 111692 20750 111694 20802
rect 111746 20750 111748 20802
rect 111356 20578 111412 20590
rect 111692 20580 111748 20750
rect 111356 20526 111358 20578
rect 111410 20526 111412 20578
rect 111356 20020 111412 20526
rect 111580 20524 111692 20580
rect 111580 20242 111636 20524
rect 111692 20514 111748 20524
rect 112364 20802 112420 20814
rect 112364 20750 112366 20802
rect 112418 20750 112420 20802
rect 111996 20412 112260 20422
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 111996 20346 112260 20356
rect 111580 20190 111582 20242
rect 111634 20190 111636 20242
rect 111580 20178 111636 20190
rect 112364 20188 112420 20750
rect 114828 20578 114884 20590
rect 114828 20526 114830 20578
rect 114882 20526 114884 20578
rect 114828 20188 114884 20526
rect 112364 20132 112532 20188
rect 112476 20066 112532 20076
rect 113372 20132 113428 20142
rect 114828 20132 114996 20188
rect 113372 20038 113428 20076
rect 110908 19908 110964 19918
rect 110908 19814 110964 19852
rect 110796 19730 110852 19740
rect 111356 19348 111412 19964
rect 111916 20018 111972 20030
rect 111916 19966 111918 20018
rect 111970 19966 111972 20018
rect 111916 19908 111972 19966
rect 112364 20020 112420 20030
rect 112364 19926 112420 19964
rect 112588 20018 112644 20030
rect 112588 19966 112590 20018
rect 112642 19966 112644 20018
rect 112476 19908 112532 19918
rect 111972 19852 112308 19908
rect 111916 19842 111972 19852
rect 112252 19348 112308 19852
rect 112476 19814 112532 19852
rect 112588 19684 112644 19966
rect 112924 20018 112980 20030
rect 112924 19966 112926 20018
rect 112978 19966 112980 20018
rect 112924 19908 112980 19966
rect 112924 19842 112980 19852
rect 113260 20018 113316 20030
rect 113260 19966 113262 20018
rect 113314 19966 113316 20018
rect 112644 19628 112756 19684
rect 112588 19618 112644 19628
rect 112364 19348 112420 19358
rect 112252 19346 112420 19348
rect 112252 19294 112366 19346
rect 112418 19294 112420 19346
rect 112252 19292 112420 19294
rect 111356 19282 111412 19292
rect 109788 19180 109956 19236
rect 109452 19142 109508 19180
rect 109116 18508 109284 18564
rect 108668 18450 108948 18452
rect 108668 18398 108670 18450
rect 108722 18398 108894 18450
rect 108946 18398 108948 18450
rect 108668 18396 108948 18398
rect 109228 18452 109284 18508
rect 109340 18452 109396 18462
rect 109228 18450 109396 18452
rect 109228 18398 109342 18450
rect 109394 18398 109396 18450
rect 109228 18396 109396 18398
rect 108668 18386 108724 18396
rect 108892 18386 108948 18396
rect 109116 18340 109172 18350
rect 109116 18246 109172 18284
rect 109340 18228 109396 18396
rect 109564 18452 109620 18462
rect 109564 18450 109732 18452
rect 109564 18398 109566 18450
rect 109618 18398 109732 18450
rect 109564 18396 109732 18398
rect 109564 18386 109620 18396
rect 109340 18162 109396 18172
rect 109116 17666 109172 17678
rect 109116 17614 109118 17666
rect 109170 17614 109172 17666
rect 108892 17444 108948 17454
rect 109116 17444 109172 17614
rect 108892 17442 109172 17444
rect 108892 17390 108894 17442
rect 108946 17390 109172 17442
rect 108892 17388 109172 17390
rect 109228 17668 109284 17678
rect 108780 16882 108836 16894
rect 108780 16830 108782 16882
rect 108834 16830 108836 16882
rect 108780 16772 108836 16830
rect 108892 16884 108948 17388
rect 108892 16818 108948 16828
rect 109228 16882 109284 17612
rect 109228 16830 109230 16882
rect 109282 16830 109284 16882
rect 108780 16706 108836 16716
rect 108556 16156 108724 16212
rect 108108 16044 108388 16100
rect 107772 15764 107828 15774
rect 107548 15540 107604 15550
rect 107492 15538 107604 15540
rect 107492 15486 107550 15538
rect 107602 15486 107604 15538
rect 107492 15484 107604 15486
rect 107436 15446 107492 15484
rect 107548 15474 107604 15484
rect 107100 15138 107156 15148
rect 107660 15204 107716 15214
rect 106988 14478 106990 14530
rect 107042 14478 107044 14530
rect 106988 14466 107044 14478
rect 107660 14530 107716 15148
rect 107772 15148 107828 15708
rect 107884 15540 107940 16044
rect 108332 15988 108388 16044
rect 108556 16098 108612 16156
rect 108556 16046 108558 16098
rect 108610 16046 108612 16098
rect 108556 16034 108612 16046
rect 108668 16100 108724 16156
rect 109228 16100 109284 16830
rect 109564 17444 109620 17454
rect 109564 16884 109620 17388
rect 109676 17108 109732 18396
rect 109788 18340 109844 18350
rect 109788 17666 109844 18284
rect 109788 17614 109790 17666
rect 109842 17614 109844 17666
rect 109788 17602 109844 17614
rect 109788 17108 109844 17118
rect 109676 17106 109844 17108
rect 109676 17054 109790 17106
rect 109842 17054 109844 17106
rect 109676 17052 109844 17054
rect 109788 17042 109844 17052
rect 109900 17106 109956 19180
rect 110236 19170 110292 19180
rect 112364 19236 112420 19292
rect 112364 19170 112420 19180
rect 112700 19234 112756 19628
rect 112700 19182 112702 19234
rect 112754 19182 112756 19234
rect 112700 19170 112756 19182
rect 113148 19236 113204 19246
rect 113148 19122 113204 19180
rect 113148 19070 113150 19122
rect 113202 19070 113204 19122
rect 113148 19058 113204 19070
rect 112812 19010 112868 19022
rect 112812 18958 112814 19010
rect 112866 18958 112868 19010
rect 111996 18844 112260 18854
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 111996 18778 112260 18788
rect 112812 18676 112868 18958
rect 112364 18620 112868 18676
rect 112924 19010 112980 19022
rect 112924 18958 112926 19010
rect 112978 18958 112980 19010
rect 111020 18452 111076 18462
rect 111020 18338 111076 18396
rect 111692 18452 111748 18462
rect 111692 18358 111748 18396
rect 112140 18452 112196 18462
rect 111020 18286 111022 18338
rect 111074 18286 111076 18338
rect 111020 17892 111076 18286
rect 111916 18340 111972 18350
rect 111916 18246 111972 18284
rect 112140 18228 112196 18396
rect 112364 18450 112420 18620
rect 112364 18398 112366 18450
rect 112418 18398 112420 18450
rect 112364 18386 112420 18398
rect 112140 18162 112196 18172
rect 112812 18340 112868 18350
rect 111020 17826 111076 17836
rect 112252 17444 112308 17482
rect 112308 17388 112420 17444
rect 112252 17378 112308 17388
rect 111996 17276 112260 17286
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 111996 17210 112260 17220
rect 109900 17054 109902 17106
rect 109954 17054 109956 17106
rect 109900 17042 109956 17054
rect 109676 16884 109732 16894
rect 109564 16882 109732 16884
rect 109564 16830 109678 16882
rect 109730 16830 109732 16882
rect 109564 16828 109732 16830
rect 109676 16818 109732 16828
rect 111916 16884 111972 16894
rect 112140 16884 112196 16894
rect 111972 16882 112196 16884
rect 111972 16830 112142 16882
rect 112194 16830 112196 16882
rect 111972 16828 112196 16830
rect 111916 16790 111972 16828
rect 112140 16818 112196 16828
rect 108668 16044 109284 16100
rect 108332 15932 108500 15988
rect 107884 15474 107940 15484
rect 107996 15874 108052 15886
rect 107996 15822 107998 15874
rect 108050 15822 108052 15874
rect 107996 15314 108052 15822
rect 108108 15874 108164 15886
rect 108108 15822 108110 15874
rect 108162 15822 108164 15874
rect 108108 15764 108164 15822
rect 108444 15876 108500 15932
rect 108892 15876 108948 15886
rect 108444 15874 108948 15876
rect 108444 15822 108894 15874
rect 108946 15822 108948 15874
rect 108444 15820 108948 15822
rect 108108 15708 108388 15764
rect 108220 15538 108276 15550
rect 108220 15486 108222 15538
rect 108274 15486 108276 15538
rect 107996 15262 107998 15314
rect 108050 15262 108052 15314
rect 107996 15250 108052 15262
rect 108108 15314 108164 15326
rect 108108 15262 108110 15314
rect 108162 15262 108164 15314
rect 108108 15148 108164 15262
rect 107772 15092 108164 15148
rect 107660 14478 107662 14530
rect 107714 14478 107716 14530
rect 107212 14420 107268 14430
rect 107212 13970 107268 14364
rect 107212 13918 107214 13970
rect 107266 13918 107268 13970
rect 107212 13906 107268 13918
rect 107660 13746 107716 14478
rect 108108 14530 108164 14542
rect 108108 14478 108110 14530
rect 108162 14478 108164 14530
rect 108108 14308 108164 14478
rect 108108 14242 108164 14252
rect 107660 13694 107662 13746
rect 107714 13694 107716 13746
rect 107548 13636 107604 13646
rect 107548 12962 107604 13580
rect 107660 13076 107716 13694
rect 108220 13746 108276 15486
rect 108332 14084 108388 15708
rect 108444 15426 108500 15820
rect 108892 15810 108948 15820
rect 108780 15540 108836 15550
rect 108780 15446 108836 15484
rect 109228 15538 109284 16044
rect 110236 16772 110292 16782
rect 110236 16098 110292 16716
rect 110236 16046 110238 16098
rect 110290 16046 110292 16098
rect 110236 16034 110292 16046
rect 112364 16098 112420 17388
rect 112364 16046 112366 16098
rect 112418 16046 112420 16098
rect 112364 16034 112420 16046
rect 112588 17108 112644 17118
rect 109228 15486 109230 15538
rect 109282 15486 109284 15538
rect 109228 15474 109284 15486
rect 110348 15874 110404 15886
rect 110348 15822 110350 15874
rect 110402 15822 110404 15874
rect 108444 15374 108446 15426
rect 108498 15374 108500 15426
rect 108444 14420 108500 15374
rect 108892 15428 108948 15438
rect 108892 15334 108948 15372
rect 109004 15314 109060 15326
rect 109004 15262 109006 15314
rect 109058 15262 109060 15314
rect 109004 14644 109060 15262
rect 109788 15204 109844 15214
rect 109788 15110 109844 15148
rect 109004 14578 109060 14588
rect 108444 14354 108500 14364
rect 108332 14018 108388 14028
rect 108220 13694 108222 13746
rect 108274 13694 108276 13746
rect 108220 13682 108276 13694
rect 109004 13636 109060 13646
rect 107660 13010 107716 13020
rect 108108 13524 108164 13534
rect 107548 12910 107550 12962
rect 107602 12910 107604 12962
rect 107548 12898 107604 12910
rect 106988 12740 107044 12750
rect 106988 12290 107044 12684
rect 107660 12740 107716 12750
rect 107660 12404 107716 12684
rect 107884 12740 107940 12750
rect 107884 12646 107940 12684
rect 107548 12348 107716 12404
rect 108108 12404 108164 13468
rect 108668 13300 108724 13310
rect 108220 13076 108276 13086
rect 108220 12982 108276 13020
rect 108668 13074 108724 13244
rect 108668 13022 108670 13074
rect 108722 13022 108724 13074
rect 108668 13010 108724 13022
rect 108892 13188 108948 13198
rect 108668 12404 108724 12414
rect 108108 12348 108276 12404
rect 106988 12238 106990 12290
rect 107042 12238 107044 12290
rect 106988 12226 107044 12238
rect 107436 12290 107492 12302
rect 107436 12238 107438 12290
rect 107490 12238 107492 12290
rect 107324 12180 107380 12190
rect 107324 12086 107380 12124
rect 106988 11172 107044 11182
rect 106988 11170 107268 11172
rect 106988 11118 106990 11170
rect 107042 11118 107268 11170
rect 106988 11116 107268 11118
rect 106988 11106 107044 11116
rect 106876 10892 107044 10948
rect 106428 9716 106484 9726
rect 106652 9716 106708 10668
rect 106764 9828 106820 9838
rect 106764 9826 106932 9828
rect 106764 9774 106766 9826
rect 106818 9774 106932 9826
rect 106764 9772 106932 9774
rect 106764 9762 106820 9772
rect 106428 9714 106708 9716
rect 106428 9662 106430 9714
rect 106482 9662 106708 9714
rect 106428 9660 106708 9662
rect 106204 9268 106260 9278
rect 106204 8930 106260 9212
rect 106204 8878 106206 8930
rect 106258 8878 106260 8930
rect 106204 8866 106260 8878
rect 106428 8820 106484 9660
rect 106428 8754 106484 8764
rect 106764 9602 106820 9614
rect 106764 9550 106766 9602
rect 106818 9550 106820 9602
rect 105980 8652 106148 8708
rect 105980 8260 106036 8652
rect 106764 8484 106820 9550
rect 106316 8428 106820 8484
rect 106204 8372 106260 8382
rect 106092 8260 106148 8270
rect 105980 8258 106148 8260
rect 105980 8206 106094 8258
rect 106146 8206 106148 8258
rect 105980 8204 106148 8206
rect 106092 8194 106148 8204
rect 105588 7420 105812 7476
rect 105532 7382 105588 7420
rect 105756 6916 105812 7420
rect 105756 6850 105812 6860
rect 106204 7028 106260 8316
rect 106316 7586 106372 8428
rect 106540 8260 106596 8270
rect 106540 8258 106708 8260
rect 106540 8206 106542 8258
rect 106594 8206 106708 8258
rect 106540 8204 106708 8206
rect 106540 8194 106596 8204
rect 106316 7534 106318 7586
rect 106370 7534 106372 7586
rect 106316 7522 106372 7534
rect 106428 8034 106484 8046
rect 106428 7982 106430 8034
rect 106482 7982 106484 8034
rect 105420 6626 105476 6636
rect 106092 6580 106148 6590
rect 106204 6580 106260 6972
rect 106092 6578 106260 6580
rect 106092 6526 106094 6578
rect 106146 6526 106260 6578
rect 106092 6524 106260 6526
rect 106092 6514 106148 6524
rect 104748 5506 104804 5516
rect 104860 6020 104916 6030
rect 103964 3714 104020 3724
rect 103964 3556 104020 3566
rect 103964 3462 104020 3500
rect 104524 3388 104580 5068
rect 104636 5010 104692 5022
rect 104636 4958 104638 5010
rect 104690 4958 104692 5010
rect 104636 4004 104692 4958
rect 104636 3938 104692 3948
rect 104748 4450 104804 4462
rect 104748 4398 104750 4450
rect 104802 4398 104804 4450
rect 104748 3666 104804 4398
rect 104748 3614 104750 3666
rect 104802 3614 104804 3666
rect 104748 3602 104804 3614
rect 104860 3388 104916 5964
rect 105420 6020 105476 6030
rect 105756 6020 105812 6030
rect 105420 6018 105812 6020
rect 105420 5966 105422 6018
rect 105474 5966 105758 6018
rect 105810 5966 105812 6018
rect 105420 5964 105812 5966
rect 105420 5954 105476 5964
rect 105756 5954 105812 5964
rect 104412 3332 104580 3388
rect 104636 3332 104916 3388
rect 105644 4676 105700 4686
rect 105644 4338 105700 4620
rect 105868 4564 105924 4574
rect 105868 4470 105924 4508
rect 105644 4286 105646 4338
rect 105698 4286 105700 4338
rect 104412 2884 104468 3332
rect 104412 2818 104468 2828
rect 104636 800 104692 3332
rect 105644 2772 105700 4286
rect 106428 4338 106484 7982
rect 106540 6916 106596 6926
rect 106540 6466 106596 6860
rect 106540 6414 106542 6466
rect 106594 6414 106596 6466
rect 106540 6402 106596 6414
rect 106652 6690 106708 8204
rect 106652 6638 106654 6690
rect 106706 6638 106708 6690
rect 106652 6468 106708 6638
rect 106652 6402 106708 6412
rect 106876 6132 106932 9772
rect 106988 8036 107044 10892
rect 107100 10052 107156 10062
rect 107100 9826 107156 9996
rect 107100 9774 107102 9826
rect 107154 9774 107156 9826
rect 107100 9762 107156 9774
rect 106988 7970 107044 7980
rect 107212 6580 107268 11116
rect 107436 9268 107492 12238
rect 107548 11956 107604 12348
rect 107996 12292 108052 12302
rect 107996 12198 108052 12236
rect 107660 12180 107716 12190
rect 107660 12178 107828 12180
rect 107660 12126 107662 12178
rect 107714 12126 107828 12178
rect 107660 12124 107828 12126
rect 107660 12114 107716 12124
rect 107548 11900 107716 11956
rect 107548 11284 107604 11294
rect 107548 11190 107604 11228
rect 107660 10052 107716 11900
rect 107772 11394 107828 12124
rect 108108 12178 108164 12190
rect 108108 12126 108110 12178
rect 108162 12126 108164 12178
rect 107996 11956 108052 11966
rect 107772 11342 107774 11394
rect 107826 11342 107828 11394
rect 107772 11330 107828 11342
rect 107884 11954 108052 11956
rect 107884 11902 107998 11954
rect 108050 11902 108052 11954
rect 107884 11900 108052 11902
rect 107436 9202 107492 9212
rect 107548 9996 107716 10052
rect 107212 6514 107268 6524
rect 107436 8484 107492 8494
rect 107436 6468 107492 8428
rect 107436 6402 107492 6412
rect 107548 6802 107604 9996
rect 107660 9826 107716 9838
rect 107660 9774 107662 9826
rect 107714 9774 107716 9826
rect 107660 8372 107716 9774
rect 107884 9156 107940 11900
rect 107996 11890 108052 11900
rect 108108 11956 108164 12126
rect 108108 11890 108164 11900
rect 108108 11282 108164 11294
rect 108108 11230 108110 11282
rect 108162 11230 108164 11282
rect 107996 11170 108052 11182
rect 107996 11118 107998 11170
rect 108050 11118 108052 11170
rect 107996 10164 108052 11118
rect 107996 10098 108052 10108
rect 107884 9090 107940 9100
rect 107996 9828 108052 9838
rect 107884 8484 107940 8494
rect 107996 8484 108052 9772
rect 107940 8428 108052 8484
rect 107884 8418 107940 8428
rect 107660 8306 107716 8316
rect 107660 8036 107716 8046
rect 107660 7942 107716 7980
rect 107884 8036 107940 8046
rect 107884 7942 107940 7980
rect 107548 6750 107550 6802
rect 107602 6750 107604 6802
rect 106876 6066 106932 6076
rect 106764 5012 106820 5022
rect 106764 4918 106820 4956
rect 106428 4286 106430 4338
rect 106482 4286 106484 4338
rect 106428 4274 106484 4286
rect 107324 4900 107380 4910
rect 105644 2706 105700 2716
rect 105980 4116 106036 4126
rect 105980 800 106036 4060
rect 107212 4116 107268 4126
rect 107212 4022 107268 4060
rect 106876 3444 106932 3482
rect 106876 2884 106932 3388
rect 107324 3442 107380 4844
rect 107324 3390 107326 3442
rect 107378 3390 107380 3442
rect 107324 3378 107380 3390
rect 107436 4788 107492 4798
rect 107548 4788 107604 6750
rect 107884 6020 107940 6030
rect 107884 5926 107940 5964
rect 107660 5012 107716 5022
rect 107660 4918 107716 4956
rect 107548 4732 107716 4788
rect 107436 3220 107492 4732
rect 107548 4228 107604 4238
rect 107548 3554 107604 4172
rect 107548 3502 107550 3554
rect 107602 3502 107604 3554
rect 107548 3490 107604 3502
rect 107548 3332 107604 3342
rect 107660 3332 107716 4732
rect 108108 4340 108164 11230
rect 108220 9826 108276 12348
rect 108556 12292 108612 12302
rect 108556 12198 108612 12236
rect 108444 12178 108500 12190
rect 108444 12126 108446 12178
rect 108498 12126 108500 12178
rect 108444 11956 108500 12126
rect 108444 11890 108500 11900
rect 108556 12068 108612 12078
rect 108556 11954 108612 12012
rect 108556 11902 108558 11954
rect 108610 11902 108612 11954
rect 108556 11890 108612 11902
rect 108668 11844 108724 12348
rect 108556 11732 108724 11788
rect 108556 11394 108612 11732
rect 108556 11342 108558 11394
rect 108610 11342 108612 11394
rect 108220 9774 108222 9826
rect 108274 9774 108276 9826
rect 108220 9762 108276 9774
rect 108332 10164 108388 10174
rect 108332 9154 108388 10108
rect 108332 9102 108334 9154
rect 108386 9102 108388 9154
rect 108332 9090 108388 9102
rect 108556 8372 108612 11342
rect 108780 11284 108836 11294
rect 108780 10612 108836 11228
rect 108780 10546 108836 10556
rect 108892 9828 108948 13132
rect 108780 9772 108948 9828
rect 108780 8596 108836 9772
rect 109004 9716 109060 13580
rect 110348 13524 110404 15822
rect 112476 15876 112532 15886
rect 112476 15782 112532 15820
rect 111996 15708 112260 15718
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 111996 15642 112260 15652
rect 112588 14980 112644 17052
rect 112812 16882 112868 18284
rect 112924 17108 112980 18958
rect 113260 18452 113316 19966
rect 113484 20020 113540 20030
rect 113932 20020 113988 20030
rect 113484 20018 113988 20020
rect 113484 19966 113486 20018
rect 113538 19966 113934 20018
rect 113986 19966 113988 20018
rect 113484 19964 113988 19966
rect 113484 19796 113540 19964
rect 113932 19954 113988 19964
rect 113484 19730 113540 19740
rect 114940 19908 114996 20132
rect 114044 19348 114100 19358
rect 114044 19254 114100 19292
rect 114156 19012 114212 19022
rect 114156 18918 114212 18956
rect 114940 18562 114996 19852
rect 114940 18510 114942 18562
rect 114994 18510 114996 18562
rect 114940 18498 114996 18510
rect 113260 18386 113316 18396
rect 117964 18340 118020 18350
rect 115052 18228 115108 18238
rect 115052 18134 115108 18172
rect 112924 17042 112980 17052
rect 115276 17108 115332 17118
rect 115332 17052 115668 17108
rect 115276 17014 115332 17052
rect 115612 16994 115668 17052
rect 115612 16942 115614 16994
rect 115666 16942 115668 16994
rect 115612 16930 115668 16942
rect 112812 16830 112814 16882
rect 112866 16830 112868 16882
rect 112812 16818 112868 16830
rect 115724 16658 115780 16670
rect 115724 16606 115726 16658
rect 115778 16606 115780 16658
rect 114940 15876 114996 15886
rect 114940 15148 114996 15820
rect 115724 15148 115780 16606
rect 114940 15092 115108 15148
rect 115724 15092 115892 15148
rect 112588 14914 112644 14924
rect 110572 14644 110628 14654
rect 110628 14588 110740 14644
rect 110572 14550 110628 14588
rect 110460 14308 110516 14318
rect 110460 13972 110516 14252
rect 110572 13972 110628 13982
rect 110460 13970 110628 13972
rect 110460 13918 110574 13970
rect 110626 13918 110628 13970
rect 110460 13916 110628 13918
rect 110572 13906 110628 13916
rect 110348 13458 110404 13468
rect 109116 13188 109172 13198
rect 109116 13074 109172 13132
rect 109116 13022 109118 13074
rect 109170 13022 109172 13074
rect 109116 13010 109172 13022
rect 110348 13076 110404 13086
rect 109564 12964 109620 12974
rect 109564 12870 109620 12908
rect 110012 12964 110068 12974
rect 109676 12740 109732 12750
rect 109340 12404 109396 12414
rect 109340 12310 109396 12348
rect 109452 12178 109508 12190
rect 109452 12126 109454 12178
rect 109506 12126 109508 12178
rect 109340 11954 109396 11966
rect 109340 11902 109342 11954
rect 109394 11902 109396 11954
rect 109340 11620 109396 11902
rect 109116 11564 109396 11620
rect 109116 11172 109172 11564
rect 109452 11508 109508 12126
rect 109452 11442 109508 11452
rect 109228 11396 109284 11406
rect 109228 11394 109396 11396
rect 109228 11342 109230 11394
rect 109282 11342 109396 11394
rect 109228 11340 109396 11342
rect 109228 11330 109284 11340
rect 109116 11116 109284 11172
rect 109228 10164 109284 11116
rect 109116 10108 109284 10164
rect 109116 10052 109172 10108
rect 109116 9986 109172 9996
rect 109228 9940 109284 9950
rect 109228 9846 109284 9884
rect 109004 9660 109172 9716
rect 108780 8530 108836 8540
rect 108892 9602 108948 9614
rect 108892 9550 108894 9602
rect 108946 9550 108948 9602
rect 108892 8484 108948 9550
rect 109004 9044 109060 9054
rect 109004 8950 109060 8988
rect 108892 8428 109060 8484
rect 108556 8306 108612 8316
rect 108892 8036 108948 8046
rect 108444 7812 108500 7822
rect 108444 7362 108500 7756
rect 108892 7586 108948 7980
rect 108892 7534 108894 7586
rect 108946 7534 108948 7586
rect 108892 7522 108948 7534
rect 109004 7364 109060 8428
rect 108444 7310 108446 7362
rect 108498 7310 108500 7362
rect 108444 7140 108500 7310
rect 108444 7074 108500 7084
rect 108892 7308 109060 7364
rect 108780 6132 108836 6142
rect 108780 6038 108836 6076
rect 108108 4274 108164 4284
rect 108556 5348 108612 5358
rect 108332 3892 108388 3902
rect 108332 3442 108388 3836
rect 108332 3390 108334 3442
rect 108386 3390 108388 3442
rect 108332 3378 108388 3390
rect 107604 3276 107716 3332
rect 108556 3332 108612 5292
rect 108780 5236 108836 5246
rect 108668 5234 108836 5236
rect 108668 5182 108782 5234
rect 108834 5182 108836 5234
rect 108668 5180 108836 5182
rect 108668 3554 108724 5180
rect 108780 5170 108836 5180
rect 108668 3502 108670 3554
rect 108722 3502 108724 3554
rect 108668 3490 108724 3502
rect 108892 3556 108948 7308
rect 109004 7140 109060 7150
rect 109004 6130 109060 7084
rect 109004 6078 109006 6130
rect 109058 6078 109060 6130
rect 109004 6066 109060 6078
rect 109116 6018 109172 9660
rect 109116 5966 109118 6018
rect 109170 5966 109172 6018
rect 109116 5954 109172 5966
rect 109228 6468 109284 6478
rect 109228 4340 109284 6412
rect 109340 5796 109396 11340
rect 109452 11172 109508 11182
rect 109452 11170 109620 11172
rect 109452 11118 109454 11170
rect 109506 11118 109620 11170
rect 109452 11116 109620 11118
rect 109452 11106 109508 11116
rect 109452 10724 109508 10734
rect 109452 10630 109508 10668
rect 109564 7476 109620 11116
rect 109676 10722 109732 12684
rect 109900 12068 109956 12078
rect 109900 11974 109956 12012
rect 110012 11844 110068 12908
rect 110348 12402 110404 13020
rect 110684 12962 110740 14588
rect 111468 14308 111524 14318
rect 111468 13858 111524 14252
rect 111996 14140 112260 14150
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 111996 14074 112260 14084
rect 111468 13806 111470 13858
rect 111522 13806 111524 13858
rect 111468 13794 111524 13806
rect 112028 13636 112084 13646
rect 111804 13634 112084 13636
rect 111804 13582 112030 13634
rect 112082 13582 112084 13634
rect 111804 13580 112084 13582
rect 110684 12910 110686 12962
rect 110738 12910 110740 12962
rect 110684 12898 110740 12910
rect 111132 13524 111188 13534
rect 110796 12740 110852 12750
rect 110348 12350 110350 12402
rect 110402 12350 110404 12402
rect 110348 12338 110404 12350
rect 110460 12738 110852 12740
rect 110460 12686 110798 12738
rect 110850 12686 110852 12738
rect 110460 12684 110852 12686
rect 110012 11778 110068 11788
rect 109900 11732 109956 11742
rect 109900 11394 109956 11676
rect 109900 11342 109902 11394
rect 109954 11342 109956 11394
rect 109900 11330 109956 11342
rect 110124 11170 110180 11182
rect 110124 11118 110126 11170
rect 110178 11118 110180 11170
rect 109676 10670 109678 10722
rect 109730 10670 109732 10722
rect 109676 10658 109732 10670
rect 109788 10834 109844 10846
rect 109788 10782 109790 10834
rect 109842 10782 109844 10834
rect 109676 9604 109732 9614
rect 109676 9042 109732 9548
rect 109676 8990 109678 9042
rect 109730 8990 109732 9042
rect 109676 8484 109732 8990
rect 109676 8418 109732 8428
rect 109564 7410 109620 7420
rect 109676 6692 109732 6702
rect 109788 6692 109844 10782
rect 110012 10724 110068 10734
rect 110012 10630 110068 10668
rect 109900 10612 109956 10622
rect 109900 8820 109956 10556
rect 110124 9604 110180 11118
rect 110348 10498 110404 10510
rect 110348 10446 110350 10498
rect 110402 10446 110404 10498
rect 110348 10388 110404 10446
rect 110124 9538 110180 9548
rect 110236 10052 110292 10062
rect 109900 8754 109956 8764
rect 110236 8148 110292 9996
rect 109676 6690 109844 6692
rect 109676 6638 109678 6690
rect 109730 6638 109844 6690
rect 109676 6636 109844 6638
rect 110012 8146 110292 8148
rect 110012 8094 110238 8146
rect 110290 8094 110292 8146
rect 110012 8092 110292 8094
rect 109676 6626 109732 6636
rect 109452 5796 109508 5806
rect 109340 5794 109508 5796
rect 109340 5742 109454 5794
rect 109506 5742 109508 5794
rect 109340 5740 109508 5742
rect 109452 5730 109508 5740
rect 109564 5572 109620 5582
rect 109340 4340 109396 4350
rect 109228 4338 109396 4340
rect 109228 4286 109342 4338
rect 109394 4286 109396 4338
rect 109228 4284 109396 4286
rect 109340 4274 109396 4284
rect 109564 4226 109620 5516
rect 110012 4788 110068 8092
rect 110236 8082 110292 8092
rect 110236 7364 110292 7374
rect 110236 7270 110292 7308
rect 110348 7140 110404 10332
rect 110236 7084 110404 7140
rect 110236 6804 110292 7084
rect 110236 6738 110292 6748
rect 110348 6692 110404 6702
rect 110348 6598 110404 6636
rect 110124 5236 110180 5246
rect 110124 5142 110180 5180
rect 110012 4722 110068 4732
rect 110124 4676 110180 4686
rect 109564 4174 109566 4226
rect 109618 4174 109620 4226
rect 109564 4162 109620 4174
rect 109676 4338 109732 4350
rect 109676 4286 109678 4338
rect 109730 4286 109732 4338
rect 109228 4114 109284 4126
rect 109228 4062 109230 4114
rect 109282 4062 109284 4114
rect 109004 3556 109060 3566
rect 108892 3554 109060 3556
rect 108892 3502 109006 3554
rect 109058 3502 109060 3554
rect 108892 3500 109060 3502
rect 109004 3490 109060 3500
rect 109228 3556 109284 4062
rect 109228 3490 109284 3500
rect 109676 3892 109732 4286
rect 108556 3276 108724 3332
rect 107548 3266 107604 3276
rect 106876 2818 106932 2828
rect 107324 3164 107492 3220
rect 107324 800 107380 3164
rect 108668 800 108724 3276
rect 109676 3220 109732 3836
rect 110124 3780 110180 4620
rect 110124 3714 110180 3724
rect 110460 3668 110516 12684
rect 110796 12674 110852 12684
rect 110908 12628 110964 12638
rect 110796 12516 110852 12526
rect 110796 12402 110852 12460
rect 110796 12350 110798 12402
rect 110850 12350 110852 12402
rect 110796 12338 110852 12350
rect 110684 11282 110740 11294
rect 110684 11230 110686 11282
rect 110738 11230 110740 11282
rect 110572 10948 110628 10958
rect 110572 10612 110628 10892
rect 110572 10546 110628 10556
rect 110684 9156 110740 11230
rect 110796 11170 110852 11182
rect 110796 11118 110798 11170
rect 110850 11118 110852 11170
rect 110796 10388 110852 11118
rect 110908 11172 110964 12572
rect 111020 11508 111076 11518
rect 111020 11394 111076 11452
rect 111020 11342 111022 11394
rect 111074 11342 111076 11394
rect 111020 11330 111076 11342
rect 110908 11116 111076 11172
rect 110908 10836 110964 10846
rect 110908 10742 110964 10780
rect 111020 10388 111076 11116
rect 110796 10322 110852 10332
rect 110908 10332 111076 10388
rect 110684 9100 110852 9156
rect 110572 8930 110628 8942
rect 110572 8878 110574 8930
rect 110626 8878 110628 8930
rect 110572 8708 110628 8878
rect 110572 8642 110628 8652
rect 110684 8932 110740 8942
rect 110684 8596 110740 8876
rect 110684 8484 110740 8540
rect 110572 8428 110740 8484
rect 110572 7698 110628 8428
rect 110684 8260 110740 8270
rect 110684 8166 110740 8204
rect 110572 7646 110574 7698
rect 110626 7646 110628 7698
rect 110572 7634 110628 7646
rect 110572 7476 110628 7486
rect 110572 5796 110628 7420
rect 110796 7252 110852 9100
rect 110908 8146 110964 10332
rect 111132 8708 111188 13468
rect 111580 13522 111636 13534
rect 111580 13470 111582 13522
rect 111634 13470 111636 13522
rect 111244 12740 111300 12750
rect 111244 12646 111300 12684
rect 111580 12292 111636 13470
rect 111692 12852 111748 12862
rect 111692 12758 111748 12796
rect 111580 12236 111748 12292
rect 111580 12066 111636 12078
rect 111580 12014 111582 12066
rect 111634 12014 111636 12066
rect 111580 11954 111636 12014
rect 111580 11902 111582 11954
rect 111634 11902 111636 11954
rect 111580 11732 111636 11902
rect 111580 11666 111636 11676
rect 111468 11282 111524 11294
rect 111468 11230 111470 11282
rect 111522 11230 111524 11282
rect 111468 11060 111524 11230
rect 111356 11004 111524 11060
rect 111580 11170 111636 11182
rect 111580 11118 111582 11170
rect 111634 11118 111636 11170
rect 111356 10052 111412 11004
rect 111580 10836 111636 11118
rect 111244 9996 111412 10052
rect 111468 10780 111636 10836
rect 111244 9828 111300 9996
rect 111468 9940 111524 10780
rect 111468 9874 111524 9884
rect 111580 10612 111636 10622
rect 111244 8932 111300 9772
rect 111356 9714 111412 9726
rect 111356 9662 111358 9714
rect 111410 9662 111412 9714
rect 111356 9156 111412 9662
rect 111356 9090 111412 9100
rect 111580 9044 111636 10556
rect 111692 9268 111748 12236
rect 111804 11396 111860 13580
rect 112028 13570 112084 13580
rect 112140 12964 112196 12974
rect 112140 12870 112196 12908
rect 112700 12852 112756 12862
rect 111996 12572 112260 12582
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 111996 12506 112260 12516
rect 112700 12404 112756 12796
rect 113036 12740 113092 12750
rect 113820 12740 113876 12750
rect 113036 12738 113316 12740
rect 113036 12686 113038 12738
rect 113090 12686 113316 12738
rect 113036 12684 113316 12686
rect 113036 12674 113092 12684
rect 112700 12338 112756 12348
rect 112028 12068 112084 12078
rect 112028 12066 112420 12068
rect 112028 12014 112030 12066
rect 112082 12014 112420 12066
rect 112028 12012 112420 12014
rect 112028 12002 112084 12012
rect 112140 11396 112196 11406
rect 111804 11340 111972 11396
rect 111916 11284 111972 11340
rect 112140 11302 112196 11340
rect 111916 11218 111972 11228
rect 111804 11170 111860 11182
rect 111804 11118 111806 11170
rect 111858 11118 111860 11170
rect 111804 10164 111860 11118
rect 111996 11004 112260 11014
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 111996 10938 112260 10948
rect 112140 10498 112196 10510
rect 112140 10446 112142 10498
rect 112194 10446 112196 10498
rect 112140 10276 112196 10446
rect 112140 10210 112196 10220
rect 111804 10098 111860 10108
rect 112028 10052 112084 10062
rect 112364 10052 112420 12012
rect 112476 12066 112532 12078
rect 112476 12014 112478 12066
rect 112530 12014 112532 12066
rect 112476 11956 112532 12014
rect 112924 12068 112980 12078
rect 112924 11974 112980 12012
rect 112476 11890 112532 11900
rect 112588 11954 112644 11966
rect 112588 11902 112590 11954
rect 112642 11902 112644 11954
rect 112588 11506 112644 11902
rect 112588 11454 112590 11506
rect 112642 11454 112644 11506
rect 112588 11442 112644 11454
rect 112700 11618 112756 11630
rect 112700 11566 112702 11618
rect 112754 11566 112756 11618
rect 112700 10612 112756 11566
rect 112084 9996 112420 10052
rect 112588 10610 112756 10612
rect 112588 10558 112702 10610
rect 112754 10558 112756 10610
rect 112588 10556 112756 10558
rect 112028 9986 112084 9996
rect 112588 9940 112644 10556
rect 112700 10546 112756 10556
rect 112812 11508 112868 11518
rect 112140 9884 112644 9940
rect 112140 9826 112196 9884
rect 112140 9774 112142 9826
rect 112194 9774 112196 9826
rect 112140 9762 112196 9774
rect 111996 9436 112260 9446
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 111996 9370 112260 9380
rect 111692 9202 111748 9212
rect 111468 9042 111636 9044
rect 111468 8990 111582 9042
rect 111634 8990 111636 9042
rect 111468 8988 111636 8990
rect 111244 8876 111412 8932
rect 111132 8652 111300 8708
rect 111132 8484 111188 8494
rect 110908 8094 110910 8146
rect 110962 8094 110964 8146
rect 110908 8082 110964 8094
rect 111020 8146 111076 8158
rect 111020 8094 111022 8146
rect 111074 8094 111076 8146
rect 111020 8036 111076 8094
rect 110908 7924 110964 7934
rect 110908 7698 110964 7868
rect 110908 7646 110910 7698
rect 110962 7646 110964 7698
rect 110908 7634 110964 7646
rect 111020 7252 111076 7980
rect 110796 7196 111076 7252
rect 110796 6468 110852 7196
rect 110908 6692 110964 6702
rect 111132 6692 111188 8428
rect 111244 7028 111300 8652
rect 111356 8596 111412 8876
rect 111356 8530 111412 8540
rect 111356 8370 111412 8382
rect 111356 8318 111358 8370
rect 111410 8318 111412 8370
rect 111356 8148 111412 8318
rect 111356 8082 111412 8092
rect 111468 7698 111524 8988
rect 111580 8978 111636 8988
rect 112364 9044 112420 9884
rect 112476 9714 112532 9726
rect 112476 9662 112478 9714
rect 112530 9662 112532 9714
rect 112476 9604 112532 9662
rect 112476 9538 112532 9548
rect 112700 9714 112756 9726
rect 112700 9662 112702 9714
rect 112754 9662 112756 9714
rect 112476 9268 112532 9278
rect 112700 9268 112756 9662
rect 112532 9212 112644 9268
rect 112476 9202 112532 9212
rect 112364 8978 112420 8988
rect 112140 8930 112196 8942
rect 112140 8878 112142 8930
rect 112194 8878 112196 8930
rect 112140 8260 112196 8878
rect 112476 8708 112532 8718
rect 112140 8194 112196 8204
rect 112364 8484 112420 8494
rect 112476 8484 112532 8652
rect 112588 8596 112644 9212
rect 112700 9202 112756 9212
rect 112812 9044 112868 11452
rect 113036 11172 113092 11182
rect 113036 11078 113092 11116
rect 113260 10276 113316 12684
rect 113820 12404 113876 12684
rect 113484 12402 113876 12404
rect 113484 12350 113822 12402
rect 113874 12350 113876 12402
rect 113484 12348 113876 12350
rect 113372 12066 113428 12078
rect 113372 12014 113374 12066
rect 113426 12014 113428 12066
rect 113372 11954 113428 12014
rect 113372 11902 113374 11954
rect 113426 11902 113428 11954
rect 113372 11890 113428 11902
rect 113484 11618 113540 12348
rect 113820 12338 113876 12348
rect 113484 11566 113486 11618
rect 113538 11566 113540 11618
rect 113484 11506 113540 11566
rect 114380 11618 114436 11630
rect 114380 11566 114382 11618
rect 114434 11566 114436 11618
rect 114380 11508 114436 11566
rect 113484 11454 113486 11506
rect 113538 11454 113540 11506
rect 113484 11442 113540 11454
rect 114268 11506 114436 11508
rect 114268 11454 114382 11506
rect 114434 11454 114436 11506
rect 114268 11452 114436 11454
rect 114044 11170 114100 11182
rect 114044 11118 114046 11170
rect 114098 11118 114100 11170
rect 113372 10500 113428 10510
rect 113372 10498 113652 10500
rect 113372 10446 113374 10498
rect 113426 10446 113652 10498
rect 113372 10444 113652 10446
rect 113372 10434 113428 10444
rect 113260 10220 113540 10276
rect 113148 10164 113204 10174
rect 113204 10108 113316 10164
rect 113148 10098 113204 10108
rect 113148 9826 113204 9838
rect 113148 9774 113150 9826
rect 113202 9774 113204 9826
rect 112924 9602 112980 9614
rect 112924 9550 112926 9602
rect 112978 9550 112980 9602
rect 112924 9380 112980 9550
rect 113148 9492 113204 9774
rect 113148 9426 113204 9436
rect 112924 9314 112980 9324
rect 113148 9156 113204 9166
rect 113036 9154 113204 9156
rect 113036 9102 113150 9154
rect 113202 9102 113204 9154
rect 113036 9100 113204 9102
rect 112924 9044 112980 9054
rect 112812 9042 112980 9044
rect 112812 8990 112926 9042
rect 112978 8990 112980 9042
rect 112812 8988 112980 8990
rect 112924 8978 112980 8988
rect 113036 9044 113092 9100
rect 113148 9090 113204 9100
rect 113036 8978 113092 8988
rect 113260 9042 113316 10108
rect 113260 8990 113262 9042
rect 113314 8990 113316 9042
rect 113260 8978 113316 8990
rect 113372 9714 113428 9726
rect 113372 9662 113374 9714
rect 113426 9662 113428 9714
rect 113372 9604 113428 9662
rect 113372 9044 113428 9548
rect 113484 9380 113540 10220
rect 113596 9604 113652 10444
rect 113708 9940 113764 9950
rect 113708 9826 113764 9884
rect 113708 9774 113710 9826
rect 113762 9774 113764 9826
rect 113708 9762 113764 9774
rect 113932 9716 113988 9726
rect 113932 9622 113988 9660
rect 113708 9604 113764 9614
rect 113596 9602 113764 9604
rect 113596 9550 113710 9602
rect 113762 9550 113764 9602
rect 113596 9548 113764 9550
rect 113708 9538 113764 9548
rect 113820 9492 113876 9502
rect 113484 9324 113764 9380
rect 113484 9044 113540 9054
rect 113372 8988 113484 9044
rect 113484 8950 113540 8988
rect 112588 8540 113092 8596
rect 112476 8428 112644 8484
rect 111996 7868 112260 7878
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 111996 7802 112260 7812
rect 111468 7646 111470 7698
rect 111522 7646 111524 7698
rect 111468 7634 111524 7646
rect 112028 7362 112084 7374
rect 112028 7310 112030 7362
rect 112082 7310 112084 7362
rect 112028 7028 112084 7310
rect 112364 7364 112420 8428
rect 112476 7364 112532 7374
rect 112364 7362 112532 7364
rect 112364 7310 112478 7362
rect 112530 7310 112532 7362
rect 112364 7308 112532 7310
rect 111244 6972 111748 7028
rect 110908 6690 111188 6692
rect 110908 6638 110910 6690
rect 110962 6638 111188 6690
rect 110908 6636 111188 6638
rect 110908 6626 110964 6636
rect 111356 6580 111412 6590
rect 111244 6578 111412 6580
rect 111244 6526 111358 6578
rect 111410 6526 111412 6578
rect 111244 6524 111412 6526
rect 110796 6412 110964 6468
rect 110684 6020 110740 6030
rect 110684 5926 110740 5964
rect 110572 5740 110852 5796
rect 110796 4562 110852 5740
rect 110796 4510 110798 4562
rect 110850 4510 110852 4562
rect 110796 4498 110852 4510
rect 110908 4564 110964 6412
rect 111244 5572 111300 6524
rect 111356 6514 111412 6524
rect 111356 6020 111412 6030
rect 111356 5926 111412 5964
rect 111244 5506 111300 5516
rect 111580 5908 111636 5918
rect 110908 4450 110964 4508
rect 111356 5236 111412 5246
rect 111356 5010 111412 5180
rect 111356 4958 111358 5010
rect 111410 4958 111412 5010
rect 111356 4564 111412 4958
rect 111356 4498 111412 4508
rect 110908 4398 110910 4450
rect 110962 4398 110964 4450
rect 110908 4386 110964 4398
rect 110572 4340 110628 4350
rect 111580 4340 111636 5852
rect 110572 4246 110628 4284
rect 111356 4284 111636 4340
rect 110460 3602 110516 3612
rect 109676 3154 109732 3164
rect 110012 3330 110068 3342
rect 110012 3278 110014 3330
rect 110066 3278 110068 3330
rect 110012 800 110068 3278
rect 111356 800 111412 4284
rect 111692 4228 111748 6972
rect 112028 6962 112084 6972
rect 112364 6580 112420 6618
rect 112364 6514 112420 6524
rect 111804 6466 111860 6478
rect 111804 6414 111806 6466
rect 111858 6414 111860 6466
rect 111804 5348 111860 6414
rect 112364 6356 112420 6366
rect 111996 6300 112260 6310
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 111996 6234 112260 6244
rect 111804 5282 111860 5292
rect 112364 5236 112420 6300
rect 112364 5170 112420 5180
rect 111916 5124 111972 5134
rect 111916 5030 111972 5068
rect 111804 4900 111860 4910
rect 111804 4806 111860 4844
rect 111996 4732 112260 4742
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 111996 4666 112260 4676
rect 111692 4162 111748 4172
rect 112252 4228 112308 4238
rect 112252 4134 112308 4172
rect 112476 3388 112532 7308
rect 112588 4900 112644 8428
rect 112924 6580 112980 6590
rect 112588 4338 112644 4844
rect 112588 4286 112590 4338
rect 112642 4286 112644 4338
rect 112588 4274 112644 4286
rect 112700 6020 112756 6030
rect 111468 3332 112532 3388
rect 111468 2996 111524 3332
rect 111996 3164 112260 3174
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 111996 3098 112260 3108
rect 111468 2930 111524 2940
rect 112700 800 112756 5964
rect 112924 5908 112980 6524
rect 112924 5842 112980 5852
rect 113036 5234 113092 8540
rect 113484 8372 113540 8382
rect 113484 8278 113540 8316
rect 113708 6580 113764 9324
rect 113820 8036 113876 9436
rect 113932 9044 113988 9054
rect 113932 8950 113988 8988
rect 113820 7970 113876 7980
rect 114044 7812 114100 11118
rect 114156 9940 114212 9950
rect 114156 9826 114212 9884
rect 114156 9774 114158 9826
rect 114210 9774 114212 9826
rect 114156 9762 114212 9774
rect 114156 9156 114212 9166
rect 114156 9062 114212 9100
rect 114268 8260 114324 11452
rect 114380 11442 114436 11452
rect 114828 11618 114884 11630
rect 114828 11566 114830 11618
rect 114882 11566 114884 11618
rect 114828 11506 114884 11566
rect 114828 11454 114830 11506
rect 114882 11454 114884 11506
rect 114828 11442 114884 11454
rect 114380 10500 114436 10510
rect 114380 9714 114436 10444
rect 114828 10388 114884 10398
rect 114492 9828 114548 9838
rect 114492 9734 114548 9772
rect 114380 9662 114382 9714
rect 114434 9662 114436 9714
rect 114380 9650 114436 9662
rect 114828 9266 114884 10332
rect 114828 9214 114830 9266
rect 114882 9214 114884 9266
rect 114828 9202 114884 9214
rect 114604 9042 114660 9054
rect 114604 8990 114606 9042
rect 114658 8990 114660 9042
rect 114268 8166 114324 8204
rect 114380 8930 114436 8942
rect 114380 8878 114382 8930
rect 114434 8878 114436 8930
rect 114044 7746 114100 7756
rect 114380 7588 114436 8878
rect 114604 8372 114660 8990
rect 114604 8306 114660 8316
rect 114604 8146 114660 8158
rect 114940 8148 114996 8158
rect 114604 8094 114606 8146
rect 114658 8094 114660 8146
rect 114604 7924 114660 8094
rect 114828 8146 114996 8148
rect 114828 8094 114942 8146
rect 114994 8094 114996 8146
rect 114828 8092 114996 8094
rect 114604 7858 114660 7868
rect 114716 8034 114772 8046
rect 114716 7982 114718 8034
rect 114770 7982 114772 8034
rect 114604 7588 114660 7598
rect 114380 7586 114660 7588
rect 114380 7534 114606 7586
rect 114658 7534 114660 7586
rect 114380 7532 114660 7534
rect 114604 7522 114660 7532
rect 114716 7476 114772 7982
rect 114828 8036 114884 8092
rect 114940 8082 114996 8092
rect 114828 7970 114884 7980
rect 114716 7410 114772 7420
rect 115052 7140 115108 15092
rect 115500 10500 115556 10510
rect 115500 10406 115556 10444
rect 115612 9828 115668 9838
rect 115668 9772 115780 9828
rect 115612 9734 115668 9772
rect 115276 9602 115332 9614
rect 115276 9550 115278 9602
rect 115330 9550 115332 9602
rect 115276 9156 115332 9550
rect 115500 9604 115556 9614
rect 115388 9268 115444 9278
rect 115388 9174 115444 9212
rect 115276 9090 115332 9100
rect 115164 9042 115220 9054
rect 115164 8990 115166 9042
rect 115218 8990 115220 9042
rect 115164 8708 115220 8990
rect 115164 8652 115444 8708
rect 115388 8370 115444 8652
rect 115500 8484 115556 9548
rect 115500 8418 115556 8428
rect 115612 9154 115668 9166
rect 115612 9102 115614 9154
rect 115666 9102 115668 9154
rect 115388 8318 115390 8370
rect 115442 8318 115444 8370
rect 115388 8306 115444 8318
rect 115276 8260 115332 8270
rect 115276 7474 115332 8204
rect 115612 8148 115668 9102
rect 115724 9154 115780 9772
rect 115724 9102 115726 9154
rect 115778 9102 115780 9154
rect 115724 9090 115780 9102
rect 115612 8082 115668 8092
rect 115276 7422 115278 7474
rect 115330 7422 115332 7474
rect 115276 7410 115332 7422
rect 115724 7588 115780 7598
rect 115052 7074 115108 7084
rect 115612 7364 115668 7374
rect 113708 6514 113764 6524
rect 114268 6804 114324 6814
rect 113484 6356 113540 6366
rect 113484 6018 113540 6300
rect 114268 6132 114324 6748
rect 114716 6580 114772 6590
rect 114716 6486 114772 6524
rect 115500 6580 115556 6590
rect 115500 6486 115556 6524
rect 114268 6066 114324 6076
rect 114380 6468 114436 6478
rect 114380 6130 114436 6412
rect 114380 6078 114382 6130
rect 114434 6078 114436 6130
rect 114380 6066 114436 6078
rect 115164 6132 115220 6142
rect 113484 5966 113486 6018
rect 113538 5966 113540 6018
rect 113484 5954 113540 5966
rect 115164 6018 115220 6076
rect 115164 5966 115166 6018
rect 115218 5966 115220 6018
rect 115164 5954 115220 5966
rect 115612 5348 115668 7308
rect 113036 5182 113038 5234
rect 113090 5182 113092 5234
rect 113036 5170 113092 5182
rect 115276 5292 115668 5348
rect 113260 5122 113316 5134
rect 113260 5070 113262 5122
rect 113314 5070 113316 5122
rect 113260 4900 113316 5070
rect 113820 5010 113876 5022
rect 113820 4958 113822 5010
rect 113874 4958 113876 5010
rect 113036 4564 113092 4574
rect 113036 4450 113092 4508
rect 113036 4398 113038 4450
rect 113090 4398 113092 4450
rect 113036 4386 113092 4398
rect 113260 4340 113316 4844
rect 112924 3668 112980 3678
rect 112924 3574 112980 3612
rect 113260 3554 113316 4284
rect 113260 3502 113262 3554
rect 113314 3502 113316 3554
rect 113260 3490 113316 3502
rect 113372 4898 113428 4910
rect 113372 4846 113374 4898
rect 113426 4846 113428 4898
rect 113372 3108 113428 4846
rect 113820 4564 113876 4958
rect 113708 3444 113764 3454
rect 113820 3444 113876 4508
rect 113708 3442 113876 3444
rect 113708 3390 113710 3442
rect 113762 3390 113876 3442
rect 113708 3388 113876 3390
rect 113932 4562 113988 4574
rect 113932 4510 113934 4562
rect 113986 4510 113988 4562
rect 113708 3378 113764 3388
rect 113372 3042 113428 3052
rect 113932 2772 113988 4510
rect 115164 4228 115220 4238
rect 115164 4134 115220 4172
rect 115276 3554 115332 5292
rect 115500 4562 115556 4574
rect 115500 4510 115502 4562
rect 115554 4510 115556 4562
rect 115388 4340 115444 4350
rect 115388 4246 115444 4284
rect 115276 3502 115278 3554
rect 115330 3502 115332 3554
rect 115276 3490 115332 3502
rect 113932 2706 113988 2716
rect 114044 3444 114100 3454
rect 114044 800 114100 3388
rect 114604 3332 114660 3342
rect 114604 3238 114660 3276
rect 115052 3330 115108 3342
rect 115052 3278 115054 3330
rect 115106 3278 115108 3330
rect 115052 2660 115108 3278
rect 115500 2996 115556 4510
rect 115500 2930 115556 2940
rect 115724 2772 115780 7532
rect 115836 5236 115892 15092
rect 116060 11620 116116 11630
rect 115948 10500 116004 10510
rect 115948 10406 116004 10444
rect 116060 10050 116116 11564
rect 117292 10724 117348 10734
rect 117348 10668 117460 10724
rect 117292 10658 117348 10668
rect 116060 9998 116062 10050
rect 116114 9998 116116 10050
rect 116060 9938 116116 9998
rect 116060 9886 116062 9938
rect 116114 9886 116116 9938
rect 116060 9874 116116 9886
rect 116396 10498 116452 10510
rect 116396 10446 116398 10498
rect 116450 10446 116452 10498
rect 115948 9716 116004 9726
rect 115948 9266 116004 9660
rect 116396 9604 116452 10446
rect 117068 10052 117124 10062
rect 117068 10050 117236 10052
rect 117068 9998 117070 10050
rect 117122 9998 117236 10050
rect 117068 9996 117236 9998
rect 117068 9986 117124 9996
rect 116396 9538 116452 9548
rect 116508 9602 116564 9614
rect 116508 9550 116510 9602
rect 116562 9550 116564 9602
rect 115948 9214 115950 9266
rect 116002 9214 116004 9266
rect 115948 9202 116004 9214
rect 116172 9156 116228 9166
rect 116172 9062 116228 9100
rect 116284 9042 116340 9054
rect 116284 8990 116286 9042
rect 116338 8990 116340 9042
rect 116284 8820 116340 8990
rect 116284 8754 116340 8764
rect 116396 7588 116452 7598
rect 116396 7494 116452 7532
rect 116284 6916 116340 6926
rect 116172 5236 116228 5246
rect 115836 5234 116228 5236
rect 115836 5182 116174 5234
rect 116226 5182 116228 5234
rect 115836 5180 116228 5182
rect 116172 5170 116228 5180
rect 115948 4900 116004 4910
rect 115948 4450 116004 4844
rect 115948 4398 115950 4450
rect 116002 4398 116004 4450
rect 115948 4386 116004 4398
rect 116172 3556 116228 3566
rect 116284 3556 116340 6860
rect 116508 5908 116564 9550
rect 116956 9604 117012 9614
rect 116956 9602 117124 9604
rect 116956 9550 116958 9602
rect 117010 9550 117124 9602
rect 116956 9548 117124 9550
rect 116956 9538 117012 9548
rect 116732 8930 116788 8942
rect 116732 8878 116734 8930
rect 116786 8878 116788 8930
rect 116732 8260 116788 8878
rect 116732 8194 116788 8204
rect 116620 8146 116676 8158
rect 116620 8094 116622 8146
rect 116674 8094 116676 8146
rect 116620 7028 116676 8094
rect 116620 6972 116788 7028
rect 116508 5852 116676 5908
rect 116396 5572 116452 5582
rect 116396 5122 116452 5516
rect 116396 5070 116398 5122
rect 116450 5070 116452 5122
rect 116396 5058 116452 5070
rect 116620 4004 116676 5852
rect 116732 5796 116788 6972
rect 116844 6802 116900 6814
rect 116844 6750 116846 6802
rect 116898 6750 116900 6802
rect 116844 6020 116900 6750
rect 116844 5954 116900 5964
rect 116956 5796 117012 5806
rect 116732 5794 117012 5796
rect 116732 5742 116958 5794
rect 117010 5742 117012 5794
rect 116732 5740 117012 5742
rect 116956 5730 117012 5740
rect 117068 5796 117124 9548
rect 117180 9266 117236 9996
rect 117180 9214 117182 9266
rect 117234 9214 117236 9266
rect 117180 9202 117236 9214
rect 117180 8820 117236 8830
rect 117180 8258 117236 8764
rect 117180 8206 117182 8258
rect 117234 8206 117236 8258
rect 117180 6690 117236 8206
rect 117292 8036 117348 8046
rect 117292 7942 117348 7980
rect 117404 7812 117460 10668
rect 117628 8932 117684 8942
rect 117628 8838 117684 8876
rect 117964 8708 118020 18284
rect 118412 14980 118468 14990
rect 118468 14924 118580 14980
rect 118412 14914 118468 14924
rect 118300 10836 118356 10846
rect 118356 10780 118468 10836
rect 118300 10770 118356 10780
rect 118076 8932 118132 8942
rect 118076 8930 118244 8932
rect 118076 8878 118078 8930
rect 118130 8878 118244 8930
rect 118076 8876 118244 8878
rect 118076 8866 118132 8876
rect 117964 8652 118132 8708
rect 117628 8482 117684 8494
rect 117628 8430 117630 8482
rect 117682 8430 117684 8482
rect 117516 8372 117572 8382
rect 117516 8258 117572 8316
rect 117516 8206 117518 8258
rect 117570 8206 117572 8258
rect 117516 8194 117572 8206
rect 117292 7756 117460 7812
rect 117292 6914 117348 7756
rect 117404 7364 117460 7374
rect 117404 7270 117460 7308
rect 117292 6862 117294 6914
rect 117346 6862 117348 6914
rect 117292 6850 117348 6862
rect 117180 6638 117182 6690
rect 117234 6638 117236 6690
rect 117180 6626 117236 6638
rect 117292 6468 117348 6478
rect 117292 6374 117348 6412
rect 117628 6132 117684 8430
rect 117852 8034 117908 8046
rect 117852 7982 117854 8034
rect 117906 7982 117908 8034
rect 117740 7474 117796 7486
rect 117740 7422 117742 7474
rect 117794 7422 117796 7474
rect 117740 7364 117796 7422
rect 117740 7298 117796 7308
rect 117852 6804 117908 7982
rect 117852 6738 117908 6748
rect 117964 7028 118020 7038
rect 117628 6066 117684 6076
rect 117852 5908 117908 5918
rect 117068 5730 117124 5740
rect 117628 5794 117684 5806
rect 117628 5742 117630 5794
rect 117682 5742 117684 5794
rect 117628 5684 117684 5742
rect 117628 5618 117684 5628
rect 117852 5572 117908 5852
rect 117740 5516 117852 5572
rect 116956 5010 117012 5022
rect 116956 4958 116958 5010
rect 117010 4958 117012 5010
rect 116956 4900 117012 4958
rect 116956 4834 117012 4844
rect 116620 3938 116676 3948
rect 116732 4676 116788 4686
rect 116172 3554 116340 3556
rect 116172 3502 116174 3554
rect 116226 3502 116340 3554
rect 116172 3500 116340 3502
rect 116172 3490 116228 3500
rect 115052 2594 115108 2604
rect 115388 2716 115780 2772
rect 115388 800 115444 2716
rect 116732 800 116788 4620
rect 117740 4338 117796 5516
rect 117852 5506 117908 5516
rect 117852 4900 117908 4910
rect 117852 4806 117908 4844
rect 117740 4286 117742 4338
rect 117794 4286 117796 4338
rect 117740 4274 117796 4286
rect 117852 4338 117908 4350
rect 117852 4286 117854 4338
rect 117906 4286 117908 4338
rect 117852 4004 117908 4286
rect 117964 4226 118020 6972
rect 118076 5906 118132 8652
rect 118188 8482 118244 8876
rect 118188 8430 118190 8482
rect 118242 8430 118244 8482
rect 118188 8418 118244 8430
rect 118300 8260 118356 8270
rect 118300 8166 118356 8204
rect 118188 7364 118244 7374
rect 118188 7270 118244 7308
rect 118412 7140 118468 10780
rect 118188 7084 118468 7140
rect 118188 6802 118244 7084
rect 118188 6750 118190 6802
rect 118242 6750 118244 6802
rect 118188 6738 118244 6750
rect 118076 5854 118078 5906
rect 118130 5854 118132 5906
rect 118076 5842 118132 5854
rect 118524 5572 118580 14924
rect 119756 14532 119812 55022
rect 125132 32788 125188 55916
rect 127356 55692 127620 55702
rect 127412 55636 127460 55692
rect 127516 55636 127564 55692
rect 127356 55626 127620 55636
rect 127708 55468 127764 56030
rect 131516 56082 131572 56094
rect 131516 56030 131518 56082
rect 131570 56030 131572 56082
rect 131516 55468 131572 56030
rect 127484 55412 127764 55468
rect 131180 55412 131572 55468
rect 127260 55298 127316 55310
rect 127260 55246 127262 55298
rect 127314 55246 127316 55298
rect 126812 55188 126868 55198
rect 126812 54404 126868 55132
rect 127260 55188 127316 55246
rect 127260 55122 127316 55132
rect 127484 55186 127540 55412
rect 127484 55134 127486 55186
rect 127538 55134 127540 55186
rect 127484 55122 127540 55134
rect 126812 54338 126868 54348
rect 131180 55074 131236 55412
rect 135100 55410 135156 56252
rect 135324 56242 135380 56252
rect 138908 56308 138964 59200
rect 142716 57092 142772 59200
rect 142716 57026 142772 57036
rect 144508 57092 144564 57102
rect 142716 56476 142980 56486
rect 142772 56420 142820 56476
rect 142876 56420 142924 56476
rect 142716 56410 142980 56420
rect 138908 56242 138964 56252
rect 140140 56308 140196 56318
rect 140140 56214 140196 56252
rect 144508 56194 144564 57036
rect 146524 56308 146580 59200
rect 146748 56308 146804 56318
rect 146524 56306 146804 56308
rect 146524 56254 146750 56306
rect 146802 56254 146804 56306
rect 146524 56252 146804 56254
rect 144508 56142 144510 56194
rect 144562 56142 144564 56194
rect 144508 56130 144564 56142
rect 139244 56082 139300 56094
rect 139244 56030 139246 56082
rect 139298 56030 139300 56082
rect 135772 55972 135828 55982
rect 135772 55878 135828 55916
rect 136892 55972 136948 55982
rect 135100 55358 135102 55410
rect 135154 55358 135156 55410
rect 135100 55346 135156 55358
rect 131180 55022 131182 55074
rect 131234 55022 131236 55074
rect 127356 54124 127620 54134
rect 127412 54068 127460 54124
rect 127516 54068 127564 54124
rect 127356 54058 127620 54068
rect 127356 52556 127620 52566
rect 127412 52500 127460 52556
rect 127516 52500 127564 52556
rect 127356 52490 127620 52500
rect 127356 50988 127620 50998
rect 127412 50932 127460 50988
rect 127516 50932 127564 50988
rect 127356 50922 127620 50932
rect 127356 49420 127620 49430
rect 127412 49364 127460 49420
rect 127516 49364 127564 49420
rect 127356 49354 127620 49364
rect 127356 47852 127620 47862
rect 127412 47796 127460 47852
rect 127516 47796 127564 47852
rect 127356 47786 127620 47796
rect 127356 46284 127620 46294
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127356 46218 127620 46228
rect 127356 44716 127620 44726
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127356 44650 127620 44660
rect 127356 43148 127620 43158
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127356 43082 127620 43092
rect 127356 41580 127620 41590
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127356 41514 127620 41524
rect 127356 40012 127620 40022
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127356 39946 127620 39956
rect 127356 38444 127620 38454
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127356 38378 127620 38388
rect 127356 36876 127620 36886
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127356 36810 127620 36820
rect 127356 35308 127620 35318
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127356 35242 127620 35252
rect 127356 33740 127620 33750
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127356 33674 127620 33684
rect 125132 32722 125188 32732
rect 127356 32172 127620 32182
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127356 32106 127620 32116
rect 127356 30604 127620 30614
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127356 30538 127620 30548
rect 127356 29036 127620 29046
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127356 28970 127620 28980
rect 127356 27468 127620 27478
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127356 27402 127620 27412
rect 127356 25900 127620 25910
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127356 25834 127620 25844
rect 127356 24332 127620 24342
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127356 24266 127620 24276
rect 127356 22764 127620 22774
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127356 22698 127620 22708
rect 127356 21196 127620 21206
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127356 21130 127620 21140
rect 127356 19628 127620 19638
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127356 19562 127620 19572
rect 119756 14466 119812 14476
rect 120092 18228 120148 18238
rect 119532 13972 119588 13982
rect 118636 8930 118692 8942
rect 118636 8878 118638 8930
rect 118690 8878 118692 8930
rect 118636 6468 118692 8878
rect 118748 8260 118804 8270
rect 118748 7700 118804 8204
rect 119196 8036 119252 8046
rect 118748 7606 118804 7644
rect 118860 8034 119252 8036
rect 118860 7982 119198 8034
rect 119250 7982 119252 8034
rect 118860 7980 119252 7982
rect 118636 6402 118692 6412
rect 118636 5684 118692 5694
rect 118636 5590 118692 5628
rect 118524 4340 118580 5516
rect 118748 5012 118804 5022
rect 118860 5012 118916 7980
rect 119196 7970 119252 7980
rect 119420 7364 119476 7374
rect 119308 7362 119476 7364
rect 119308 7310 119422 7362
rect 119474 7310 119476 7362
rect 119308 7308 119476 7310
rect 118748 5010 118916 5012
rect 118748 4958 118750 5010
rect 118802 4958 118916 5010
rect 118748 4956 118916 4958
rect 119084 6020 119140 6030
rect 118748 4676 118804 4956
rect 118748 4610 118804 4620
rect 117964 4174 117966 4226
rect 118018 4174 118020 4226
rect 117964 4162 118020 4174
rect 118300 4284 118580 4340
rect 118300 4004 118356 4284
rect 118412 4116 118468 4126
rect 118412 4022 118468 4060
rect 117852 3948 118356 4004
rect 118076 3668 118132 3678
rect 117628 3444 117684 3482
rect 117628 3378 117684 3388
rect 118076 800 118132 3612
rect 119084 3554 119140 5964
rect 119308 5124 119364 7308
rect 119420 7298 119476 7308
rect 119420 5796 119476 5806
rect 119420 5702 119476 5740
rect 119308 5058 119364 5068
rect 119084 3502 119086 3554
rect 119138 3502 119140 3554
rect 119084 3490 119140 3502
rect 119420 4004 119476 4014
rect 118860 3444 118916 3482
rect 118860 3378 118916 3388
rect 119420 800 119476 3948
rect 119532 3444 119588 13916
rect 119868 7700 119924 7710
rect 119868 7606 119924 7644
rect 119644 5908 119700 5918
rect 119644 5814 119700 5852
rect 119980 5908 120036 5918
rect 120092 5908 120148 18172
rect 127356 18060 127620 18070
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127356 17994 127620 18004
rect 127356 16492 127620 16502
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127356 16426 127620 16436
rect 127356 14924 127620 14934
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127356 14858 127620 14868
rect 131180 14420 131236 55022
rect 136892 27748 136948 55916
rect 139020 55298 139076 55310
rect 139020 55246 139022 55298
rect 139074 55246 139076 55298
rect 138348 55188 138404 55198
rect 138348 55094 138404 55132
rect 139020 55188 139076 55246
rect 139020 55122 139076 55132
rect 139244 55186 139300 56030
rect 142940 56082 142996 56094
rect 142940 56030 142942 56082
rect 142994 56030 142996 56082
rect 142940 55468 142996 56030
rect 139244 55134 139246 55186
rect 139298 55134 139300 55186
rect 139244 55122 139300 55134
rect 142604 55412 142996 55468
rect 146748 55468 146804 56252
rect 150332 56308 150388 59200
rect 150332 56242 150388 56252
rect 151564 56308 151620 56318
rect 151564 56214 151620 56252
rect 154140 56308 154196 59200
rect 154140 56242 154196 56252
rect 155372 56308 155428 56318
rect 155372 56214 155428 56252
rect 150780 56082 150836 56094
rect 150780 56030 150782 56082
rect 150834 56030 150836 56082
rect 147196 55972 147252 55982
rect 147196 55878 147252 55916
rect 149772 55970 149828 55982
rect 149772 55918 149774 55970
rect 149826 55918 149828 55970
rect 146748 55412 146916 55468
rect 136892 27682 136948 27692
rect 142604 55074 142660 55412
rect 146860 55410 146916 55412
rect 146860 55358 146862 55410
rect 146914 55358 146916 55410
rect 146860 55346 146916 55358
rect 149772 55412 149828 55918
rect 149772 55346 149828 55356
rect 150780 55412 150836 56030
rect 154588 56082 154644 56094
rect 154588 56030 154590 56082
rect 154642 56030 154644 56082
rect 154588 55468 154644 56030
rect 158076 55692 158340 55702
rect 158132 55636 158180 55692
rect 158236 55636 158284 55692
rect 158076 55626 158340 55636
rect 150780 55346 150836 55356
rect 154028 55412 154644 55468
rect 142604 55022 142606 55074
rect 142658 55022 142660 55074
rect 142604 16212 142660 55022
rect 154028 55074 154084 55412
rect 154028 55022 154030 55074
rect 154082 55022 154084 55074
rect 142716 54908 142980 54918
rect 142772 54852 142820 54908
rect 142876 54852 142924 54908
rect 142716 54842 142980 54852
rect 142716 53340 142980 53350
rect 142772 53284 142820 53340
rect 142876 53284 142924 53340
rect 142716 53274 142980 53284
rect 142716 51772 142980 51782
rect 142772 51716 142820 51772
rect 142876 51716 142924 51772
rect 142716 51706 142980 51716
rect 142716 50204 142980 50214
rect 142772 50148 142820 50204
rect 142876 50148 142924 50204
rect 142716 50138 142980 50148
rect 142716 48636 142980 48646
rect 142772 48580 142820 48636
rect 142876 48580 142924 48636
rect 142716 48570 142980 48580
rect 142716 47068 142980 47078
rect 142772 47012 142820 47068
rect 142876 47012 142924 47068
rect 142716 47002 142980 47012
rect 142716 45500 142980 45510
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142716 45434 142980 45444
rect 142716 43932 142980 43942
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142716 43866 142980 43876
rect 142716 42364 142980 42374
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142716 42298 142980 42308
rect 142716 40796 142980 40806
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142716 40730 142980 40740
rect 142716 39228 142980 39238
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142716 39162 142980 39172
rect 142716 37660 142980 37670
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142716 37594 142980 37604
rect 142716 36092 142980 36102
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142716 36026 142980 36036
rect 142716 34524 142980 34534
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142716 34458 142980 34468
rect 142716 32956 142980 32966
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142716 32890 142980 32900
rect 142716 31388 142980 31398
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142716 31322 142980 31332
rect 142716 29820 142980 29830
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142716 29754 142980 29764
rect 142716 28252 142980 28262
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142716 28186 142980 28196
rect 142716 26684 142980 26694
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142716 26618 142980 26628
rect 142716 25116 142980 25126
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142716 25050 142980 25060
rect 142716 23548 142980 23558
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142716 23482 142980 23492
rect 142716 21980 142980 21990
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142716 21914 142980 21924
rect 142716 20412 142980 20422
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142716 20346 142980 20356
rect 142716 18844 142980 18854
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142716 18778 142980 18788
rect 142716 17276 142980 17286
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142716 17210 142980 17220
rect 142604 16146 142660 16156
rect 154028 16100 154084 55022
rect 158076 54124 158340 54134
rect 158132 54068 158180 54124
rect 158236 54068 158284 54124
rect 158076 54058 158340 54068
rect 158076 52556 158340 52566
rect 158132 52500 158180 52556
rect 158236 52500 158284 52556
rect 158076 52490 158340 52500
rect 158076 50988 158340 50998
rect 158132 50932 158180 50988
rect 158236 50932 158284 50988
rect 158076 50922 158340 50932
rect 158076 49420 158340 49430
rect 158132 49364 158180 49420
rect 158236 49364 158284 49420
rect 158076 49354 158340 49364
rect 158076 47852 158340 47862
rect 158132 47796 158180 47852
rect 158236 47796 158284 47852
rect 158076 47786 158340 47796
rect 158076 46284 158340 46294
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158076 46218 158340 46228
rect 158076 44716 158340 44726
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158076 44650 158340 44660
rect 158076 43148 158340 43158
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158076 43082 158340 43092
rect 158076 41580 158340 41590
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158076 41514 158340 41524
rect 158076 40012 158340 40022
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158076 39946 158340 39956
rect 158076 38444 158340 38454
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158076 38378 158340 38388
rect 158076 36876 158340 36886
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158076 36810 158340 36820
rect 158076 35308 158340 35318
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158076 35242 158340 35252
rect 158076 33740 158340 33750
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158076 33674 158340 33684
rect 158076 32172 158340 32182
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158076 32106 158340 32116
rect 158076 30604 158340 30614
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158076 30538 158340 30548
rect 158076 29036 158340 29046
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158076 28970 158340 28980
rect 158076 27468 158340 27478
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158076 27402 158340 27412
rect 158076 25900 158340 25910
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158076 25834 158340 25844
rect 158076 24332 158340 24342
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158076 24266 158340 24276
rect 158076 22764 158340 22774
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158076 22698 158340 22708
rect 158076 21196 158340 21206
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158076 21130 158340 21140
rect 158076 19628 158340 19638
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158076 19562 158340 19572
rect 158076 18060 158340 18070
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158076 17994 158340 18004
rect 158076 16492 158340 16502
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158076 16426 158340 16436
rect 154028 16034 154084 16044
rect 142716 15708 142980 15718
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142716 15642 142980 15652
rect 158076 14924 158340 14934
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158076 14858 158340 14868
rect 131180 14354 131236 14364
rect 142716 14140 142980 14150
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142716 14074 142980 14084
rect 127356 13356 127620 13366
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127356 13290 127620 13300
rect 158076 13356 158340 13366
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158076 13290 158340 13300
rect 121772 12852 121828 12862
rect 121772 8372 121828 12796
rect 142716 12572 142980 12582
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142716 12506 142980 12516
rect 145516 12068 145572 12078
rect 122668 11956 122724 11966
rect 122668 9268 122724 11900
rect 127356 11788 127620 11798
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127356 11722 127620 11732
rect 142716 11004 142980 11014
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142716 10938 142980 10948
rect 127356 10220 127620 10230
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127356 10154 127620 10164
rect 142716 9436 142980 9446
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142716 9370 142980 9380
rect 122668 9202 122724 9212
rect 137900 9268 137956 9278
rect 121772 8306 121828 8316
rect 126476 9156 126532 9166
rect 121324 7812 121380 7822
rect 120316 7588 120372 7598
rect 120316 7494 120372 7532
rect 119980 5906 120148 5908
rect 119980 5854 119982 5906
rect 120034 5854 120148 5906
rect 119980 5852 120148 5854
rect 120316 6578 120372 6590
rect 120316 6526 120318 6578
rect 120370 6526 120372 6578
rect 119980 5842 120036 5852
rect 120316 5460 120372 6526
rect 120876 6466 120932 6478
rect 120876 6414 120878 6466
rect 120930 6414 120932 6466
rect 120316 5394 120372 5404
rect 120652 5906 120708 5918
rect 120652 5854 120654 5906
rect 120706 5854 120708 5906
rect 120540 5236 120596 5246
rect 119756 5234 120596 5236
rect 119756 5182 120542 5234
rect 120594 5182 120596 5234
rect 119756 5180 120596 5182
rect 119756 4450 119812 5180
rect 120540 5170 120596 5180
rect 119756 4398 119758 4450
rect 119810 4398 119812 4450
rect 119756 4386 119812 4398
rect 119756 4116 119812 4126
rect 119756 3554 119812 4060
rect 119756 3502 119758 3554
rect 119810 3502 119812 3554
rect 119756 3490 119812 3502
rect 120652 3556 120708 5854
rect 120764 4228 120820 4238
rect 120764 4134 120820 4172
rect 120652 3490 120708 3500
rect 119532 3378 119588 3388
rect 120764 3444 120820 3454
rect 120764 800 120820 3388
rect 120876 2884 120932 6414
rect 121212 6018 121268 6030
rect 121212 5966 121214 6018
rect 121266 5966 121268 6018
rect 120988 5906 121044 5918
rect 120988 5854 120990 5906
rect 121042 5854 121044 5906
rect 120988 5236 121044 5854
rect 121100 5236 121156 5246
rect 120988 5234 121156 5236
rect 120988 5182 121102 5234
rect 121154 5182 121156 5234
rect 120988 5180 121156 5182
rect 121100 5170 121156 5180
rect 121100 4450 121156 4462
rect 121100 4398 121102 4450
rect 121154 4398 121156 4450
rect 121100 4228 121156 4398
rect 121212 4452 121268 5966
rect 121212 4386 121268 4396
rect 121324 4228 121380 7756
rect 122668 7476 122724 7486
rect 121660 6466 121716 6478
rect 121660 6414 121662 6466
rect 121714 6414 121716 6466
rect 121660 6020 121716 6414
rect 122556 6466 122612 6478
rect 122556 6414 122558 6466
rect 122610 6414 122612 6466
rect 121660 5964 122388 6020
rect 121660 5794 121716 5806
rect 122220 5796 122276 5806
rect 121660 5742 121662 5794
rect 121714 5742 121716 5794
rect 121660 5572 121716 5742
rect 121660 5506 121716 5516
rect 121772 5794 122276 5796
rect 121772 5742 122222 5794
rect 122274 5742 122276 5794
rect 121772 5740 122276 5742
rect 121772 5012 121828 5740
rect 122220 5730 122276 5740
rect 121436 4956 121828 5012
rect 122108 5012 122164 5022
rect 122332 5012 122388 5964
rect 122108 5010 122388 5012
rect 122108 4958 122110 5010
rect 122162 4958 122388 5010
rect 122108 4956 122388 4958
rect 121436 4450 121492 4956
rect 121436 4398 121438 4450
rect 121490 4398 121492 4450
rect 121436 4386 121492 4398
rect 121100 4172 121380 4228
rect 121884 4226 121940 4238
rect 121884 4174 121886 4226
rect 121938 4174 121940 4226
rect 121884 3780 121940 4174
rect 122108 4004 122164 4956
rect 122556 4676 122612 6414
rect 122108 3938 122164 3948
rect 122332 4226 122388 4238
rect 122332 4174 122334 4226
rect 122386 4174 122388 4226
rect 122332 3892 122388 4174
rect 122332 3826 122388 3836
rect 121884 3714 121940 3724
rect 120988 3668 121044 3678
rect 120988 3574 121044 3612
rect 122108 3668 122164 3678
rect 120876 2818 120932 2828
rect 122108 800 122164 3612
rect 122556 3444 122612 4620
rect 122556 3378 122612 3388
rect 122668 3442 122724 7420
rect 123788 6466 123844 6478
rect 123788 6414 123790 6466
rect 123842 6414 123844 6466
rect 123228 6018 123284 6030
rect 123228 5966 123230 6018
rect 123282 5966 123284 6018
rect 122892 5460 122948 5470
rect 122892 4562 122948 5404
rect 123228 5234 123284 5966
rect 123788 5908 123844 6414
rect 125804 6466 125860 6478
rect 125804 6414 125806 6466
rect 125858 6414 125860 6466
rect 125804 6244 125860 6414
rect 125468 6188 125860 6244
rect 124348 6020 124404 6030
rect 124348 6018 124964 6020
rect 124348 5966 124350 6018
rect 124402 5966 124964 6018
rect 124348 5964 124964 5966
rect 124348 5954 124404 5964
rect 124012 5908 124068 5918
rect 123788 5906 124068 5908
rect 123788 5854 124014 5906
rect 124066 5854 124068 5906
rect 123788 5852 124068 5854
rect 123228 5182 123230 5234
rect 123282 5182 123284 5234
rect 123228 5170 123284 5182
rect 122892 4510 122894 4562
rect 122946 4510 122948 4562
rect 122892 4498 122948 4510
rect 122780 4452 122836 4462
rect 122780 4358 122836 4396
rect 122892 4228 122948 4238
rect 122892 3554 122948 4172
rect 124012 4116 124068 5852
rect 124796 5012 124852 5022
rect 124572 4452 124628 4462
rect 124572 4338 124628 4396
rect 124572 4286 124574 4338
rect 124626 4286 124628 4338
rect 124572 4274 124628 4286
rect 122892 3502 122894 3554
rect 122946 3502 122948 3554
rect 122892 3490 122948 3502
rect 123452 4060 124068 4116
rect 122668 3390 122670 3442
rect 122722 3390 122724 3442
rect 122668 3378 122724 3390
rect 123452 800 123508 4060
rect 124572 3668 124628 3678
rect 124572 3574 124628 3612
rect 123564 3556 123620 3566
rect 123564 3462 123620 3500
rect 124796 800 124852 4956
rect 124908 4338 124964 5964
rect 125244 5010 125300 5022
rect 125244 4958 125246 5010
rect 125298 4958 125300 5010
rect 125244 4676 125300 4958
rect 125468 5012 125524 6188
rect 125580 6018 125636 6030
rect 125580 5966 125582 6018
rect 125634 5966 125636 6018
rect 125580 5460 125636 5966
rect 125580 5404 125972 5460
rect 125916 5346 125972 5404
rect 125916 5294 125918 5346
rect 125970 5294 125972 5346
rect 125916 5282 125972 5294
rect 125580 5012 125636 5022
rect 125468 4956 125580 5012
rect 125580 4946 125636 4956
rect 125244 4610 125300 4620
rect 126140 4564 126196 4574
rect 126028 4452 126084 4462
rect 126140 4452 126196 4508
rect 126028 4450 126196 4452
rect 126028 4398 126030 4450
rect 126082 4398 126196 4450
rect 126028 4396 126196 4398
rect 126028 4386 126084 4396
rect 124908 4286 124910 4338
rect 124962 4286 124964 4338
rect 124908 4274 124964 4286
rect 126140 3668 126196 3678
rect 126140 800 126196 3612
rect 126476 3442 126532 9100
rect 127356 8652 127620 8662
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127356 8586 127620 8596
rect 128828 8372 128884 8382
rect 127356 7084 127620 7094
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127356 7018 127620 7028
rect 126588 5794 126644 5806
rect 126588 5742 126590 5794
rect 126642 5742 126644 5794
rect 126588 3556 126644 5742
rect 127708 5794 127764 5806
rect 127708 5742 127710 5794
rect 127762 5742 127764 5794
rect 127148 5684 127204 5694
rect 126700 3556 126756 3566
rect 126588 3554 126756 3556
rect 126588 3502 126702 3554
rect 126754 3502 126756 3554
rect 126588 3500 126756 3502
rect 127148 3556 127204 5628
rect 127356 5516 127620 5526
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127356 5450 127620 5460
rect 127708 4564 127764 5742
rect 128044 5012 128100 5022
rect 128044 4918 128100 4956
rect 128828 5010 128884 8316
rect 134092 6468 134148 6478
rect 128828 4958 128830 5010
rect 128882 4958 128884 5010
rect 128828 4946 128884 4958
rect 129164 5122 129220 5134
rect 129164 5070 129166 5122
rect 129218 5070 129220 5122
rect 127708 4508 127988 4564
rect 127260 4452 127316 4462
rect 127260 4358 127316 4396
rect 127932 4452 127988 4508
rect 127596 4340 127652 4350
rect 127820 4340 127876 4350
rect 127596 4338 127876 4340
rect 127596 4286 127598 4338
rect 127650 4286 127822 4338
rect 127874 4286 127876 4338
rect 127596 4284 127876 4286
rect 127596 4274 127652 4284
rect 127820 4274 127876 4284
rect 127356 3948 127620 3958
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127356 3882 127620 3892
rect 127372 3556 127428 3566
rect 127148 3554 127428 3556
rect 127148 3502 127374 3554
rect 127426 3502 127428 3554
rect 127148 3500 127428 3502
rect 126700 3490 126756 3500
rect 127372 3490 127428 3500
rect 127932 3444 127988 4396
rect 129164 4228 129220 5070
rect 132300 5122 132356 5134
rect 132300 5070 132302 5122
rect 132354 5070 132356 5122
rect 131180 4788 131236 4798
rect 129948 4452 130004 4462
rect 129948 4358 130004 4396
rect 129164 4162 129220 4172
rect 130732 4228 130788 4238
rect 130732 4134 130788 4172
rect 128380 3668 128436 3678
rect 128380 3574 128436 3612
rect 126476 3390 126478 3442
rect 126530 3390 126532 3442
rect 126476 3378 126532 3390
rect 127484 3388 127988 3444
rect 128828 3556 128884 3566
rect 127484 800 127540 3388
rect 128828 800 128884 3500
rect 130396 3556 130452 3566
rect 130396 3462 130452 3500
rect 131180 3554 131236 4732
rect 131740 4450 131796 4462
rect 131740 4398 131742 4450
rect 131794 4398 131796 4450
rect 131180 3502 131182 3554
rect 131234 3502 131236 3554
rect 131180 3490 131236 3502
rect 131516 4340 131572 4350
rect 130172 3444 130228 3454
rect 130172 800 130228 3388
rect 131516 800 131572 4284
rect 131740 3556 131796 4398
rect 132300 4340 132356 5070
rect 133868 5012 133924 5022
rect 133532 5010 133924 5012
rect 133532 4958 133870 5010
rect 133922 4958 133924 5010
rect 133532 4956 133924 4958
rect 133532 4898 133588 4956
rect 133868 4946 133924 4956
rect 133532 4846 133534 4898
rect 133586 4846 133588 4898
rect 132524 4564 132580 4574
rect 132524 4470 132580 4508
rect 132300 4274 132356 4284
rect 132748 4340 132804 4350
rect 132748 4246 132804 4284
rect 131740 3490 131796 3500
rect 132748 3444 132804 3454
rect 132748 3350 132804 3388
rect 132860 924 133140 980
rect 132860 800 132916 924
rect 99596 700 100100 756
rect 100576 0 100688 800
rect 101920 0 102032 800
rect 103264 0 103376 800
rect 104608 0 104720 800
rect 105952 0 106064 800
rect 107296 0 107408 800
rect 108640 0 108752 800
rect 109984 0 110096 800
rect 111328 0 111440 800
rect 112672 0 112784 800
rect 114016 0 114128 800
rect 115360 0 115472 800
rect 116704 0 116816 800
rect 118048 0 118160 800
rect 119392 0 119504 800
rect 120736 0 120848 800
rect 122080 0 122192 800
rect 123424 0 123536 800
rect 124768 0 124880 800
rect 126112 0 126224 800
rect 127456 0 127568 800
rect 128800 0 128912 800
rect 130144 0 130256 800
rect 131488 0 131600 800
rect 132832 0 132944 800
rect 133084 756 133140 924
rect 133532 756 133588 4846
rect 134092 3442 134148 6412
rect 136220 5348 136276 5358
rect 134988 5236 135044 5246
rect 134316 5234 135044 5236
rect 134316 5182 134990 5234
rect 135042 5182 135044 5234
rect 134316 5180 135044 5182
rect 134092 3390 134094 3442
rect 134146 3390 134148 3442
rect 134092 3378 134148 3390
rect 134204 3668 134260 3678
rect 134204 800 134260 3612
rect 134316 3554 134372 5180
rect 134988 5170 135044 5180
rect 135772 5124 135828 5134
rect 135772 4450 135828 5068
rect 135772 4398 135774 4450
rect 135826 4398 135828 4450
rect 135772 4386 135828 4398
rect 135996 4898 136052 4910
rect 135996 4846 135998 4898
rect 136050 4846 136052 4898
rect 135548 4338 135604 4350
rect 135548 4286 135550 4338
rect 135602 4286 135604 4338
rect 135100 4228 135156 4238
rect 134316 3502 134318 3554
rect 134370 3502 134372 3554
rect 134316 3490 134372 3502
rect 134988 4226 135156 4228
rect 134988 4174 135102 4226
rect 135154 4174 135156 4226
rect 134988 4172 135156 4174
rect 134988 3554 135044 4172
rect 135100 4162 135156 4172
rect 135548 4228 135604 4286
rect 135996 4228 136052 4846
rect 136220 4450 136276 5292
rect 137340 5236 137396 5246
rect 136220 4398 136222 4450
rect 136274 4398 136276 4450
rect 136220 4386 136276 4398
rect 136892 4452 136948 4462
rect 135548 4172 136052 4228
rect 134988 3502 134990 3554
rect 135042 3502 135044 3554
rect 134988 2996 135044 3502
rect 134988 2930 135044 2940
rect 135548 800 135604 4172
rect 136108 3668 136164 3678
rect 136108 3574 136164 3612
rect 136892 800 136948 4396
rect 137340 4338 137396 5180
rect 137452 5122 137508 5134
rect 137452 5070 137454 5122
rect 137506 5070 137508 5122
rect 137452 4452 137508 5070
rect 137676 4452 137732 4462
rect 137788 4452 137844 4462
rect 137452 4396 137676 4452
rect 137732 4450 137844 4452
rect 137732 4398 137790 4450
rect 137842 4398 137844 4450
rect 137732 4396 137844 4398
rect 137676 4386 137732 4396
rect 137788 4386 137844 4396
rect 137340 4286 137342 4338
rect 137394 4286 137396 4338
rect 137340 4274 137396 4286
rect 137900 3442 137956 9212
rect 142716 7868 142980 7878
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142716 7802 142980 7812
rect 141036 7700 141092 7710
rect 138908 5794 138964 5806
rect 138908 5742 138910 5794
rect 138962 5742 138964 5794
rect 138908 5460 138964 5742
rect 138908 5394 138964 5404
rect 139020 5682 139076 5694
rect 139020 5630 139022 5682
rect 139074 5630 139076 5682
rect 138236 5124 138292 5134
rect 138236 5030 138292 5068
rect 138348 4900 138404 4910
rect 138348 4806 138404 4844
rect 139020 4340 139076 5630
rect 140140 5236 140196 5246
rect 140140 5142 140196 5180
rect 139020 4274 139076 4284
rect 138908 4228 138964 4238
rect 139580 4228 139636 4238
rect 138236 4226 138964 4228
rect 138236 4174 138910 4226
rect 138962 4174 138964 4226
rect 138236 4172 138964 4174
rect 138236 3554 138292 4172
rect 138908 4162 138964 4172
rect 139244 4226 139636 4228
rect 139244 4174 139582 4226
rect 139634 4174 139636 4226
rect 139244 4172 139636 4174
rect 138236 3502 138238 3554
rect 138290 3502 138292 3554
rect 138236 3490 138292 3502
rect 138348 3668 138404 3678
rect 137900 3390 137902 3442
rect 137954 3390 137956 3442
rect 137900 3378 137956 3390
rect 138348 980 138404 3612
rect 139244 3556 139300 4172
rect 139580 4162 139636 4172
rect 140924 3780 140980 3790
rect 139804 3668 139860 3678
rect 139804 3574 139860 3612
rect 139244 3462 139300 3500
rect 139580 3556 139636 3566
rect 138236 924 138404 980
rect 138236 800 138292 924
rect 139580 800 139636 3500
rect 140924 800 140980 3724
rect 141036 3444 141092 7644
rect 142716 6300 142980 6310
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142716 6234 142980 6244
rect 143836 5794 143892 5806
rect 143836 5742 143838 5794
rect 143890 5742 143892 5794
rect 142940 5460 142996 5470
rect 142996 5404 143108 5460
rect 142940 5394 142996 5404
rect 142044 5348 142100 5358
rect 141708 5124 141764 5134
rect 141372 5010 141428 5022
rect 141372 4958 141374 5010
rect 141426 4958 141428 5010
rect 141372 4450 141428 4958
rect 141372 4398 141374 4450
rect 141426 4398 141428 4450
rect 141372 4386 141428 4398
rect 141484 4900 141540 4910
rect 141484 4338 141540 4844
rect 141484 4286 141486 4338
rect 141538 4286 141540 4338
rect 141484 4274 141540 4286
rect 141708 4338 141764 5068
rect 141708 4286 141710 4338
rect 141762 4286 141764 4338
rect 141708 4274 141764 4286
rect 141932 4340 141988 4350
rect 141932 4246 141988 4284
rect 142044 4338 142100 5292
rect 142044 4286 142046 4338
rect 142098 4286 142100 4338
rect 142044 4274 142100 4286
rect 142156 5236 142212 5246
rect 142044 3556 142100 3566
rect 142156 3556 142212 5180
rect 142940 5236 142996 5246
rect 142940 5142 142996 5180
rect 142716 5122 142772 5134
rect 142716 5070 142718 5122
rect 142770 5070 142772 5122
rect 142716 4900 142772 5070
rect 142492 4844 142716 4900
rect 142492 3780 142548 4844
rect 142716 4834 142772 4844
rect 142716 4732 142980 4742
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142716 4666 142980 4676
rect 142828 4564 142884 4574
rect 143052 4564 143108 5404
rect 142828 4562 143108 4564
rect 142828 4510 142830 4562
rect 142882 4510 143108 4562
rect 142828 4508 143108 4510
rect 142828 4498 142884 4508
rect 143052 4340 143108 4350
rect 142492 3714 142548 3724
rect 142604 4228 142660 4238
rect 142044 3554 142212 3556
rect 142044 3502 142046 3554
rect 142098 3502 142212 3554
rect 142044 3500 142212 3502
rect 142268 3668 142324 3678
rect 142044 3490 142100 3500
rect 141036 3378 141092 3388
rect 141708 3444 141764 3454
rect 141708 3350 141764 3388
rect 142268 800 142324 3612
rect 142604 3556 142660 4172
rect 142380 3554 142660 3556
rect 142380 3502 142606 3554
rect 142658 3502 142660 3554
rect 142380 3500 142660 3502
rect 142380 3108 142436 3500
rect 142604 3490 142660 3500
rect 143052 3556 143108 4284
rect 143612 4228 143668 4238
rect 143612 4134 143668 4172
rect 143612 3668 143668 3678
rect 143612 3574 143668 3612
rect 143052 3490 143108 3500
rect 143836 3444 143892 5742
rect 144172 5796 144228 5806
rect 144172 5794 144340 5796
rect 144172 5742 144174 5794
rect 144226 5742 144340 5794
rect 144172 5740 144340 5742
rect 144172 5730 144228 5740
rect 143948 5010 144004 5022
rect 143948 4958 143950 5010
rect 144002 4958 144004 5010
rect 143948 4900 144004 4958
rect 143948 4834 144004 4844
rect 144172 4450 144228 4462
rect 144172 4398 144174 4450
rect 144226 4398 144228 4450
rect 144172 3444 144228 4398
rect 144284 4340 144340 5740
rect 144732 5124 144788 5134
rect 144732 5010 144788 5068
rect 144732 4958 144734 5010
rect 144786 4958 144788 5010
rect 144732 4946 144788 4958
rect 145068 5010 145124 5022
rect 145068 4958 145070 5010
rect 145122 4958 145124 5010
rect 144284 4274 144340 4284
rect 143612 3388 144228 3444
rect 144956 4228 145012 4238
rect 145068 4228 145124 4958
rect 145292 4228 145348 4238
rect 145068 4226 145348 4228
rect 145068 4174 145294 4226
rect 145346 4174 145348 4226
rect 145068 4172 145348 4174
rect 142716 3164 142980 3174
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142716 3098 142980 3108
rect 142380 3042 142436 3052
rect 143612 800 143668 3388
rect 144956 800 145012 4172
rect 145292 4162 145348 4172
rect 145516 3442 145572 12012
rect 158076 11788 158340 11798
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158076 11722 158340 11732
rect 158076 10220 158340 10230
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158076 10154 158340 10164
rect 158076 8652 158340 8662
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158076 8586 158340 8596
rect 158076 7084 158340 7094
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158076 7018 158340 7028
rect 158076 5516 158340 5526
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158076 5450 158340 5460
rect 147868 5348 147924 5358
rect 147644 5124 147700 5134
rect 146188 4226 146244 4238
rect 146188 4174 146190 4226
rect 146242 4174 146244 4226
rect 146188 3668 146244 4174
rect 147532 4228 147588 4238
rect 147532 4134 147588 4172
rect 145964 3612 146580 3668
rect 145852 3556 145908 3566
rect 145852 3462 145908 3500
rect 145516 3390 145518 3442
rect 145570 3390 145572 3442
rect 145516 3378 145572 3390
rect 145964 2772 146020 3612
rect 146524 3554 146580 3612
rect 146524 3502 146526 3554
rect 146578 3502 146580 3554
rect 146524 3490 146580 3502
rect 145964 2706 146020 2716
rect 146300 3444 146356 3454
rect 146300 800 146356 3388
rect 147532 3444 147588 3454
rect 147532 3330 147588 3388
rect 147532 3278 147534 3330
rect 147586 3278 147588 3330
rect 147532 3266 147588 3278
rect 147644 800 147700 5068
rect 147868 4898 147924 5292
rect 150668 5236 150724 5246
rect 149996 5234 150724 5236
rect 149996 5182 150670 5234
rect 150722 5182 150724 5234
rect 149996 5180 150724 5182
rect 148092 5124 148148 5134
rect 148092 5030 148148 5068
rect 149212 5122 149268 5134
rect 149212 5070 149214 5122
rect 149266 5070 149268 5122
rect 149212 5012 149268 5070
rect 149548 5012 149604 5022
rect 147868 4846 147870 4898
rect 147922 4846 147924 4898
rect 147868 4834 147924 4846
rect 148988 5010 149604 5012
rect 148988 4958 149550 5010
rect 149602 4958 149604 5010
rect 148988 4956 149604 4958
rect 148876 4450 148932 4462
rect 148876 4398 148878 4450
rect 148930 4398 148932 4450
rect 147868 4228 147924 4238
rect 147756 4226 147924 4228
rect 147756 4174 147870 4226
rect 147922 4174 147924 4226
rect 147756 4172 147924 4174
rect 147756 3556 147812 4172
rect 147868 4162 147924 4172
rect 148876 4228 148932 4398
rect 148876 4162 148932 4172
rect 147756 3490 147812 3500
rect 148988 800 149044 4956
rect 149548 4946 149604 4956
rect 149772 5012 149828 5022
rect 149660 4450 149716 4462
rect 149660 4398 149662 4450
rect 149714 4398 149716 4450
rect 149660 1652 149716 4398
rect 149772 3666 149828 4956
rect 149996 4562 150052 5180
rect 150668 5170 150724 5180
rect 149996 4510 149998 4562
rect 150050 4510 150052 4562
rect 149996 4498 150052 4510
rect 158076 3948 158340 3958
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158076 3882 158340 3892
rect 149772 3614 149774 3666
rect 149826 3614 149828 3666
rect 149772 3556 149828 3614
rect 149772 3490 149828 3500
rect 150332 3668 150388 3678
rect 149660 1586 149716 1596
rect 150332 800 150388 3612
rect 151564 3668 151620 3678
rect 151564 3574 151620 3612
rect 150556 3556 150612 3566
rect 150556 3462 150612 3500
rect 133084 700 133588 756
rect 134176 0 134288 800
rect 135520 0 135632 800
rect 136864 0 136976 800
rect 138208 0 138320 800
rect 139552 0 139664 800
rect 140896 0 141008 800
rect 142240 0 142352 800
rect 143584 0 143696 800
rect 144928 0 145040 800
rect 146272 0 146384 800
rect 147616 0 147728 800
rect 148960 0 149072 800
rect 150304 0 150416 800
<< via2 >>
rect 6188 56194 6244 56196
rect 6188 56142 6190 56194
rect 6190 56142 6242 56194
rect 6242 56142 6244 56194
rect 6188 56140 6244 56142
rect 9212 56140 9268 56196
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 28476 56252 28532 56308
rect 29708 56306 29764 56308
rect 29708 56254 29710 56306
rect 29710 56254 29762 56306
rect 29762 56254 29764 56306
rect 29708 56252 29764 56254
rect 19852 55916 19908 55972
rect 20972 55970 21028 55972
rect 20972 55918 20974 55970
rect 20974 55918 21026 55970
rect 21026 55918 21028 55970
rect 20972 55916 21028 55918
rect 27916 55916 27972 55972
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 51324 56252 51380 56308
rect 52556 56306 52612 56308
rect 52556 56254 52558 56306
rect 52558 56254 52610 56306
rect 52610 56254 52612 56306
rect 52556 56252 52612 56254
rect 50092 56028 50148 56084
rect 42700 55916 42756 55972
rect 43820 55970 43876 55972
rect 43820 55918 43822 55970
rect 43822 55918 43874 55970
rect 43874 55918 43876 55970
rect 43820 55916 43876 55918
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 26908 27692 26964 27748
rect 24444 26796 24500 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 25788 26796 25844 26852
rect 25340 26572 25396 26628
rect 23436 25506 23492 25508
rect 23436 25454 23438 25506
rect 23438 25454 23490 25506
rect 23490 25454 23492 25506
rect 23436 25452 23492 25454
rect 24780 26290 24836 26292
rect 24780 26238 24782 26290
rect 24782 26238 24834 26290
rect 24834 26238 24836 26290
rect 24780 26236 24836 26238
rect 26348 26850 26404 26852
rect 26348 26798 26350 26850
rect 26350 26798 26402 26850
rect 26402 26798 26404 26850
rect 26348 26796 26404 26798
rect 26684 26572 26740 26628
rect 26012 26514 26068 26516
rect 26012 26462 26014 26514
rect 26014 26462 26066 26514
rect 26066 26462 26068 26514
rect 26012 26460 26068 26462
rect 25564 26290 25620 26292
rect 25564 26238 25566 26290
rect 25566 26238 25618 26290
rect 25618 26238 25620 26290
rect 25564 26236 25620 26238
rect 24556 25452 24612 25508
rect 23436 25228 23492 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 27020 26572 27076 26628
rect 27132 26514 27188 26516
rect 27132 26462 27134 26514
rect 27134 26462 27186 26514
rect 27186 26462 27188 26514
rect 27132 26460 27188 26462
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 21084 21756 21140 21812
rect 22540 23042 22596 23044
rect 22540 22990 22542 23042
rect 22542 22990 22594 23042
rect 22594 22990 22596 23042
rect 22540 22988 22596 22990
rect 23324 22988 23380 23044
rect 21868 21756 21924 21812
rect 21868 21474 21924 21476
rect 21868 21422 21870 21474
rect 21870 21422 21922 21474
rect 21922 21422 21924 21474
rect 21868 21420 21924 21422
rect 21980 20860 22036 20916
rect 23324 21420 23380 21476
rect 23772 22876 23828 22932
rect 23660 22258 23716 22260
rect 23660 22206 23662 22258
rect 23662 22206 23714 22258
rect 23714 22206 23716 22258
rect 23660 22204 23716 22206
rect 23884 22258 23940 22260
rect 23884 22206 23886 22258
rect 23886 22206 23938 22258
rect 23938 22206 23940 22258
rect 23884 22204 23940 22206
rect 26908 24556 26964 24612
rect 24668 23324 24724 23380
rect 25340 23378 25396 23380
rect 25340 23326 25342 23378
rect 25342 23326 25394 23378
rect 25394 23326 25396 23378
rect 25340 23324 25396 23326
rect 25340 22930 25396 22932
rect 25340 22878 25342 22930
rect 25342 22878 25394 22930
rect 25394 22878 25396 22930
rect 25340 22876 25396 22878
rect 25452 22316 25508 22372
rect 24780 22204 24836 22260
rect 23996 21644 24052 21700
rect 23996 21308 24052 21364
rect 23884 21196 23940 21252
rect 24444 21308 24500 21364
rect 23660 20972 23716 21028
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 21980 20188 22036 20244
rect 19852 19906 19908 19908
rect 19852 19854 19854 19906
rect 19854 19854 19906 19906
rect 19906 19854 19908 19906
rect 19852 19852 19908 19854
rect 24220 21196 24276 21252
rect 23324 20188 23380 20244
rect 23884 20300 23940 20356
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19180 18508 19236 18564
rect 21532 18508 21588 18564
rect 22764 19852 22820 19908
rect 23436 19180 23492 19236
rect 22876 18620 22932 18676
rect 22428 18508 22484 18564
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 9212 17052 9268 17108
rect 19628 17106 19684 17108
rect 19628 17054 19630 17106
rect 19630 17054 19682 17106
rect 19682 17054 19684 17106
rect 19628 17052 19684 17054
rect 20188 17052 20244 17108
rect 19292 16716 19348 16772
rect 20300 16770 20356 16772
rect 20300 16718 20302 16770
rect 20302 16718 20354 16770
rect 20354 16718 20356 16770
rect 20300 16716 20356 16718
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 17948 16098 18004 16100
rect 17948 16046 17950 16098
rect 17950 16046 18002 16098
rect 18002 16046 18004 16098
rect 17948 16044 18004 16046
rect 9212 15932 9268 15988
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 18620 15484 18676 15540
rect 19628 15260 19684 15316
rect 17164 14252 17220 14308
rect 17836 13020 17892 13076
rect 19068 13468 19124 13524
rect 18620 12684 18676 12740
rect 15596 12348 15652 12404
rect 18172 12402 18228 12404
rect 18172 12350 18174 12402
rect 18174 12350 18226 12402
rect 18226 12350 18228 12402
rect 18172 12348 18228 12350
rect 20748 16210 20804 16212
rect 20748 16158 20750 16210
rect 20750 16158 20802 16210
rect 20802 16158 20804 16210
rect 20748 16156 20804 16158
rect 20412 16044 20468 16100
rect 22764 17666 22820 17668
rect 22764 17614 22766 17666
rect 22766 17614 22818 17666
rect 22818 17614 22820 17666
rect 22764 17612 22820 17614
rect 23996 20188 24052 20244
rect 23884 19234 23940 19236
rect 23884 19182 23886 19234
rect 23886 19182 23938 19234
rect 23938 19182 23940 19234
rect 23884 19180 23940 19182
rect 23324 17836 23380 17892
rect 23772 17836 23828 17892
rect 23548 17724 23604 17780
rect 24108 17666 24164 17668
rect 24108 17614 24110 17666
rect 24110 17614 24162 17666
rect 24162 17614 24164 17666
rect 24108 17612 24164 17614
rect 22652 17164 22708 17220
rect 21644 16994 21700 16996
rect 21644 16942 21646 16994
rect 21646 16942 21698 16994
rect 21698 16942 21700 16994
rect 21644 16940 21700 16942
rect 21644 16098 21700 16100
rect 21644 16046 21646 16098
rect 21646 16046 21698 16098
rect 21698 16046 21700 16098
rect 21644 16044 21700 16046
rect 20748 15538 20804 15540
rect 20748 15486 20750 15538
rect 20750 15486 20802 15538
rect 20802 15486 20804 15538
rect 20748 15484 20804 15486
rect 20972 15484 21028 15540
rect 20636 15314 20692 15316
rect 20636 15262 20638 15314
rect 20638 15262 20690 15314
rect 20690 15262 20692 15314
rect 20636 15260 20692 15262
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20412 14306 20468 14308
rect 20412 14254 20414 14306
rect 20414 14254 20466 14306
rect 20466 14254 20468 14306
rect 20412 14252 20468 14254
rect 20076 13916 20132 13972
rect 19740 13468 19796 13524
rect 20076 13244 20132 13300
rect 19852 13074 19908 13076
rect 19852 13022 19854 13074
rect 19854 13022 19906 13074
rect 19906 13022 19908 13074
rect 19852 13020 19908 13022
rect 17724 12124 17780 12180
rect 18172 11116 18228 11172
rect 16940 10668 16996 10724
rect 15932 7756 15988 7812
rect 17500 10610 17556 10612
rect 17500 10558 17502 10610
rect 17502 10558 17554 10610
rect 17554 10558 17556 10610
rect 17500 10556 17556 10558
rect 18956 12402 19012 12404
rect 18956 12350 18958 12402
rect 18958 12350 19010 12402
rect 19010 12350 19012 12402
rect 18956 12348 19012 12350
rect 20412 13522 20468 13524
rect 20412 13470 20414 13522
rect 20414 13470 20466 13522
rect 20466 13470 20468 13522
rect 20412 13468 20468 13470
rect 19628 12684 19684 12740
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19628 12178 19684 12180
rect 19628 12126 19630 12178
rect 19630 12126 19682 12178
rect 19682 12126 19684 12178
rect 19628 12124 19684 12126
rect 18956 12066 19012 12068
rect 18956 12014 18958 12066
rect 18958 12014 19010 12066
rect 19010 12014 19012 12066
rect 18956 12012 19012 12014
rect 19180 11954 19236 11956
rect 19180 11902 19182 11954
rect 19182 11902 19234 11954
rect 19234 11902 19236 11954
rect 19180 11900 19236 11902
rect 18956 11228 19012 11284
rect 19740 11676 19796 11732
rect 19404 11282 19460 11284
rect 19404 11230 19406 11282
rect 19406 11230 19458 11282
rect 19458 11230 19460 11282
rect 19404 11228 19460 11230
rect 18508 10556 18564 10612
rect 19964 12066 20020 12068
rect 19964 12014 19966 12066
rect 19966 12014 20018 12066
rect 20018 12014 20020 12066
rect 19964 12012 20020 12014
rect 20076 11452 20132 11508
rect 20300 11618 20356 11620
rect 20300 11566 20302 11618
rect 20302 11566 20354 11618
rect 20354 11566 20356 11618
rect 20300 11564 20356 11566
rect 20524 11394 20580 11396
rect 20524 11342 20526 11394
rect 20526 11342 20578 11394
rect 20578 11342 20580 11394
rect 20524 11340 20580 11342
rect 20188 11170 20244 11172
rect 20188 11118 20190 11170
rect 20190 11118 20242 11170
rect 20242 11118 20244 11170
rect 20188 11116 20244 11118
rect 18844 9938 18900 9940
rect 18844 9886 18846 9938
rect 18846 9886 18898 9938
rect 18898 9886 18900 9938
rect 18844 9884 18900 9886
rect 16940 7756 16996 7812
rect 18060 8146 18116 8148
rect 18060 8094 18062 8146
rect 18062 8094 18114 8146
rect 18114 8094 18116 8146
rect 18060 8092 18116 8094
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 20300 11004 20356 11060
rect 20972 13468 21028 13524
rect 21420 13244 21476 13300
rect 21868 13468 21924 13524
rect 22204 15426 22260 15428
rect 22204 15374 22206 15426
rect 22206 15374 22258 15426
rect 22258 15374 22260 15426
rect 22204 15372 22260 15374
rect 22428 15314 22484 15316
rect 22428 15262 22430 15314
rect 22430 15262 22482 15314
rect 22482 15262 22484 15314
rect 22428 15260 22484 15262
rect 22764 16716 22820 16772
rect 22764 15538 22820 15540
rect 22764 15486 22766 15538
rect 22766 15486 22818 15538
rect 22818 15486 22820 15538
rect 22764 15484 22820 15486
rect 22876 16156 22932 16212
rect 23324 15484 23380 15540
rect 22652 14252 22708 14308
rect 20972 12178 21028 12180
rect 20972 12126 20974 12178
rect 20974 12126 21026 12178
rect 21026 12126 21028 12178
rect 20972 12124 21028 12126
rect 21308 11788 21364 11844
rect 21532 12290 21588 12292
rect 21532 12238 21534 12290
rect 21534 12238 21586 12290
rect 21586 12238 21588 12290
rect 21532 12236 21588 12238
rect 21420 11676 21476 11732
rect 21196 11564 21252 11620
rect 20748 11452 20804 11508
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20188 9212 20244 9268
rect 20188 8428 20244 8484
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 17388 6972 17444 7028
rect 18508 6972 18564 7028
rect 16828 6524 16884 6580
rect 18396 6076 18452 6132
rect 16380 5234 16436 5236
rect 16380 5182 16382 5234
rect 16382 5182 16434 5234
rect 16434 5182 16436 5234
rect 16380 5180 16436 5182
rect 16604 5180 16660 5236
rect 11340 5068 11396 5124
rect 13804 4450 13860 4452
rect 13804 4398 13806 4450
rect 13806 4398 13858 4450
rect 13858 4398 13860 4450
rect 13804 4396 13860 4398
rect 15484 4450 15540 4452
rect 15484 4398 15486 4450
rect 15486 4398 15538 4450
rect 15538 4398 15540 4450
rect 15484 4396 15540 4398
rect 11900 3612 11956 3668
rect 13356 3666 13412 3668
rect 13356 3614 13358 3666
rect 13358 3614 13410 3666
rect 13410 3614 13412 3666
rect 13356 3612 13412 3614
rect 15484 4114 15540 4116
rect 15484 4062 15486 4114
rect 15486 4062 15538 4114
rect 15538 4062 15540 4114
rect 15484 4060 15540 4062
rect 14588 3388 14644 3444
rect 17500 5516 17556 5572
rect 17052 5068 17108 5124
rect 17836 4956 17892 5012
rect 16828 4450 16884 4452
rect 16828 4398 16830 4450
rect 16830 4398 16882 4450
rect 16882 4398 16884 4450
rect 16828 4396 16884 4398
rect 16156 3612 16212 3668
rect 15708 2828 15764 2884
rect 17052 3666 17108 3668
rect 17052 3614 17054 3666
rect 17054 3614 17106 3666
rect 17106 3614 17108 3666
rect 17052 3612 17108 3614
rect 17836 4060 17892 4116
rect 16268 3388 16324 3444
rect 17500 3442 17556 3444
rect 17500 3390 17502 3442
rect 17502 3390 17554 3442
rect 17554 3390 17556 3442
rect 17500 3388 17556 3390
rect 17948 3612 18004 3668
rect 18060 3442 18116 3444
rect 18060 3390 18062 3442
rect 18062 3390 18114 3442
rect 18114 3390 18116 3442
rect 18060 3388 18116 3390
rect 17836 2492 17892 2548
rect 18620 6636 18676 6692
rect 20076 6972 20132 7028
rect 19628 6466 19684 6468
rect 19628 6414 19630 6466
rect 19630 6414 19682 6466
rect 19682 6414 19684 6466
rect 19628 6412 19684 6414
rect 21420 11004 21476 11060
rect 21756 12178 21812 12180
rect 21756 12126 21758 12178
rect 21758 12126 21810 12178
rect 21810 12126 21812 12178
rect 21756 12124 21812 12126
rect 22428 12290 22484 12292
rect 22428 12238 22430 12290
rect 22430 12238 22482 12290
rect 22482 12238 22484 12290
rect 22428 12236 22484 12238
rect 22204 12178 22260 12180
rect 22204 12126 22206 12178
rect 22206 12126 22258 12178
rect 22258 12126 22260 12178
rect 22204 12124 22260 12126
rect 22876 12178 22932 12180
rect 22876 12126 22878 12178
rect 22878 12126 22930 12178
rect 22930 12126 22932 12178
rect 22876 12124 22932 12126
rect 22204 11788 22260 11844
rect 21644 11282 21700 11284
rect 21644 11230 21646 11282
rect 21646 11230 21698 11282
rect 21698 11230 21700 11282
rect 21644 11228 21700 11230
rect 21644 11004 21700 11060
rect 20972 10556 21028 10612
rect 21420 10610 21476 10612
rect 21420 10558 21422 10610
rect 21422 10558 21474 10610
rect 21474 10558 21476 10610
rect 21420 10556 21476 10558
rect 22092 11004 22148 11060
rect 22092 10610 22148 10612
rect 22092 10558 22094 10610
rect 22094 10558 22146 10610
rect 22146 10558 22148 10610
rect 22092 10556 22148 10558
rect 21532 9938 21588 9940
rect 21532 9886 21534 9938
rect 21534 9886 21586 9938
rect 21586 9886 21588 9938
rect 21532 9884 21588 9886
rect 20748 9602 20804 9604
rect 20748 9550 20750 9602
rect 20750 9550 20802 9602
rect 20802 9550 20804 9602
rect 20748 9548 20804 9550
rect 20972 9266 21028 9268
rect 20972 9214 20974 9266
rect 20974 9214 21026 9266
rect 21026 9214 21028 9266
rect 20972 9212 21028 9214
rect 20412 8930 20468 8932
rect 20412 8878 20414 8930
rect 20414 8878 20466 8930
rect 20466 8878 20468 8930
rect 20412 8876 20468 8878
rect 21756 9154 21812 9156
rect 21756 9102 21758 9154
rect 21758 9102 21810 9154
rect 21810 9102 21812 9154
rect 21756 9100 21812 9102
rect 21756 8316 21812 8372
rect 21420 8204 21476 8260
rect 20412 8146 20468 8148
rect 20412 8094 20414 8146
rect 20414 8094 20466 8146
rect 20466 8094 20468 8146
rect 20412 8092 20468 8094
rect 21532 7980 21588 8036
rect 21980 9324 22036 9380
rect 22540 11676 22596 11732
rect 22876 11116 22932 11172
rect 22204 9100 22260 9156
rect 22988 10780 23044 10836
rect 23324 12348 23380 12404
rect 23660 10444 23716 10500
rect 22428 9154 22484 9156
rect 22428 9102 22430 9154
rect 22430 9102 22482 9154
rect 22482 9102 22484 9154
rect 22428 9100 22484 9102
rect 22316 8876 22372 8932
rect 22540 8316 22596 8372
rect 21644 7868 21700 7924
rect 20524 7362 20580 7364
rect 20524 7310 20526 7362
rect 20526 7310 20578 7362
rect 20578 7310 20580 7362
rect 20524 7308 20580 7310
rect 21308 7196 21364 7252
rect 19068 5628 19124 5684
rect 19180 5292 19236 5348
rect 18844 4956 18900 5012
rect 18620 4898 18676 4900
rect 18620 4846 18622 4898
rect 18622 4846 18674 4898
rect 18674 4846 18676 4898
rect 18620 4844 18676 4846
rect 18732 3666 18788 3668
rect 18732 3614 18734 3666
rect 18734 3614 18786 3666
rect 18786 3614 18788 3666
rect 18732 3612 18788 3614
rect 19292 5234 19348 5236
rect 19292 5182 19294 5234
rect 19294 5182 19346 5234
rect 19346 5182 19348 5234
rect 19292 5180 19348 5182
rect 18956 4450 19012 4452
rect 18956 4398 18958 4450
rect 18958 4398 19010 4450
rect 19010 4398 19012 4450
rect 18956 4396 19012 4398
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20412 6524 20468 6580
rect 21084 6412 21140 6468
rect 20300 5292 20356 5348
rect 20300 5010 20356 5012
rect 20300 4958 20302 5010
rect 20302 4958 20354 5010
rect 20354 4958 20356 5010
rect 20300 4956 20356 4958
rect 21532 5404 21588 5460
rect 21308 5122 21364 5124
rect 21308 5070 21310 5122
rect 21310 5070 21362 5122
rect 21362 5070 21364 5122
rect 21308 5068 21364 5070
rect 20636 4844 20692 4900
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 22764 7980 22820 8036
rect 24556 20914 24612 20916
rect 24556 20862 24558 20914
rect 24558 20862 24610 20914
rect 24610 20862 24612 20914
rect 24556 20860 24612 20862
rect 24332 20076 24388 20132
rect 24332 19180 24388 19236
rect 24668 20300 24724 20356
rect 24444 18620 24500 18676
rect 24780 18620 24836 18676
rect 24556 17778 24612 17780
rect 24556 17726 24558 17778
rect 24558 17726 24610 17778
rect 24610 17726 24612 17778
rect 24556 17724 24612 17726
rect 27020 22428 27076 22484
rect 26684 22316 26740 22372
rect 26236 21868 26292 21924
rect 26012 21644 26068 21700
rect 25900 21532 25956 21588
rect 25004 20972 25060 21028
rect 25900 20860 25956 20916
rect 26684 21586 26740 21588
rect 26684 21534 26686 21586
rect 26686 21534 26738 21586
rect 26738 21534 26740 21586
rect 26684 21532 26740 21534
rect 27244 24556 27300 24612
rect 28476 55020 28532 55076
rect 29372 55074 29428 55076
rect 29372 55022 29374 55074
rect 29374 55022 29426 55074
rect 29426 55022 29428 55074
rect 29372 55020 29428 55022
rect 28364 26572 28420 26628
rect 28364 24892 28420 24948
rect 27244 23100 27300 23156
rect 27132 20972 27188 21028
rect 26460 20130 26516 20132
rect 26460 20078 26462 20130
rect 26462 20078 26514 20130
rect 26514 20078 26516 20130
rect 26460 20076 26516 20078
rect 26236 20018 26292 20020
rect 26236 19966 26238 20018
rect 26238 19966 26290 20018
rect 26290 19966 26292 20018
rect 26236 19964 26292 19966
rect 25340 19068 25396 19124
rect 27020 19404 27076 19460
rect 27804 23772 27860 23828
rect 27804 23100 27860 23156
rect 28140 22428 28196 22484
rect 28028 22258 28084 22260
rect 28028 22206 28030 22258
rect 28030 22206 28082 22258
rect 28082 22206 28084 22258
rect 28028 22204 28084 22206
rect 27692 21980 27748 22036
rect 27580 21026 27636 21028
rect 27580 20974 27582 21026
rect 27582 20974 27634 21026
rect 27634 20974 27636 21026
rect 27580 20972 27636 20974
rect 28140 22092 28196 22148
rect 27916 20300 27972 20356
rect 25340 18562 25396 18564
rect 25340 18510 25342 18562
rect 25342 18510 25394 18562
rect 25394 18510 25396 18562
rect 25340 18508 25396 18510
rect 26460 18562 26516 18564
rect 26460 18510 26462 18562
rect 26462 18510 26514 18562
rect 26514 18510 26516 18562
rect 26460 18508 26516 18510
rect 24892 16716 24948 16772
rect 24892 16098 24948 16100
rect 24892 16046 24894 16098
rect 24894 16046 24946 16098
rect 24946 16046 24948 16098
rect 24892 16044 24948 16046
rect 27356 17836 27412 17892
rect 25788 15484 25844 15540
rect 25228 15426 25284 15428
rect 25228 15374 25230 15426
rect 25230 15374 25282 15426
rect 25282 15374 25284 15426
rect 25228 15372 25284 15374
rect 24556 15260 24612 15316
rect 25340 15314 25396 15316
rect 25340 15262 25342 15314
rect 25342 15262 25394 15314
rect 25394 15262 25396 15314
rect 25340 15260 25396 15262
rect 26124 15484 26180 15540
rect 23996 12402 24052 12404
rect 23996 12350 23998 12402
rect 23998 12350 24050 12402
rect 24050 12350 24052 12402
rect 23996 12348 24052 12350
rect 24220 13244 24276 13300
rect 24668 13020 24724 13076
rect 24780 12348 24836 12404
rect 23884 11788 23940 11844
rect 24556 12178 24612 12180
rect 24556 12126 24558 12178
rect 24558 12126 24610 12178
rect 24610 12126 24612 12178
rect 24556 12124 24612 12126
rect 23884 10834 23940 10836
rect 23884 10782 23886 10834
rect 23886 10782 23938 10834
rect 23938 10782 23940 10834
rect 23884 10780 23940 10782
rect 23772 9212 23828 9268
rect 24668 11788 24724 11844
rect 24332 11340 24388 11396
rect 25228 14140 25284 14196
rect 25676 14252 25732 14308
rect 24892 11676 24948 11732
rect 25004 14028 25060 14084
rect 27132 16604 27188 16660
rect 27804 19068 27860 19124
rect 27804 17388 27860 17444
rect 26684 15260 26740 15316
rect 25788 14140 25844 14196
rect 26124 13244 26180 13300
rect 25004 12684 25060 12740
rect 25452 13074 25508 13076
rect 25452 13022 25454 13074
rect 25454 13022 25506 13074
rect 25506 13022 25508 13074
rect 25452 13020 25508 13022
rect 25340 12178 25396 12180
rect 25340 12126 25342 12178
rect 25342 12126 25394 12178
rect 25394 12126 25396 12178
rect 25340 12124 25396 12126
rect 26684 14252 26740 14308
rect 27356 13634 27412 13636
rect 27356 13582 27358 13634
rect 27358 13582 27410 13634
rect 27410 13582 27412 13634
rect 27356 13580 27412 13582
rect 27356 13356 27412 13412
rect 26684 13244 26740 13300
rect 25788 12348 25844 12404
rect 25564 12236 25620 12292
rect 26236 12290 26292 12292
rect 26236 12238 26238 12290
rect 26238 12238 26290 12290
rect 26290 12238 26292 12290
rect 26236 12236 26292 12238
rect 25452 12012 25508 12068
rect 25228 11900 25284 11956
rect 25340 11170 25396 11172
rect 25340 11118 25342 11170
rect 25342 11118 25394 11170
rect 25394 11118 25396 11170
rect 25340 11116 25396 11118
rect 24444 10444 24500 10500
rect 24220 10386 24276 10388
rect 24220 10334 24222 10386
rect 24222 10334 24274 10386
rect 24274 10334 24276 10386
rect 24220 10332 24276 10334
rect 25228 10386 25284 10388
rect 25228 10334 25230 10386
rect 25230 10334 25282 10386
rect 25282 10334 25284 10386
rect 25228 10332 25284 10334
rect 25116 9938 25172 9940
rect 25116 9886 25118 9938
rect 25118 9886 25170 9938
rect 25170 9886 25172 9938
rect 25116 9884 25172 9886
rect 25564 10386 25620 10388
rect 25564 10334 25566 10386
rect 25566 10334 25618 10386
rect 25618 10334 25620 10386
rect 25564 10332 25620 10334
rect 27132 12684 27188 12740
rect 26460 11788 26516 11844
rect 26796 11900 26852 11956
rect 22316 7420 22372 7476
rect 23436 8204 23492 8260
rect 23212 7474 23268 7476
rect 23212 7422 23214 7474
rect 23214 7422 23266 7474
rect 23266 7422 23268 7474
rect 23212 7420 23268 7422
rect 22876 7308 22932 7364
rect 22540 7084 22596 7140
rect 21756 6578 21812 6580
rect 21756 6526 21758 6578
rect 21758 6526 21810 6578
rect 21810 6526 21812 6578
rect 21756 6524 21812 6526
rect 21868 5906 21924 5908
rect 21868 5854 21870 5906
rect 21870 5854 21922 5906
rect 21922 5854 21924 5906
rect 21868 5852 21924 5854
rect 22316 5404 22372 5460
rect 22764 6972 22820 7028
rect 22540 6636 22596 6692
rect 21868 5292 21924 5348
rect 21756 5180 21812 5236
rect 22652 6748 22708 6804
rect 22876 6524 22932 6580
rect 23436 6972 23492 7028
rect 24444 8876 24500 8932
rect 23884 8258 23940 8260
rect 23884 8206 23886 8258
rect 23886 8206 23938 8258
rect 23938 8206 23940 8258
rect 23884 8204 23940 8206
rect 24332 7868 24388 7924
rect 23324 6076 23380 6132
rect 22092 4284 22148 4340
rect 22876 4396 22932 4452
rect 20188 3612 20244 3668
rect 19740 3442 19796 3444
rect 19740 3390 19742 3442
rect 19742 3390 19794 3442
rect 19794 3390 19796 3442
rect 19740 3388 19796 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 20972 3666 21028 3668
rect 20972 3614 20974 3666
rect 20974 3614 21026 3666
rect 21026 3614 21028 3666
rect 20972 3612 21028 3614
rect 21308 3388 21364 3444
rect 23436 6524 23492 6580
rect 23212 5852 23268 5908
rect 23548 5180 23604 5236
rect 23660 6524 23716 6580
rect 23212 4956 23268 5012
rect 23324 4508 23380 4564
rect 24668 7980 24724 8036
rect 24556 7698 24612 7700
rect 24556 7646 24558 7698
rect 24558 7646 24610 7698
rect 24610 7646 24612 7698
rect 24556 7644 24612 7646
rect 24668 7586 24724 7588
rect 24668 7534 24670 7586
rect 24670 7534 24722 7586
rect 24722 7534 24724 7586
rect 24668 7532 24724 7534
rect 24556 7308 24612 7364
rect 23996 6524 24052 6580
rect 24332 6972 24388 7028
rect 24780 7196 24836 7252
rect 26124 10780 26180 10836
rect 26572 10610 26628 10612
rect 26572 10558 26574 10610
rect 26574 10558 26626 10610
rect 26626 10558 26628 10610
rect 26572 10556 26628 10558
rect 26236 10444 26292 10500
rect 27132 11954 27188 11956
rect 27132 11902 27134 11954
rect 27134 11902 27186 11954
rect 27186 11902 27188 11954
rect 27132 11900 27188 11902
rect 26908 11788 26964 11844
rect 27244 10780 27300 10836
rect 27020 10498 27076 10500
rect 27020 10446 27022 10498
rect 27022 10446 27074 10498
rect 27074 10446 27076 10498
rect 27020 10444 27076 10446
rect 26796 10332 26852 10388
rect 26124 9548 26180 9604
rect 25228 8540 25284 8596
rect 24780 6412 24836 6468
rect 23772 3836 23828 3892
rect 24108 4338 24164 4340
rect 24108 4286 24110 4338
rect 24110 4286 24162 4338
rect 24162 4286 24164 4338
rect 24108 4284 24164 4286
rect 25228 5628 25284 5684
rect 25564 7756 25620 7812
rect 25452 7196 25508 7252
rect 26012 8652 26068 8708
rect 25788 8204 25844 8260
rect 25676 7420 25732 7476
rect 25788 7644 25844 7700
rect 25900 7532 25956 7588
rect 25900 6524 25956 6580
rect 25900 5628 25956 5684
rect 25676 4956 25732 5012
rect 25676 4508 25732 4564
rect 24444 4338 24500 4340
rect 24444 4286 24446 4338
rect 24446 4286 24498 4338
rect 24498 4286 24500 4338
rect 24444 4284 24500 4286
rect 25228 4172 25284 4228
rect 26236 7756 26292 7812
rect 26236 6748 26292 6804
rect 27692 12124 27748 12180
rect 27580 11900 27636 11956
rect 27692 11788 27748 11844
rect 28588 20802 28644 20804
rect 28588 20750 28590 20802
rect 28590 20750 28642 20802
rect 28642 20750 28644 20802
rect 28588 20748 28644 20750
rect 28588 19906 28644 19908
rect 28588 19854 28590 19906
rect 28590 19854 28642 19906
rect 28642 19854 28644 19906
rect 28588 19852 28644 19854
rect 28476 19404 28532 19460
rect 51548 56082 51604 56084
rect 51548 56030 51550 56082
rect 51550 56030 51602 56082
rect 51602 56030 51604 56082
rect 51548 56028 51604 56030
rect 62748 56252 62804 56308
rect 63980 56306 64036 56308
rect 63980 56254 63982 56306
rect 63982 56254 64034 56306
rect 64034 56254 64036 56306
rect 63980 56252 64036 56254
rect 61292 56028 61348 56084
rect 43708 55020 43764 55076
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 37884 30828 37940 30884
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 32844 30268 32900 30324
rect 29820 27692 29876 27748
rect 29708 27580 29764 27636
rect 29372 22540 29428 22596
rect 29372 22370 29428 22372
rect 29372 22318 29374 22370
rect 29374 22318 29426 22370
rect 29426 22318 29428 22370
rect 29372 22316 29428 22318
rect 29036 22258 29092 22260
rect 29036 22206 29038 22258
rect 29038 22206 29090 22258
rect 29090 22206 29092 22258
rect 29036 22204 29092 22206
rect 29148 22092 29204 22148
rect 29820 21756 29876 21812
rect 29372 20802 29428 20804
rect 29372 20750 29374 20802
rect 29374 20750 29426 20802
rect 29426 20750 29428 20802
rect 29372 20748 29428 20750
rect 29148 20300 29204 20356
rect 28700 18396 28756 18452
rect 28700 17612 28756 17668
rect 28812 19068 28868 19124
rect 27916 16604 27972 16660
rect 28812 16156 28868 16212
rect 28476 15036 28532 15092
rect 29036 15260 29092 15316
rect 29260 18844 29316 18900
rect 29596 18396 29652 18452
rect 32620 28028 32676 28084
rect 30940 27970 30996 27972
rect 30940 27918 30942 27970
rect 30942 27918 30994 27970
rect 30994 27918 30996 27970
rect 30940 27916 30996 27918
rect 31612 27916 31668 27972
rect 30156 27746 30212 27748
rect 30156 27694 30158 27746
rect 30158 27694 30210 27746
rect 30210 27694 30212 27746
rect 30156 27692 30212 27694
rect 30716 27580 30772 27636
rect 31388 27020 31444 27076
rect 30268 26290 30324 26292
rect 30268 26238 30270 26290
rect 30270 26238 30322 26290
rect 30322 26238 30324 26290
rect 30268 26236 30324 26238
rect 30940 26290 30996 26292
rect 30940 26238 30942 26290
rect 30942 26238 30994 26290
rect 30994 26238 30996 26290
rect 30940 26236 30996 26238
rect 31724 27804 31780 27860
rect 31724 27074 31780 27076
rect 31724 27022 31726 27074
rect 31726 27022 31778 27074
rect 31778 27022 31780 27074
rect 31724 27020 31780 27022
rect 31836 26572 31892 26628
rect 30492 26012 30548 26068
rect 31836 26012 31892 26068
rect 31388 24946 31444 24948
rect 31388 24894 31390 24946
rect 31390 24894 31442 24946
rect 31442 24894 31444 24946
rect 31388 24892 31444 24894
rect 31276 24834 31332 24836
rect 31276 24782 31278 24834
rect 31278 24782 31330 24834
rect 31330 24782 31332 24834
rect 31276 24780 31332 24782
rect 30492 24610 30548 24612
rect 30492 24558 30494 24610
rect 30494 24558 30546 24610
rect 30546 24558 30548 24610
rect 30492 24556 30548 24558
rect 31948 25506 32004 25508
rect 31948 25454 31950 25506
rect 31950 25454 32002 25506
rect 32002 25454 32004 25506
rect 31948 25452 32004 25454
rect 31836 24780 31892 24836
rect 30492 23660 30548 23716
rect 31164 23660 31220 23716
rect 31500 22540 31556 22596
rect 30716 21644 30772 21700
rect 30044 21474 30100 21476
rect 30044 21422 30046 21474
rect 30046 21422 30098 21474
rect 30098 21422 30100 21474
rect 30044 21420 30100 21422
rect 30044 20802 30100 20804
rect 30044 20750 30046 20802
rect 30046 20750 30098 20802
rect 30098 20750 30100 20802
rect 30044 20748 30100 20750
rect 30268 19964 30324 20020
rect 29596 15874 29652 15876
rect 29596 15822 29598 15874
rect 29598 15822 29650 15874
rect 29650 15822 29652 15874
rect 29596 15820 29652 15822
rect 30940 20018 30996 20020
rect 30940 19966 30942 20018
rect 30942 19966 30994 20018
rect 30994 19966 30996 20018
rect 30940 19964 30996 19966
rect 31164 19906 31220 19908
rect 31164 19854 31166 19906
rect 31166 19854 31218 19906
rect 31218 19854 31220 19906
rect 31164 19852 31220 19854
rect 30268 19122 30324 19124
rect 30268 19070 30270 19122
rect 30270 19070 30322 19122
rect 30322 19070 30324 19122
rect 30268 19068 30324 19070
rect 31052 18956 31108 19012
rect 30268 18450 30324 18452
rect 30268 18398 30270 18450
rect 30270 18398 30322 18450
rect 30322 18398 30324 18450
rect 30268 18396 30324 18398
rect 30492 18450 30548 18452
rect 30492 18398 30494 18450
rect 30494 18398 30546 18450
rect 30546 18398 30548 18450
rect 30492 18396 30548 18398
rect 32620 24722 32676 24724
rect 32620 24670 32622 24722
rect 32622 24670 32674 24722
rect 32674 24670 32676 24722
rect 32620 24668 32676 24670
rect 32060 24556 32116 24612
rect 32172 23772 32228 23828
rect 31836 22428 31892 22484
rect 32732 22482 32788 22484
rect 32732 22430 32734 22482
rect 32734 22430 32786 22482
rect 32786 22430 32788 22482
rect 32732 22428 32788 22430
rect 31612 21698 31668 21700
rect 31612 21646 31614 21698
rect 31614 21646 31666 21698
rect 31666 21646 31668 21698
rect 31612 21644 31668 21646
rect 31724 20076 31780 20132
rect 31612 19852 31668 19908
rect 31948 19740 32004 19796
rect 31836 19180 31892 19236
rect 32284 20130 32340 20132
rect 32284 20078 32286 20130
rect 32286 20078 32338 20130
rect 32338 20078 32340 20130
rect 32284 20076 32340 20078
rect 32396 19852 32452 19908
rect 32172 19740 32228 19796
rect 31388 18508 31444 18564
rect 31836 18284 31892 18340
rect 30828 17442 30884 17444
rect 30828 17390 30830 17442
rect 30830 17390 30882 17442
rect 30882 17390 30884 17442
rect 30828 17388 30884 17390
rect 29932 16828 29988 16884
rect 29820 16098 29876 16100
rect 29820 16046 29822 16098
rect 29822 16046 29874 16098
rect 29874 16046 29876 16098
rect 29820 16044 29876 16046
rect 30380 16716 30436 16772
rect 30492 16098 30548 16100
rect 30492 16046 30494 16098
rect 30494 16046 30546 16098
rect 30546 16046 30548 16098
rect 30492 16044 30548 16046
rect 30380 15708 30436 15764
rect 29148 14418 29204 14420
rect 29148 14366 29150 14418
rect 29150 14366 29202 14418
rect 29202 14366 29204 14418
rect 29148 14364 29204 14366
rect 29708 14306 29764 14308
rect 29708 14254 29710 14306
rect 29710 14254 29762 14306
rect 29762 14254 29764 14306
rect 29708 14252 29764 14254
rect 28252 13356 28308 13412
rect 28140 11564 28196 11620
rect 28364 12684 28420 12740
rect 29148 12348 29204 12404
rect 29932 12850 29988 12852
rect 29932 12798 29934 12850
rect 29934 12798 29986 12850
rect 29986 12798 29988 12850
rect 29932 12796 29988 12798
rect 29596 12572 29652 12628
rect 29708 12290 29764 12292
rect 29708 12238 29710 12290
rect 29710 12238 29762 12290
rect 29762 12238 29764 12290
rect 29708 12236 29764 12238
rect 28812 12124 28868 12180
rect 28364 11788 28420 11844
rect 27020 8988 27076 9044
rect 26572 8034 26628 8036
rect 26572 7982 26574 8034
rect 26574 7982 26626 8034
rect 26626 7982 26628 8034
rect 26572 7980 26628 7982
rect 26460 6300 26516 6356
rect 27132 8876 27188 8932
rect 28028 10892 28084 10948
rect 28476 11564 28532 11620
rect 28028 10610 28084 10612
rect 28028 10558 28030 10610
rect 28030 10558 28082 10610
rect 28082 10558 28084 10610
rect 28028 10556 28084 10558
rect 27916 9436 27972 9492
rect 27804 8876 27860 8932
rect 27804 8428 27860 8484
rect 28028 8316 28084 8372
rect 26684 6188 26740 6244
rect 26908 6412 26964 6468
rect 26796 6076 26852 6132
rect 26348 5852 26404 5908
rect 24668 3948 24724 4004
rect 26236 4060 26292 4116
rect 26460 4620 26516 4676
rect 23548 3052 23604 3108
rect 24892 3330 24948 3332
rect 24892 3278 24894 3330
rect 24894 3278 24946 3330
rect 24946 3278 24948 3330
rect 24892 3276 24948 3278
rect 24556 3164 24612 3220
rect 23100 2940 23156 2996
rect 27244 7586 27300 7588
rect 27244 7534 27246 7586
rect 27246 7534 27298 7586
rect 27298 7534 27300 7586
rect 27244 7532 27300 7534
rect 28476 9436 28532 9492
rect 28364 8876 28420 8932
rect 28252 8316 28308 8372
rect 28364 7980 28420 8036
rect 28140 6690 28196 6692
rect 28140 6638 28142 6690
rect 28142 6638 28194 6690
rect 28194 6638 28196 6690
rect 28140 6636 28196 6638
rect 27580 6466 27636 6468
rect 27580 6414 27582 6466
rect 27582 6414 27634 6466
rect 27634 6414 27636 6466
rect 27580 6412 27636 6414
rect 27356 6300 27412 6356
rect 27244 6018 27300 6020
rect 27244 5966 27246 6018
rect 27246 5966 27298 6018
rect 27298 5966 27300 6018
rect 27244 5964 27300 5966
rect 27356 5852 27412 5908
rect 28476 7420 28532 7476
rect 28700 11506 28756 11508
rect 28700 11454 28702 11506
rect 28702 11454 28754 11506
rect 28754 11454 28756 11506
rect 28700 11452 28756 11454
rect 28700 8146 28756 8148
rect 28700 8094 28702 8146
rect 28702 8094 28754 8146
rect 28754 8094 28756 8146
rect 28700 8092 28756 8094
rect 28924 11452 28980 11508
rect 28924 10668 28980 10724
rect 29932 11340 29988 11396
rect 29260 11170 29316 11172
rect 29260 11118 29262 11170
rect 29262 11118 29314 11170
rect 29314 11118 29316 11170
rect 29260 11116 29316 11118
rect 28924 9100 28980 9156
rect 29372 9772 29428 9828
rect 29260 9100 29316 9156
rect 29932 11170 29988 11172
rect 29932 11118 29934 11170
rect 29934 11118 29986 11170
rect 29986 11118 29988 11170
rect 29932 11116 29988 11118
rect 29932 10668 29988 10724
rect 30156 14364 30212 14420
rect 30492 13916 30548 13972
rect 30380 13746 30436 13748
rect 30380 13694 30382 13746
rect 30382 13694 30434 13746
rect 30434 13694 30436 13746
rect 30380 13692 30436 13694
rect 30268 13634 30324 13636
rect 30268 13582 30270 13634
rect 30270 13582 30322 13634
rect 30322 13582 30324 13634
rect 30268 13580 30324 13582
rect 31164 17052 31220 17108
rect 30716 16882 30772 16884
rect 30716 16830 30718 16882
rect 30718 16830 30770 16882
rect 30770 16830 30772 16882
rect 30716 16828 30772 16830
rect 31052 16716 31108 16772
rect 31500 16828 31556 16884
rect 31836 16882 31892 16884
rect 31836 16830 31838 16882
rect 31838 16830 31890 16882
rect 31890 16830 31892 16882
rect 31836 16828 31892 16830
rect 32060 18620 32116 18676
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 36876 29036 36932 29092
rect 33404 28028 33460 28084
rect 33180 27804 33236 27860
rect 34188 27916 34244 27972
rect 35756 27916 35812 27972
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34636 26348 34692 26404
rect 35644 26962 35700 26964
rect 35644 26910 35646 26962
rect 35646 26910 35698 26962
rect 35698 26910 35700 26962
rect 35644 26908 35700 26910
rect 35868 27804 35924 27860
rect 35532 26290 35588 26292
rect 35532 26238 35534 26290
rect 35534 26238 35586 26290
rect 35586 26238 35588 26290
rect 35532 26236 35588 26238
rect 34748 26012 34804 26068
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 33964 25394 34020 25396
rect 33964 25342 33966 25394
rect 33966 25342 34018 25394
rect 34018 25342 34020 25394
rect 33964 25340 34020 25342
rect 34860 25506 34916 25508
rect 34860 25454 34862 25506
rect 34862 25454 34914 25506
rect 34914 25454 34916 25506
rect 34860 25452 34916 25454
rect 33628 25282 33684 25284
rect 33628 25230 33630 25282
rect 33630 25230 33682 25282
rect 33682 25230 33684 25282
rect 33628 25228 33684 25230
rect 34748 24722 34804 24724
rect 34748 24670 34750 24722
rect 34750 24670 34802 24722
rect 34802 24670 34804 24722
rect 34748 24668 34804 24670
rect 33068 23660 33124 23716
rect 34076 23266 34132 23268
rect 34076 23214 34078 23266
rect 34078 23214 34130 23266
rect 34130 23214 34132 23266
rect 34076 23212 34132 23214
rect 33516 23100 33572 23156
rect 33404 21698 33460 21700
rect 33404 21646 33406 21698
rect 33406 21646 33458 21698
rect 33458 21646 33460 21698
rect 33404 21644 33460 21646
rect 35196 25730 35252 25732
rect 35196 25678 35198 25730
rect 35198 25678 35250 25730
rect 35250 25678 35252 25730
rect 35196 25676 35252 25678
rect 35756 26124 35812 26180
rect 35756 25788 35812 25844
rect 35308 24834 35364 24836
rect 35308 24782 35310 24834
rect 35310 24782 35362 24834
rect 35362 24782 35364 24834
rect 35308 24780 35364 24782
rect 35756 24780 35812 24836
rect 34972 23996 35028 24052
rect 34188 23100 34244 23156
rect 34412 23714 34468 23716
rect 34412 23662 34414 23714
rect 34414 23662 34466 23714
rect 34466 23662 34468 23714
rect 34412 23660 34468 23662
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 33740 22316 33796 22372
rect 33628 21420 33684 21476
rect 33404 20018 33460 20020
rect 33404 19966 33406 20018
rect 33406 19966 33458 20018
rect 33458 19966 33460 20018
rect 33404 19964 33460 19966
rect 32956 18956 33012 19012
rect 33628 19852 33684 19908
rect 33628 19292 33684 19348
rect 33180 18620 33236 18676
rect 32172 16716 32228 16772
rect 31052 16044 31108 16100
rect 31836 16098 31892 16100
rect 31836 16046 31838 16098
rect 31838 16046 31890 16098
rect 31890 16046 31892 16098
rect 31836 16044 31892 16046
rect 31052 15874 31108 15876
rect 31052 15822 31054 15874
rect 31054 15822 31106 15874
rect 31106 15822 31108 15874
rect 31052 15820 31108 15822
rect 31052 14252 31108 14308
rect 35644 23436 35700 23492
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34412 21698 34468 21700
rect 34412 21646 34414 21698
rect 34414 21646 34466 21698
rect 34466 21646 34468 21698
rect 34412 21644 34468 21646
rect 34636 21532 34692 21588
rect 34412 21420 34468 21476
rect 33852 20018 33908 20020
rect 33852 19966 33854 20018
rect 33854 19966 33906 20018
rect 33906 19966 33908 20018
rect 33852 19964 33908 19966
rect 34188 20130 34244 20132
rect 34188 20078 34190 20130
rect 34190 20078 34242 20130
rect 34242 20078 34244 20130
rect 34188 20076 34244 20078
rect 34076 19740 34132 19796
rect 33852 19234 33908 19236
rect 33852 19182 33854 19234
rect 33854 19182 33906 19234
rect 33906 19182 33908 19234
rect 33852 19180 33908 19182
rect 32620 17948 32676 18004
rect 32396 16882 32452 16884
rect 32396 16830 32398 16882
rect 32398 16830 32450 16882
rect 32450 16830 32452 16882
rect 32396 16828 32452 16830
rect 33180 17612 33236 17668
rect 33516 18226 33572 18228
rect 33516 18174 33518 18226
rect 33518 18174 33570 18226
rect 33570 18174 33572 18226
rect 33516 18172 33572 18174
rect 33628 17948 33684 18004
rect 33740 18338 33796 18340
rect 33740 18286 33742 18338
rect 33742 18286 33794 18338
rect 33794 18286 33796 18338
rect 33740 18284 33796 18286
rect 33404 16322 33460 16324
rect 33404 16270 33406 16322
rect 33406 16270 33458 16322
rect 33458 16270 33460 16322
rect 33404 16268 33460 16270
rect 32508 16098 32564 16100
rect 32508 16046 32510 16098
rect 32510 16046 32562 16098
rect 32562 16046 32564 16098
rect 32508 16044 32564 16046
rect 34300 19180 34356 19236
rect 36540 26402 36596 26404
rect 36540 26350 36542 26402
rect 36542 26350 36594 26402
rect 36594 26350 36596 26402
rect 36540 26348 36596 26350
rect 36316 25730 36372 25732
rect 36316 25678 36318 25730
rect 36318 25678 36370 25730
rect 36370 25678 36372 25730
rect 36316 25676 36372 25678
rect 36652 26178 36708 26180
rect 36652 26126 36654 26178
rect 36654 26126 36706 26178
rect 36706 26126 36708 26178
rect 36652 26124 36708 26126
rect 36764 26066 36820 26068
rect 36764 26014 36766 26066
rect 36766 26014 36818 26066
rect 36818 26014 36820 26066
rect 36764 26012 36820 26014
rect 36092 25228 36148 25284
rect 37436 26236 37492 26292
rect 37772 26124 37828 26180
rect 37548 26012 37604 26068
rect 36988 25228 37044 25284
rect 36204 24668 36260 24724
rect 36988 24780 37044 24836
rect 37100 24668 37156 24724
rect 36988 24556 37044 24612
rect 36316 24498 36372 24500
rect 36316 24446 36318 24498
rect 36318 24446 36370 24498
rect 36370 24446 36372 24498
rect 36316 24444 36372 24446
rect 37436 24498 37492 24500
rect 37436 24446 37438 24498
rect 37438 24446 37490 24498
rect 37490 24446 37492 24498
rect 37436 24444 37492 24446
rect 37548 23884 37604 23940
rect 37436 23548 37492 23604
rect 36428 23212 36484 23268
rect 36428 22482 36484 22484
rect 36428 22430 36430 22482
rect 36430 22430 36482 22482
rect 36482 22430 36484 22482
rect 36428 22428 36484 22430
rect 36988 22764 37044 22820
rect 35644 21532 35700 21588
rect 37212 22204 37268 22260
rect 35532 21420 35588 21476
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34860 20300 34916 20356
rect 36652 21474 36708 21476
rect 36652 21422 36654 21474
rect 36654 21422 36706 21474
rect 36706 21422 36708 21474
rect 36652 21420 36708 21422
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 36092 19964 36148 20020
rect 35868 19906 35924 19908
rect 35868 19854 35870 19906
rect 35870 19854 35922 19906
rect 35922 19854 35924 19906
rect 35868 19852 35924 19854
rect 35532 18508 35588 18564
rect 34524 17666 34580 17668
rect 34524 17614 34526 17666
rect 34526 17614 34578 17666
rect 34578 17614 34580 17666
rect 34524 17612 34580 17614
rect 33740 16828 33796 16884
rect 34748 18450 34804 18452
rect 34748 18398 34750 18450
rect 34750 18398 34802 18450
rect 34802 18398 34804 18450
rect 34748 18396 34804 18398
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35644 17724 35700 17780
rect 34860 17442 34916 17444
rect 34860 17390 34862 17442
rect 34862 17390 34914 17442
rect 34914 17390 34916 17442
rect 34860 17388 34916 17390
rect 36204 18172 36260 18228
rect 36204 17948 36260 18004
rect 35980 16828 36036 16884
rect 34636 16716 34692 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34972 16268 35028 16324
rect 31948 15036 32004 15092
rect 30828 12962 30884 12964
rect 30828 12910 30830 12962
rect 30830 12910 30882 12962
rect 30882 12910 30884 12962
rect 30828 12908 30884 12910
rect 30268 12178 30324 12180
rect 30268 12126 30270 12178
rect 30270 12126 30322 12178
rect 30322 12126 30324 12178
rect 30268 12124 30324 12126
rect 30268 11564 30324 11620
rect 29708 10332 29764 10388
rect 29260 8764 29316 8820
rect 29036 8652 29092 8708
rect 28700 7756 28756 7812
rect 29484 9042 29540 9044
rect 29484 8990 29486 9042
rect 29486 8990 29538 9042
rect 29538 8990 29540 9042
rect 29484 8988 29540 8990
rect 29484 8370 29540 8372
rect 29484 8318 29486 8370
rect 29486 8318 29538 8370
rect 29538 8318 29540 8370
rect 29484 8316 29540 8318
rect 28812 7644 28868 7700
rect 28588 6860 28644 6916
rect 28364 6412 28420 6468
rect 27132 4396 27188 4452
rect 28028 4732 28084 4788
rect 27804 4172 27860 4228
rect 28140 4620 28196 4676
rect 28812 6972 28868 7028
rect 29148 7474 29204 7476
rect 29148 7422 29150 7474
rect 29150 7422 29202 7474
rect 29202 7422 29204 7474
rect 29148 7420 29204 7422
rect 29260 6972 29316 7028
rect 29260 6802 29316 6804
rect 29260 6750 29262 6802
rect 29262 6750 29314 6802
rect 29314 6750 29316 6802
rect 29260 6748 29316 6750
rect 29148 6412 29204 6468
rect 28924 6300 28980 6356
rect 28812 4956 28868 5012
rect 28924 5964 28980 6020
rect 28700 4732 28756 4788
rect 28476 4396 28532 4452
rect 29484 7084 29540 7140
rect 29596 6972 29652 7028
rect 29484 6914 29540 6916
rect 29484 6862 29486 6914
rect 29486 6862 29538 6914
rect 29538 6862 29540 6914
rect 29484 6860 29540 6862
rect 29596 5964 29652 6020
rect 29484 5122 29540 5124
rect 29484 5070 29486 5122
rect 29486 5070 29538 5122
rect 29538 5070 29540 5122
rect 29484 5068 29540 5070
rect 29148 4450 29204 4452
rect 29148 4398 29150 4450
rect 29150 4398 29202 4450
rect 29202 4398 29204 4450
rect 29148 4396 29204 4398
rect 28924 3948 28980 4004
rect 28700 3554 28756 3556
rect 28700 3502 28702 3554
rect 28702 3502 28754 3554
rect 28754 3502 28756 3554
rect 28700 3500 28756 3502
rect 29932 9826 29988 9828
rect 29932 9774 29934 9826
rect 29934 9774 29986 9826
rect 29986 9774 29988 9826
rect 29932 9772 29988 9774
rect 30940 12850 30996 12852
rect 30940 12798 30942 12850
rect 30942 12798 30994 12850
rect 30994 12798 30996 12850
rect 30940 12796 30996 12798
rect 30604 12572 30660 12628
rect 30940 12124 30996 12180
rect 31164 13858 31220 13860
rect 31164 13806 31166 13858
rect 31166 13806 31218 13858
rect 31218 13806 31220 13858
rect 31164 13804 31220 13806
rect 31500 13804 31556 13860
rect 31388 13692 31444 13748
rect 31500 13244 31556 13300
rect 31724 13356 31780 13412
rect 31052 12460 31108 12516
rect 30828 11340 30884 11396
rect 30492 9996 30548 10052
rect 30044 9042 30100 9044
rect 30044 8990 30046 9042
rect 30046 8990 30098 9042
rect 30098 8990 30100 9042
rect 30044 8988 30100 8990
rect 29932 8258 29988 8260
rect 29932 8206 29934 8258
rect 29934 8206 29986 8258
rect 29986 8206 29988 8258
rect 29932 8204 29988 8206
rect 30044 7756 30100 7812
rect 29932 6578 29988 6580
rect 29932 6526 29934 6578
rect 29934 6526 29986 6578
rect 29986 6526 29988 6578
rect 29932 6524 29988 6526
rect 29820 6076 29876 6132
rect 30604 9548 30660 9604
rect 30268 8764 30324 8820
rect 30940 10556 30996 10612
rect 31948 13186 32004 13188
rect 31948 13134 31950 13186
rect 31950 13134 32002 13186
rect 32002 13134 32004 13186
rect 31948 13132 32004 13134
rect 32508 14252 32564 14308
rect 32172 13356 32228 13412
rect 32284 13132 32340 13188
rect 32060 12684 32116 12740
rect 32508 12962 32564 12964
rect 32508 12910 32510 12962
rect 32510 12910 32562 12962
rect 32562 12910 32564 12962
rect 32508 12908 32564 12910
rect 34412 15874 34468 15876
rect 34412 15822 34414 15874
rect 34414 15822 34466 15874
rect 34466 15822 34468 15874
rect 34412 15820 34468 15822
rect 34860 15484 34916 15540
rect 33964 15372 34020 15428
rect 33516 14252 33572 14308
rect 33516 13634 33572 13636
rect 33516 13582 33518 13634
rect 33518 13582 33570 13634
rect 33570 13582 33572 13634
rect 33516 13580 33572 13582
rect 32844 12850 32900 12852
rect 32844 12798 32846 12850
rect 32846 12798 32898 12850
rect 32898 12798 32900 12850
rect 32844 12796 32900 12798
rect 32060 12012 32116 12068
rect 31388 10780 31444 10836
rect 31052 9548 31108 9604
rect 30716 8988 30772 9044
rect 30156 6860 30212 6916
rect 30268 8428 30324 8484
rect 30492 8316 30548 8372
rect 30828 8428 30884 8484
rect 30716 8258 30772 8260
rect 30716 8206 30718 8258
rect 30718 8206 30770 8258
rect 30770 8206 30772 8258
rect 30716 8204 30772 8206
rect 31052 7586 31108 7588
rect 31052 7534 31054 7586
rect 31054 7534 31106 7586
rect 31106 7534 31108 7586
rect 31052 7532 31108 7534
rect 30492 6972 30548 7028
rect 30604 6914 30660 6916
rect 30604 6862 30606 6914
rect 30606 6862 30658 6914
rect 30658 6862 30660 6914
rect 30604 6860 30660 6862
rect 30044 5964 30100 6020
rect 30828 6802 30884 6804
rect 30828 6750 30830 6802
rect 30830 6750 30882 6802
rect 30882 6750 30884 6802
rect 30828 6748 30884 6750
rect 30492 6636 30548 6692
rect 30604 6524 30660 6580
rect 29820 4732 29876 4788
rect 30716 4956 30772 5012
rect 29820 4338 29876 4340
rect 29820 4286 29822 4338
rect 29822 4286 29874 4338
rect 29874 4286 29876 4338
rect 29820 4284 29876 4286
rect 30604 4226 30660 4228
rect 30604 4174 30606 4226
rect 30606 4174 30658 4226
rect 30658 4174 30660 4226
rect 30604 4172 30660 4174
rect 31052 3500 31108 3556
rect 31612 10722 31668 10724
rect 31612 10670 31614 10722
rect 31614 10670 31666 10722
rect 31666 10670 31668 10722
rect 31612 10668 31668 10670
rect 31388 7756 31444 7812
rect 31388 7196 31444 7252
rect 31948 10444 32004 10500
rect 32844 12236 32900 12292
rect 34300 15036 34356 15092
rect 35532 15484 35588 15540
rect 35644 15820 35700 15876
rect 35868 15484 35924 15540
rect 36092 15874 36148 15876
rect 36092 15822 36094 15874
rect 36094 15822 36146 15874
rect 36146 15822 36148 15874
rect 36092 15820 36148 15822
rect 36428 16210 36484 16212
rect 36428 16158 36430 16210
rect 36430 16158 36482 16210
rect 36482 16158 36484 16210
rect 36428 16156 36484 16158
rect 35644 15314 35700 15316
rect 35644 15262 35646 15314
rect 35646 15262 35698 15314
rect 35698 15262 35700 15314
rect 35644 15260 35700 15262
rect 36316 15426 36372 15428
rect 36316 15374 36318 15426
rect 36318 15374 36370 15426
rect 36370 15374 36372 15426
rect 36316 15372 36372 15374
rect 36204 15314 36260 15316
rect 36204 15262 36206 15314
rect 36206 15262 36258 15314
rect 36258 15262 36260 15314
rect 36204 15260 36260 15262
rect 37548 20690 37604 20692
rect 37548 20638 37550 20690
rect 37550 20638 37602 20690
rect 37602 20638 37604 20690
rect 37548 20636 37604 20638
rect 37100 19852 37156 19908
rect 37324 19292 37380 19348
rect 37548 19234 37604 19236
rect 37548 19182 37550 19234
rect 37550 19182 37602 19234
rect 37602 19182 37604 19234
rect 37548 19180 37604 19182
rect 36876 16828 36932 16884
rect 37772 17052 37828 17108
rect 49644 55074 49700 55076
rect 49644 55022 49646 55074
rect 49646 55022 49698 55074
rect 49698 55022 49700 55074
rect 49644 55020 49700 55022
rect 50988 55020 51044 55076
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 59948 55074 60004 55076
rect 59948 55022 59950 55074
rect 59950 55022 60002 55074
rect 60002 55022 60004 55074
rect 59948 55020 60004 55022
rect 60956 55298 61012 55300
rect 60956 55246 60958 55298
rect 60958 55246 61010 55298
rect 61010 55246 61012 55298
rect 60956 55244 61012 55246
rect 62972 56082 63028 56084
rect 62972 56030 62974 56082
rect 62974 56030 63026 56082
rect 63026 56030 63028 56082
rect 62972 56028 63028 56030
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 70364 56252 70420 56308
rect 71596 56306 71652 56308
rect 71596 56254 71598 56306
rect 71598 56254 71650 56306
rect 71650 56254 71652 56306
rect 71596 56252 71652 56254
rect 67116 56194 67172 56196
rect 67116 56142 67118 56194
rect 67118 56142 67170 56194
rect 67170 56142 67172 56194
rect 67116 56140 67172 56142
rect 68012 56140 68068 56196
rect 61740 55244 61796 55300
rect 60508 55020 60564 55076
rect 62188 55298 62244 55300
rect 62188 55246 62190 55298
rect 62190 55246 62242 55298
rect 62242 55246 62244 55298
rect 62188 55244 62244 55246
rect 62972 55244 63028 55300
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 46844 31948 46900 32004
rect 43372 28812 43428 28868
rect 38556 26684 38612 26740
rect 38332 26572 38388 26628
rect 38332 26402 38388 26404
rect 38332 26350 38334 26402
rect 38334 26350 38386 26402
rect 38386 26350 38388 26402
rect 38332 26348 38388 26350
rect 37996 26236 38052 26292
rect 38444 26236 38500 26292
rect 37996 25340 38052 25396
rect 39452 26402 39508 26404
rect 39452 26350 39454 26402
rect 39454 26350 39506 26402
rect 39506 26350 39508 26402
rect 39452 26348 39508 26350
rect 39004 26124 39060 26180
rect 38780 25452 38836 25508
rect 38220 25282 38276 25284
rect 38220 25230 38222 25282
rect 38222 25230 38274 25282
rect 38274 25230 38276 25282
rect 38220 25228 38276 25230
rect 38444 24892 38500 24948
rect 38892 25340 38948 25396
rect 39900 26962 39956 26964
rect 39900 26910 39902 26962
rect 39902 26910 39954 26962
rect 39954 26910 39956 26962
rect 39900 26908 39956 26910
rect 40124 26908 40180 26964
rect 39900 26460 39956 26516
rect 39788 26290 39844 26292
rect 39788 26238 39790 26290
rect 39790 26238 39842 26290
rect 39842 26238 39844 26290
rect 39788 26236 39844 26238
rect 39676 26124 39732 26180
rect 38556 24444 38612 24500
rect 38332 23436 38388 23492
rect 37996 22764 38052 22820
rect 39564 25506 39620 25508
rect 39564 25454 39566 25506
rect 39566 25454 39618 25506
rect 39618 25454 39620 25506
rect 39564 25452 39620 25454
rect 40796 26962 40852 26964
rect 40796 26910 40798 26962
rect 40798 26910 40850 26962
rect 40850 26910 40852 26962
rect 40796 26908 40852 26910
rect 40572 26684 40628 26740
rect 40236 26348 40292 26404
rect 40124 25282 40180 25284
rect 40124 25230 40126 25282
rect 40126 25230 40178 25282
rect 40178 25230 40180 25282
rect 40124 25228 40180 25230
rect 41916 26514 41972 26516
rect 41916 26462 41918 26514
rect 41918 26462 41970 26514
rect 41970 26462 41972 26514
rect 41916 26460 41972 26462
rect 42028 26402 42084 26404
rect 42028 26350 42030 26402
rect 42030 26350 42082 26402
rect 42082 26350 42084 26402
rect 42028 26348 42084 26350
rect 42588 26402 42644 26404
rect 42588 26350 42590 26402
rect 42590 26350 42642 26402
rect 42642 26350 42644 26402
rect 42588 26348 42644 26350
rect 43260 26402 43316 26404
rect 43260 26350 43262 26402
rect 43262 26350 43314 26402
rect 43314 26350 43316 26402
rect 43260 26348 43316 26350
rect 41468 26290 41524 26292
rect 41468 26238 41470 26290
rect 41470 26238 41522 26290
rect 41522 26238 41524 26290
rect 41468 26236 41524 26238
rect 42812 26236 42868 26292
rect 41356 26178 41412 26180
rect 41356 26126 41358 26178
rect 41358 26126 41410 26178
rect 41410 26126 41412 26178
rect 41356 26124 41412 26126
rect 40348 25452 40404 25508
rect 40460 25394 40516 25396
rect 40460 25342 40462 25394
rect 40462 25342 40514 25394
rect 40514 25342 40516 25394
rect 40460 25340 40516 25342
rect 39452 25004 39508 25060
rect 40236 24668 40292 24724
rect 39564 23938 39620 23940
rect 39564 23886 39566 23938
rect 39566 23886 39618 23938
rect 39618 23886 39620 23938
rect 39564 23884 39620 23886
rect 40012 23772 40068 23828
rect 40460 23826 40516 23828
rect 40460 23774 40462 23826
rect 40462 23774 40514 23826
rect 40514 23774 40516 23826
rect 40460 23772 40516 23774
rect 39452 23714 39508 23716
rect 39452 23662 39454 23714
rect 39454 23662 39506 23714
rect 39506 23662 39508 23714
rect 39452 23660 39508 23662
rect 38556 23548 38612 23604
rect 41244 25506 41300 25508
rect 41244 25454 41246 25506
rect 41246 25454 41298 25506
rect 41298 25454 41300 25506
rect 41244 25452 41300 25454
rect 41020 25282 41076 25284
rect 41020 25230 41022 25282
rect 41022 25230 41074 25282
rect 41074 25230 41076 25282
rect 41020 25228 41076 25230
rect 41132 24668 41188 24724
rect 40796 23436 40852 23492
rect 41132 23324 41188 23380
rect 41020 23266 41076 23268
rect 41020 23214 41022 23266
rect 41022 23214 41074 23266
rect 41074 23214 41076 23266
rect 41020 23212 41076 23214
rect 40796 22988 40852 23044
rect 39788 22428 39844 22484
rect 40348 22482 40404 22484
rect 40348 22430 40350 22482
rect 40350 22430 40402 22482
rect 40402 22430 40404 22482
rect 40348 22428 40404 22430
rect 39116 22258 39172 22260
rect 39116 22206 39118 22258
rect 39118 22206 39170 22258
rect 39170 22206 39172 22258
rect 39116 22204 39172 22206
rect 38444 20636 38500 20692
rect 40012 20188 40068 20244
rect 38108 20076 38164 20132
rect 38444 20130 38500 20132
rect 38444 20078 38446 20130
rect 38446 20078 38498 20130
rect 38498 20078 38500 20130
rect 38444 20076 38500 20078
rect 39004 20076 39060 20132
rect 37996 19906 38052 19908
rect 37996 19854 37998 19906
rect 37998 19854 38050 19906
rect 38050 19854 38052 19906
rect 37996 19852 38052 19854
rect 39004 19906 39060 19908
rect 39004 19854 39006 19906
rect 39006 19854 39058 19906
rect 39058 19854 39060 19906
rect 39004 19852 39060 19854
rect 38220 19292 38276 19348
rect 39116 19404 39172 19460
rect 37996 19234 38052 19236
rect 37996 19182 37998 19234
rect 37998 19182 38050 19234
rect 38050 19182 38052 19234
rect 37996 19180 38052 19182
rect 39900 19180 39956 19236
rect 36988 16156 37044 16212
rect 37212 16828 37268 16884
rect 36988 15820 37044 15876
rect 39452 17612 39508 17668
rect 39004 17500 39060 17556
rect 38220 17388 38276 17444
rect 39564 17554 39620 17556
rect 39564 17502 39566 17554
rect 39566 17502 39618 17554
rect 39618 17502 39620 17554
rect 39564 17500 39620 17502
rect 39228 17442 39284 17444
rect 39228 17390 39230 17442
rect 39230 17390 39282 17442
rect 39282 17390 39284 17442
rect 39228 17388 39284 17390
rect 39004 17276 39060 17332
rect 38220 16604 38276 16660
rect 37660 15708 37716 15764
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34412 14306 34468 14308
rect 34412 14254 34414 14306
rect 34414 14254 34466 14306
rect 34466 14254 34468 14306
rect 34412 14252 34468 14254
rect 34636 13746 34692 13748
rect 34636 13694 34638 13746
rect 34638 13694 34690 13746
rect 34690 13694 34692 13746
rect 34636 13692 34692 13694
rect 34300 13580 34356 13636
rect 34188 13522 34244 13524
rect 34188 13470 34190 13522
rect 34190 13470 34242 13522
rect 34242 13470 34244 13522
rect 34188 13468 34244 13470
rect 33964 12908 34020 12964
rect 33852 12684 33908 12740
rect 34300 11116 34356 11172
rect 32508 10668 32564 10724
rect 33404 10722 33460 10724
rect 33404 10670 33406 10722
rect 33406 10670 33458 10722
rect 33458 10670 33460 10722
rect 33404 10668 33460 10670
rect 33068 10610 33124 10612
rect 33068 10558 33070 10610
rect 33070 10558 33122 10610
rect 33122 10558 33124 10610
rect 33068 10556 33124 10558
rect 32956 10444 33012 10500
rect 32284 9884 32340 9940
rect 31836 8764 31892 8820
rect 31500 5740 31556 5796
rect 31612 8428 31668 8484
rect 31276 3836 31332 3892
rect 31724 6860 31780 6916
rect 32508 9042 32564 9044
rect 32508 8990 32510 9042
rect 32510 8990 32562 9042
rect 32562 8990 32564 9042
rect 32508 8988 32564 8990
rect 32172 8316 32228 8372
rect 32620 8258 32676 8260
rect 32620 8206 32622 8258
rect 32622 8206 32674 8258
rect 32674 8206 32676 8258
rect 32620 8204 32676 8206
rect 32956 9660 33012 9716
rect 33068 9436 33124 9492
rect 32732 8092 32788 8148
rect 32172 7868 32228 7924
rect 32284 7532 32340 7588
rect 31836 5516 31892 5572
rect 31836 4732 31892 4788
rect 32060 6188 32116 6244
rect 32060 6018 32116 6020
rect 32060 5966 32062 6018
rect 32062 5966 32114 6018
rect 32114 5966 32116 6018
rect 32060 5964 32116 5966
rect 32620 7474 32676 7476
rect 32620 7422 32622 7474
rect 32622 7422 32674 7474
rect 32674 7422 32676 7474
rect 32620 7420 32676 7422
rect 33404 9884 33460 9940
rect 33516 9826 33572 9828
rect 33516 9774 33518 9826
rect 33518 9774 33570 9826
rect 33570 9774 33572 9826
rect 33516 9772 33572 9774
rect 33404 8204 33460 8260
rect 33180 6524 33236 6580
rect 33516 8092 33572 8148
rect 33852 8092 33908 8148
rect 32956 5292 33012 5348
rect 33180 4956 33236 5012
rect 32060 4844 32116 4900
rect 32060 4450 32116 4452
rect 32060 4398 32062 4450
rect 32062 4398 32114 4450
rect 32114 4398 32116 4450
rect 32060 4396 32116 4398
rect 32172 4172 32228 4228
rect 33180 3948 33236 4004
rect 31612 1596 31668 1652
rect 33292 3164 33348 3220
rect 33404 4060 33460 4116
rect 33852 6972 33908 7028
rect 34188 10444 34244 10500
rect 34076 9548 34132 9604
rect 34076 7756 34132 7812
rect 34636 11564 34692 11620
rect 35308 13916 35364 13972
rect 35084 13468 35140 13524
rect 35756 14364 35812 14420
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 34972 12796 35028 12852
rect 35084 12572 35140 12628
rect 35532 12124 35588 12180
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35532 11564 35588 11620
rect 35084 11228 35140 11284
rect 35420 11340 35476 11396
rect 35084 10556 35140 10612
rect 35868 13916 35924 13972
rect 35756 13468 35812 13524
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35308 9714 35364 9716
rect 35308 9662 35310 9714
rect 35310 9662 35362 9714
rect 35362 9662 35364 9714
rect 35308 9660 35364 9662
rect 35196 9548 35252 9604
rect 35644 10332 35700 10388
rect 34524 9212 34580 9268
rect 34076 7084 34132 7140
rect 34076 6188 34132 6244
rect 33964 4508 34020 4564
rect 34748 8988 34804 9044
rect 34636 8092 34692 8148
rect 34636 6748 34692 6804
rect 33740 4226 33796 4228
rect 33740 4174 33742 4226
rect 33742 4174 33794 4226
rect 33794 4174 33796 4226
rect 33740 4172 33796 4174
rect 34636 5964 34692 6020
rect 34636 4732 34692 4788
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34860 4732 34916 4788
rect 35308 5180 35364 5236
rect 34860 4508 34916 4564
rect 34636 4396 34692 4452
rect 34972 4284 35028 4340
rect 35644 8204 35700 8260
rect 35756 11004 35812 11060
rect 37996 15314 38052 15316
rect 37996 15262 37998 15314
rect 37998 15262 38050 15314
rect 38050 15262 38052 15314
rect 37996 15260 38052 15262
rect 37100 14530 37156 14532
rect 37100 14478 37102 14530
rect 37102 14478 37154 14530
rect 37154 14478 37156 14530
rect 37100 14476 37156 14478
rect 37324 14476 37380 14532
rect 37100 14252 37156 14308
rect 36652 13692 36708 13748
rect 35980 11452 36036 11508
rect 37100 13692 37156 13748
rect 36764 13634 36820 13636
rect 36764 13582 36766 13634
rect 36766 13582 36818 13634
rect 36818 13582 36820 13634
rect 36764 13580 36820 13582
rect 36652 12908 36708 12964
rect 37100 13468 37156 13524
rect 36988 12850 37044 12852
rect 36988 12798 36990 12850
rect 36990 12798 37042 12850
rect 37042 12798 37044 12850
rect 36988 12796 37044 12798
rect 36540 12012 36596 12068
rect 36092 11170 36148 11172
rect 36092 11118 36094 11170
rect 36094 11118 36146 11170
rect 36146 11118 36148 11170
rect 36092 11116 36148 11118
rect 35980 9996 36036 10052
rect 35868 8764 35924 8820
rect 36316 10444 36372 10500
rect 36988 11788 37044 11844
rect 37436 14252 37492 14308
rect 37436 13468 37492 13524
rect 37548 13580 37604 13636
rect 37212 11788 37268 11844
rect 37324 12348 37380 12404
rect 36988 10892 37044 10948
rect 36540 10780 36596 10836
rect 37884 12796 37940 12852
rect 37660 12178 37716 12180
rect 37660 12126 37662 12178
rect 37662 12126 37714 12178
rect 37714 12126 37716 12178
rect 37660 12124 37716 12126
rect 38668 16882 38724 16884
rect 38668 16830 38670 16882
rect 38670 16830 38722 16882
rect 38722 16830 38724 16882
rect 38668 16828 38724 16830
rect 38332 16268 38388 16324
rect 38332 15708 38388 15764
rect 38332 15538 38388 15540
rect 38332 15486 38334 15538
rect 38334 15486 38386 15538
rect 38386 15486 38388 15538
rect 38332 15484 38388 15486
rect 39004 15202 39060 15204
rect 39004 15150 39006 15202
rect 39006 15150 39058 15202
rect 39058 15150 39060 15202
rect 39004 15148 39060 15150
rect 38444 14418 38500 14420
rect 38444 14366 38446 14418
rect 38446 14366 38498 14418
rect 38498 14366 38500 14418
rect 38444 14364 38500 14366
rect 39564 14252 39620 14308
rect 38220 13916 38276 13972
rect 38108 13692 38164 13748
rect 38108 13132 38164 13188
rect 38332 12962 38388 12964
rect 38332 12910 38334 12962
rect 38334 12910 38386 12962
rect 38386 12910 38388 12962
rect 38332 12908 38388 12910
rect 37996 11340 38052 11396
rect 37660 11282 37716 11284
rect 37660 11230 37662 11282
rect 37662 11230 37714 11282
rect 37714 11230 37716 11282
rect 37660 11228 37716 11230
rect 37548 11004 37604 11060
rect 38332 10892 38388 10948
rect 36988 10498 37044 10500
rect 36988 10446 36990 10498
rect 36990 10446 37042 10498
rect 37042 10446 37044 10498
rect 36988 10444 37044 10446
rect 37100 9996 37156 10052
rect 36428 9436 36484 9492
rect 36988 9436 37044 9492
rect 36988 8428 37044 8484
rect 37548 9660 37604 9716
rect 37772 9660 37828 9716
rect 37100 8370 37156 8372
rect 37100 8318 37102 8370
rect 37102 8318 37154 8370
rect 37154 8318 37156 8370
rect 37100 8316 37156 8318
rect 37212 8092 37268 8148
rect 35756 5852 35812 5908
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34972 3554 35028 3556
rect 34972 3502 34974 3554
rect 34974 3502 35026 3554
rect 35026 3502 35028 3554
rect 34972 3500 35028 3502
rect 33628 3052 33684 3108
rect 33516 2604 33572 2660
rect 36428 6748 36484 6804
rect 36092 4956 36148 5012
rect 37660 8370 37716 8372
rect 37660 8318 37662 8370
rect 37662 8318 37714 8370
rect 37714 8318 37716 8370
rect 37660 8316 37716 8318
rect 37884 8764 37940 8820
rect 37660 6748 37716 6804
rect 37548 6636 37604 6692
rect 37436 6412 37492 6468
rect 37324 6188 37380 6244
rect 37548 6018 37604 6020
rect 37548 5966 37550 6018
rect 37550 5966 37602 6018
rect 37602 5966 37604 6018
rect 37548 5964 37604 5966
rect 39452 14028 39508 14084
rect 38780 13132 38836 13188
rect 38444 10220 38500 10276
rect 38556 11340 38612 11396
rect 38780 10892 38836 10948
rect 39004 11282 39060 11284
rect 39004 11230 39006 11282
rect 39006 11230 39058 11282
rect 39058 11230 39060 11282
rect 39004 11228 39060 11230
rect 39228 12124 39284 12180
rect 38668 10556 38724 10612
rect 38332 9772 38388 9828
rect 38332 9100 38388 9156
rect 38220 8540 38276 8596
rect 38556 9772 38612 9828
rect 38668 9714 38724 9716
rect 38668 9662 38670 9714
rect 38670 9662 38722 9714
rect 38722 9662 38724 9714
rect 38668 9660 38724 9662
rect 38556 9548 38612 9604
rect 38668 9154 38724 9156
rect 38668 9102 38670 9154
rect 38670 9102 38722 9154
rect 38722 9102 38724 9154
rect 38668 9100 38724 9102
rect 38108 6524 38164 6580
rect 36988 5740 37044 5796
rect 36764 5628 36820 5684
rect 37324 5740 37380 5796
rect 38220 5964 38276 6020
rect 37212 5180 37268 5236
rect 36876 4844 36932 4900
rect 36316 4172 36372 4228
rect 36204 3612 36260 3668
rect 35980 3554 36036 3556
rect 35980 3502 35982 3554
rect 35982 3502 36034 3554
rect 36034 3502 36036 3554
rect 35980 3500 36036 3502
rect 37436 4956 37492 5012
rect 35756 1036 35812 1092
rect 38556 6636 38612 6692
rect 38332 5852 38388 5908
rect 38444 5740 38500 5796
rect 38332 5180 38388 5236
rect 39004 8540 39060 8596
rect 39564 13916 39620 13972
rect 39676 14140 39732 14196
rect 39900 14028 39956 14084
rect 40236 19516 40292 19572
rect 41468 22652 41524 22708
rect 42252 23772 42308 23828
rect 41916 23436 41972 23492
rect 41804 22988 41860 23044
rect 42028 23378 42084 23380
rect 42028 23326 42030 23378
rect 42030 23326 42082 23378
rect 42082 23326 42084 23378
rect 42028 23324 42084 23326
rect 42140 23266 42196 23268
rect 42140 23214 42142 23266
rect 42142 23214 42194 23266
rect 42194 23214 42196 23266
rect 42140 23212 42196 23214
rect 41916 22876 41972 22932
rect 41468 21474 41524 21476
rect 41468 21422 41470 21474
rect 41470 21422 41522 21474
rect 41522 21422 41524 21474
rect 41468 21420 41524 21422
rect 41692 20860 41748 20916
rect 41916 22428 41972 22484
rect 41020 19516 41076 19572
rect 41020 18396 41076 18452
rect 40236 17500 40292 17556
rect 41020 17554 41076 17556
rect 41020 17502 41022 17554
rect 41022 17502 41074 17554
rect 41074 17502 41076 17554
rect 41020 17500 41076 17502
rect 41580 19068 41636 19124
rect 42588 23772 42644 23828
rect 42364 23266 42420 23268
rect 42364 23214 42366 23266
rect 42366 23214 42418 23266
rect 42418 23214 42420 23266
rect 42364 23212 42420 23214
rect 43148 25340 43204 25396
rect 45164 29372 45220 29428
rect 46172 29426 46228 29428
rect 46172 29374 46174 29426
rect 46174 29374 46226 29426
rect 46226 29374 46228 29426
rect 46172 29372 46228 29374
rect 46060 29260 46116 29316
rect 46732 28364 46788 28420
rect 46060 27916 46116 27972
rect 45052 27746 45108 27748
rect 45052 27694 45054 27746
rect 45054 27694 45106 27746
rect 45106 27694 45108 27746
rect 45052 27692 45108 27694
rect 44828 27634 44884 27636
rect 44828 27582 44830 27634
rect 44830 27582 44882 27634
rect 44882 27582 44884 27634
rect 44828 27580 44884 27582
rect 45052 27356 45108 27412
rect 43596 26236 43652 26292
rect 44268 26290 44324 26292
rect 44268 26238 44270 26290
rect 44270 26238 44322 26290
rect 44322 26238 44324 26290
rect 44268 26236 44324 26238
rect 44604 26236 44660 26292
rect 44044 25676 44100 25732
rect 43820 25394 43876 25396
rect 43820 25342 43822 25394
rect 43822 25342 43874 25394
rect 43874 25342 43876 25394
rect 43820 25340 43876 25342
rect 43708 25228 43764 25284
rect 44716 26124 44772 26180
rect 44828 25676 44884 25732
rect 45164 25900 45220 25956
rect 44604 25340 44660 25396
rect 45724 27580 45780 27636
rect 45724 27132 45780 27188
rect 45948 27580 46004 27636
rect 45836 26908 45892 26964
rect 45388 26572 45444 26628
rect 45276 25564 45332 25620
rect 45388 25506 45444 25508
rect 45388 25454 45390 25506
rect 45390 25454 45442 25506
rect 45442 25454 45444 25506
rect 45388 25452 45444 25454
rect 45164 25228 45220 25284
rect 45052 24892 45108 24948
rect 45500 24780 45556 24836
rect 43820 23996 43876 24052
rect 44492 23884 44548 23940
rect 44604 23772 44660 23828
rect 44828 24332 44884 24388
rect 42812 23548 42868 23604
rect 43372 23548 43428 23604
rect 43708 23436 43764 23492
rect 45388 23996 45444 24052
rect 45164 23772 45220 23828
rect 45052 23436 45108 23492
rect 42588 22652 42644 22708
rect 42700 22540 42756 22596
rect 42028 21586 42084 21588
rect 42028 21534 42030 21586
rect 42030 21534 42082 21586
rect 42082 21534 42084 21586
rect 42028 21532 42084 21534
rect 42028 19516 42084 19572
rect 42140 19404 42196 19460
rect 41804 18396 41860 18452
rect 42364 19292 42420 19348
rect 41916 18284 41972 18340
rect 42588 18620 42644 18676
rect 42812 19122 42868 19124
rect 42812 19070 42814 19122
rect 42814 19070 42866 19122
rect 42866 19070 42868 19122
rect 42812 19068 42868 19070
rect 43484 22876 43540 22932
rect 43372 22204 43428 22260
rect 43708 22652 43764 22708
rect 46172 27692 46228 27748
rect 46172 27020 46228 27076
rect 46732 27132 46788 27188
rect 46508 25900 46564 25956
rect 46396 24946 46452 24948
rect 46396 24894 46398 24946
rect 46398 24894 46450 24946
rect 46450 24894 46452 24946
rect 46396 24892 46452 24894
rect 46620 25228 46676 25284
rect 46508 24780 46564 24836
rect 45388 23548 45444 23604
rect 45276 23154 45332 23156
rect 45276 23102 45278 23154
rect 45278 23102 45330 23154
rect 45330 23102 45332 23154
rect 45276 23100 45332 23102
rect 45388 22146 45444 22148
rect 45388 22094 45390 22146
rect 45390 22094 45442 22146
rect 45442 22094 45444 22146
rect 45388 22092 45444 22094
rect 43932 21196 43988 21252
rect 44044 20636 44100 20692
rect 44268 20748 44324 20804
rect 45388 20636 45444 20692
rect 43260 19516 43316 19572
rect 43372 19292 43428 19348
rect 43148 19068 43204 19124
rect 43148 18338 43204 18340
rect 43148 18286 43150 18338
rect 43150 18286 43202 18338
rect 43202 18286 43204 18338
rect 43148 18284 43204 18286
rect 42364 17724 42420 17780
rect 41580 17612 41636 17668
rect 40908 16210 40964 16212
rect 40908 16158 40910 16210
rect 40910 16158 40962 16210
rect 40962 16158 40964 16210
rect 40908 16156 40964 16158
rect 40572 16098 40628 16100
rect 40572 16046 40574 16098
rect 40574 16046 40626 16098
rect 40626 16046 40628 16098
rect 40572 16044 40628 16046
rect 40348 15874 40404 15876
rect 40348 15822 40350 15874
rect 40350 15822 40402 15874
rect 40402 15822 40404 15874
rect 40348 15820 40404 15822
rect 40796 15708 40852 15764
rect 41356 16268 41412 16324
rect 41692 16156 41748 16212
rect 42140 16268 42196 16324
rect 41804 16044 41860 16100
rect 41692 15708 41748 15764
rect 42140 14700 42196 14756
rect 39452 11452 39508 11508
rect 39564 11788 39620 11844
rect 39340 11282 39396 11284
rect 39340 11230 39342 11282
rect 39342 11230 39394 11282
rect 39394 11230 39396 11282
rect 39340 11228 39396 11230
rect 39676 10722 39732 10724
rect 39676 10670 39678 10722
rect 39678 10670 39730 10722
rect 39730 10670 39732 10722
rect 39676 10668 39732 10670
rect 39452 9996 39508 10052
rect 39340 9548 39396 9604
rect 39676 9266 39732 9268
rect 39676 9214 39678 9266
rect 39678 9214 39730 9266
rect 39730 9214 39732 9266
rect 39676 9212 39732 9214
rect 39116 8428 39172 8484
rect 39228 8316 39284 8372
rect 39004 7084 39060 7140
rect 39004 6860 39060 6916
rect 39228 7196 39284 7252
rect 39340 7084 39396 7140
rect 39564 8652 39620 8708
rect 39340 6860 39396 6916
rect 39004 6524 39060 6580
rect 39228 6412 39284 6468
rect 39116 6076 39172 6132
rect 39564 7868 39620 7924
rect 39564 6972 39620 7028
rect 39676 6748 39732 6804
rect 39788 8540 39844 8596
rect 39564 6690 39620 6692
rect 39564 6638 39566 6690
rect 39566 6638 39618 6690
rect 39618 6638 39620 6690
rect 39564 6636 39620 6638
rect 39452 6300 39508 6356
rect 40012 12124 40068 12180
rect 40124 14028 40180 14084
rect 43372 18620 43428 18676
rect 43708 19180 43764 19236
rect 45388 18956 45444 19012
rect 44268 18396 44324 18452
rect 43260 16380 43316 16436
rect 42812 16268 42868 16324
rect 42364 14588 42420 14644
rect 41020 13746 41076 13748
rect 41020 13694 41022 13746
rect 41022 13694 41074 13746
rect 41074 13694 41076 13746
rect 41020 13692 41076 13694
rect 41692 13692 41748 13748
rect 40348 13634 40404 13636
rect 40348 13582 40350 13634
rect 40350 13582 40402 13634
rect 40402 13582 40404 13634
rect 40348 13580 40404 13582
rect 40684 13468 40740 13524
rect 40908 12178 40964 12180
rect 40908 12126 40910 12178
rect 40910 12126 40962 12178
rect 40962 12126 40964 12178
rect 40908 12124 40964 12126
rect 40124 11564 40180 11620
rect 40348 11954 40404 11956
rect 40348 11902 40350 11954
rect 40350 11902 40402 11954
rect 40402 11902 40404 11954
rect 40348 11900 40404 11902
rect 40236 11452 40292 11508
rect 40012 11340 40068 11396
rect 40236 11116 40292 11172
rect 40124 10892 40180 10948
rect 40012 9660 40068 9716
rect 39900 8092 39956 8148
rect 39900 7474 39956 7476
rect 39900 7422 39902 7474
rect 39902 7422 39954 7474
rect 39954 7422 39956 7474
rect 39900 7420 39956 7422
rect 40236 10332 40292 10388
rect 40572 10444 40628 10500
rect 40460 9884 40516 9940
rect 41244 11282 41300 11284
rect 41244 11230 41246 11282
rect 41246 11230 41298 11282
rect 41298 11230 41300 11282
rect 41244 11228 41300 11230
rect 40796 9996 40852 10052
rect 40908 9884 40964 9940
rect 40908 9660 40964 9716
rect 40348 8428 40404 8484
rect 40236 7698 40292 7700
rect 40236 7646 40238 7698
rect 40238 7646 40290 7698
rect 40290 7646 40292 7698
rect 40236 7644 40292 7646
rect 40012 7196 40068 7252
rect 40124 6412 40180 6468
rect 39900 5906 39956 5908
rect 39900 5854 39902 5906
rect 39902 5854 39954 5906
rect 39954 5854 39956 5906
rect 39900 5852 39956 5854
rect 40012 5628 40068 5684
rect 38892 5180 38948 5236
rect 39900 5234 39956 5236
rect 39900 5182 39902 5234
rect 39902 5182 39954 5234
rect 39954 5182 39956 5234
rect 39900 5180 39956 5182
rect 39452 4732 39508 4788
rect 39116 4620 39172 4676
rect 39340 4562 39396 4564
rect 39340 4510 39342 4562
rect 39342 4510 39394 4562
rect 39394 4510 39396 4562
rect 39340 4508 39396 4510
rect 39004 4060 39060 4116
rect 38556 3500 38612 3556
rect 38444 2492 38500 2548
rect 38780 3388 38836 3444
rect 40236 6076 40292 6132
rect 40236 5906 40292 5908
rect 40236 5854 40238 5906
rect 40238 5854 40290 5906
rect 40290 5854 40292 5906
rect 40236 5852 40292 5854
rect 40236 5628 40292 5684
rect 40236 5068 40292 5124
rect 41356 10610 41412 10612
rect 41356 10558 41358 10610
rect 41358 10558 41410 10610
rect 41410 10558 41412 10610
rect 41356 10556 41412 10558
rect 41132 10498 41188 10500
rect 41132 10446 41134 10498
rect 41134 10446 41186 10498
rect 41186 10446 41188 10498
rect 41132 10444 41188 10446
rect 41356 9884 41412 9940
rect 40572 6860 40628 6916
rect 40684 6076 40740 6132
rect 41132 7644 41188 7700
rect 41580 10386 41636 10388
rect 41580 10334 41582 10386
rect 41582 10334 41634 10386
rect 41634 10334 41636 10386
rect 41580 10332 41636 10334
rect 42588 14028 42644 14084
rect 42140 13970 42196 13972
rect 42140 13918 42142 13970
rect 42142 13918 42194 13970
rect 42194 13918 42196 13970
rect 42140 13916 42196 13918
rect 42812 13020 42868 13076
rect 41804 12348 41860 12404
rect 42364 12290 42420 12292
rect 42364 12238 42366 12290
rect 42366 12238 42418 12290
rect 42418 12238 42420 12290
rect 42364 12236 42420 12238
rect 41916 12178 41972 12180
rect 41916 12126 41918 12178
rect 41918 12126 41970 12178
rect 41970 12126 41972 12178
rect 41916 12124 41972 12126
rect 43148 12460 43204 12516
rect 42812 11788 42868 11844
rect 42924 11900 42980 11956
rect 41692 9884 41748 9940
rect 41356 8652 41412 8708
rect 41356 8258 41412 8260
rect 41356 8206 41358 8258
rect 41358 8206 41410 8258
rect 41410 8206 41412 8258
rect 41356 8204 41412 8206
rect 41020 7250 41076 7252
rect 41020 7198 41022 7250
rect 41022 7198 41074 7250
rect 41074 7198 41076 7250
rect 41020 7196 41076 7198
rect 41020 6972 41076 7028
rect 41132 6636 41188 6692
rect 41580 7420 41636 7476
rect 41580 6690 41636 6692
rect 41580 6638 41582 6690
rect 41582 6638 41634 6690
rect 41634 6638 41636 6690
rect 41580 6636 41636 6638
rect 41020 5964 41076 6020
rect 40908 5906 40964 5908
rect 40908 5854 40910 5906
rect 40910 5854 40962 5906
rect 40962 5854 40964 5906
rect 40908 5852 40964 5854
rect 41468 6076 41524 6132
rect 40796 4844 40852 4900
rect 41132 5292 41188 5348
rect 41244 5180 41300 5236
rect 41356 5068 41412 5124
rect 41468 4844 41524 4900
rect 41468 4396 41524 4452
rect 40796 3666 40852 3668
rect 40796 3614 40798 3666
rect 40798 3614 40850 3666
rect 40850 3614 40852 3666
rect 40796 3612 40852 3614
rect 40460 2828 40516 2884
rect 41916 10780 41972 10836
rect 42140 10722 42196 10724
rect 42140 10670 42142 10722
rect 42142 10670 42194 10722
rect 42194 10670 42196 10722
rect 42140 10668 42196 10670
rect 42476 11340 42532 11396
rect 42700 11564 42756 11620
rect 42588 11282 42644 11284
rect 42588 11230 42590 11282
rect 42590 11230 42642 11282
rect 42642 11230 42644 11282
rect 42588 11228 42644 11230
rect 43036 11676 43092 11732
rect 42588 10834 42644 10836
rect 42588 10782 42590 10834
rect 42590 10782 42642 10834
rect 42642 10782 42644 10834
rect 42588 10780 42644 10782
rect 42812 11452 42868 11508
rect 42476 10444 42532 10500
rect 42252 10108 42308 10164
rect 42028 8204 42084 8260
rect 41804 6636 41860 6692
rect 41916 5964 41972 6020
rect 41692 4226 41748 4228
rect 41692 4174 41694 4226
rect 41694 4174 41746 4226
rect 41746 4174 41748 4226
rect 41692 4172 41748 4174
rect 42252 6524 42308 6580
rect 42364 6300 42420 6356
rect 42252 5122 42308 5124
rect 42252 5070 42254 5122
rect 42254 5070 42306 5122
rect 42306 5070 42308 5122
rect 42252 5068 42308 5070
rect 42140 3948 42196 4004
rect 41804 3388 41860 3444
rect 42588 4956 42644 5012
rect 42588 4562 42644 4564
rect 42588 4510 42590 4562
rect 42590 4510 42642 4562
rect 42642 4510 42644 4562
rect 42588 4508 42644 4510
rect 42812 7980 42868 8036
rect 42812 5794 42868 5796
rect 42812 5742 42814 5794
rect 42814 5742 42866 5794
rect 42866 5742 42868 5794
rect 42812 5740 42868 5742
rect 43036 10892 43092 10948
rect 43036 10108 43092 10164
rect 43148 10386 43204 10388
rect 43148 10334 43150 10386
rect 43150 10334 43202 10386
rect 43202 10334 43204 10386
rect 43148 10332 43204 10334
rect 43820 15820 43876 15876
rect 46732 24108 46788 24164
rect 46060 23996 46116 24052
rect 46732 23938 46788 23940
rect 46732 23886 46734 23938
rect 46734 23886 46786 23938
rect 46786 23886 46788 23938
rect 46732 23884 46788 23886
rect 46284 23826 46340 23828
rect 46284 23774 46286 23826
rect 46286 23774 46338 23826
rect 46338 23774 46340 23826
rect 46284 23772 46340 23774
rect 46396 23660 46452 23716
rect 45612 21644 45668 21700
rect 46284 23548 46340 23604
rect 45612 20860 45668 20916
rect 45836 20860 45892 20916
rect 45948 20802 46004 20804
rect 45948 20750 45950 20802
rect 45950 20750 46002 20802
rect 46002 20750 46004 20802
rect 45948 20748 46004 20750
rect 45612 20188 45668 20244
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 48300 30940 48356 30996
rect 47292 29314 47348 29316
rect 47292 29262 47294 29314
rect 47294 29262 47346 29314
rect 47346 29262 47348 29314
rect 47292 29260 47348 29262
rect 46956 23266 47012 23268
rect 46956 23214 46958 23266
rect 46958 23214 47010 23266
rect 47010 23214 47012 23266
rect 46956 23212 47012 23214
rect 46620 21698 46676 21700
rect 46620 21646 46622 21698
rect 46622 21646 46674 21698
rect 46674 21646 46676 21698
rect 46620 21644 46676 21646
rect 47964 26908 48020 26964
rect 47852 26796 47908 26852
rect 47292 25676 47348 25732
rect 47740 25228 47796 25284
rect 48076 26236 48132 26292
rect 48188 25788 48244 25844
rect 48076 25676 48132 25732
rect 47180 24108 47236 24164
rect 47628 23996 47684 24052
rect 47292 23938 47348 23940
rect 47292 23886 47294 23938
rect 47294 23886 47346 23938
rect 47346 23886 47348 23938
rect 47292 23884 47348 23886
rect 47180 23436 47236 23492
rect 47628 23100 47684 23156
rect 47852 23212 47908 23268
rect 47404 22764 47460 22820
rect 47180 22540 47236 22596
rect 47068 22482 47124 22484
rect 47068 22430 47070 22482
rect 47070 22430 47122 22482
rect 47122 22430 47124 22482
rect 47068 22428 47124 22430
rect 46844 22092 46900 22148
rect 46844 21644 46900 21700
rect 46732 20748 46788 20804
rect 46844 20690 46900 20692
rect 46844 20638 46846 20690
rect 46846 20638 46898 20690
rect 46898 20638 46900 20690
rect 46844 20636 46900 20638
rect 48188 22988 48244 23044
rect 48076 22764 48132 22820
rect 47068 21474 47124 21476
rect 47068 21422 47070 21474
rect 47070 21422 47122 21474
rect 47122 21422 47124 21474
rect 47068 21420 47124 21422
rect 47404 21084 47460 21140
rect 47740 20860 47796 20916
rect 47068 20578 47124 20580
rect 47068 20526 47070 20578
rect 47070 20526 47122 20578
rect 47122 20526 47124 20578
rect 47068 20524 47124 20526
rect 46284 19628 46340 19684
rect 46060 19180 46116 19236
rect 46284 18956 46340 19012
rect 46844 18732 46900 18788
rect 45724 17836 45780 17892
rect 44268 15538 44324 15540
rect 44268 15486 44270 15538
rect 44270 15486 44322 15538
rect 44322 15486 44324 15538
rect 44268 15484 44324 15486
rect 45276 15484 45332 15540
rect 45836 17666 45892 17668
rect 45836 17614 45838 17666
rect 45838 17614 45890 17666
rect 45890 17614 45892 17666
rect 45836 17612 45892 17614
rect 46284 17612 46340 17668
rect 45724 17164 45780 17220
rect 46172 17164 46228 17220
rect 45948 16994 46004 16996
rect 45948 16942 45950 16994
rect 45950 16942 46002 16994
rect 46002 16942 46004 16994
rect 45948 16940 46004 16942
rect 46060 16828 46116 16884
rect 44940 14476 44996 14532
rect 44492 14028 44548 14084
rect 43932 13074 43988 13076
rect 43932 13022 43934 13074
rect 43934 13022 43986 13074
rect 43986 13022 43988 13074
rect 43932 13020 43988 13022
rect 45388 14700 45444 14756
rect 45164 13356 45220 13412
rect 44828 12796 44884 12852
rect 45836 12796 45892 12852
rect 43820 12402 43876 12404
rect 43820 12350 43822 12402
rect 43822 12350 43874 12402
rect 43874 12350 43876 12402
rect 43820 12348 43876 12350
rect 43708 11954 43764 11956
rect 43708 11902 43710 11954
rect 43710 11902 43762 11954
rect 43762 11902 43764 11954
rect 43708 11900 43764 11902
rect 43596 11788 43652 11844
rect 43596 10556 43652 10612
rect 43372 8988 43428 9044
rect 42924 5628 42980 5684
rect 42924 5180 42980 5236
rect 43036 8316 43092 8372
rect 43148 6524 43204 6580
rect 42924 3554 42980 3556
rect 42924 3502 42926 3554
rect 42926 3502 42978 3554
rect 42978 3502 42980 3554
rect 42924 3500 42980 3502
rect 43372 5964 43428 6020
rect 43596 10108 43652 10164
rect 44044 12012 44100 12068
rect 43932 11004 43988 11060
rect 44940 11228 44996 11284
rect 44156 11004 44212 11060
rect 43932 10108 43988 10164
rect 44268 10610 44324 10612
rect 44268 10558 44270 10610
rect 44270 10558 44322 10610
rect 44322 10558 44324 10610
rect 44268 10556 44324 10558
rect 44156 10220 44212 10276
rect 43820 9996 43876 10052
rect 43820 8316 43876 8372
rect 43260 5234 43316 5236
rect 43260 5182 43262 5234
rect 43262 5182 43314 5234
rect 43314 5182 43316 5234
rect 43260 5180 43316 5182
rect 43148 3276 43204 3332
rect 42476 2268 42532 2324
rect 42252 924 42308 980
rect 44156 9772 44212 9828
rect 44604 10610 44660 10612
rect 44604 10558 44606 10610
rect 44606 10558 44658 10610
rect 44658 10558 44660 10610
rect 44604 10556 44660 10558
rect 44716 10444 44772 10500
rect 44492 9996 44548 10052
rect 44716 9996 44772 10052
rect 45836 12460 45892 12516
rect 45612 12402 45668 12404
rect 45612 12350 45614 12402
rect 45614 12350 45666 12402
rect 45666 12350 45668 12402
rect 45612 12348 45668 12350
rect 45612 11788 45668 11844
rect 45836 11788 45892 11844
rect 46508 18396 46564 18452
rect 46956 17164 47012 17220
rect 46508 16940 46564 16996
rect 46508 16156 46564 16212
rect 47292 20188 47348 20244
rect 47292 17666 47348 17668
rect 47292 17614 47294 17666
rect 47294 17614 47346 17666
rect 47346 17614 47348 17666
rect 47292 17612 47348 17614
rect 48188 21420 48244 21476
rect 49756 30716 49812 30772
rect 49308 29932 49364 29988
rect 49084 29314 49140 29316
rect 49084 29262 49086 29314
rect 49086 29262 49138 29314
rect 49138 29262 49140 29314
rect 49084 29260 49140 29262
rect 49420 29036 49476 29092
rect 49308 28924 49364 28980
rect 48188 20690 48244 20692
rect 48188 20638 48190 20690
rect 48190 20638 48242 20690
rect 48242 20638 48244 20690
rect 48188 20636 48244 20638
rect 48524 28476 48580 28532
rect 49420 28588 49476 28644
rect 48860 27634 48916 27636
rect 48860 27582 48862 27634
rect 48862 27582 48914 27634
rect 48914 27582 48916 27634
rect 48860 27580 48916 27582
rect 48636 27468 48692 27524
rect 48748 26962 48804 26964
rect 48748 26910 48750 26962
rect 48750 26910 48802 26962
rect 48802 26910 48804 26962
rect 48748 26908 48804 26910
rect 48860 26514 48916 26516
rect 48860 26462 48862 26514
rect 48862 26462 48914 26514
rect 48914 26462 48916 26514
rect 48860 26460 48916 26462
rect 49420 27020 49476 27076
rect 48860 26236 48916 26292
rect 48636 26012 48692 26068
rect 48636 24892 48692 24948
rect 48972 26012 49028 26068
rect 49084 26124 49140 26180
rect 48972 25618 49028 25620
rect 48972 25566 48974 25618
rect 48974 25566 49026 25618
rect 49026 25566 49028 25618
rect 48972 25564 49028 25566
rect 49420 26348 49476 26404
rect 49196 24556 49252 24612
rect 48636 23548 48692 23604
rect 49420 24108 49476 24164
rect 49084 22876 49140 22932
rect 48748 21644 48804 21700
rect 48860 21474 48916 21476
rect 48860 21422 48862 21474
rect 48862 21422 48914 21474
rect 48914 21422 48916 21474
rect 48860 21420 48916 21422
rect 48748 21196 48804 21252
rect 47964 20076 48020 20132
rect 47516 18284 47572 18340
rect 47740 18450 47796 18452
rect 47740 18398 47742 18450
rect 47742 18398 47794 18450
rect 47794 18398 47796 18450
rect 47740 18396 47796 18398
rect 49084 19852 49140 19908
rect 48188 18620 48244 18676
rect 48076 18396 48132 18452
rect 48972 19234 49028 19236
rect 48972 19182 48974 19234
rect 48974 19182 49026 19234
rect 49026 19182 49028 19234
rect 48972 19180 49028 19182
rect 49644 28530 49700 28532
rect 49644 28478 49646 28530
rect 49646 28478 49698 28530
rect 49698 28478 49700 28530
rect 49644 28476 49700 28478
rect 49644 27858 49700 27860
rect 49644 27806 49646 27858
rect 49646 27806 49698 27858
rect 49698 27806 49700 27858
rect 49644 27804 49700 27806
rect 51100 29932 51156 29988
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50988 29260 51044 29316
rect 50540 29036 50596 29092
rect 49868 28476 49924 28532
rect 49980 28418 50036 28420
rect 49980 28366 49982 28418
rect 49982 28366 50034 28418
rect 50034 28366 50036 28418
rect 49980 28364 50036 28366
rect 50316 28028 50372 28084
rect 50316 27858 50372 27860
rect 50316 27806 50318 27858
rect 50318 27806 50370 27858
rect 50370 27806 50372 27858
rect 50316 27804 50372 27806
rect 50092 27580 50148 27636
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50540 28028 50596 28084
rect 50988 28476 51044 28532
rect 49756 27244 49812 27300
rect 50428 27244 50484 27300
rect 50204 26908 50260 26964
rect 49756 26572 49812 26628
rect 49644 26402 49700 26404
rect 49644 26350 49646 26402
rect 49646 26350 49698 26402
rect 49698 26350 49700 26402
rect 49644 26348 49700 26350
rect 49644 25676 49700 25732
rect 49532 23042 49588 23044
rect 49532 22990 49534 23042
rect 49534 22990 49586 23042
rect 49586 22990 49588 23042
rect 49532 22988 49588 22990
rect 49532 22764 49588 22820
rect 49196 19628 49252 19684
rect 49084 19068 49140 19124
rect 49196 19180 49252 19236
rect 48412 18732 48468 18788
rect 48860 18450 48916 18452
rect 48860 18398 48862 18450
rect 48862 18398 48914 18450
rect 48914 18398 48916 18450
rect 48860 18396 48916 18398
rect 48300 18060 48356 18116
rect 48412 17948 48468 18004
rect 47404 17164 47460 17220
rect 47292 16716 47348 16772
rect 47628 16994 47684 16996
rect 47628 16942 47630 16994
rect 47630 16942 47682 16994
rect 47682 16942 47684 16994
rect 47628 16940 47684 16942
rect 47852 16882 47908 16884
rect 47852 16830 47854 16882
rect 47854 16830 47906 16882
rect 47906 16830 47908 16882
rect 47852 16828 47908 16830
rect 48076 16882 48132 16884
rect 48076 16830 48078 16882
rect 48078 16830 48130 16882
rect 48130 16830 48132 16882
rect 48076 16828 48132 16830
rect 48300 16492 48356 16548
rect 48860 17666 48916 17668
rect 48860 17614 48862 17666
rect 48862 17614 48914 17666
rect 48914 17614 48916 17666
rect 48860 17612 48916 17614
rect 49868 26124 49924 26180
rect 50764 27634 50820 27636
rect 50764 27582 50766 27634
rect 50766 27582 50818 27634
rect 50818 27582 50820 27634
rect 50764 27580 50820 27582
rect 50988 27580 51044 27636
rect 51996 30380 52052 30436
rect 51772 29314 51828 29316
rect 51772 29262 51774 29314
rect 51774 29262 51826 29314
rect 51826 29262 51828 29314
rect 51772 29260 51828 29262
rect 51436 28028 51492 28084
rect 51100 27468 51156 27524
rect 50988 27244 51044 27300
rect 51772 27746 51828 27748
rect 51772 27694 51774 27746
rect 51774 27694 51826 27746
rect 51826 27694 51828 27746
rect 51772 27692 51828 27694
rect 51212 27244 51268 27300
rect 51548 27468 51604 27524
rect 50652 26796 50708 26852
rect 51436 27074 51492 27076
rect 51436 27022 51438 27074
rect 51438 27022 51490 27074
rect 51490 27022 51492 27074
rect 51436 27020 51492 27022
rect 50988 26684 51044 26740
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50092 25506 50148 25508
rect 50092 25454 50094 25506
rect 50094 25454 50146 25506
rect 50146 25454 50148 25506
rect 50092 25452 50148 25454
rect 49868 24610 49924 24612
rect 49868 24558 49870 24610
rect 49870 24558 49922 24610
rect 49922 24558 49924 24610
rect 49868 24556 49924 24558
rect 49868 22428 49924 22484
rect 50316 26460 50372 26516
rect 50764 26460 50820 26516
rect 50652 26348 50708 26404
rect 50876 26290 50932 26292
rect 50876 26238 50878 26290
rect 50878 26238 50930 26290
rect 50930 26238 50932 26290
rect 50876 26236 50932 26238
rect 50876 26012 50932 26068
rect 50764 25564 50820 25620
rect 50540 25506 50596 25508
rect 50540 25454 50542 25506
rect 50542 25454 50594 25506
rect 50594 25454 50596 25506
rect 50540 25452 50596 25454
rect 50316 25394 50372 25396
rect 50316 25342 50318 25394
rect 50318 25342 50370 25394
rect 50370 25342 50372 25394
rect 50316 25340 50372 25342
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50764 24892 50820 24948
rect 51100 25452 51156 25508
rect 51772 27298 51828 27300
rect 51772 27246 51774 27298
rect 51774 27246 51826 27298
rect 51826 27246 51828 27298
rect 51772 27244 51828 27246
rect 54796 30210 54852 30212
rect 54796 30158 54798 30210
rect 54798 30158 54850 30210
rect 54850 30158 54852 30210
rect 54796 30156 54852 30158
rect 52780 29986 52836 29988
rect 52780 29934 52782 29986
rect 52782 29934 52834 29986
rect 52834 29934 52836 29986
rect 52780 29932 52836 29934
rect 54124 29986 54180 29988
rect 54124 29934 54126 29986
rect 54126 29934 54178 29986
rect 54178 29934 54180 29986
rect 54124 29932 54180 29934
rect 52108 29484 52164 29540
rect 54572 29538 54628 29540
rect 54572 29486 54574 29538
rect 54574 29486 54626 29538
rect 54626 29486 54628 29538
rect 54572 29484 54628 29486
rect 53900 29314 53956 29316
rect 53900 29262 53902 29314
rect 53902 29262 53954 29314
rect 53954 29262 53956 29314
rect 53900 29260 53956 29262
rect 53788 29036 53844 29092
rect 53004 28642 53060 28644
rect 53004 28590 53006 28642
rect 53006 28590 53058 28642
rect 53058 28590 53060 28642
rect 53004 28588 53060 28590
rect 53452 28642 53508 28644
rect 53452 28590 53454 28642
rect 53454 28590 53506 28642
rect 53506 28590 53508 28642
rect 53452 28588 53508 28590
rect 53228 27858 53284 27860
rect 53228 27806 53230 27858
rect 53230 27806 53282 27858
rect 53282 27806 53284 27858
rect 53228 27804 53284 27806
rect 51996 27244 52052 27300
rect 52108 27580 52164 27636
rect 52668 27580 52724 27636
rect 51884 26684 51940 26740
rect 52108 26066 52164 26068
rect 52108 26014 52110 26066
rect 52110 26014 52162 26066
rect 52162 26014 52164 26066
rect 52108 26012 52164 26014
rect 51660 25676 51716 25732
rect 51324 25004 51380 25060
rect 51548 24892 51604 24948
rect 52108 25340 52164 25396
rect 50428 24722 50484 24724
rect 50428 24670 50430 24722
rect 50430 24670 50482 24722
rect 50482 24670 50484 24722
rect 50428 24668 50484 24670
rect 50204 24108 50260 24164
rect 50428 24162 50484 24164
rect 50428 24110 50430 24162
rect 50430 24110 50482 24162
rect 50482 24110 50484 24162
rect 50428 24108 50484 24110
rect 51212 24556 51268 24612
rect 51660 24610 51716 24612
rect 51660 24558 51662 24610
rect 51662 24558 51714 24610
rect 51714 24558 51716 24610
rect 51660 24556 51716 24558
rect 50988 24220 51044 24276
rect 50764 23938 50820 23940
rect 50764 23886 50766 23938
rect 50766 23886 50818 23938
rect 50818 23886 50820 23938
rect 50764 23884 50820 23886
rect 52556 24498 52612 24500
rect 52556 24446 52558 24498
rect 52558 24446 52610 24498
rect 52610 24446 52612 24498
rect 52556 24444 52612 24446
rect 51548 24108 51604 24164
rect 51772 23938 51828 23940
rect 51772 23886 51774 23938
rect 51774 23886 51826 23938
rect 51826 23886 51828 23938
rect 51772 23884 51828 23886
rect 50316 23212 50372 23268
rect 50204 22204 50260 22260
rect 50204 21756 50260 21812
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50876 23100 50932 23156
rect 50652 22876 50708 22932
rect 50876 22876 50932 22932
rect 50540 22764 50596 22820
rect 51324 23660 51380 23716
rect 51212 23548 51268 23604
rect 51436 23548 51492 23604
rect 51324 22988 51380 23044
rect 51548 23436 51604 23492
rect 51996 23660 52052 23716
rect 51660 23324 51716 23380
rect 51772 23548 51828 23604
rect 51324 22594 51380 22596
rect 51324 22542 51326 22594
rect 51326 22542 51378 22594
rect 51378 22542 51380 22594
rect 51324 22540 51380 22542
rect 51548 22428 51604 22484
rect 50988 22370 51044 22372
rect 50988 22318 50990 22370
rect 50990 22318 51042 22370
rect 51042 22318 51044 22370
rect 50988 22316 51044 22318
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50204 21026 50260 21028
rect 50204 20974 50206 21026
rect 50206 20974 50258 21026
rect 50258 20974 50260 21026
rect 50204 20972 50260 20974
rect 49532 19010 49588 19012
rect 49532 18958 49534 19010
rect 49534 18958 49586 19010
rect 49586 18958 49588 19010
rect 49532 18956 49588 18958
rect 49980 19010 50036 19012
rect 49980 18958 49982 19010
rect 49982 18958 50034 19010
rect 50034 18958 50036 19010
rect 49980 18956 50036 18958
rect 49756 18620 49812 18676
rect 49420 18284 49476 18340
rect 49308 18060 49364 18116
rect 49532 17666 49588 17668
rect 49532 17614 49534 17666
rect 49534 17614 49586 17666
rect 49586 17614 49588 17666
rect 49532 17612 49588 17614
rect 49868 17554 49924 17556
rect 49868 17502 49870 17554
rect 49870 17502 49922 17554
rect 49922 17502 49924 17554
rect 49868 17500 49924 17502
rect 48412 17052 48468 17108
rect 49868 17106 49924 17108
rect 49868 17054 49870 17106
rect 49870 17054 49922 17106
rect 49922 17054 49924 17106
rect 49868 17052 49924 17054
rect 48524 16940 48580 16996
rect 47180 15820 47236 15876
rect 47404 15874 47460 15876
rect 47404 15822 47406 15874
rect 47406 15822 47458 15874
rect 47458 15822 47460 15874
rect 47404 15820 47460 15822
rect 46396 14924 46452 14980
rect 48076 15708 48132 15764
rect 46396 13970 46452 13972
rect 46396 13918 46398 13970
rect 46398 13918 46450 13970
rect 46450 13918 46452 13970
rect 46396 13916 46452 13918
rect 46396 12460 46452 12516
rect 45164 11116 45220 11172
rect 44828 9884 44884 9940
rect 45164 9938 45220 9940
rect 45164 9886 45166 9938
rect 45166 9886 45218 9938
rect 45218 9886 45220 9938
rect 45164 9884 45220 9886
rect 45836 11170 45892 11172
rect 45836 11118 45838 11170
rect 45838 11118 45890 11170
rect 45890 11118 45892 11170
rect 45836 11116 45892 11118
rect 46172 12178 46228 12180
rect 46172 12126 46174 12178
rect 46174 12126 46226 12178
rect 46226 12126 46228 12178
rect 46172 12124 46228 12126
rect 46060 10780 46116 10836
rect 45500 9996 45556 10052
rect 44716 9100 44772 9156
rect 45500 9660 45556 9716
rect 44380 8204 44436 8260
rect 45052 8258 45108 8260
rect 45052 8206 45054 8258
rect 45054 8206 45106 8258
rect 45106 8206 45108 8258
rect 45052 8204 45108 8206
rect 43708 7532 43764 7588
rect 43708 6636 43764 6692
rect 44156 6578 44212 6580
rect 44156 6526 44158 6578
rect 44158 6526 44210 6578
rect 44210 6526 44212 6578
rect 44156 6524 44212 6526
rect 43932 6412 43988 6468
rect 43596 4956 43652 5012
rect 44940 7644 44996 7700
rect 44380 6748 44436 6804
rect 45500 9324 45556 9380
rect 45276 8316 45332 8372
rect 45276 8034 45332 8036
rect 45276 7982 45278 8034
rect 45278 7982 45330 8034
rect 45330 7982 45332 8034
rect 45276 7980 45332 7982
rect 47180 14812 47236 14868
rect 46956 12348 47012 12404
rect 46620 12178 46676 12180
rect 46620 12126 46622 12178
rect 46622 12126 46674 12178
rect 46674 12126 46676 12178
rect 46620 12124 46676 12126
rect 46732 10610 46788 10612
rect 46732 10558 46734 10610
rect 46734 10558 46786 10610
rect 46786 10558 46788 10610
rect 46732 10556 46788 10558
rect 46732 10332 46788 10388
rect 45948 9714 46004 9716
rect 45948 9662 45950 9714
rect 45950 9662 46002 9714
rect 46002 9662 46004 9714
rect 45948 9660 46004 9662
rect 45836 9436 45892 9492
rect 46396 9324 46452 9380
rect 46732 9996 46788 10052
rect 45612 9212 45668 9268
rect 46284 9100 46340 9156
rect 45612 8428 45668 8484
rect 45724 8258 45780 8260
rect 45724 8206 45726 8258
rect 45726 8206 45778 8258
rect 45778 8206 45780 8258
rect 45724 8204 45780 8206
rect 44940 6972 44996 7028
rect 44380 6578 44436 6580
rect 44380 6526 44382 6578
rect 44382 6526 44434 6578
rect 44434 6526 44436 6578
rect 44380 6524 44436 6526
rect 44268 6412 44324 6468
rect 44604 6412 44660 6468
rect 43932 4732 43988 4788
rect 44044 6300 44100 6356
rect 43708 4226 43764 4228
rect 43708 4174 43710 4226
rect 43710 4174 43762 4226
rect 43762 4174 43764 4226
rect 43708 4172 43764 4174
rect 44604 4396 44660 4452
rect 45052 6748 45108 6804
rect 45388 6524 45444 6580
rect 45388 6188 45444 6244
rect 45276 5852 45332 5908
rect 45388 5516 45444 5572
rect 45836 7084 45892 7140
rect 46284 6972 46340 7028
rect 45948 6690 46004 6692
rect 45948 6638 45950 6690
rect 45950 6638 46002 6690
rect 46002 6638 46004 6690
rect 45948 6636 46004 6638
rect 46396 6636 46452 6692
rect 46508 9100 46564 9156
rect 46732 7644 46788 7700
rect 45612 5346 45668 5348
rect 45612 5294 45614 5346
rect 45614 5294 45666 5346
rect 45666 5294 45668 5346
rect 45612 5292 45668 5294
rect 46508 4508 46564 4564
rect 47180 12460 47236 12516
rect 47292 12684 47348 12740
rect 47516 12460 47572 12516
rect 48636 16098 48692 16100
rect 48636 16046 48638 16098
rect 48638 16046 48690 16098
rect 48690 16046 48692 16098
rect 48636 16044 48692 16046
rect 48188 15820 48244 15876
rect 48300 15484 48356 15540
rect 48860 16716 48916 16772
rect 49532 16828 49588 16884
rect 49868 16492 49924 16548
rect 49644 16268 49700 16324
rect 49196 15820 49252 15876
rect 48972 15708 49028 15764
rect 48860 15538 48916 15540
rect 48860 15486 48862 15538
rect 48862 15486 48914 15538
rect 48914 15486 48916 15538
rect 48860 15484 48916 15486
rect 49756 16044 49812 16100
rect 49420 15538 49476 15540
rect 49420 15486 49422 15538
rect 49422 15486 49474 15538
rect 49474 15486 49476 15538
rect 49420 15484 49476 15486
rect 51548 22092 51604 22148
rect 51660 21980 51716 22036
rect 51884 22988 51940 23044
rect 51100 21698 51156 21700
rect 51100 21646 51102 21698
rect 51102 21646 51154 21698
rect 51154 21646 51156 21698
rect 51100 21644 51156 21646
rect 51212 21586 51268 21588
rect 51212 21534 51214 21586
rect 51214 21534 51266 21586
rect 51266 21534 51268 21586
rect 51212 21532 51268 21534
rect 51324 21420 51380 21476
rect 51324 20802 51380 20804
rect 51324 20750 51326 20802
rect 51326 20750 51378 20802
rect 51378 20750 51380 20802
rect 51324 20748 51380 20750
rect 50764 20578 50820 20580
rect 50764 20526 50766 20578
rect 50766 20526 50818 20578
rect 50818 20526 50820 20578
rect 50764 20524 50820 20526
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50204 20076 50260 20132
rect 50876 19964 50932 20020
rect 51772 21532 51828 21588
rect 51660 20860 51716 20916
rect 51772 21196 51828 21252
rect 51660 20690 51716 20692
rect 51660 20638 51662 20690
rect 51662 20638 51714 20690
rect 51714 20638 51716 20690
rect 51660 20636 51716 20638
rect 50204 19628 50260 19684
rect 52332 23660 52388 23716
rect 52220 23436 52276 23492
rect 53340 27020 53396 27076
rect 53676 26796 53732 26852
rect 53116 26402 53172 26404
rect 53116 26350 53118 26402
rect 53118 26350 53170 26402
rect 53170 26350 53172 26402
rect 53116 26348 53172 26350
rect 52892 26012 52948 26068
rect 52780 25564 52836 25620
rect 53004 25506 53060 25508
rect 53004 25454 53006 25506
rect 53006 25454 53058 25506
rect 53058 25454 53060 25506
rect 53004 25452 53060 25454
rect 52780 24108 52836 24164
rect 52892 23548 52948 23604
rect 52668 23324 52724 23380
rect 52780 23436 52836 23492
rect 52556 23100 52612 23156
rect 52108 22988 52164 23044
rect 52332 23042 52388 23044
rect 52332 22990 52334 23042
rect 52334 22990 52386 23042
rect 52386 22990 52388 23042
rect 52332 22988 52388 22990
rect 52220 22540 52276 22596
rect 52332 22092 52388 22148
rect 52444 22876 52500 22932
rect 52108 21980 52164 22036
rect 51996 21756 52052 21812
rect 51436 19740 51492 19796
rect 51324 19292 51380 19348
rect 50092 18396 50148 18452
rect 50316 18956 50372 19012
rect 51436 18956 51492 19012
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50092 17388 50148 17444
rect 50204 17052 50260 17108
rect 50988 18396 51044 18452
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 51212 17948 51268 18004
rect 50988 17554 51044 17556
rect 50988 17502 50990 17554
rect 50990 17502 51042 17554
rect 51042 17502 51044 17554
rect 50988 17500 51044 17502
rect 51100 17276 51156 17332
rect 50316 16940 50372 16996
rect 50876 16940 50932 16996
rect 49980 15484 50036 15540
rect 50204 16828 50260 16884
rect 51324 17164 51380 17220
rect 51100 16828 51156 16884
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 49196 14700 49252 14756
rect 48188 13634 48244 13636
rect 48188 13582 48190 13634
rect 48190 13582 48242 13634
rect 48242 13582 48244 13634
rect 48188 13580 48244 13582
rect 48076 13522 48132 13524
rect 48076 13470 48078 13522
rect 48078 13470 48130 13522
rect 48130 13470 48132 13522
rect 48076 13468 48132 13470
rect 48076 13132 48132 13188
rect 48524 12738 48580 12740
rect 48524 12686 48526 12738
rect 48526 12686 48578 12738
rect 48578 12686 48580 12738
rect 48524 12684 48580 12686
rect 47964 12402 48020 12404
rect 47964 12350 47966 12402
rect 47966 12350 48018 12402
rect 48018 12350 48020 12402
rect 47964 12348 48020 12350
rect 47852 11676 47908 11732
rect 47292 9436 47348 9492
rect 47068 8316 47124 8372
rect 46956 7980 47012 8036
rect 47180 7196 47236 7252
rect 47292 7084 47348 7140
rect 47180 4620 47236 4676
rect 47292 6636 47348 6692
rect 47628 11340 47684 11396
rect 47740 10220 47796 10276
rect 47516 9660 47572 9716
rect 47628 9996 47684 10052
rect 47964 10108 48020 10164
rect 47404 4956 47460 5012
rect 47628 7308 47684 7364
rect 47852 6748 47908 6804
rect 47740 5292 47796 5348
rect 48524 11394 48580 11396
rect 48524 11342 48526 11394
rect 48526 11342 48578 11394
rect 48578 11342 48580 11394
rect 48524 11340 48580 11342
rect 48188 11282 48244 11284
rect 48188 11230 48190 11282
rect 48190 11230 48242 11282
rect 48242 11230 48244 11282
rect 48188 11228 48244 11230
rect 48748 12290 48804 12292
rect 48748 12238 48750 12290
rect 48750 12238 48802 12290
rect 48802 12238 48804 12290
rect 48748 12236 48804 12238
rect 48860 12124 48916 12180
rect 48860 11228 48916 11284
rect 48300 9266 48356 9268
rect 48300 9214 48302 9266
rect 48302 9214 48354 9266
rect 48354 9214 48356 9266
rect 48300 9212 48356 9214
rect 48188 9100 48244 9156
rect 48524 10108 48580 10164
rect 49084 12178 49140 12180
rect 49084 12126 49086 12178
rect 49086 12126 49138 12178
rect 49138 12126 49140 12178
rect 49084 12124 49140 12126
rect 49084 11676 49140 11732
rect 49420 13132 49476 13188
rect 50764 15484 50820 15540
rect 49644 12908 49700 12964
rect 49308 12850 49364 12852
rect 49308 12798 49310 12850
rect 49310 12798 49362 12850
rect 49362 12798 49364 12850
rect 49308 12796 49364 12798
rect 49308 12236 49364 12292
rect 49756 13020 49812 13076
rect 49532 12738 49588 12740
rect 49532 12686 49534 12738
rect 49534 12686 49586 12738
rect 49586 12686 49588 12738
rect 49532 12684 49588 12686
rect 49308 11900 49364 11956
rect 49196 10780 49252 10836
rect 49196 10610 49252 10612
rect 49196 10558 49198 10610
rect 49198 10558 49250 10610
rect 49250 10558 49252 10610
rect 49196 10556 49252 10558
rect 48636 10220 48692 10276
rect 48972 9884 49028 9940
rect 49196 9826 49252 9828
rect 49196 9774 49198 9826
rect 49198 9774 49250 9826
rect 49250 9774 49252 9826
rect 49196 9772 49252 9774
rect 49756 12290 49812 12292
rect 49756 12238 49758 12290
rect 49758 12238 49810 12290
rect 49810 12238 49812 12290
rect 49756 12236 49812 12238
rect 49868 12124 49924 12180
rect 50316 14364 50372 14420
rect 50204 13970 50260 13972
rect 50204 13918 50206 13970
rect 50206 13918 50258 13970
rect 50258 13918 50260 13970
rect 50204 13916 50260 13918
rect 50876 15372 50932 15428
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50316 13020 50372 13076
rect 52108 20914 52164 20916
rect 52108 20862 52110 20914
rect 52110 20862 52162 20914
rect 52162 20862 52164 20914
rect 52108 20860 52164 20862
rect 52108 20636 52164 20692
rect 51884 19964 51940 20020
rect 51772 19740 51828 19796
rect 51996 19852 52052 19908
rect 52332 21196 52388 21252
rect 52220 19964 52276 20020
rect 52220 19292 52276 19348
rect 52892 23154 52948 23156
rect 52892 23102 52894 23154
rect 52894 23102 52946 23154
rect 52946 23102 52948 23154
rect 52892 23100 52948 23102
rect 52668 22370 52724 22372
rect 52668 22318 52670 22370
rect 52670 22318 52722 22370
rect 52722 22318 52724 22370
rect 52668 22316 52724 22318
rect 52892 21810 52948 21812
rect 52892 21758 52894 21810
rect 52894 21758 52946 21810
rect 52946 21758 52948 21810
rect 52892 21756 52948 21758
rect 53116 22988 53172 23044
rect 53340 25506 53396 25508
rect 53340 25454 53342 25506
rect 53342 25454 53394 25506
rect 53394 25454 53396 25506
rect 53340 25452 53396 25454
rect 53564 24444 53620 24500
rect 53900 28700 53956 28756
rect 54348 28588 54404 28644
rect 53900 26572 53956 26628
rect 53900 26348 53956 26404
rect 54348 27858 54404 27860
rect 54348 27806 54350 27858
rect 54350 27806 54402 27858
rect 54402 27806 54404 27858
rect 54348 27804 54404 27806
rect 55020 29538 55076 29540
rect 55020 29486 55022 29538
rect 55022 29486 55074 29538
rect 55074 29486 55076 29538
rect 55020 29484 55076 29486
rect 55244 29260 55300 29316
rect 55468 29932 55524 29988
rect 54908 28924 54964 28980
rect 55132 28924 55188 28980
rect 55356 28476 55412 28532
rect 55132 27804 55188 27860
rect 55020 27074 55076 27076
rect 55020 27022 55022 27074
rect 55022 27022 55074 27074
rect 55074 27022 55076 27074
rect 55020 27020 55076 27022
rect 54124 26796 54180 26852
rect 54572 26572 54628 26628
rect 54460 26348 54516 26404
rect 54012 25564 54068 25620
rect 53900 24220 53956 24276
rect 53900 23996 53956 24052
rect 54460 25394 54516 25396
rect 54460 25342 54462 25394
rect 54462 25342 54514 25394
rect 54514 25342 54516 25394
rect 54460 25340 54516 25342
rect 54236 25282 54292 25284
rect 54236 25230 54238 25282
rect 54238 25230 54290 25282
rect 54290 25230 54292 25282
rect 54236 25228 54292 25230
rect 54124 24220 54180 24276
rect 53340 23154 53396 23156
rect 53340 23102 53342 23154
rect 53342 23102 53394 23154
rect 53394 23102 53396 23154
rect 53340 23100 53396 23102
rect 53676 23436 53732 23492
rect 53564 22876 53620 22932
rect 53900 23212 53956 23268
rect 53788 22652 53844 22708
rect 54012 23154 54068 23156
rect 54012 23102 54014 23154
rect 54014 23102 54066 23154
rect 54066 23102 54068 23154
rect 54012 23100 54068 23102
rect 52668 21644 52724 21700
rect 52556 21532 52612 21588
rect 52556 20860 52612 20916
rect 53676 21756 53732 21812
rect 53340 20748 53396 20804
rect 53676 21084 53732 21140
rect 52892 20578 52948 20580
rect 52892 20526 52894 20578
rect 52894 20526 52946 20578
rect 52946 20526 52948 20578
rect 52892 20524 52948 20526
rect 52780 20412 52836 20468
rect 53004 20130 53060 20132
rect 53004 20078 53006 20130
rect 53006 20078 53058 20130
rect 53058 20078 53060 20130
rect 53004 20076 53060 20078
rect 53340 20188 53396 20244
rect 52892 19628 52948 19684
rect 52444 19516 52500 19572
rect 51996 19234 52052 19236
rect 51996 19182 51998 19234
rect 51998 19182 52050 19234
rect 52050 19182 52052 19234
rect 51996 19180 52052 19182
rect 51772 18338 51828 18340
rect 51772 18286 51774 18338
rect 51774 18286 51826 18338
rect 51826 18286 51828 18338
rect 51772 18284 51828 18286
rect 51660 18172 51716 18228
rect 52668 18450 52724 18452
rect 52668 18398 52670 18450
rect 52670 18398 52722 18450
rect 52722 18398 52724 18450
rect 52668 18396 52724 18398
rect 53116 19628 53172 19684
rect 53340 19404 53396 19460
rect 54348 22876 54404 22932
rect 53564 20188 53620 20244
rect 53564 19628 53620 19684
rect 53564 19122 53620 19124
rect 53564 19070 53566 19122
rect 53566 19070 53618 19122
rect 53618 19070 53620 19122
rect 53564 19068 53620 19070
rect 53116 18956 53172 19012
rect 53004 18284 53060 18340
rect 52892 18226 52948 18228
rect 52892 18174 52894 18226
rect 52894 18174 52946 18226
rect 52946 18174 52948 18226
rect 52892 18172 52948 18174
rect 52780 18060 52836 18116
rect 53340 18060 53396 18116
rect 51660 17500 51716 17556
rect 52444 17500 52500 17556
rect 51884 17164 51940 17220
rect 52332 17276 52388 17332
rect 51772 15372 51828 15428
rect 51100 13468 51156 13524
rect 50988 13356 51044 13412
rect 50876 12796 50932 12852
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50764 12236 50820 12292
rect 50204 12124 50260 12180
rect 49532 11282 49588 11284
rect 49532 11230 49534 11282
rect 49534 11230 49586 11282
rect 49586 11230 49588 11282
rect 49532 11228 49588 11230
rect 49644 11452 49700 11508
rect 49420 9324 49476 9380
rect 49532 11004 49588 11060
rect 48412 8428 48468 8484
rect 48300 7980 48356 8036
rect 48188 7532 48244 7588
rect 48188 7362 48244 7364
rect 48188 7310 48190 7362
rect 48190 7310 48242 7362
rect 48242 7310 48244 7362
rect 48188 7308 48244 7310
rect 48300 6076 48356 6132
rect 48076 5010 48132 5012
rect 48076 4958 48078 5010
rect 48078 4958 48130 5010
rect 48130 4958 48132 5010
rect 48076 4956 48132 4958
rect 47964 4732 48020 4788
rect 47628 4284 47684 4340
rect 48860 8370 48916 8372
rect 48860 8318 48862 8370
rect 48862 8318 48914 8370
rect 48914 8318 48916 8370
rect 48860 8316 48916 8318
rect 48636 6802 48692 6804
rect 48636 6750 48638 6802
rect 48638 6750 48690 6802
rect 48690 6750 48692 6802
rect 48636 6748 48692 6750
rect 48860 6860 48916 6916
rect 50092 11676 50148 11732
rect 51100 12178 51156 12180
rect 51100 12126 51102 12178
rect 51102 12126 51154 12178
rect 51154 12126 51156 12178
rect 51100 12124 51156 12126
rect 50316 11004 50372 11060
rect 49756 9826 49812 9828
rect 49756 9774 49758 9826
rect 49758 9774 49810 9826
rect 49810 9774 49812 9826
rect 49756 9772 49812 9774
rect 49756 9548 49812 9604
rect 49756 8876 49812 8932
rect 50204 10610 50260 10612
rect 50204 10558 50206 10610
rect 50206 10558 50258 10610
rect 50258 10558 50260 10610
rect 50204 10556 50260 10558
rect 50204 10332 50260 10388
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50316 10108 50372 10164
rect 50092 9212 50148 9268
rect 49420 8258 49476 8260
rect 49420 8206 49422 8258
rect 49422 8206 49474 8258
rect 49474 8206 49476 8258
rect 49420 8204 49476 8206
rect 49532 8092 49588 8148
rect 49308 7420 49364 7476
rect 49196 6690 49252 6692
rect 49196 6638 49198 6690
rect 49198 6638 49250 6690
rect 49250 6638 49252 6690
rect 49196 6636 49252 6638
rect 48748 6300 48804 6356
rect 48860 6524 48916 6580
rect 49756 8316 49812 8372
rect 49756 7980 49812 8036
rect 49644 6524 49700 6580
rect 49756 7420 49812 7476
rect 50316 9548 50372 9604
rect 48860 5906 48916 5908
rect 48860 5854 48862 5906
rect 48862 5854 48914 5906
rect 48914 5854 48916 5906
rect 48860 5852 48916 5854
rect 48748 5234 48804 5236
rect 48748 5182 48750 5234
rect 48750 5182 48802 5234
rect 48802 5182 48804 5234
rect 48748 5180 48804 5182
rect 48748 4338 48804 4340
rect 48748 4286 48750 4338
rect 48750 4286 48802 4338
rect 48802 4286 48804 4338
rect 48748 4284 48804 4286
rect 48076 2940 48132 2996
rect 49644 5740 49700 5796
rect 49196 5628 49252 5684
rect 49308 4450 49364 4452
rect 49308 4398 49310 4450
rect 49310 4398 49362 4450
rect 49362 4398 49364 4450
rect 49308 4396 49364 4398
rect 49868 7362 49924 7364
rect 49868 7310 49870 7362
rect 49870 7310 49922 7362
rect 49922 7310 49924 7362
rect 49868 7308 49924 7310
rect 50092 6860 50148 6916
rect 49980 6578 50036 6580
rect 49980 6526 49982 6578
rect 49982 6526 50034 6578
rect 50034 6526 50036 6578
rect 49980 6524 50036 6526
rect 50540 9826 50596 9828
rect 50540 9774 50542 9826
rect 50542 9774 50594 9826
rect 50594 9774 50596 9826
rect 50540 9772 50596 9774
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50988 9436 51044 9492
rect 50764 9380 50820 9382
rect 51212 9042 51268 9044
rect 51212 8990 51214 9042
rect 51214 8990 51266 9042
rect 51266 8990 51268 9042
rect 51212 8988 51268 8990
rect 50540 8204 50596 8260
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50652 7698 50708 7700
rect 50652 7646 50654 7698
rect 50654 7646 50706 7698
rect 50706 7646 50708 7698
rect 50652 7644 50708 7646
rect 50540 6412 50596 6468
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 51100 8764 51156 8820
rect 50988 6748 51044 6804
rect 51324 8652 51380 8708
rect 50876 4956 50932 5012
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 49420 2716 49476 2772
rect 48860 1484 48916 1540
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 51660 15036 51716 15092
rect 52220 15036 52276 15092
rect 52108 13804 52164 13860
rect 51772 11452 51828 11508
rect 51660 11340 51716 11396
rect 51548 10892 51604 10948
rect 52220 12348 52276 12404
rect 52108 11564 52164 11620
rect 51996 10780 52052 10836
rect 51660 9714 51716 9716
rect 51660 9662 51662 9714
rect 51662 9662 51714 9714
rect 51714 9662 51716 9714
rect 51660 9660 51716 9662
rect 51548 8652 51604 8708
rect 51548 8316 51604 8372
rect 51548 6860 51604 6916
rect 51660 6300 51716 6356
rect 51548 5740 51604 5796
rect 51884 10498 51940 10500
rect 51884 10446 51886 10498
rect 51886 10446 51938 10498
rect 51938 10446 51940 10498
rect 51884 10444 51940 10446
rect 51884 9772 51940 9828
rect 51996 9436 52052 9492
rect 52332 9548 52388 9604
rect 51884 8652 51940 8708
rect 52332 8428 52388 8484
rect 52892 17612 52948 17668
rect 52556 17052 52612 17108
rect 52780 16044 52836 16100
rect 52892 16492 52948 16548
rect 54348 20802 54404 20804
rect 54348 20750 54350 20802
rect 54350 20750 54402 20802
rect 54402 20750 54404 20802
rect 54348 20748 54404 20750
rect 54124 20188 54180 20244
rect 53900 19906 53956 19908
rect 53900 19854 53902 19906
rect 53902 19854 53954 19906
rect 53954 19854 53956 19906
rect 53900 19852 53956 19854
rect 54012 19122 54068 19124
rect 54012 19070 54014 19122
rect 54014 19070 54066 19122
rect 54066 19070 54068 19122
rect 54012 19068 54068 19070
rect 53900 16940 53956 16996
rect 54012 17724 54068 17780
rect 53676 16492 53732 16548
rect 52668 15874 52724 15876
rect 52668 15822 52670 15874
rect 52670 15822 52722 15874
rect 52722 15822 52724 15874
rect 52668 15820 52724 15822
rect 52668 15372 52724 15428
rect 52892 15148 52948 15204
rect 52780 14588 52836 14644
rect 52668 13746 52724 13748
rect 52668 13694 52670 13746
rect 52670 13694 52722 13746
rect 52722 13694 52724 13746
rect 52668 13692 52724 13694
rect 53116 15036 53172 15092
rect 54124 15874 54180 15876
rect 54124 15822 54126 15874
rect 54126 15822 54178 15874
rect 54178 15822 54180 15874
rect 54124 15820 54180 15822
rect 54124 15538 54180 15540
rect 54124 15486 54126 15538
rect 54126 15486 54178 15538
rect 54178 15486 54180 15538
rect 54124 15484 54180 15486
rect 54236 15202 54292 15204
rect 54236 15150 54238 15202
rect 54238 15150 54290 15202
rect 54290 15150 54292 15202
rect 54236 15148 54292 15150
rect 54684 23996 54740 24052
rect 54684 23266 54740 23268
rect 54684 23214 54686 23266
rect 54686 23214 54738 23266
rect 54738 23214 54740 23266
rect 54684 23212 54740 23214
rect 55132 23548 55188 23604
rect 55020 23154 55076 23156
rect 55020 23102 55022 23154
rect 55022 23102 55074 23154
rect 55074 23102 55076 23154
rect 55020 23100 55076 23102
rect 55020 22540 55076 22596
rect 55356 24722 55412 24724
rect 55356 24670 55358 24722
rect 55358 24670 55410 24722
rect 55410 24670 55412 24722
rect 55356 24668 55412 24670
rect 55244 23212 55300 23268
rect 55356 23660 55412 23716
rect 55804 29036 55860 29092
rect 55916 30156 55972 30212
rect 55692 28700 55748 28756
rect 55580 27970 55636 27972
rect 55580 27918 55582 27970
rect 55582 27918 55634 27970
rect 55634 27918 55636 27970
rect 55580 27916 55636 27918
rect 55916 28642 55972 28644
rect 55916 28590 55918 28642
rect 55918 28590 55970 28642
rect 55970 28590 55972 28642
rect 55916 28588 55972 28590
rect 55692 26290 55748 26292
rect 55692 26238 55694 26290
rect 55694 26238 55746 26290
rect 55746 26238 55748 26290
rect 55692 26236 55748 26238
rect 55916 26402 55972 26404
rect 55916 26350 55918 26402
rect 55918 26350 55970 26402
rect 55970 26350 55972 26402
rect 55916 26348 55972 26350
rect 60956 31948 61012 32004
rect 56588 29260 56644 29316
rect 56812 29148 56868 29204
rect 56476 28924 56532 28980
rect 56364 28028 56420 28084
rect 56924 28588 56980 28644
rect 57820 28700 57876 28756
rect 57036 28364 57092 28420
rect 57148 27916 57204 27972
rect 56924 26572 56980 26628
rect 56028 25116 56084 25172
rect 56140 26236 56196 26292
rect 55804 24946 55860 24948
rect 55804 24894 55806 24946
rect 55806 24894 55858 24946
rect 55858 24894 55860 24946
rect 55804 24892 55860 24894
rect 55916 24834 55972 24836
rect 55916 24782 55918 24834
rect 55918 24782 55970 24834
rect 55970 24782 55972 24834
rect 55916 24780 55972 24782
rect 57820 28418 57876 28420
rect 57820 28366 57822 28418
rect 57822 28366 57874 28418
rect 57874 28366 57876 28418
rect 57820 28364 57876 28366
rect 58492 28700 58548 28756
rect 59388 28924 59444 28980
rect 58044 28418 58100 28420
rect 58044 28366 58046 28418
rect 58046 28366 58098 28418
rect 58098 28366 58100 28418
rect 58044 28364 58100 28366
rect 59052 28364 59108 28420
rect 58828 27804 58884 27860
rect 57820 27634 57876 27636
rect 57820 27582 57822 27634
rect 57822 27582 57874 27634
rect 57874 27582 57876 27634
rect 57820 27580 57876 27582
rect 57708 27020 57764 27076
rect 57148 26290 57204 26292
rect 57148 26238 57150 26290
rect 57150 26238 57202 26290
rect 57202 26238 57204 26290
rect 57148 26236 57204 26238
rect 56812 25452 56868 25508
rect 55692 23660 55748 23716
rect 55692 23324 55748 23380
rect 55804 23212 55860 23268
rect 57148 25116 57204 25172
rect 57036 24834 57092 24836
rect 57036 24782 57038 24834
rect 57038 24782 57090 24834
rect 57090 24782 57092 24834
rect 57036 24780 57092 24782
rect 56924 24668 56980 24724
rect 56476 23548 56532 23604
rect 55804 22652 55860 22708
rect 55468 22428 55524 22484
rect 54908 21308 54964 21364
rect 54796 20802 54852 20804
rect 54796 20750 54798 20802
rect 54798 20750 54850 20802
rect 54850 20750 54852 20802
rect 54796 20748 54852 20750
rect 54684 20636 54740 20692
rect 55132 21084 55188 21140
rect 55132 19404 55188 19460
rect 54684 17836 54740 17892
rect 55356 19122 55412 19124
rect 55356 19070 55358 19122
rect 55358 19070 55410 19122
rect 55410 19070 55412 19122
rect 55356 19068 55412 19070
rect 55244 17724 55300 17780
rect 55804 21868 55860 21924
rect 56028 21084 56084 21140
rect 55916 20636 55972 20692
rect 55692 19122 55748 19124
rect 55692 19070 55694 19122
rect 55694 19070 55746 19122
rect 55746 19070 55748 19122
rect 55692 19068 55748 19070
rect 56028 18956 56084 19012
rect 55916 18396 55972 18452
rect 56924 23154 56980 23156
rect 56924 23102 56926 23154
rect 56926 23102 56978 23154
rect 56978 23102 56980 23154
rect 56924 23100 56980 23102
rect 55580 17612 55636 17668
rect 57148 23884 57204 23940
rect 57036 22652 57092 22708
rect 57036 22482 57092 22484
rect 57036 22430 57038 22482
rect 57038 22430 57090 22482
rect 57090 22430 57092 22482
rect 57036 22428 57092 22430
rect 57148 22092 57204 22148
rect 56588 21868 56644 21924
rect 58044 27020 58100 27076
rect 58156 26572 58212 26628
rect 58716 26348 58772 26404
rect 58044 26236 58100 26292
rect 59388 28700 59444 28756
rect 59052 27132 59108 27188
rect 57708 24722 57764 24724
rect 57708 24670 57710 24722
rect 57710 24670 57762 24722
rect 57762 24670 57764 24722
rect 57708 24668 57764 24670
rect 57708 23996 57764 24052
rect 57372 21756 57428 21812
rect 57820 23266 57876 23268
rect 57820 23214 57822 23266
rect 57822 23214 57874 23266
rect 57874 23214 57876 23266
rect 57820 23212 57876 23214
rect 58156 25340 58212 25396
rect 58492 24892 58548 24948
rect 58268 24834 58324 24836
rect 58268 24782 58270 24834
rect 58270 24782 58322 24834
rect 58322 24782 58324 24834
rect 58268 24780 58324 24782
rect 58828 24668 58884 24724
rect 58604 24050 58660 24052
rect 58604 23998 58606 24050
rect 58606 23998 58658 24050
rect 58658 23998 58660 24050
rect 58604 23996 58660 23998
rect 58380 23772 58436 23828
rect 57932 23100 57988 23156
rect 58268 23324 58324 23380
rect 58380 22204 58436 22260
rect 57372 21196 57428 21252
rect 57484 20860 57540 20916
rect 58268 20914 58324 20916
rect 58268 20862 58270 20914
rect 58270 20862 58322 20914
rect 58322 20862 58324 20914
rect 58268 20860 58324 20862
rect 56588 19180 56644 19236
rect 57484 20524 57540 20580
rect 58604 22146 58660 22148
rect 58604 22094 58606 22146
rect 58606 22094 58658 22146
rect 58658 22094 58660 22146
rect 58604 22092 58660 22094
rect 59388 27356 59444 27412
rect 59836 27858 59892 27860
rect 59836 27806 59838 27858
rect 59838 27806 59890 27858
rect 59890 27806 59892 27858
rect 59836 27804 59892 27806
rect 59500 26908 59556 26964
rect 59612 26012 59668 26068
rect 59500 25506 59556 25508
rect 59500 25454 59502 25506
rect 59502 25454 59554 25506
rect 59554 25454 59556 25506
rect 59500 25452 59556 25454
rect 59164 25116 59220 25172
rect 60620 27858 60676 27860
rect 60620 27806 60622 27858
rect 60622 27806 60674 27858
rect 60674 27806 60676 27858
rect 60620 27804 60676 27806
rect 60508 27356 60564 27412
rect 60844 27468 60900 27524
rect 62076 29820 62132 29876
rect 61068 27858 61124 27860
rect 61068 27806 61070 27858
rect 61070 27806 61122 27858
rect 61122 27806 61124 27858
rect 61068 27804 61124 27806
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 81276 56474 81332 56476
rect 81276 56422 81278 56474
rect 81278 56422 81330 56474
rect 81330 56422 81332 56474
rect 81276 56420 81332 56422
rect 81380 56474 81436 56476
rect 81380 56422 81382 56474
rect 81382 56422 81434 56474
rect 81434 56422 81436 56474
rect 81380 56420 81436 56422
rect 81484 56474 81540 56476
rect 81484 56422 81486 56474
rect 81486 56422 81538 56474
rect 81538 56422 81540 56474
rect 81484 56420 81540 56422
rect 81788 56252 81844 56308
rect 83020 56306 83076 56308
rect 83020 56254 83022 56306
rect 83022 56254 83074 56306
rect 83074 56254 83076 56306
rect 83020 56252 83076 56254
rect 69804 55298 69860 55300
rect 69804 55246 69806 55298
rect 69806 55246 69858 55298
rect 69858 55246 69860 55298
rect 69804 55244 69860 55246
rect 70140 55132 70196 55188
rect 71036 55298 71092 55300
rect 71036 55246 71038 55298
rect 71038 55246 71090 55298
rect 71090 55246 71092 55298
rect 71036 55244 71092 55246
rect 70700 55186 70756 55188
rect 70700 55134 70702 55186
rect 70702 55134 70754 55186
rect 70754 55134 70756 55186
rect 70700 55132 70756 55134
rect 71484 55186 71540 55188
rect 71484 55134 71486 55186
rect 71486 55134 71538 55186
rect 71538 55134 71540 55186
rect 71484 55132 71540 55134
rect 74620 30940 74676 30996
rect 74060 30828 74116 30884
rect 68012 30492 68068 30548
rect 69468 30716 69524 30772
rect 62972 29820 63028 29876
rect 60508 26684 60564 26740
rect 61180 27244 61236 27300
rect 59500 24892 59556 24948
rect 59164 23042 59220 23044
rect 59164 22990 59166 23042
rect 59166 22990 59218 23042
rect 59218 22990 59220 23042
rect 59164 22988 59220 22990
rect 60508 25452 60564 25508
rect 60284 24892 60340 24948
rect 59948 23212 60004 23268
rect 60060 23772 60116 23828
rect 58940 22764 58996 22820
rect 59836 23154 59892 23156
rect 59836 23102 59838 23154
rect 59838 23102 59890 23154
rect 59890 23102 59892 23154
rect 59836 23100 59892 23102
rect 58828 21756 58884 21812
rect 59052 22652 59108 22708
rect 59052 21868 59108 21924
rect 59836 22428 59892 22484
rect 61628 27186 61684 27188
rect 61628 27134 61630 27186
rect 61630 27134 61682 27186
rect 61682 27134 61684 27186
rect 61628 27132 61684 27134
rect 61852 26962 61908 26964
rect 61852 26910 61854 26962
rect 61854 26910 61906 26962
rect 61906 26910 61908 26962
rect 61852 26908 61908 26910
rect 61292 26796 61348 26852
rect 63196 28028 63252 28084
rect 62748 27468 62804 27524
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 68236 28812 68292 28868
rect 63644 28028 63700 28084
rect 63756 27970 63812 27972
rect 63756 27918 63758 27970
rect 63758 27918 63810 27970
rect 63810 27918 63812 27970
rect 63756 27916 63812 27918
rect 64764 28082 64820 28084
rect 64764 28030 64766 28082
rect 64766 28030 64818 28082
rect 64818 28030 64820 28082
rect 64764 28028 64820 28030
rect 65660 28028 65716 28084
rect 65324 27970 65380 27972
rect 65324 27918 65326 27970
rect 65326 27918 65378 27970
rect 65378 27918 65380 27970
rect 65324 27916 65380 27918
rect 65100 27858 65156 27860
rect 65100 27806 65102 27858
rect 65102 27806 65154 27858
rect 65154 27806 65156 27858
rect 65100 27804 65156 27806
rect 66108 28140 66164 28196
rect 67676 28364 67732 28420
rect 65996 27916 66052 27972
rect 65884 27858 65940 27860
rect 65884 27806 65886 27858
rect 65886 27806 65938 27858
rect 65938 27806 65940 27858
rect 65884 27804 65940 27806
rect 66220 27858 66276 27860
rect 66220 27806 66222 27858
rect 66222 27806 66274 27858
rect 66274 27806 66276 27858
rect 66220 27804 66276 27806
rect 63308 27580 63364 27636
rect 63644 27186 63700 27188
rect 63644 27134 63646 27186
rect 63646 27134 63698 27186
rect 63698 27134 63700 27186
rect 63644 27132 63700 27134
rect 63196 27020 63252 27076
rect 63980 27074 64036 27076
rect 63980 27022 63982 27074
rect 63982 27022 64034 27074
rect 64034 27022 64036 27074
rect 63980 27020 64036 27022
rect 64764 27020 64820 27076
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 66444 27186 66500 27188
rect 66444 27134 66446 27186
rect 66446 27134 66498 27186
rect 66498 27134 66500 27186
rect 66444 27132 66500 27134
rect 61964 26796 62020 26852
rect 61180 26236 61236 26292
rect 62636 26684 62692 26740
rect 61964 26236 62020 26292
rect 60956 26012 61012 26068
rect 60732 25282 60788 25284
rect 60732 25230 60734 25282
rect 60734 25230 60786 25282
rect 60786 25230 60788 25282
rect 60732 25228 60788 25230
rect 60284 23154 60340 23156
rect 60284 23102 60286 23154
rect 60286 23102 60338 23154
rect 60338 23102 60340 23154
rect 60284 23100 60340 23102
rect 61516 26012 61572 26068
rect 61180 25900 61236 25956
rect 62188 25788 62244 25844
rect 60956 24108 61012 24164
rect 60396 22988 60452 23044
rect 59388 22146 59444 22148
rect 59388 22094 59390 22146
rect 59390 22094 59442 22146
rect 59442 22094 59444 22146
rect 59388 22092 59444 22094
rect 58828 20578 58884 20580
rect 58828 20526 58830 20578
rect 58830 20526 58882 20578
rect 58882 20526 58884 20578
rect 58828 20524 58884 20526
rect 58268 19516 58324 19572
rect 57484 19292 57540 19348
rect 58268 19122 58324 19124
rect 58268 19070 58270 19122
rect 58270 19070 58322 19122
rect 58322 19070 58324 19122
rect 58268 19068 58324 19070
rect 58156 18844 58212 18900
rect 56812 18284 56868 18340
rect 56252 17948 56308 18004
rect 55020 16940 55076 16996
rect 55692 16828 55748 16884
rect 55916 16380 55972 16436
rect 56588 18226 56644 18228
rect 56588 18174 56590 18226
rect 56590 18174 56642 18226
rect 56642 18174 56644 18226
rect 56588 18172 56644 18174
rect 56140 17778 56196 17780
rect 56140 17726 56142 17778
rect 56142 17726 56194 17778
rect 56194 17726 56196 17778
rect 56140 17724 56196 17726
rect 56700 17612 56756 17668
rect 56812 17500 56868 17556
rect 57820 18338 57876 18340
rect 57820 18286 57822 18338
rect 57822 18286 57874 18338
rect 57874 18286 57876 18338
rect 57820 18284 57876 18286
rect 57372 18172 57428 18228
rect 57260 18060 57316 18116
rect 57260 17164 57316 17220
rect 57596 17276 57652 17332
rect 56700 17106 56756 17108
rect 56700 17054 56702 17106
rect 56702 17054 56754 17106
rect 56754 17054 56756 17106
rect 56700 17052 56756 17054
rect 56588 16828 56644 16884
rect 57036 16882 57092 16884
rect 57036 16830 57038 16882
rect 57038 16830 57090 16882
rect 57090 16830 57092 16882
rect 57036 16828 57092 16830
rect 56028 16268 56084 16324
rect 56588 16380 56644 16436
rect 57484 16098 57540 16100
rect 57484 16046 57486 16098
rect 57486 16046 57538 16098
rect 57538 16046 57540 16098
rect 57484 16044 57540 16046
rect 56252 15708 56308 15764
rect 55132 15538 55188 15540
rect 55132 15486 55134 15538
rect 55134 15486 55186 15538
rect 55186 15486 55188 15538
rect 55132 15484 55188 15486
rect 54012 14812 54068 14868
rect 53116 13804 53172 13860
rect 52780 12572 52836 12628
rect 53004 12962 53060 12964
rect 53004 12910 53006 12962
rect 53006 12910 53058 12962
rect 53058 12910 53060 12962
rect 53004 12908 53060 12910
rect 54572 14306 54628 14308
rect 54572 14254 54574 14306
rect 54574 14254 54626 14306
rect 54626 14254 54628 14306
rect 54572 14252 54628 14254
rect 54348 12962 54404 12964
rect 54348 12910 54350 12962
rect 54350 12910 54402 12962
rect 54402 12910 54404 12962
rect 54348 12908 54404 12910
rect 52892 12124 52948 12180
rect 52668 11900 52724 11956
rect 52780 11506 52836 11508
rect 52780 11454 52782 11506
rect 52782 11454 52834 11506
rect 52834 11454 52836 11506
rect 52780 11452 52836 11454
rect 53004 11394 53060 11396
rect 53004 11342 53006 11394
rect 53006 11342 53058 11394
rect 53058 11342 53060 11394
rect 53004 11340 53060 11342
rect 53452 12572 53508 12628
rect 53564 12460 53620 12516
rect 53452 12348 53508 12404
rect 52444 9884 52500 9940
rect 53340 10332 53396 10388
rect 52556 9266 52612 9268
rect 52556 9214 52558 9266
rect 52558 9214 52610 9266
rect 52610 9214 52612 9266
rect 52556 9212 52612 9214
rect 52780 9042 52836 9044
rect 52780 8990 52782 9042
rect 52782 8990 52834 9042
rect 52834 8990 52836 9042
rect 52780 8988 52836 8990
rect 52780 8204 52836 8260
rect 51996 7868 52052 7924
rect 52220 7644 52276 7700
rect 51884 7308 51940 7364
rect 52108 6802 52164 6804
rect 52108 6750 52110 6802
rect 52110 6750 52162 6802
rect 52162 6750 52164 6802
rect 52108 6748 52164 6750
rect 52108 6412 52164 6468
rect 51884 6018 51940 6020
rect 51884 5966 51886 6018
rect 51886 5966 51938 6018
rect 51938 5966 51940 6018
rect 51884 5964 51940 5966
rect 51548 4732 51604 4788
rect 51212 4396 51268 4452
rect 51884 4338 51940 4340
rect 51884 4286 51886 4338
rect 51886 4286 51938 4338
rect 51938 4286 51940 4338
rect 51884 4284 51940 4286
rect 51548 3442 51604 3444
rect 51548 3390 51550 3442
rect 51550 3390 51602 3442
rect 51602 3390 51604 3442
rect 51548 3388 51604 3390
rect 51996 2828 52052 2884
rect 52332 7308 52388 7364
rect 52332 7084 52388 7140
rect 52556 7474 52612 7476
rect 52556 7422 52558 7474
rect 52558 7422 52610 7474
rect 52610 7422 52612 7474
rect 52556 7420 52612 7422
rect 52444 6412 52500 6468
rect 52556 6076 52612 6132
rect 52668 6636 52724 6692
rect 53004 8146 53060 8148
rect 53004 8094 53006 8146
rect 53006 8094 53058 8146
rect 53058 8094 53060 8146
rect 53004 8092 53060 8094
rect 53228 8316 53284 8372
rect 53228 8146 53284 8148
rect 53228 8094 53230 8146
rect 53230 8094 53282 8146
rect 53282 8094 53284 8146
rect 53228 8092 53284 8094
rect 53116 7980 53172 8036
rect 52892 6748 52948 6804
rect 53004 7308 53060 7364
rect 52780 5964 52836 6020
rect 53564 11900 53620 11956
rect 53900 11900 53956 11956
rect 53788 11564 53844 11620
rect 54124 11282 54180 11284
rect 54124 11230 54126 11282
rect 54126 11230 54178 11282
rect 54178 11230 54180 11282
rect 54124 11228 54180 11230
rect 54012 10780 54068 10836
rect 54460 12572 54516 12628
rect 54684 12460 54740 12516
rect 54460 10834 54516 10836
rect 54460 10782 54462 10834
rect 54462 10782 54514 10834
rect 54514 10782 54516 10834
rect 54460 10780 54516 10782
rect 53788 10722 53844 10724
rect 53788 10670 53790 10722
rect 53790 10670 53842 10722
rect 53842 10670 53844 10722
rect 53788 10668 53844 10670
rect 53676 10556 53732 10612
rect 53452 7308 53508 7364
rect 53340 6748 53396 6804
rect 54572 10556 54628 10612
rect 58380 18620 58436 18676
rect 58604 18562 58660 18564
rect 58604 18510 58606 18562
rect 58606 18510 58658 18562
rect 58658 18510 58660 18562
rect 58604 18508 58660 18510
rect 58492 18284 58548 18340
rect 59052 20860 59108 20916
rect 59052 20412 59108 20468
rect 59164 19964 59220 20020
rect 59052 19516 59108 19572
rect 59836 22258 59892 22260
rect 59836 22206 59838 22258
rect 59838 22206 59890 22258
rect 59890 22206 59892 22258
rect 59836 22204 59892 22206
rect 60060 21868 60116 21924
rect 59500 21586 59556 21588
rect 59500 21534 59502 21586
rect 59502 21534 59554 21586
rect 59554 21534 59556 21586
rect 59500 21532 59556 21534
rect 59388 20802 59444 20804
rect 59388 20750 59390 20802
rect 59390 20750 59442 20802
rect 59442 20750 59444 20802
rect 59388 20748 59444 20750
rect 60956 23826 61012 23828
rect 60956 23774 60958 23826
rect 60958 23774 61010 23826
rect 61010 23774 61012 23826
rect 60956 23772 61012 23774
rect 61068 22988 61124 23044
rect 61628 25228 61684 25284
rect 64204 26850 64260 26852
rect 64204 26798 64206 26850
rect 64206 26798 64258 26850
rect 64258 26798 64260 26850
rect 64204 26796 64260 26798
rect 64428 26684 64484 26740
rect 63644 26572 63700 26628
rect 63756 26460 63812 26516
rect 63196 26290 63252 26292
rect 63196 26238 63198 26290
rect 63198 26238 63250 26290
rect 63250 26238 63252 26290
rect 63196 26236 63252 26238
rect 65436 26684 65492 26740
rect 67004 26460 67060 26516
rect 67452 26684 67508 26740
rect 67900 26962 67956 26964
rect 67900 26910 67902 26962
rect 67902 26910 67954 26962
rect 67954 26910 67956 26962
rect 67900 26908 67956 26910
rect 67788 26796 67844 26852
rect 67564 26572 67620 26628
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 64988 25452 65044 25508
rect 62860 24946 62916 24948
rect 62860 24894 62862 24946
rect 62862 24894 62914 24946
rect 62914 24894 62916 24946
rect 62860 24892 62916 24894
rect 64316 24892 64372 24948
rect 61404 23324 61460 23380
rect 60956 22092 61012 22148
rect 60844 21810 60900 21812
rect 60844 21758 60846 21810
rect 60846 21758 60898 21810
rect 60898 21758 60900 21810
rect 60844 21756 60900 21758
rect 59948 20914 60004 20916
rect 59948 20862 59950 20914
rect 59950 20862 60002 20914
rect 60002 20862 60004 20914
rect 59948 20860 60004 20862
rect 60508 20914 60564 20916
rect 60508 20862 60510 20914
rect 60510 20862 60562 20914
rect 60562 20862 60564 20914
rect 60508 20860 60564 20862
rect 59724 20748 59780 20804
rect 60620 20802 60676 20804
rect 60620 20750 60622 20802
rect 60622 20750 60674 20802
rect 60674 20750 60676 20802
rect 60620 20748 60676 20750
rect 59388 20524 59444 20580
rect 59724 20412 59780 20468
rect 60956 21532 61012 21588
rect 60956 20802 61012 20804
rect 60956 20750 60958 20802
rect 60958 20750 61010 20802
rect 61010 20750 61012 20802
rect 60956 20748 61012 20750
rect 60732 20188 60788 20244
rect 62524 20188 62580 20244
rect 60060 20076 60116 20132
rect 59836 19740 59892 19796
rect 59276 19404 59332 19460
rect 59388 19516 59444 19572
rect 58716 17106 58772 17108
rect 58716 17054 58718 17106
rect 58718 17054 58770 17106
rect 58770 17054 58772 17106
rect 58716 17052 58772 17054
rect 58940 17554 58996 17556
rect 58940 17502 58942 17554
rect 58942 17502 58994 17554
rect 58994 17502 58996 17554
rect 58940 17500 58996 17502
rect 58828 16828 58884 16884
rect 59164 16828 59220 16884
rect 59276 16044 59332 16100
rect 60956 20130 61012 20132
rect 60956 20078 60958 20130
rect 60958 20078 61010 20130
rect 61010 20078 61012 20130
rect 60956 20076 61012 20078
rect 60172 19964 60228 20020
rect 60172 18956 60228 19012
rect 60732 19068 60788 19124
rect 60620 18732 60676 18788
rect 59724 18508 59780 18564
rect 59500 18450 59556 18452
rect 59500 18398 59502 18450
rect 59502 18398 59554 18450
rect 59554 18398 59556 18450
rect 59500 18396 59556 18398
rect 59724 18226 59780 18228
rect 59724 18174 59726 18226
rect 59726 18174 59778 18226
rect 59778 18174 59780 18226
rect 59724 18172 59780 18174
rect 59500 17554 59556 17556
rect 59500 17502 59502 17554
rect 59502 17502 59554 17554
rect 59554 17502 59556 17554
rect 59500 17500 59556 17502
rect 59948 17276 60004 17332
rect 60396 17276 60452 17332
rect 62412 19180 62468 19236
rect 62300 19122 62356 19124
rect 62300 19070 62302 19122
rect 62302 19070 62354 19122
rect 62354 19070 62356 19122
rect 62300 19068 62356 19070
rect 61180 18508 61236 18564
rect 61292 19010 61348 19012
rect 61292 18958 61294 19010
rect 61294 18958 61346 19010
rect 61346 18958 61348 19010
rect 61292 18956 61348 18958
rect 60732 18284 60788 18340
rect 61068 18396 61124 18452
rect 60620 18172 60676 18228
rect 61068 18060 61124 18116
rect 61964 18284 62020 18340
rect 60732 16882 60788 16884
rect 60732 16830 60734 16882
rect 60734 16830 60786 16882
rect 60786 16830 60788 16882
rect 60732 16828 60788 16830
rect 60956 16882 61012 16884
rect 60956 16830 60958 16882
rect 60958 16830 61010 16882
rect 61010 16830 61012 16882
rect 60956 16828 61012 16830
rect 60620 16156 60676 16212
rect 59388 15484 59444 15540
rect 58156 14924 58212 14980
rect 55132 13746 55188 13748
rect 55132 13694 55134 13746
rect 55134 13694 55186 13746
rect 55186 13694 55188 13746
rect 55132 13692 55188 13694
rect 55244 13580 55300 13636
rect 55132 12236 55188 12292
rect 54908 12178 54964 12180
rect 54908 12126 54910 12178
rect 54910 12126 54962 12178
rect 54962 12126 54964 12178
rect 54908 12124 54964 12126
rect 54796 10444 54852 10500
rect 55916 12908 55972 12964
rect 56028 12402 56084 12404
rect 56028 12350 56030 12402
rect 56030 12350 56082 12402
rect 56082 12350 56084 12402
rect 56028 12348 56084 12350
rect 55916 12124 55972 12180
rect 55580 11228 55636 11284
rect 55468 10834 55524 10836
rect 55468 10782 55470 10834
rect 55470 10782 55522 10834
rect 55522 10782 55524 10834
rect 55468 10780 55524 10782
rect 55916 10892 55972 10948
rect 55132 10220 55188 10276
rect 53900 10108 53956 10164
rect 53340 6412 53396 6468
rect 52668 5906 52724 5908
rect 52668 5854 52670 5906
rect 52670 5854 52722 5906
rect 52722 5854 52724 5906
rect 52668 5852 52724 5854
rect 52780 5404 52836 5460
rect 52780 5010 52836 5012
rect 52780 4958 52782 5010
rect 52782 4958 52834 5010
rect 52834 4958 52836 5010
rect 52780 4956 52836 4958
rect 53004 4844 53060 4900
rect 53340 6018 53396 6020
rect 53340 5966 53342 6018
rect 53342 5966 53394 6018
rect 53394 5966 53396 6018
rect 53340 5964 53396 5966
rect 53340 5292 53396 5348
rect 53676 5122 53732 5124
rect 53676 5070 53678 5122
rect 53678 5070 53730 5122
rect 53730 5070 53732 5122
rect 53676 5068 53732 5070
rect 55020 9996 55076 10052
rect 54348 9154 54404 9156
rect 54348 9102 54350 9154
rect 54350 9102 54402 9154
rect 54402 9102 54404 9154
rect 54348 9100 54404 9102
rect 55692 9772 55748 9828
rect 55804 9884 55860 9940
rect 55244 9660 55300 9716
rect 56812 13746 56868 13748
rect 56812 13694 56814 13746
rect 56814 13694 56866 13746
rect 56866 13694 56868 13746
rect 56812 13692 56868 13694
rect 56700 13634 56756 13636
rect 56700 13582 56702 13634
rect 56702 13582 56754 13634
rect 56754 13582 56756 13634
rect 56700 13580 56756 13582
rect 56812 12796 56868 12852
rect 56588 10780 56644 10836
rect 57036 12684 57092 12740
rect 57036 12348 57092 12404
rect 57148 13580 57204 13636
rect 56924 12178 56980 12180
rect 56924 12126 56926 12178
rect 56926 12126 56978 12178
rect 56978 12126 56980 12178
rect 56924 12124 56980 12126
rect 57036 12012 57092 12068
rect 57596 13692 57652 13748
rect 57708 12850 57764 12852
rect 57708 12798 57710 12850
rect 57710 12798 57762 12850
rect 57762 12798 57764 12850
rect 57708 12796 57764 12798
rect 58044 13634 58100 13636
rect 58044 13582 58046 13634
rect 58046 13582 58098 13634
rect 58098 13582 58100 13634
rect 58044 13580 58100 13582
rect 57260 12348 57316 12404
rect 57484 11340 57540 11396
rect 58044 11900 58100 11956
rect 57148 11004 57204 11060
rect 56924 10668 56980 10724
rect 56140 10610 56196 10612
rect 56140 10558 56142 10610
rect 56142 10558 56194 10610
rect 56194 10558 56196 10610
rect 56140 10556 56196 10558
rect 56700 9996 56756 10052
rect 56028 9714 56084 9716
rect 56028 9662 56030 9714
rect 56030 9662 56082 9714
rect 56082 9662 56084 9714
rect 56028 9660 56084 9662
rect 56140 9602 56196 9604
rect 56140 9550 56142 9602
rect 56142 9550 56194 9602
rect 56194 9550 56196 9602
rect 56140 9548 56196 9550
rect 56812 9548 56868 9604
rect 55356 8876 55412 8932
rect 55244 8428 55300 8484
rect 53900 7532 53956 7588
rect 54012 7474 54068 7476
rect 54012 7422 54014 7474
rect 54014 7422 54066 7474
rect 54066 7422 54068 7474
rect 54012 7420 54068 7422
rect 54684 8092 54740 8148
rect 54460 7980 54516 8036
rect 54684 7308 54740 7364
rect 54124 6524 54180 6580
rect 54348 6636 54404 6692
rect 54236 5852 54292 5908
rect 54684 6300 54740 6356
rect 53116 3388 53172 3444
rect 54908 5122 54964 5124
rect 54908 5070 54910 5122
rect 54910 5070 54962 5122
rect 54962 5070 54964 5122
rect 54908 5068 54964 5070
rect 55020 4956 55076 5012
rect 55916 9154 55972 9156
rect 55916 9102 55918 9154
rect 55918 9102 55970 9154
rect 55970 9102 55972 9154
rect 55916 9100 55972 9102
rect 55692 8540 55748 8596
rect 55580 8428 55636 8484
rect 58380 12460 58436 12516
rect 57260 10610 57316 10612
rect 57260 10558 57262 10610
rect 57262 10558 57314 10610
rect 57314 10558 57316 10610
rect 57260 10556 57316 10558
rect 57708 10332 57764 10388
rect 57932 10498 57988 10500
rect 57932 10446 57934 10498
rect 57934 10446 57986 10498
rect 57986 10446 57988 10498
rect 57932 10444 57988 10446
rect 57932 9996 57988 10052
rect 56140 9042 56196 9044
rect 56140 8990 56142 9042
rect 56142 8990 56194 9042
rect 56194 8990 56196 9042
rect 56140 8988 56196 8990
rect 56588 8764 56644 8820
rect 56812 8540 56868 8596
rect 56028 8428 56084 8484
rect 56700 8428 56756 8484
rect 56028 7644 56084 7700
rect 55692 7474 55748 7476
rect 55692 7422 55694 7474
rect 55694 7422 55746 7474
rect 55746 7422 55748 7474
rect 55692 7420 55748 7422
rect 55468 7084 55524 7140
rect 55580 6300 55636 6356
rect 55692 4284 55748 4340
rect 55804 6524 55860 6580
rect 56476 7644 56532 7700
rect 56140 7308 56196 7364
rect 56028 6412 56084 6468
rect 53788 3164 53844 3220
rect 56924 8428 56980 8484
rect 56588 7586 56644 7588
rect 56588 7534 56590 7586
rect 56590 7534 56642 7586
rect 56642 7534 56644 7586
rect 56588 7532 56644 7534
rect 57148 9100 57204 9156
rect 58268 11228 58324 11284
rect 58716 15036 58772 15092
rect 60508 15708 60564 15764
rect 58604 13468 58660 13524
rect 59276 13356 59332 13412
rect 58716 12124 58772 12180
rect 58716 11506 58772 11508
rect 58716 11454 58718 11506
rect 58718 11454 58770 11506
rect 58770 11454 58772 11506
rect 58716 11452 58772 11454
rect 58828 12684 58884 12740
rect 58828 11004 58884 11060
rect 58156 9826 58212 9828
rect 58156 9774 58158 9826
rect 58158 9774 58210 9826
rect 58210 9774 58212 9826
rect 58156 9772 58212 9774
rect 58268 9602 58324 9604
rect 58268 9550 58270 9602
rect 58270 9550 58322 9602
rect 58322 9550 58324 9602
rect 58268 9548 58324 9550
rect 57036 7868 57092 7924
rect 56812 7084 56868 7140
rect 56476 5516 56532 5572
rect 56700 6972 56756 7028
rect 57036 6972 57092 7028
rect 56812 6018 56868 6020
rect 56812 5966 56814 6018
rect 56814 5966 56866 6018
rect 56866 5966 56868 6018
rect 56812 5964 56868 5966
rect 56588 5180 56644 5236
rect 56588 4844 56644 4900
rect 56700 4450 56756 4452
rect 56700 4398 56702 4450
rect 56702 4398 56754 4450
rect 56754 4398 56756 4450
rect 56700 4396 56756 4398
rect 57036 5404 57092 5460
rect 57036 5234 57092 5236
rect 57036 5182 57038 5234
rect 57038 5182 57090 5234
rect 57090 5182 57092 5234
rect 57036 5180 57092 5182
rect 57260 7698 57316 7700
rect 57260 7646 57262 7698
rect 57262 7646 57314 7698
rect 57314 7646 57316 7698
rect 57260 7644 57316 7646
rect 57484 6524 57540 6580
rect 57596 8428 57652 8484
rect 57708 6802 57764 6804
rect 57708 6750 57710 6802
rect 57710 6750 57762 6802
rect 57762 6750 57764 6802
rect 57708 6748 57764 6750
rect 57708 5794 57764 5796
rect 57708 5742 57710 5794
rect 57710 5742 57762 5794
rect 57762 5742 57764 5794
rect 57708 5740 57764 5742
rect 57260 5292 57316 5348
rect 57148 4956 57204 5012
rect 57596 3612 57652 3668
rect 56140 1260 56196 1316
rect 58380 6748 58436 6804
rect 59500 13074 59556 13076
rect 59500 13022 59502 13074
rect 59502 13022 59554 13074
rect 59554 13022 59556 13074
rect 59500 13020 59556 13022
rect 59276 10834 59332 10836
rect 59276 10782 59278 10834
rect 59278 10782 59330 10834
rect 59330 10782 59332 10834
rect 59276 10780 59332 10782
rect 59052 10444 59108 10500
rect 58716 10108 58772 10164
rect 59276 10386 59332 10388
rect 59276 10334 59278 10386
rect 59278 10334 59330 10386
rect 59330 10334 59332 10386
rect 59276 10332 59332 10334
rect 59388 9884 59444 9940
rect 59948 13244 60004 13300
rect 59836 12908 59892 12964
rect 59836 12012 59892 12068
rect 60060 13132 60116 13188
rect 59836 11564 59892 11620
rect 59948 11116 60004 11172
rect 60060 11452 60116 11508
rect 59052 9548 59108 9604
rect 59164 9154 59220 9156
rect 59164 9102 59166 9154
rect 59166 9102 59218 9154
rect 59218 9102 59220 9154
rect 59164 9100 59220 9102
rect 58716 7644 58772 7700
rect 58492 6412 58548 6468
rect 58940 4956 58996 5012
rect 59052 3666 59108 3668
rect 59052 3614 59054 3666
rect 59054 3614 59106 3666
rect 59106 3614 59108 3666
rect 59052 3612 59108 3614
rect 59948 9826 60004 9828
rect 59948 9774 59950 9826
rect 59950 9774 60002 9826
rect 60002 9774 60004 9826
rect 59948 9772 60004 9774
rect 59724 9548 59780 9604
rect 59500 8146 59556 8148
rect 59500 8094 59502 8146
rect 59502 8094 59554 8146
rect 59554 8094 59556 8146
rect 59500 8092 59556 8094
rect 59836 9436 59892 9492
rect 59836 7644 59892 7700
rect 60620 14700 60676 14756
rect 61964 17164 62020 17220
rect 61068 16268 61124 16324
rect 61404 16828 61460 16884
rect 61404 15708 61460 15764
rect 60732 14476 60788 14532
rect 61628 15260 61684 15316
rect 60508 13468 60564 13524
rect 60732 13244 60788 13300
rect 60620 13132 60676 13188
rect 62076 16828 62132 16884
rect 62188 17276 62244 17332
rect 62860 17724 62916 17780
rect 62412 16882 62468 16884
rect 62412 16830 62414 16882
rect 62414 16830 62466 16882
rect 62466 16830 62468 16882
rect 62412 16828 62468 16830
rect 62748 17164 62804 17220
rect 62076 16322 62132 16324
rect 62076 16270 62078 16322
rect 62078 16270 62130 16322
rect 62130 16270 62132 16322
rect 62076 16268 62132 16270
rect 62188 15372 62244 15428
rect 61404 14530 61460 14532
rect 61404 14478 61406 14530
rect 61406 14478 61458 14530
rect 61458 14478 61460 14530
rect 61404 14476 61460 14478
rect 61628 14530 61684 14532
rect 61628 14478 61630 14530
rect 61630 14478 61682 14530
rect 61682 14478 61684 14530
rect 61628 14476 61684 14478
rect 61068 14028 61124 14084
rect 60956 13244 61012 13300
rect 61068 13356 61124 13412
rect 61516 13356 61572 13412
rect 61628 13468 61684 13524
rect 61404 13244 61460 13300
rect 60620 12796 60676 12852
rect 60508 12460 60564 12516
rect 60844 12460 60900 12516
rect 61292 12290 61348 12292
rect 61292 12238 61294 12290
rect 61294 12238 61346 12290
rect 61346 12238 61348 12290
rect 61292 12236 61348 12238
rect 60732 11452 60788 11508
rect 60508 11282 60564 11284
rect 60508 11230 60510 11282
rect 60510 11230 60562 11282
rect 60562 11230 60564 11282
rect 60508 11228 60564 11230
rect 60396 9996 60452 10052
rect 60844 10780 60900 10836
rect 60844 9660 60900 9716
rect 60732 9100 60788 9156
rect 60284 7532 60340 7588
rect 59948 5068 60004 5124
rect 60284 5964 60340 6020
rect 59388 1596 59444 1652
rect 59276 1148 59332 1204
rect 60508 7084 60564 7140
rect 61068 9714 61124 9716
rect 61068 9662 61070 9714
rect 61070 9662 61122 9714
rect 61122 9662 61124 9714
rect 61068 9660 61124 9662
rect 61740 13186 61796 13188
rect 61740 13134 61742 13186
rect 61742 13134 61794 13186
rect 61794 13134 61796 13186
rect 61740 13132 61796 13134
rect 61292 10332 61348 10388
rect 61516 12460 61572 12516
rect 61740 12236 61796 12292
rect 61628 11452 61684 11508
rect 62076 14924 62132 14980
rect 62188 14476 62244 14532
rect 62076 14028 62132 14084
rect 61964 13916 62020 13972
rect 61964 11452 62020 11508
rect 61852 11340 61908 11396
rect 62524 14476 62580 14532
rect 62524 13858 62580 13860
rect 62524 13806 62526 13858
rect 62526 13806 62578 13858
rect 62578 13806 62580 13858
rect 62524 13804 62580 13806
rect 64764 24834 64820 24836
rect 64764 24782 64766 24834
rect 64766 24782 64818 24834
rect 64818 24782 64820 24834
rect 64764 24780 64820 24782
rect 64428 24220 64484 24276
rect 63084 23042 63140 23044
rect 63084 22990 63086 23042
rect 63086 22990 63138 23042
rect 63138 22990 63140 23042
rect 63084 22988 63140 22990
rect 63308 20972 63364 21028
rect 63868 22764 63924 22820
rect 63420 18620 63476 18676
rect 63532 22316 63588 22372
rect 63084 18338 63140 18340
rect 63084 18286 63086 18338
rect 63086 18286 63138 18338
rect 63138 18286 63140 18338
rect 63084 18284 63140 18286
rect 62748 14812 62804 14868
rect 62860 16716 62916 16772
rect 63420 16882 63476 16884
rect 63420 16830 63422 16882
rect 63422 16830 63474 16882
rect 63474 16830 63476 16882
rect 63420 16828 63476 16830
rect 63084 16268 63140 16324
rect 63196 15314 63252 15316
rect 63196 15262 63198 15314
rect 63198 15262 63250 15314
rect 63250 15262 63252 15314
rect 63196 15260 63252 15262
rect 63084 15148 63140 15204
rect 63868 22092 63924 22148
rect 63644 21756 63700 21812
rect 64092 21084 64148 21140
rect 64764 22764 64820 22820
rect 65436 24892 65492 24948
rect 65772 24556 65828 24612
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 67788 24668 67844 24724
rect 68012 25116 68068 25172
rect 67788 24050 67844 24052
rect 67788 23998 67790 24050
rect 67790 23998 67842 24050
rect 67842 23998 67844 24050
rect 67788 23996 67844 23998
rect 68012 23772 68068 23828
rect 65324 22764 65380 22820
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 63868 19740 63924 19796
rect 64428 20860 64484 20916
rect 64092 20412 64148 20468
rect 64652 20748 64708 20804
rect 64204 19234 64260 19236
rect 64204 19182 64206 19234
rect 64206 19182 64258 19234
rect 64258 19182 64260 19234
rect 64204 19180 64260 19182
rect 64204 18508 64260 18564
rect 64652 19180 64708 19236
rect 64540 19068 64596 19124
rect 64316 17948 64372 18004
rect 64764 18620 64820 18676
rect 63868 17666 63924 17668
rect 63868 17614 63870 17666
rect 63870 17614 63922 17666
rect 63922 17614 63924 17666
rect 63868 17612 63924 17614
rect 63756 17052 63812 17108
rect 64540 17106 64596 17108
rect 64540 17054 64542 17106
rect 64542 17054 64594 17106
rect 64594 17054 64596 17106
rect 64540 17052 64596 17054
rect 64540 16828 64596 16884
rect 62860 14924 62916 14980
rect 62860 14028 62916 14084
rect 62748 13244 62804 13300
rect 62076 11340 62132 11396
rect 61628 11116 61684 11172
rect 61964 11170 62020 11172
rect 61964 11118 61966 11170
rect 61966 11118 62018 11170
rect 62018 11118 62020 11170
rect 61964 11116 62020 11118
rect 61964 10892 62020 10948
rect 61180 9548 61236 9604
rect 61180 9266 61236 9268
rect 61180 9214 61182 9266
rect 61182 9214 61234 9266
rect 61234 9214 61236 9266
rect 61180 9212 61236 9214
rect 62188 10668 62244 10724
rect 62076 10332 62132 10388
rect 61740 9324 61796 9380
rect 61852 8988 61908 9044
rect 62076 8988 62132 9044
rect 61740 8316 61796 8372
rect 60844 7362 60900 7364
rect 60844 7310 60846 7362
rect 60846 7310 60898 7362
rect 60898 7310 60900 7362
rect 60844 7308 60900 7310
rect 60844 7084 60900 7140
rect 60732 6690 60788 6692
rect 60732 6638 60734 6690
rect 60734 6638 60786 6690
rect 60786 6638 60788 6690
rect 60732 6636 60788 6638
rect 60620 6018 60676 6020
rect 60620 5966 60622 6018
rect 60622 5966 60674 6018
rect 60674 5966 60676 6018
rect 60620 5964 60676 5966
rect 61068 7308 61124 7364
rect 61068 6914 61124 6916
rect 61068 6862 61070 6914
rect 61070 6862 61122 6914
rect 61122 6862 61124 6914
rect 61068 6860 61124 6862
rect 60396 4956 60452 5012
rect 61292 7532 61348 7588
rect 61516 7084 61572 7140
rect 61180 6524 61236 6580
rect 61852 8204 61908 8260
rect 61964 7532 62020 7588
rect 61852 7084 61908 7140
rect 62412 10780 62468 10836
rect 63308 15036 63364 15092
rect 63644 15372 63700 15428
rect 63756 15314 63812 15316
rect 63756 15262 63758 15314
rect 63758 15262 63810 15314
rect 63810 15262 63812 15314
rect 63756 15260 63812 15262
rect 63644 14476 63700 14532
rect 63756 14588 63812 14644
rect 63756 13970 63812 13972
rect 63756 13918 63758 13970
rect 63758 13918 63810 13970
rect 63810 13918 63812 13970
rect 63756 13916 63812 13918
rect 63420 13074 63476 13076
rect 63420 13022 63422 13074
rect 63422 13022 63474 13074
rect 63474 13022 63476 13074
rect 63420 13020 63476 13022
rect 63868 13020 63924 13076
rect 63084 12124 63140 12180
rect 62972 11788 63028 11844
rect 62524 9826 62580 9828
rect 62524 9774 62526 9826
rect 62526 9774 62578 9826
rect 62578 9774 62580 9826
rect 62524 9772 62580 9774
rect 62860 10780 62916 10836
rect 62972 10668 63028 10724
rect 63084 10556 63140 10612
rect 62412 9266 62468 9268
rect 62412 9214 62414 9266
rect 62414 9214 62466 9266
rect 62466 9214 62468 9266
rect 62412 9212 62468 9214
rect 61740 6412 61796 6468
rect 62300 8540 62356 8596
rect 63084 9772 63140 9828
rect 63420 10556 63476 10612
rect 63420 9826 63476 9828
rect 63420 9774 63422 9826
rect 63422 9774 63474 9826
rect 63474 9774 63476 9826
rect 63420 9772 63476 9774
rect 62860 9602 62916 9604
rect 62860 9550 62862 9602
rect 62862 9550 62914 9602
rect 62914 9550 62916 9602
rect 62860 9548 62916 9550
rect 62748 9042 62804 9044
rect 62748 8990 62750 9042
rect 62750 8990 62802 9042
rect 62802 8990 62804 9042
rect 62748 8988 62804 8990
rect 63420 9042 63476 9044
rect 63420 8990 63422 9042
rect 63422 8990 63474 9042
rect 63474 8990 63476 9042
rect 63420 8988 63476 8990
rect 62636 8540 62692 8596
rect 62524 7756 62580 7812
rect 63420 8316 63476 8372
rect 62860 7644 62916 7700
rect 63196 6748 63252 6804
rect 63308 7308 63364 7364
rect 62188 6412 62244 6468
rect 63084 6412 63140 6468
rect 61516 4620 61572 4676
rect 61404 2492 61460 2548
rect 61964 5068 62020 5124
rect 61740 4956 61796 5012
rect 62524 4396 62580 4452
rect 61740 3442 61796 3444
rect 61740 3390 61742 3442
rect 61742 3390 61794 3442
rect 61794 3390 61796 3442
rect 61740 3388 61796 3390
rect 63420 7084 63476 7140
rect 63532 7756 63588 7812
rect 63308 4060 63364 4116
rect 64988 19740 65044 19796
rect 65212 20802 65268 20804
rect 65212 20750 65214 20802
rect 65214 20750 65266 20802
rect 65266 20750 65268 20802
rect 65212 20748 65268 20750
rect 65324 20076 65380 20132
rect 65436 22540 65492 22596
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 66556 20860 66612 20916
rect 64540 14812 64596 14868
rect 65436 19628 65492 19684
rect 65100 18620 65156 18676
rect 65100 17612 65156 17668
rect 64764 14140 64820 14196
rect 64428 13746 64484 13748
rect 64428 13694 64430 13746
rect 64430 13694 64482 13746
rect 64482 13694 64484 13746
rect 64428 13692 64484 13694
rect 64092 13020 64148 13076
rect 63980 10556 64036 10612
rect 64204 11340 64260 11396
rect 64316 11004 64372 11060
rect 64204 9714 64260 9716
rect 64204 9662 64206 9714
rect 64206 9662 64258 9714
rect 64258 9662 64260 9714
rect 64204 9660 64260 9662
rect 63980 8930 64036 8932
rect 63980 8878 63982 8930
rect 63982 8878 64034 8930
rect 64034 8878 64036 8930
rect 63980 8876 64036 8878
rect 63980 8428 64036 8484
rect 63868 5852 63924 5908
rect 63644 4844 63700 4900
rect 64316 9548 64372 9604
rect 66220 19740 66276 19796
rect 66332 20412 66388 20468
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 65772 19068 65828 19124
rect 66892 20076 66948 20132
rect 66780 19346 66836 19348
rect 66780 19294 66782 19346
rect 66782 19294 66834 19346
rect 66834 19294 66836 19346
rect 66780 19292 66836 19294
rect 69356 28418 69412 28420
rect 69356 28366 69358 28418
rect 69358 28366 69410 28418
rect 69410 28366 69412 28418
rect 69356 28364 69412 28366
rect 68460 27020 68516 27076
rect 68796 26572 68852 26628
rect 68348 26402 68404 26404
rect 68348 26350 68350 26402
rect 68350 26350 68402 26402
rect 68402 26350 68404 26402
rect 68348 26348 68404 26350
rect 69132 26572 69188 26628
rect 68908 25228 68964 25284
rect 68684 25116 68740 25172
rect 68908 24946 68964 24948
rect 68908 24894 68910 24946
rect 68910 24894 68962 24946
rect 68962 24894 68964 24946
rect 68908 24892 68964 24894
rect 68348 24722 68404 24724
rect 68348 24670 68350 24722
rect 68350 24670 68402 24722
rect 68402 24670 68404 24722
rect 68348 24668 68404 24670
rect 68908 24668 68964 24724
rect 69020 23996 69076 24052
rect 68796 23826 68852 23828
rect 68796 23774 68798 23826
rect 68798 23774 68850 23826
rect 68850 23774 68852 23826
rect 68796 23772 68852 23774
rect 73388 30492 73444 30548
rect 72716 28364 72772 28420
rect 70364 27858 70420 27860
rect 70364 27806 70366 27858
rect 70366 27806 70418 27858
rect 70418 27806 70420 27858
rect 70364 27804 70420 27806
rect 70700 27580 70756 27636
rect 69580 27186 69636 27188
rect 69580 27134 69582 27186
rect 69582 27134 69634 27186
rect 69634 27134 69636 27186
rect 69580 27132 69636 27134
rect 70140 27356 70196 27412
rect 69468 26348 69524 26404
rect 69244 25116 69300 25172
rect 69468 25228 69524 25284
rect 69356 25004 69412 25060
rect 69244 24050 69300 24052
rect 69244 23998 69246 24050
rect 69246 23998 69298 24050
rect 69298 23998 69300 24050
rect 69244 23996 69300 23998
rect 69580 25116 69636 25172
rect 69468 24610 69524 24612
rect 69468 24558 69470 24610
rect 69470 24558 69522 24610
rect 69522 24558 69524 24610
rect 69468 24556 69524 24558
rect 69356 23826 69412 23828
rect 69356 23774 69358 23826
rect 69358 23774 69410 23826
rect 69410 23774 69412 23826
rect 69356 23772 69412 23774
rect 68572 23436 68628 23492
rect 68012 20972 68068 21028
rect 69804 26908 69860 26964
rect 70364 27074 70420 27076
rect 70364 27022 70366 27074
rect 70366 27022 70418 27074
rect 70418 27022 70420 27074
rect 70364 27020 70420 27022
rect 71372 28028 71428 28084
rect 71148 27356 71204 27412
rect 71596 27298 71652 27300
rect 71596 27246 71598 27298
rect 71598 27246 71650 27298
rect 71650 27246 71652 27298
rect 71596 27244 71652 27246
rect 71708 27074 71764 27076
rect 71708 27022 71710 27074
rect 71710 27022 71762 27074
rect 71762 27022 71764 27074
rect 71708 27020 71764 27022
rect 72380 27244 72436 27300
rect 70252 26796 70308 26852
rect 71260 26962 71316 26964
rect 71260 26910 71262 26962
rect 71262 26910 71314 26962
rect 71314 26910 71316 26962
rect 71260 26908 71316 26910
rect 70476 26572 70532 26628
rect 70476 25564 70532 25620
rect 70700 25506 70756 25508
rect 70700 25454 70702 25506
rect 70702 25454 70754 25506
rect 70754 25454 70756 25506
rect 70700 25452 70756 25454
rect 69916 25394 69972 25396
rect 69916 25342 69918 25394
rect 69918 25342 69970 25394
rect 69970 25342 69972 25394
rect 69916 25340 69972 25342
rect 70028 25228 70084 25284
rect 70588 25282 70644 25284
rect 70588 25230 70590 25282
rect 70590 25230 70642 25282
rect 70642 25230 70644 25282
rect 70588 25228 70644 25230
rect 70364 25116 70420 25172
rect 70364 24722 70420 24724
rect 70364 24670 70366 24722
rect 70366 24670 70418 24722
rect 70418 24670 70420 24722
rect 70364 24668 70420 24670
rect 71260 24892 71316 24948
rect 71148 24834 71204 24836
rect 71148 24782 71150 24834
rect 71150 24782 71202 24834
rect 71202 24782 71204 24834
rect 71148 24780 71204 24782
rect 71708 26514 71764 26516
rect 71708 26462 71710 26514
rect 71710 26462 71762 26514
rect 71762 26462 71764 26514
rect 71708 26460 71764 26462
rect 72156 26460 72212 26516
rect 73276 27074 73332 27076
rect 73276 27022 73278 27074
rect 73278 27022 73330 27074
rect 73330 27022 73332 27074
rect 73276 27020 73332 27022
rect 73948 27580 74004 27636
rect 73612 27244 73668 27300
rect 73724 26962 73780 26964
rect 73724 26910 73726 26962
rect 73726 26910 73778 26962
rect 73778 26910 73780 26962
rect 73724 26908 73780 26910
rect 73948 26962 74004 26964
rect 73948 26910 73950 26962
rect 73950 26910 74002 26962
rect 74002 26910 74004 26962
rect 73948 26908 74004 26910
rect 72828 26796 72884 26852
rect 71596 25618 71652 25620
rect 71596 25566 71598 25618
rect 71598 25566 71650 25618
rect 71650 25566 71652 25618
rect 71596 25564 71652 25566
rect 71708 26124 71764 26180
rect 72828 26290 72884 26292
rect 72828 26238 72830 26290
rect 72830 26238 72882 26290
rect 72882 26238 72884 26290
rect 72828 26236 72884 26238
rect 74284 27746 74340 27748
rect 74284 27694 74286 27746
rect 74286 27694 74338 27746
rect 74338 27694 74340 27746
rect 74284 27692 74340 27694
rect 74172 27132 74228 27188
rect 74060 26796 74116 26852
rect 73948 26402 74004 26404
rect 73948 26350 73950 26402
rect 73950 26350 74002 26402
rect 74002 26350 74004 26402
rect 73948 26348 74004 26350
rect 73836 26290 73892 26292
rect 73836 26238 73838 26290
rect 73838 26238 73890 26290
rect 73890 26238 73892 26290
rect 73836 26236 73892 26238
rect 72044 25506 72100 25508
rect 72044 25454 72046 25506
rect 72046 25454 72098 25506
rect 72098 25454 72100 25506
rect 72044 25452 72100 25454
rect 72492 25004 72548 25060
rect 72716 25340 72772 25396
rect 72604 24892 72660 24948
rect 71708 24834 71764 24836
rect 71708 24782 71710 24834
rect 71710 24782 71762 24834
rect 71762 24782 71764 24834
rect 71708 24780 71764 24782
rect 71372 24444 71428 24500
rect 74396 26236 74452 26292
rect 74172 25004 74228 25060
rect 74396 24892 74452 24948
rect 73388 24668 73444 24724
rect 73052 24050 73108 24052
rect 73052 23998 73054 24050
rect 73054 23998 73106 24050
rect 73106 23998 73108 24050
rect 73052 23996 73108 23998
rect 74172 24780 74228 24836
rect 74172 23996 74228 24052
rect 72268 23100 72324 23156
rect 72492 23154 72548 23156
rect 72492 23102 72494 23154
rect 72494 23102 72546 23154
rect 72546 23102 72548 23154
rect 72492 23100 72548 23102
rect 73052 22988 73108 23044
rect 77196 29372 77252 29428
rect 81116 55186 81172 55188
rect 81116 55134 81118 55186
rect 81118 55134 81170 55186
rect 81170 55134 81172 55186
rect 81116 55132 81172 55134
rect 81564 55132 81620 55188
rect 93212 56252 93268 56308
rect 94444 56306 94500 56308
rect 94444 56254 94446 56306
rect 94446 56254 94498 56306
rect 94498 56254 94500 56306
rect 94444 56252 94500 56254
rect 97020 56252 97076 56308
rect 98252 56306 98308 56308
rect 98252 56254 98254 56306
rect 98254 56254 98306 56306
rect 98306 56254 98308 56306
rect 98252 56252 98308 56254
rect 96636 55690 96692 55692
rect 96636 55638 96638 55690
rect 96638 55638 96690 55690
rect 96690 55638 96692 55690
rect 96636 55636 96692 55638
rect 96740 55690 96796 55692
rect 96740 55638 96742 55690
rect 96742 55638 96794 55690
rect 96794 55638 96796 55690
rect 96740 55636 96796 55638
rect 96844 55690 96900 55692
rect 96844 55638 96846 55690
rect 96846 55638 96898 55690
rect 96898 55638 96900 55690
rect 96844 55636 96900 55638
rect 81276 54906 81332 54908
rect 81276 54854 81278 54906
rect 81278 54854 81330 54906
rect 81330 54854 81332 54906
rect 81276 54852 81332 54854
rect 81380 54906 81436 54908
rect 81380 54854 81382 54906
rect 81382 54854 81434 54906
rect 81434 54854 81436 54906
rect 81380 54852 81436 54854
rect 81484 54906 81540 54908
rect 81484 54854 81486 54906
rect 81486 54854 81538 54906
rect 81538 54854 81540 54906
rect 81484 54852 81540 54854
rect 81276 53338 81332 53340
rect 81276 53286 81278 53338
rect 81278 53286 81330 53338
rect 81330 53286 81332 53338
rect 81276 53284 81332 53286
rect 81380 53338 81436 53340
rect 81380 53286 81382 53338
rect 81382 53286 81434 53338
rect 81434 53286 81436 53338
rect 81380 53284 81436 53286
rect 81484 53338 81540 53340
rect 81484 53286 81486 53338
rect 81486 53286 81538 53338
rect 81538 53286 81540 53338
rect 81484 53284 81540 53286
rect 81276 51770 81332 51772
rect 81276 51718 81278 51770
rect 81278 51718 81330 51770
rect 81330 51718 81332 51770
rect 81276 51716 81332 51718
rect 81380 51770 81436 51772
rect 81380 51718 81382 51770
rect 81382 51718 81434 51770
rect 81434 51718 81436 51770
rect 81380 51716 81436 51718
rect 81484 51770 81540 51772
rect 81484 51718 81486 51770
rect 81486 51718 81538 51770
rect 81538 51718 81540 51770
rect 81484 51716 81540 51718
rect 81276 50202 81332 50204
rect 81276 50150 81278 50202
rect 81278 50150 81330 50202
rect 81330 50150 81332 50202
rect 81276 50148 81332 50150
rect 81380 50202 81436 50204
rect 81380 50150 81382 50202
rect 81382 50150 81434 50202
rect 81434 50150 81436 50202
rect 81380 50148 81436 50150
rect 81484 50202 81540 50204
rect 81484 50150 81486 50202
rect 81486 50150 81538 50202
rect 81538 50150 81540 50202
rect 81484 50148 81540 50150
rect 81276 48634 81332 48636
rect 81276 48582 81278 48634
rect 81278 48582 81330 48634
rect 81330 48582 81332 48634
rect 81276 48580 81332 48582
rect 81380 48634 81436 48636
rect 81380 48582 81382 48634
rect 81382 48582 81434 48634
rect 81434 48582 81436 48634
rect 81380 48580 81436 48582
rect 81484 48634 81540 48636
rect 81484 48582 81486 48634
rect 81486 48582 81538 48634
rect 81538 48582 81540 48634
rect 81484 48580 81540 48582
rect 81276 47066 81332 47068
rect 81276 47014 81278 47066
rect 81278 47014 81330 47066
rect 81330 47014 81332 47066
rect 81276 47012 81332 47014
rect 81380 47066 81436 47068
rect 81380 47014 81382 47066
rect 81382 47014 81434 47066
rect 81434 47014 81436 47066
rect 81380 47012 81436 47014
rect 81484 47066 81540 47068
rect 81484 47014 81486 47066
rect 81486 47014 81538 47066
rect 81538 47014 81540 47066
rect 81484 47012 81540 47014
rect 81276 45498 81332 45500
rect 81276 45446 81278 45498
rect 81278 45446 81330 45498
rect 81330 45446 81332 45498
rect 81276 45444 81332 45446
rect 81380 45498 81436 45500
rect 81380 45446 81382 45498
rect 81382 45446 81434 45498
rect 81434 45446 81436 45498
rect 81380 45444 81436 45446
rect 81484 45498 81540 45500
rect 81484 45446 81486 45498
rect 81486 45446 81538 45498
rect 81538 45446 81540 45498
rect 81484 45444 81540 45446
rect 81276 43930 81332 43932
rect 81276 43878 81278 43930
rect 81278 43878 81330 43930
rect 81330 43878 81332 43930
rect 81276 43876 81332 43878
rect 81380 43930 81436 43932
rect 81380 43878 81382 43930
rect 81382 43878 81434 43930
rect 81434 43878 81436 43930
rect 81380 43876 81436 43878
rect 81484 43930 81540 43932
rect 81484 43878 81486 43930
rect 81486 43878 81538 43930
rect 81538 43878 81540 43930
rect 81484 43876 81540 43878
rect 81276 42362 81332 42364
rect 81276 42310 81278 42362
rect 81278 42310 81330 42362
rect 81330 42310 81332 42362
rect 81276 42308 81332 42310
rect 81380 42362 81436 42364
rect 81380 42310 81382 42362
rect 81382 42310 81434 42362
rect 81434 42310 81436 42362
rect 81380 42308 81436 42310
rect 81484 42362 81540 42364
rect 81484 42310 81486 42362
rect 81486 42310 81538 42362
rect 81538 42310 81540 42362
rect 81484 42308 81540 42310
rect 81276 40794 81332 40796
rect 81276 40742 81278 40794
rect 81278 40742 81330 40794
rect 81330 40742 81332 40794
rect 81276 40740 81332 40742
rect 81380 40794 81436 40796
rect 81380 40742 81382 40794
rect 81382 40742 81434 40794
rect 81434 40742 81436 40794
rect 81380 40740 81436 40742
rect 81484 40794 81540 40796
rect 81484 40742 81486 40794
rect 81486 40742 81538 40794
rect 81538 40742 81540 40794
rect 81484 40740 81540 40742
rect 81276 39226 81332 39228
rect 81276 39174 81278 39226
rect 81278 39174 81330 39226
rect 81330 39174 81332 39226
rect 81276 39172 81332 39174
rect 81380 39226 81436 39228
rect 81380 39174 81382 39226
rect 81382 39174 81434 39226
rect 81434 39174 81436 39226
rect 81380 39172 81436 39174
rect 81484 39226 81540 39228
rect 81484 39174 81486 39226
rect 81486 39174 81538 39226
rect 81538 39174 81540 39226
rect 81484 39172 81540 39174
rect 81276 37658 81332 37660
rect 81276 37606 81278 37658
rect 81278 37606 81330 37658
rect 81330 37606 81332 37658
rect 81276 37604 81332 37606
rect 81380 37658 81436 37660
rect 81380 37606 81382 37658
rect 81382 37606 81434 37658
rect 81434 37606 81436 37658
rect 81380 37604 81436 37606
rect 81484 37658 81540 37660
rect 81484 37606 81486 37658
rect 81486 37606 81538 37658
rect 81538 37606 81540 37658
rect 81484 37604 81540 37606
rect 81276 36090 81332 36092
rect 81276 36038 81278 36090
rect 81278 36038 81330 36090
rect 81330 36038 81332 36090
rect 81276 36036 81332 36038
rect 81380 36090 81436 36092
rect 81380 36038 81382 36090
rect 81382 36038 81434 36090
rect 81434 36038 81436 36090
rect 81380 36036 81436 36038
rect 81484 36090 81540 36092
rect 81484 36038 81486 36090
rect 81486 36038 81538 36090
rect 81538 36038 81540 36090
rect 81484 36036 81540 36038
rect 81276 34522 81332 34524
rect 81276 34470 81278 34522
rect 81278 34470 81330 34522
rect 81330 34470 81332 34522
rect 81276 34468 81332 34470
rect 81380 34522 81436 34524
rect 81380 34470 81382 34522
rect 81382 34470 81434 34522
rect 81434 34470 81436 34522
rect 81380 34468 81436 34470
rect 81484 34522 81540 34524
rect 81484 34470 81486 34522
rect 81486 34470 81538 34522
rect 81538 34470 81540 34522
rect 81484 34468 81540 34470
rect 81276 32954 81332 32956
rect 81276 32902 81278 32954
rect 81278 32902 81330 32954
rect 81330 32902 81332 32954
rect 81276 32900 81332 32902
rect 81380 32954 81436 32956
rect 81380 32902 81382 32954
rect 81382 32902 81434 32954
rect 81434 32902 81436 32954
rect 81380 32900 81436 32902
rect 81484 32954 81540 32956
rect 81484 32902 81486 32954
rect 81486 32902 81538 32954
rect 81538 32902 81540 32954
rect 81484 32900 81540 32902
rect 81276 31386 81332 31388
rect 81276 31334 81278 31386
rect 81278 31334 81330 31386
rect 81330 31334 81332 31386
rect 81276 31332 81332 31334
rect 81380 31386 81436 31388
rect 81380 31334 81382 31386
rect 81382 31334 81434 31386
rect 81434 31334 81436 31386
rect 81380 31332 81436 31334
rect 81484 31386 81540 31388
rect 81484 31334 81486 31386
rect 81486 31334 81538 31386
rect 81538 31334 81540 31386
rect 81484 31332 81540 31334
rect 81276 29818 81332 29820
rect 81276 29766 81278 29818
rect 81278 29766 81330 29818
rect 81330 29766 81332 29818
rect 81276 29764 81332 29766
rect 81380 29818 81436 29820
rect 81380 29766 81382 29818
rect 81382 29766 81434 29818
rect 81434 29766 81436 29818
rect 81380 29764 81436 29766
rect 81484 29818 81540 29820
rect 81484 29766 81486 29818
rect 81486 29766 81538 29818
rect 81538 29766 81540 29818
rect 81484 29764 81540 29766
rect 83244 29372 83300 29428
rect 81276 28250 81332 28252
rect 81276 28198 81278 28250
rect 81278 28198 81330 28250
rect 81330 28198 81332 28250
rect 81276 28196 81332 28198
rect 81380 28250 81436 28252
rect 81380 28198 81382 28250
rect 81382 28198 81434 28250
rect 81434 28198 81436 28250
rect 81380 28196 81436 28198
rect 81484 28250 81540 28252
rect 81484 28198 81486 28250
rect 81486 28198 81538 28250
rect 81538 28198 81540 28250
rect 81484 28196 81540 28198
rect 77308 27804 77364 27860
rect 75852 27692 75908 27748
rect 75292 27356 75348 27412
rect 74732 27132 74788 27188
rect 75180 27186 75236 27188
rect 75180 27134 75182 27186
rect 75182 27134 75234 27186
rect 75234 27134 75236 27186
rect 75180 27132 75236 27134
rect 74956 26908 75012 26964
rect 75068 26796 75124 26852
rect 74844 25676 74900 25732
rect 74732 24892 74788 24948
rect 74844 24834 74900 24836
rect 74844 24782 74846 24834
rect 74846 24782 74898 24834
rect 74898 24782 74900 24834
rect 74844 24780 74900 24782
rect 74732 24722 74788 24724
rect 74732 24670 74734 24722
rect 74734 24670 74786 24722
rect 74786 24670 74788 24722
rect 74732 24668 74788 24670
rect 75068 23714 75124 23716
rect 75068 23662 75070 23714
rect 75070 23662 75122 23714
rect 75122 23662 75124 23714
rect 75068 23660 75124 23662
rect 77196 27580 77252 27636
rect 76188 27074 76244 27076
rect 76188 27022 76190 27074
rect 76190 27022 76242 27074
rect 76242 27022 76244 27074
rect 76188 27020 76244 27022
rect 75516 26290 75572 26292
rect 75516 26238 75518 26290
rect 75518 26238 75570 26290
rect 75570 26238 75572 26290
rect 75516 26236 75572 26238
rect 75292 24610 75348 24612
rect 75292 24558 75294 24610
rect 75294 24558 75346 24610
rect 75346 24558 75348 24610
rect 75292 24556 75348 24558
rect 75180 22876 75236 22932
rect 68908 20188 68964 20244
rect 69132 21644 69188 21700
rect 67004 19852 67060 19908
rect 67004 19234 67060 19236
rect 67004 19182 67006 19234
rect 67006 19182 67058 19234
rect 67058 19182 67060 19234
rect 67004 19180 67060 19182
rect 66556 19122 66612 19124
rect 66556 19070 66558 19122
rect 66558 19070 66610 19122
rect 66610 19070 66612 19122
rect 66556 19068 66612 19070
rect 73836 22204 73892 22260
rect 70476 21196 70532 21252
rect 74172 21586 74228 21588
rect 74172 21534 74174 21586
rect 74174 21534 74226 21586
rect 74226 21534 74228 21586
rect 74172 21532 74228 21534
rect 72828 21420 72884 21476
rect 67676 19740 67732 19796
rect 67564 19234 67620 19236
rect 67564 19182 67566 19234
rect 67566 19182 67618 19234
rect 67618 19182 67620 19234
rect 67564 19180 67620 19182
rect 66444 18508 66500 18564
rect 66556 18450 66612 18452
rect 66556 18398 66558 18450
rect 66558 18398 66610 18450
rect 66610 18398 66612 18450
rect 66556 18396 66612 18398
rect 65548 18060 65604 18116
rect 65916 18058 65972 18060
rect 65772 17948 65828 18004
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 65660 17666 65716 17668
rect 65660 17614 65662 17666
rect 65662 17614 65714 17666
rect 65714 17614 65716 17666
rect 65660 17612 65716 17614
rect 65548 16828 65604 16884
rect 65772 17500 65828 17556
rect 65324 14812 65380 14868
rect 65324 14418 65380 14420
rect 65324 14366 65326 14418
rect 65326 14366 65378 14418
rect 65378 14366 65380 14418
rect 65324 14364 65380 14366
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 66444 15932 66500 15988
rect 67340 18508 67396 18564
rect 66668 15036 66724 15092
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 66332 14924 66388 14980
rect 65548 13916 65604 13972
rect 65772 14028 65828 14084
rect 65660 13858 65716 13860
rect 65660 13806 65662 13858
rect 65662 13806 65714 13858
rect 65714 13806 65716 13858
rect 65660 13804 65716 13806
rect 64876 11676 64932 11732
rect 64540 11228 64596 11284
rect 66220 13916 66276 13972
rect 66444 14418 66500 14420
rect 66444 14366 66446 14418
rect 66446 14366 66498 14418
rect 66498 14366 66500 14418
rect 66444 14364 66500 14366
rect 66668 14140 66724 14196
rect 66780 14028 66836 14084
rect 66332 13804 66388 13860
rect 64988 11564 65044 11620
rect 64652 10892 64708 10948
rect 64988 11228 65044 11284
rect 64540 9884 64596 9940
rect 65100 11170 65156 11172
rect 65100 11118 65102 11170
rect 65102 11118 65154 11170
rect 65154 11118 65156 11170
rect 65100 11116 65156 11118
rect 64876 10556 64932 10612
rect 64764 9772 64820 9828
rect 64540 8428 64596 8484
rect 64876 9100 64932 9156
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 65996 12066 66052 12068
rect 65996 12014 65998 12066
rect 65998 12014 66050 12066
rect 66050 12014 66052 12066
rect 65996 12012 66052 12014
rect 67340 16716 67396 16772
rect 67788 17442 67844 17444
rect 67788 17390 67790 17442
rect 67790 17390 67842 17442
rect 67842 17390 67844 17442
rect 67788 17388 67844 17390
rect 67340 15036 67396 15092
rect 68572 19180 68628 19236
rect 69468 18450 69524 18452
rect 69468 18398 69470 18450
rect 69470 18398 69522 18450
rect 69522 18398 69524 18450
rect 69468 18396 69524 18398
rect 69804 18284 69860 18340
rect 69916 19852 69972 19908
rect 69692 17724 69748 17780
rect 68908 17666 68964 17668
rect 68908 17614 68910 17666
rect 68910 17614 68962 17666
rect 68962 17614 68964 17666
rect 68908 17612 68964 17614
rect 69356 17612 69412 17668
rect 68684 17554 68740 17556
rect 68684 17502 68686 17554
rect 68686 17502 68738 17554
rect 68738 17502 68740 17554
rect 68684 17500 68740 17502
rect 69580 17388 69636 17444
rect 68460 17052 68516 17108
rect 68908 16994 68964 16996
rect 68908 16942 68910 16994
rect 68910 16942 68962 16994
rect 68962 16942 68964 16994
rect 68908 16940 68964 16942
rect 68348 15932 68404 15988
rect 68460 15314 68516 15316
rect 68460 15262 68462 15314
rect 68462 15262 68514 15314
rect 68514 15262 68516 15314
rect 68460 15260 68516 15262
rect 68012 15148 68068 15204
rect 67788 14700 67844 14756
rect 67004 12796 67060 12852
rect 67116 13356 67172 13412
rect 66892 11900 66948 11956
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 66332 11676 66388 11732
rect 66220 11452 66276 11508
rect 65436 11394 65492 11396
rect 65436 11342 65438 11394
rect 65438 11342 65490 11394
rect 65490 11342 65492 11394
rect 65436 11340 65492 11342
rect 65324 9772 65380 9828
rect 65436 10892 65492 10948
rect 65212 9714 65268 9716
rect 65212 9662 65214 9714
rect 65214 9662 65266 9714
rect 65266 9662 65268 9714
rect 65212 9660 65268 9662
rect 65212 9100 65268 9156
rect 64764 8204 64820 8260
rect 64876 8876 64932 8932
rect 64764 7868 64820 7924
rect 64428 7698 64484 7700
rect 64428 7646 64430 7698
rect 64430 7646 64482 7698
rect 64482 7646 64484 7698
rect 64428 7644 64484 7646
rect 64204 6860 64260 6916
rect 64316 7532 64372 7588
rect 64652 7420 64708 7476
rect 64092 5740 64148 5796
rect 67116 12012 67172 12068
rect 66668 11676 66724 11732
rect 66556 11228 66612 11284
rect 66892 11282 66948 11284
rect 66892 11230 66894 11282
rect 66894 11230 66946 11282
rect 66946 11230 66948 11282
rect 66892 11228 66948 11230
rect 66444 11116 66500 11172
rect 67564 11676 67620 11732
rect 67564 11004 67620 11060
rect 67228 10722 67284 10724
rect 67228 10670 67230 10722
rect 67230 10670 67282 10722
rect 67282 10670 67284 10722
rect 67228 10668 67284 10670
rect 66220 10556 66276 10612
rect 65884 10332 65940 10388
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 65436 9212 65492 9268
rect 64988 8204 65044 8260
rect 65436 8988 65492 9044
rect 65324 8316 65380 8372
rect 64764 6188 64820 6244
rect 64316 4620 64372 4676
rect 63084 2940 63140 2996
rect 64540 4620 64596 4676
rect 64876 5740 64932 5796
rect 65548 8764 65604 8820
rect 66444 9436 66500 9492
rect 65660 7868 65716 7924
rect 65772 9042 65828 9044
rect 65772 8990 65774 9042
rect 65774 8990 65826 9042
rect 65826 8990 65828 9042
rect 65772 8988 65828 8990
rect 66332 9042 66388 9044
rect 66332 8990 66334 9042
rect 66334 8990 66386 9042
rect 66386 8990 66388 9042
rect 66332 8988 66388 8990
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 67004 10108 67060 10164
rect 67228 10332 67284 10388
rect 66668 9660 66724 9716
rect 67004 9324 67060 9380
rect 67116 9548 67172 9604
rect 66892 9100 66948 9156
rect 66668 8258 66724 8260
rect 66668 8206 66670 8258
rect 66670 8206 66722 8258
rect 66722 8206 66724 8258
rect 66668 8204 66724 8206
rect 67452 9826 67508 9828
rect 67452 9774 67454 9826
rect 67454 9774 67506 9826
rect 67506 9774 67508 9826
rect 67452 9772 67508 9774
rect 67228 9042 67284 9044
rect 67228 8990 67230 9042
rect 67230 8990 67282 9042
rect 67282 8990 67284 9042
rect 67228 8988 67284 8990
rect 67228 8764 67284 8820
rect 66444 7868 66500 7924
rect 65436 7420 65492 7476
rect 66220 7362 66276 7364
rect 66220 7310 66222 7362
rect 66222 7310 66274 7362
rect 66274 7310 66276 7362
rect 66220 7308 66276 7310
rect 66668 7532 66724 7588
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 65436 6860 65492 6916
rect 66332 6578 66388 6580
rect 66332 6526 66334 6578
rect 66334 6526 66386 6578
rect 66386 6526 66388 6578
rect 66332 6524 66388 6526
rect 66332 5964 66388 6020
rect 65212 5068 65268 5124
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 65772 4956 65828 5012
rect 65548 4508 65604 4564
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 65884 3724 65940 3780
rect 64876 3666 64932 3668
rect 64876 3614 64878 3666
rect 64878 3614 64930 3666
rect 64930 3614 64932 3666
rect 64876 3612 64932 3614
rect 65660 3612 65716 3668
rect 66668 7196 66724 7252
rect 66892 6578 66948 6580
rect 66892 6526 66894 6578
rect 66894 6526 66946 6578
rect 66946 6526 66948 6578
rect 66892 6524 66948 6526
rect 66780 5292 66836 5348
rect 66556 4956 66612 5012
rect 66892 3612 66948 3668
rect 67116 7644 67172 7700
rect 67228 7868 67284 7924
rect 67116 7474 67172 7476
rect 67116 7422 67118 7474
rect 67118 7422 67170 7474
rect 67170 7422 67172 7474
rect 67116 7420 67172 7422
rect 67116 5740 67172 5796
rect 67452 8540 67508 8596
rect 67452 8316 67508 8372
rect 67452 7980 67508 8036
rect 67788 11116 67844 11172
rect 67900 11004 67956 11060
rect 69132 15986 69188 15988
rect 69132 15934 69134 15986
rect 69134 15934 69186 15986
rect 69186 15934 69188 15986
rect 69132 15932 69188 15934
rect 69692 15538 69748 15540
rect 69692 15486 69694 15538
rect 69694 15486 69746 15538
rect 69746 15486 69748 15538
rect 69692 15484 69748 15486
rect 69132 15202 69188 15204
rect 69132 15150 69134 15202
rect 69134 15150 69186 15202
rect 69186 15150 69188 15202
rect 69132 15148 69188 15150
rect 71260 19404 71316 19460
rect 70700 18450 70756 18452
rect 70700 18398 70702 18450
rect 70702 18398 70754 18450
rect 70754 18398 70756 18450
rect 70700 18396 70756 18398
rect 71372 19234 71428 19236
rect 71372 19182 71374 19234
rect 71374 19182 71426 19234
rect 71426 19182 71428 19234
rect 71372 19180 71428 19182
rect 73948 21474 74004 21476
rect 73948 21422 73950 21474
rect 73950 21422 74002 21474
rect 74002 21422 74004 21474
rect 73948 21420 74004 21422
rect 73948 21196 74004 21252
rect 72044 19180 72100 19236
rect 72940 20188 72996 20244
rect 71932 18508 71988 18564
rect 69020 14588 69076 14644
rect 68684 13916 68740 13972
rect 68908 14252 68964 14308
rect 68796 13244 68852 13300
rect 70476 17666 70532 17668
rect 70476 17614 70478 17666
rect 70478 17614 70530 17666
rect 70530 17614 70532 17666
rect 70476 17612 70532 17614
rect 70924 17666 70980 17668
rect 70924 17614 70926 17666
rect 70926 17614 70978 17666
rect 70978 17614 70980 17666
rect 70924 17612 70980 17614
rect 72268 18284 72324 18340
rect 72268 17948 72324 18004
rect 71820 17666 71876 17668
rect 71820 17614 71822 17666
rect 71822 17614 71874 17666
rect 71874 17614 71876 17666
rect 71820 17612 71876 17614
rect 72492 17388 72548 17444
rect 71596 16940 71652 16996
rect 72492 16940 72548 16996
rect 72044 16604 72100 16660
rect 70588 15708 70644 15764
rect 70140 15596 70196 15652
rect 70812 15596 70868 15652
rect 70700 15314 70756 15316
rect 70700 15262 70702 15314
rect 70702 15262 70754 15314
rect 70754 15262 70756 15314
rect 70700 15260 70756 15262
rect 70028 14700 70084 14756
rect 69580 13746 69636 13748
rect 69580 13694 69582 13746
rect 69582 13694 69634 13746
rect 69634 13694 69636 13746
rect 69580 13692 69636 13694
rect 69132 13132 69188 13188
rect 68124 11452 68180 11508
rect 68012 10892 68068 10948
rect 67788 10332 67844 10388
rect 67900 10668 67956 10724
rect 67788 9938 67844 9940
rect 67788 9886 67790 9938
rect 67790 9886 67842 9938
rect 67842 9886 67844 9938
rect 67788 9884 67844 9886
rect 67900 9154 67956 9156
rect 67900 9102 67902 9154
rect 67902 9102 67954 9154
rect 67954 9102 67956 9154
rect 67900 9100 67956 9102
rect 68348 11452 68404 11508
rect 68348 10556 68404 10612
rect 68572 10498 68628 10500
rect 68572 10446 68574 10498
rect 68574 10446 68626 10498
rect 68626 10446 68628 10498
rect 68572 10444 68628 10446
rect 68236 8204 68292 8260
rect 67788 7644 67844 7700
rect 67676 6748 67732 6804
rect 67564 6636 67620 6692
rect 68236 6636 68292 6692
rect 67564 5906 67620 5908
rect 67564 5854 67566 5906
rect 67566 5854 67618 5906
rect 67618 5854 67620 5906
rect 67564 5852 67620 5854
rect 68012 6018 68068 6020
rect 68012 5966 68014 6018
rect 68014 5966 68066 6018
rect 68066 5966 68068 6018
rect 68012 5964 68068 5966
rect 67788 5122 67844 5124
rect 67788 5070 67790 5122
rect 67790 5070 67842 5122
rect 67842 5070 67844 5122
rect 67788 5068 67844 5070
rect 67228 4956 67284 5012
rect 67676 5010 67732 5012
rect 67676 4958 67678 5010
rect 67678 4958 67730 5010
rect 67730 4958 67732 5010
rect 67676 4956 67732 4958
rect 68684 8876 68740 8932
rect 68460 8540 68516 8596
rect 68460 6466 68516 6468
rect 68460 6414 68462 6466
rect 68462 6414 68514 6466
rect 68514 6414 68516 6466
rect 68460 6412 68516 6414
rect 68460 6076 68516 6132
rect 68460 5740 68516 5796
rect 68460 5346 68516 5348
rect 68460 5294 68462 5346
rect 68462 5294 68514 5346
rect 68514 5294 68516 5346
rect 68460 5292 68516 5294
rect 71260 15484 71316 15540
rect 70924 15260 70980 15316
rect 71484 15538 71540 15540
rect 71484 15486 71486 15538
rect 71486 15486 71538 15538
rect 71538 15486 71540 15538
rect 71484 15484 71540 15486
rect 72380 15484 72436 15540
rect 69804 13916 69860 13972
rect 70252 13468 70308 13524
rect 69692 12572 69748 12628
rect 69020 11170 69076 11172
rect 69020 11118 69022 11170
rect 69022 11118 69074 11170
rect 69074 11118 69076 11170
rect 69020 11116 69076 11118
rect 69132 9602 69188 9604
rect 69132 9550 69134 9602
rect 69134 9550 69186 9602
rect 69186 9550 69188 9602
rect 69132 9548 69188 9550
rect 70140 12572 70196 12628
rect 70588 13020 70644 13076
rect 70476 12178 70532 12180
rect 70476 12126 70478 12178
rect 70478 12126 70530 12178
rect 70530 12126 70532 12178
rect 70476 12124 70532 12126
rect 70140 11394 70196 11396
rect 70140 11342 70142 11394
rect 70142 11342 70194 11394
rect 70194 11342 70196 11394
rect 70140 11340 70196 11342
rect 70028 11228 70084 11284
rect 69356 10892 69412 10948
rect 69468 11004 69524 11060
rect 70252 11004 70308 11060
rect 69804 10892 69860 10948
rect 70028 10108 70084 10164
rect 69468 9548 69524 9604
rect 69020 8428 69076 8484
rect 68908 8092 68964 8148
rect 69244 8092 69300 8148
rect 69580 8930 69636 8932
rect 69580 8878 69582 8930
rect 69582 8878 69634 8930
rect 69634 8878 69636 8930
rect 69580 8876 69636 8878
rect 69916 6860 69972 6916
rect 70588 9884 70644 9940
rect 70140 9714 70196 9716
rect 70140 9662 70142 9714
rect 70142 9662 70194 9714
rect 70194 9662 70196 9714
rect 70140 9660 70196 9662
rect 70476 9714 70532 9716
rect 70476 9662 70478 9714
rect 70478 9662 70530 9714
rect 70530 9662 70532 9714
rect 70476 9660 70532 9662
rect 70364 8146 70420 8148
rect 70364 8094 70366 8146
rect 70366 8094 70418 8146
rect 70418 8094 70420 8146
rect 70364 8092 70420 8094
rect 70476 7362 70532 7364
rect 70476 7310 70478 7362
rect 70478 7310 70530 7362
rect 70530 7310 70532 7362
rect 70476 7308 70532 7310
rect 68684 5122 68740 5124
rect 68684 5070 68686 5122
rect 68686 5070 68738 5122
rect 68738 5070 68740 5122
rect 68684 5068 68740 5070
rect 69132 5906 69188 5908
rect 69132 5854 69134 5906
rect 69134 5854 69186 5906
rect 69186 5854 69188 5906
rect 69132 5852 69188 5854
rect 69244 5740 69300 5796
rect 69020 5122 69076 5124
rect 69020 5070 69022 5122
rect 69022 5070 69074 5122
rect 69074 5070 69076 5122
rect 69020 5068 69076 5070
rect 68908 4732 68964 4788
rect 69244 4284 69300 4340
rect 68572 3666 68628 3668
rect 68572 3614 68574 3666
rect 68574 3614 68626 3666
rect 68626 3614 68628 3666
rect 68572 3612 68628 3614
rect 69356 5404 69412 5460
rect 69468 5292 69524 5348
rect 69468 4732 69524 4788
rect 69692 3612 69748 3668
rect 69468 3164 69524 3220
rect 70588 6860 70644 6916
rect 71036 13746 71092 13748
rect 71036 13694 71038 13746
rect 71038 13694 71090 13746
rect 71090 13694 71092 13746
rect 71036 13692 71092 13694
rect 71260 13970 71316 13972
rect 71260 13918 71262 13970
rect 71262 13918 71314 13970
rect 71314 13918 71316 13970
rect 71260 13916 71316 13918
rect 71372 13580 71428 13636
rect 72492 15426 72548 15428
rect 72492 15374 72494 15426
rect 72494 15374 72546 15426
rect 72546 15374 72548 15426
rect 72492 15372 72548 15374
rect 72380 14642 72436 14644
rect 72380 14590 72382 14642
rect 72382 14590 72434 14642
rect 72434 14590 72436 14642
rect 72380 14588 72436 14590
rect 74172 20524 74228 20580
rect 74620 22652 74676 22708
rect 75628 24892 75684 24948
rect 75628 23938 75684 23940
rect 75628 23886 75630 23938
rect 75630 23886 75682 23938
rect 75682 23886 75684 23938
rect 75628 23884 75684 23886
rect 77644 27580 77700 27636
rect 77308 27020 77364 27076
rect 76860 26178 76916 26180
rect 76860 26126 76862 26178
rect 76862 26126 76914 26178
rect 76914 26126 76916 26178
rect 76860 26124 76916 26126
rect 78540 27132 78596 27188
rect 78876 27020 78932 27076
rect 76524 25004 76580 25060
rect 76076 23884 76132 23940
rect 75628 23100 75684 23156
rect 76860 24668 76916 24724
rect 76524 23100 76580 23156
rect 76188 23042 76244 23044
rect 76188 22990 76190 23042
rect 76190 22990 76242 23042
rect 76242 22990 76244 23042
rect 76188 22988 76244 22990
rect 75740 22652 75796 22708
rect 75628 22482 75684 22484
rect 75628 22430 75630 22482
rect 75630 22430 75682 22482
rect 75682 22430 75684 22482
rect 75628 22428 75684 22430
rect 74508 22146 74564 22148
rect 74508 22094 74510 22146
rect 74510 22094 74562 22146
rect 74562 22094 74564 22146
rect 74508 22092 74564 22094
rect 74396 20300 74452 20356
rect 74172 19794 74228 19796
rect 74172 19742 74174 19794
rect 74174 19742 74226 19794
rect 74226 19742 74228 19794
rect 74172 19740 74228 19742
rect 73724 19068 73780 19124
rect 72940 18060 72996 18116
rect 73724 18396 73780 18452
rect 73276 18172 73332 18228
rect 73724 17442 73780 17444
rect 73724 17390 73726 17442
rect 73726 17390 73778 17442
rect 73778 17390 73780 17442
rect 73724 17388 73780 17390
rect 74732 21644 74788 21700
rect 74956 21644 75012 21700
rect 74732 20524 74788 20580
rect 75180 20578 75236 20580
rect 75180 20526 75182 20578
rect 75182 20526 75234 20578
rect 75234 20526 75236 20578
rect 75180 20524 75236 20526
rect 74844 20188 74900 20244
rect 74620 20130 74676 20132
rect 74620 20078 74622 20130
rect 74622 20078 74674 20130
rect 74674 20078 74676 20130
rect 74620 20076 74676 20078
rect 76300 22204 76356 22260
rect 76412 22428 76468 22484
rect 76412 21756 76468 21812
rect 75404 21532 75460 21588
rect 75404 20636 75460 20692
rect 75516 21196 75572 21252
rect 74396 19068 74452 19124
rect 73612 16716 73668 16772
rect 73276 16604 73332 16660
rect 73052 15986 73108 15988
rect 73052 15934 73054 15986
rect 73054 15934 73106 15986
rect 73106 15934 73108 15986
rect 73052 15932 73108 15934
rect 72940 15708 72996 15764
rect 74284 17388 74340 17444
rect 74172 17276 74228 17332
rect 74172 15932 74228 15988
rect 73836 15708 73892 15764
rect 73052 15372 73108 15428
rect 74284 15426 74340 15428
rect 74284 15374 74286 15426
rect 74286 15374 74338 15426
rect 74338 15374 74340 15426
rect 74284 15372 74340 15374
rect 72492 14530 72548 14532
rect 72492 14478 72494 14530
rect 72494 14478 72546 14530
rect 72546 14478 72548 14530
rect 72492 14476 72548 14478
rect 71820 13916 71876 13972
rect 72492 13580 72548 13636
rect 72380 13522 72436 13524
rect 72380 13470 72382 13522
rect 72382 13470 72434 13522
rect 72434 13470 72436 13522
rect 72380 13468 72436 13470
rect 72940 13804 72996 13860
rect 72716 12124 72772 12180
rect 72828 12460 72884 12516
rect 71036 11564 71092 11620
rect 70924 11116 70980 11172
rect 71596 11394 71652 11396
rect 71596 11342 71598 11394
rect 71598 11342 71650 11394
rect 71650 11342 71652 11394
rect 71596 11340 71652 11342
rect 71484 11170 71540 11172
rect 71484 11118 71486 11170
rect 71486 11118 71538 11170
rect 71538 11118 71540 11170
rect 71484 11116 71540 11118
rect 71708 11116 71764 11172
rect 71932 11900 71988 11956
rect 71372 11004 71428 11060
rect 71372 10668 71428 10724
rect 72156 11340 72212 11396
rect 71932 11116 71988 11172
rect 71932 10892 71988 10948
rect 70924 9714 70980 9716
rect 70924 9662 70926 9714
rect 70926 9662 70978 9714
rect 70978 9662 70980 9714
rect 70924 9660 70980 9662
rect 71260 9548 71316 9604
rect 71148 9436 71204 9492
rect 71708 9436 71764 9492
rect 71260 9212 71316 9268
rect 71708 9266 71764 9268
rect 71708 9214 71710 9266
rect 71710 9214 71762 9266
rect 71762 9214 71764 9266
rect 71708 9212 71764 9214
rect 75292 19122 75348 19124
rect 75292 19070 75294 19122
rect 75294 19070 75346 19122
rect 75346 19070 75348 19122
rect 75292 19068 75348 19070
rect 77756 26124 77812 26180
rect 78428 24946 78484 24948
rect 78428 24894 78430 24946
rect 78430 24894 78482 24946
rect 78482 24894 78484 24946
rect 78428 24892 78484 24894
rect 78204 24722 78260 24724
rect 78204 24670 78206 24722
rect 78206 24670 78258 24722
rect 78258 24670 78260 24722
rect 78204 24668 78260 24670
rect 77532 23100 77588 23156
rect 77420 21532 77476 21588
rect 77084 20802 77140 20804
rect 77084 20750 77086 20802
rect 77086 20750 77138 20802
rect 77138 20750 77140 20802
rect 77084 20748 77140 20750
rect 78316 23212 78372 23268
rect 78428 23154 78484 23156
rect 78428 23102 78430 23154
rect 78430 23102 78482 23154
rect 78482 23102 78484 23154
rect 78428 23100 78484 23102
rect 77868 22092 77924 22148
rect 77756 20860 77812 20916
rect 74844 19010 74900 19012
rect 74844 18958 74846 19010
rect 74846 18958 74898 19010
rect 74898 18958 74900 19010
rect 74844 18956 74900 18958
rect 75068 19010 75124 19012
rect 75068 18958 75070 19010
rect 75070 18958 75122 19010
rect 75122 18958 75124 19010
rect 75068 18956 75124 18958
rect 74956 18172 75012 18228
rect 75292 16268 75348 16324
rect 74956 15932 75012 15988
rect 75180 15874 75236 15876
rect 75180 15822 75182 15874
rect 75182 15822 75234 15874
rect 75234 15822 75236 15874
rect 75180 15820 75236 15822
rect 81276 26682 81332 26684
rect 81276 26630 81278 26682
rect 81278 26630 81330 26682
rect 81330 26630 81332 26682
rect 81276 26628 81332 26630
rect 81380 26682 81436 26684
rect 81380 26630 81382 26682
rect 81382 26630 81434 26682
rect 81434 26630 81436 26682
rect 81380 26628 81436 26630
rect 81484 26682 81540 26684
rect 81484 26630 81486 26682
rect 81486 26630 81538 26682
rect 81538 26630 81540 26682
rect 81484 26628 81540 26630
rect 79660 25228 79716 25284
rect 79100 24892 79156 24948
rect 78540 21420 78596 21476
rect 77868 20412 77924 20468
rect 78092 20524 78148 20580
rect 76524 19964 76580 20020
rect 75740 18396 75796 18452
rect 75516 17052 75572 17108
rect 74620 15148 74676 15204
rect 73276 14252 73332 14308
rect 73724 13244 73780 13300
rect 72380 11228 72436 11284
rect 71932 8428 71988 8484
rect 71036 7980 71092 8036
rect 71148 7308 71204 7364
rect 71260 7420 71316 7476
rect 70700 6300 70756 6356
rect 70700 5180 70756 5236
rect 71148 6860 71204 6916
rect 71148 5010 71204 5012
rect 71148 4958 71150 5010
rect 71150 4958 71202 5010
rect 71202 4958 71204 5010
rect 71148 4956 71204 4958
rect 70476 3666 70532 3668
rect 70476 3614 70478 3666
rect 70478 3614 70530 3666
rect 70530 3614 70532 3666
rect 70476 3612 70532 3614
rect 70700 2828 70756 2884
rect 71036 4732 71092 4788
rect 70252 2380 70308 2436
rect 71708 6636 71764 6692
rect 72156 9602 72212 9604
rect 72156 9550 72158 9602
rect 72158 9550 72210 9602
rect 72210 9550 72212 9602
rect 72156 9548 72212 9550
rect 72716 11116 72772 11172
rect 72828 11004 72884 11060
rect 72492 10610 72548 10612
rect 72492 10558 72494 10610
rect 72494 10558 72546 10610
rect 72546 10558 72548 10610
rect 72492 10556 72548 10558
rect 72716 10444 72772 10500
rect 72268 8540 72324 8596
rect 72492 9436 72548 9492
rect 72716 9602 72772 9604
rect 72716 9550 72718 9602
rect 72718 9550 72770 9602
rect 72770 9550 72772 9602
rect 72716 9548 72772 9550
rect 72604 9212 72660 9268
rect 72716 9324 72772 9380
rect 73052 11394 73108 11396
rect 73052 11342 73054 11394
rect 73054 11342 73106 11394
rect 73106 11342 73108 11394
rect 73052 11340 73108 11342
rect 73388 11788 73444 11844
rect 73724 12460 73780 12516
rect 73500 11564 73556 11620
rect 74732 15036 74788 15092
rect 74284 14924 74340 14980
rect 74284 14476 74340 14532
rect 74284 14306 74340 14308
rect 74284 14254 74286 14306
rect 74286 14254 74338 14306
rect 74338 14254 74340 14306
rect 74284 14252 74340 14254
rect 74956 15260 75012 15316
rect 74844 14306 74900 14308
rect 74844 14254 74846 14306
rect 74846 14254 74898 14306
rect 74898 14254 74900 14306
rect 74844 14252 74900 14254
rect 74396 13468 74452 13524
rect 74732 13804 74788 13860
rect 74172 13074 74228 13076
rect 74172 13022 74174 13074
rect 74174 13022 74226 13074
rect 74226 13022 74228 13074
rect 74172 13020 74228 13022
rect 73948 12684 74004 12740
rect 73164 10108 73220 10164
rect 72940 9996 72996 10052
rect 73724 11228 73780 11284
rect 73612 10444 73668 10500
rect 73724 9826 73780 9828
rect 73724 9774 73726 9826
rect 73726 9774 73778 9826
rect 73778 9774 73780 9826
rect 73724 9772 73780 9774
rect 73276 9714 73332 9716
rect 73276 9662 73278 9714
rect 73278 9662 73330 9714
rect 73330 9662 73332 9714
rect 73276 9660 73332 9662
rect 72828 8652 72884 8708
rect 72940 8988 72996 9044
rect 72156 7644 72212 7700
rect 72268 7586 72324 7588
rect 72268 7534 72270 7586
rect 72270 7534 72322 7586
rect 72322 7534 72324 7586
rect 72268 7532 72324 7534
rect 72380 7420 72436 7476
rect 72492 8204 72548 8260
rect 72044 7196 72100 7252
rect 74060 9324 74116 9380
rect 74508 12796 74564 12852
rect 74508 12178 74564 12180
rect 74508 12126 74510 12178
rect 74510 12126 74562 12178
rect 74562 12126 74564 12178
rect 74508 12124 74564 12126
rect 73948 9212 74004 9268
rect 73052 8540 73108 8596
rect 73164 8316 73220 8372
rect 73612 8988 73668 9044
rect 73500 8316 73556 8372
rect 73612 8652 73668 8708
rect 72492 6748 72548 6804
rect 72604 7196 72660 7252
rect 72268 6524 72324 6580
rect 72044 6300 72100 6356
rect 71596 5122 71652 5124
rect 71596 5070 71598 5122
rect 71598 5070 71650 5122
rect 71650 5070 71652 5122
rect 71596 5068 71652 5070
rect 72044 5628 72100 5684
rect 72268 6300 72324 6356
rect 72268 5068 72324 5124
rect 72380 5852 72436 5908
rect 72604 5292 72660 5348
rect 72828 7420 72884 7476
rect 72828 7084 72884 7140
rect 72828 6578 72884 6580
rect 72828 6526 72830 6578
rect 72830 6526 72882 6578
rect 72882 6526 72884 6578
rect 72828 6524 72884 6526
rect 72940 5964 72996 6020
rect 73052 5292 73108 5348
rect 73164 7084 73220 7140
rect 72716 4956 72772 5012
rect 72828 4172 72884 4228
rect 73388 6748 73444 6804
rect 73164 4338 73220 4340
rect 73164 4286 73166 4338
rect 73166 4286 73218 4338
rect 73218 4286 73220 4338
rect 73164 4284 73220 4286
rect 73388 6018 73444 6020
rect 73388 5966 73390 6018
rect 73390 5966 73442 6018
rect 73442 5966 73444 6018
rect 73388 5964 73444 5966
rect 73612 7196 73668 7252
rect 74060 7532 74116 7588
rect 73948 7474 74004 7476
rect 73948 7422 73950 7474
rect 73950 7422 74002 7474
rect 74002 7422 74004 7474
rect 73948 7420 74004 7422
rect 73724 6524 73780 6580
rect 74172 6524 74228 6580
rect 73500 5180 73556 5236
rect 74172 5234 74228 5236
rect 74172 5182 74174 5234
rect 74174 5182 74226 5234
rect 74226 5182 74228 5234
rect 74172 5180 74228 5182
rect 74396 11394 74452 11396
rect 74396 11342 74398 11394
rect 74398 11342 74450 11394
rect 74450 11342 74452 11394
rect 74396 11340 74452 11342
rect 74508 9324 74564 9380
rect 74508 8428 74564 8484
rect 74620 8988 74676 9044
rect 74284 4620 74340 4676
rect 75740 17106 75796 17108
rect 75740 17054 75742 17106
rect 75742 17054 75794 17106
rect 75794 17054 75796 17106
rect 75740 17052 75796 17054
rect 75852 19740 75908 19796
rect 75628 15986 75684 15988
rect 75628 15934 75630 15986
rect 75630 15934 75682 15986
rect 75682 15934 75684 15986
rect 75628 15932 75684 15934
rect 75292 14588 75348 14644
rect 75068 13580 75124 13636
rect 74844 12684 74900 12740
rect 74844 11394 74900 11396
rect 74844 11342 74846 11394
rect 74846 11342 74898 11394
rect 74898 11342 74900 11394
rect 74844 11340 74900 11342
rect 74844 9884 74900 9940
rect 75628 14252 75684 14308
rect 75404 13692 75460 13748
rect 75516 13858 75572 13860
rect 75516 13806 75518 13858
rect 75518 13806 75570 13858
rect 75570 13806 75572 13858
rect 75516 13804 75572 13806
rect 75292 12738 75348 12740
rect 75292 12686 75294 12738
rect 75294 12686 75346 12738
rect 75346 12686 75348 12738
rect 75292 12684 75348 12686
rect 75292 11564 75348 11620
rect 74956 9772 75012 9828
rect 77196 20076 77252 20132
rect 76748 19906 76804 19908
rect 76748 19854 76750 19906
rect 76750 19854 76802 19906
rect 76802 19854 76804 19906
rect 76748 19852 76804 19854
rect 77756 20076 77812 20132
rect 76188 18956 76244 19012
rect 77644 19964 77700 20020
rect 78540 20524 78596 20580
rect 78316 20412 78372 20468
rect 78988 23212 79044 23268
rect 78876 22764 78932 22820
rect 80444 24892 80500 24948
rect 80668 25228 80724 25284
rect 81276 25114 81332 25116
rect 80220 23266 80276 23268
rect 80220 23214 80222 23266
rect 80222 23214 80274 23266
rect 80274 23214 80276 23266
rect 80220 23212 80276 23214
rect 79548 22764 79604 22820
rect 79324 22316 79380 22372
rect 78764 20748 78820 20804
rect 78652 20076 78708 20132
rect 76636 18172 76692 18228
rect 76300 16770 76356 16772
rect 76300 16718 76302 16770
rect 76302 16718 76354 16770
rect 76354 16718 76356 16770
rect 76300 16716 76356 16718
rect 76188 16492 76244 16548
rect 76860 18284 76916 18340
rect 77420 18060 77476 18116
rect 77196 17778 77252 17780
rect 77196 17726 77198 17778
rect 77198 17726 77250 17778
rect 77250 17726 77252 17778
rect 77196 17724 77252 17726
rect 77420 17276 77476 17332
rect 76636 16828 76692 16884
rect 76860 16882 76916 16884
rect 76860 16830 76862 16882
rect 76862 16830 76914 16882
rect 76914 16830 76916 16882
rect 76860 16828 76916 16830
rect 77644 16828 77700 16884
rect 77420 16492 77476 16548
rect 76412 16268 76468 16324
rect 77308 16268 77364 16324
rect 75852 15820 75908 15876
rect 76412 15932 76468 15988
rect 76300 15874 76356 15876
rect 76300 15822 76302 15874
rect 76302 15822 76354 15874
rect 76354 15822 76356 15874
rect 76300 15820 76356 15822
rect 76748 15820 76804 15876
rect 76636 15708 76692 15764
rect 75740 11116 75796 11172
rect 75852 12236 75908 12292
rect 75852 11004 75908 11060
rect 75068 9602 75124 9604
rect 75068 9550 75070 9602
rect 75070 9550 75122 9602
rect 75122 9550 75124 9602
rect 75068 9548 75124 9550
rect 76412 13746 76468 13748
rect 76412 13694 76414 13746
rect 76414 13694 76466 13746
rect 76466 13694 76468 13746
rect 76412 13692 76468 13694
rect 76076 11394 76132 11396
rect 76076 11342 76078 11394
rect 76078 11342 76130 11394
rect 76130 11342 76132 11394
rect 76076 11340 76132 11342
rect 76412 11788 76468 11844
rect 76300 11340 76356 11396
rect 76188 11116 76244 11172
rect 76524 11340 76580 11396
rect 76412 10332 76468 10388
rect 76972 15874 77028 15876
rect 76972 15822 76974 15874
rect 76974 15822 77026 15874
rect 77026 15822 77028 15874
rect 76972 15820 77028 15822
rect 77196 15148 77252 15204
rect 77644 16268 77700 16324
rect 77420 15820 77476 15876
rect 77084 13580 77140 13636
rect 77196 12236 77252 12292
rect 77420 12236 77476 12292
rect 77196 11564 77252 11620
rect 76972 11394 77028 11396
rect 76972 11342 76974 11394
rect 76974 11342 77026 11394
rect 77026 11342 77028 11394
rect 76972 11340 77028 11342
rect 76972 11116 77028 11172
rect 76748 11004 76804 11060
rect 76972 10834 77028 10836
rect 76972 10782 76974 10834
rect 76974 10782 77026 10834
rect 77026 10782 77028 10834
rect 76972 10780 77028 10782
rect 75964 9324 76020 9380
rect 75740 8316 75796 8372
rect 75404 8258 75460 8260
rect 75404 8206 75406 8258
rect 75406 8206 75458 8258
rect 75458 8206 75460 8258
rect 75404 8204 75460 8206
rect 75404 7980 75460 8036
rect 75516 7308 75572 7364
rect 75964 7644 76020 7700
rect 75292 5964 75348 6020
rect 75740 5068 75796 5124
rect 75516 4508 75572 4564
rect 76076 6860 76132 6916
rect 76188 5068 76244 5124
rect 76300 7196 76356 7252
rect 76412 6690 76468 6692
rect 76412 6638 76414 6690
rect 76414 6638 76466 6690
rect 76466 6638 76468 6690
rect 76412 6636 76468 6638
rect 76412 6412 76468 6468
rect 76636 8930 76692 8932
rect 76636 8878 76638 8930
rect 76638 8878 76690 8930
rect 76690 8878 76692 8930
rect 76636 8876 76692 8878
rect 77084 8764 77140 8820
rect 76972 8092 77028 8148
rect 76748 7362 76804 7364
rect 76748 7310 76750 7362
rect 76750 7310 76802 7362
rect 76802 7310 76804 7362
rect 76748 7308 76804 7310
rect 77532 10444 77588 10500
rect 77420 9324 77476 9380
rect 77532 9042 77588 9044
rect 77532 8990 77534 9042
rect 77534 8990 77586 9042
rect 77586 8990 77588 9042
rect 77532 8988 77588 8990
rect 77532 8316 77588 8372
rect 77196 7308 77252 7364
rect 77308 7532 77364 7588
rect 77308 6860 77364 6916
rect 77196 6636 77252 6692
rect 76972 6018 77028 6020
rect 76972 5966 76974 6018
rect 76974 5966 77026 6018
rect 77026 5966 77028 6018
rect 76972 5964 77028 5966
rect 77084 5292 77140 5348
rect 76524 4956 76580 5012
rect 76412 4898 76468 4900
rect 76412 4846 76414 4898
rect 76414 4846 76466 4898
rect 76466 4846 76468 4898
rect 76412 4844 76468 4846
rect 76412 4620 76468 4676
rect 74284 2492 74340 2548
rect 76076 3442 76132 3444
rect 76076 3390 76078 3442
rect 76078 3390 76130 3442
rect 76130 3390 76132 3442
rect 76076 3388 76132 3390
rect 75628 2380 75684 2436
rect 76972 4562 77028 4564
rect 76972 4510 76974 4562
rect 76974 4510 77026 4562
rect 77026 4510 77028 4562
rect 76972 4508 77028 4510
rect 76524 4284 76580 4340
rect 77196 4284 77252 4340
rect 77196 4060 77252 4116
rect 76972 3500 77028 3556
rect 77980 16210 78036 16212
rect 77980 16158 77982 16210
rect 77982 16158 78034 16210
rect 78034 16158 78036 16210
rect 77980 16156 78036 16158
rect 77980 15820 78036 15876
rect 77980 15202 78036 15204
rect 77980 15150 77982 15202
rect 77982 15150 78034 15202
rect 78034 15150 78036 15202
rect 77980 15148 78036 15150
rect 78428 16268 78484 16324
rect 78540 15484 78596 15540
rect 77868 13916 77924 13972
rect 78652 14924 78708 14980
rect 78428 13916 78484 13972
rect 78204 13468 78260 13524
rect 77868 11004 77924 11060
rect 77868 9436 77924 9492
rect 77868 9100 77924 9156
rect 78092 12684 78148 12740
rect 78540 12796 78596 12852
rect 78540 12236 78596 12292
rect 78204 11340 78260 11396
rect 78204 10834 78260 10836
rect 78204 10782 78206 10834
rect 78206 10782 78258 10834
rect 78258 10782 78260 10834
rect 78204 10780 78260 10782
rect 78204 10332 78260 10388
rect 78764 12124 78820 12180
rect 78316 8930 78372 8932
rect 78316 8878 78318 8930
rect 78318 8878 78370 8930
rect 78370 8878 78372 8930
rect 78316 8876 78372 8878
rect 78204 8540 78260 8596
rect 79548 21474 79604 21476
rect 79548 21422 79550 21474
rect 79550 21422 79602 21474
rect 79602 21422 79604 21474
rect 79548 21420 79604 21422
rect 79324 20914 79380 20916
rect 79324 20862 79326 20914
rect 79326 20862 79378 20914
rect 79378 20862 79380 20914
rect 79324 20860 79380 20862
rect 78988 18396 79044 18452
rect 79212 17948 79268 18004
rect 79212 17106 79268 17108
rect 79212 17054 79214 17106
rect 79214 17054 79266 17106
rect 79266 17054 79268 17106
rect 79212 17052 79268 17054
rect 79548 18172 79604 18228
rect 79772 17612 79828 17668
rect 80668 23660 80724 23716
rect 80780 25004 80836 25060
rect 81276 25062 81278 25114
rect 81278 25062 81330 25114
rect 81330 25062 81332 25114
rect 81276 25060 81332 25062
rect 81380 25114 81436 25116
rect 81380 25062 81382 25114
rect 81382 25062 81434 25114
rect 81434 25062 81436 25114
rect 81380 25060 81436 25062
rect 81484 25114 81540 25116
rect 81484 25062 81486 25114
rect 81486 25062 81538 25114
rect 81538 25062 81540 25114
rect 81484 25060 81540 25062
rect 81116 24834 81172 24836
rect 81116 24782 81118 24834
rect 81118 24782 81170 24834
rect 81170 24782 81172 24834
rect 81116 24780 81172 24782
rect 81900 24780 81956 24836
rect 81276 23546 81332 23548
rect 81276 23494 81278 23546
rect 81278 23494 81330 23546
rect 81330 23494 81332 23546
rect 81276 23492 81332 23494
rect 81380 23546 81436 23548
rect 81380 23494 81382 23546
rect 81382 23494 81434 23546
rect 81434 23494 81436 23546
rect 81380 23492 81436 23494
rect 81484 23546 81540 23548
rect 81484 23494 81486 23546
rect 81486 23494 81538 23546
rect 81538 23494 81540 23546
rect 81484 23492 81540 23494
rect 81564 23212 81620 23268
rect 82796 24668 82852 24724
rect 80892 22988 80948 23044
rect 80220 21810 80276 21812
rect 80220 21758 80222 21810
rect 80222 21758 80274 21810
rect 80274 21758 80276 21810
rect 80220 21756 80276 21758
rect 80444 21756 80500 21812
rect 81676 22876 81732 22932
rect 82124 22876 82180 22932
rect 81276 21978 81332 21980
rect 81276 21926 81278 21978
rect 81278 21926 81330 21978
rect 81330 21926 81332 21978
rect 81276 21924 81332 21926
rect 81380 21978 81436 21980
rect 81380 21926 81382 21978
rect 81382 21926 81434 21978
rect 81434 21926 81436 21978
rect 81380 21924 81436 21926
rect 81484 21978 81540 21980
rect 81484 21926 81486 21978
rect 81486 21926 81538 21978
rect 81538 21926 81540 21978
rect 81484 21924 81540 21926
rect 81676 21868 81732 21924
rect 81452 21756 81508 21812
rect 81116 20748 81172 20804
rect 81564 20748 81620 20804
rect 80556 20524 80612 20580
rect 79996 17666 80052 17668
rect 79996 17614 79998 17666
rect 79998 17614 80050 17666
rect 80050 17614 80052 17666
rect 79996 17612 80052 17614
rect 80444 17612 80500 17668
rect 80108 17106 80164 17108
rect 80108 17054 80110 17106
rect 80110 17054 80162 17106
rect 80162 17054 80164 17106
rect 80108 17052 80164 17054
rect 79548 16044 79604 16100
rect 79996 16940 80052 16996
rect 79100 15372 79156 15428
rect 79772 15708 79828 15764
rect 79884 16044 79940 16100
rect 79548 15538 79604 15540
rect 79548 15486 79550 15538
rect 79550 15486 79602 15538
rect 79602 15486 79604 15538
rect 79548 15484 79604 15486
rect 81564 20578 81620 20580
rect 81564 20526 81566 20578
rect 81566 20526 81618 20578
rect 81618 20526 81620 20578
rect 81564 20524 81620 20526
rect 81276 20410 81332 20412
rect 81276 20358 81278 20410
rect 81278 20358 81330 20410
rect 81330 20358 81332 20410
rect 81276 20356 81332 20358
rect 81380 20410 81436 20412
rect 81380 20358 81382 20410
rect 81382 20358 81434 20410
rect 81434 20358 81436 20410
rect 81380 20356 81436 20358
rect 81484 20410 81540 20412
rect 81484 20358 81486 20410
rect 81486 20358 81538 20410
rect 81538 20358 81540 20410
rect 81484 20356 81540 20358
rect 80892 20018 80948 20020
rect 80892 19966 80894 20018
rect 80894 19966 80946 20018
rect 80946 19966 80948 20018
rect 80892 19964 80948 19966
rect 80780 17666 80836 17668
rect 80780 17614 80782 17666
rect 80782 17614 80834 17666
rect 80834 17614 80836 17666
rect 80780 17612 80836 17614
rect 81228 19628 81284 19684
rect 81564 19740 81620 19796
rect 82236 23100 82292 23156
rect 82012 21810 82068 21812
rect 82012 21758 82014 21810
rect 82014 21758 82066 21810
rect 82066 21758 82068 21810
rect 82012 21756 82068 21758
rect 82460 22876 82516 22932
rect 82684 22988 82740 23044
rect 82684 21868 82740 21924
rect 88060 28700 88116 28756
rect 86156 26178 86212 26180
rect 86156 26126 86158 26178
rect 86158 26126 86210 26178
rect 86210 26126 86212 26178
rect 86156 26124 86212 26126
rect 86604 26178 86660 26180
rect 86604 26126 86606 26178
rect 86606 26126 86658 26178
rect 86658 26126 86660 26178
rect 86604 26124 86660 26126
rect 86940 26012 86996 26068
rect 83804 24722 83860 24724
rect 83804 24670 83806 24722
rect 83806 24670 83858 24722
rect 83858 24670 83860 24722
rect 83804 24668 83860 24670
rect 83356 23660 83412 23716
rect 84364 23660 84420 23716
rect 84588 23884 84644 23940
rect 86828 23772 86884 23828
rect 84588 23660 84644 23716
rect 83356 22988 83412 23044
rect 83580 23154 83636 23156
rect 83580 23102 83582 23154
rect 83582 23102 83634 23154
rect 83634 23102 83636 23154
rect 83580 23100 83636 23102
rect 83468 22428 83524 22484
rect 84476 23042 84532 23044
rect 84476 22990 84478 23042
rect 84478 22990 84530 23042
rect 84530 22990 84532 23042
rect 84476 22988 84532 22990
rect 86156 22988 86212 23044
rect 84028 22876 84084 22932
rect 81788 20130 81844 20132
rect 81788 20078 81790 20130
rect 81790 20078 81842 20130
rect 81842 20078 81844 20130
rect 81788 20076 81844 20078
rect 82236 20130 82292 20132
rect 82236 20078 82238 20130
rect 82238 20078 82290 20130
rect 82290 20078 82292 20130
rect 82236 20076 82292 20078
rect 81676 19628 81732 19684
rect 82012 19740 82068 19796
rect 82236 19628 82292 19684
rect 81276 18842 81332 18844
rect 81276 18790 81278 18842
rect 81278 18790 81330 18842
rect 81330 18790 81332 18842
rect 81276 18788 81332 18790
rect 81380 18842 81436 18844
rect 81380 18790 81382 18842
rect 81382 18790 81434 18842
rect 81434 18790 81436 18842
rect 81380 18788 81436 18790
rect 81484 18842 81540 18844
rect 81484 18790 81486 18842
rect 81486 18790 81538 18842
rect 81538 18790 81540 18842
rect 81484 18788 81540 18790
rect 81276 17274 81332 17276
rect 81276 17222 81278 17274
rect 81278 17222 81330 17274
rect 81330 17222 81332 17274
rect 81276 17220 81332 17222
rect 81380 17274 81436 17276
rect 81380 17222 81382 17274
rect 81382 17222 81434 17274
rect 81434 17222 81436 17274
rect 81380 17220 81436 17222
rect 81484 17274 81540 17276
rect 81484 17222 81486 17274
rect 81486 17222 81538 17274
rect 81538 17222 81540 17274
rect 81484 17220 81540 17222
rect 80892 16940 80948 16996
rect 81116 16994 81172 16996
rect 81116 16942 81118 16994
rect 81118 16942 81170 16994
rect 81170 16942 81172 16994
rect 81116 16940 81172 16942
rect 80108 15932 80164 15988
rect 82012 18172 82068 18228
rect 81900 17164 81956 17220
rect 80108 15484 80164 15540
rect 79100 14140 79156 14196
rect 79324 13634 79380 13636
rect 79324 13582 79326 13634
rect 79326 13582 79378 13634
rect 79378 13582 79380 13634
rect 79324 13580 79380 13582
rect 79100 13468 79156 13524
rect 79660 12572 79716 12628
rect 78988 11282 79044 11284
rect 78988 11230 78990 11282
rect 78990 11230 79042 11282
rect 79042 11230 79044 11282
rect 78988 11228 79044 11230
rect 78988 10780 79044 10836
rect 79100 11116 79156 11172
rect 78540 8316 78596 8372
rect 78092 7980 78148 8036
rect 77980 7532 78036 7588
rect 77644 6300 77700 6356
rect 77644 5292 77700 5348
rect 77644 3388 77700 3444
rect 77756 3612 77812 3668
rect 78428 6076 78484 6132
rect 78316 5964 78372 6020
rect 79212 8316 79268 8372
rect 78988 7532 79044 7588
rect 78652 5852 78708 5908
rect 79436 12290 79492 12292
rect 79436 12238 79438 12290
rect 79438 12238 79490 12290
rect 79490 12238 79492 12290
rect 79436 12236 79492 12238
rect 79660 12236 79716 12292
rect 79548 11788 79604 11844
rect 81340 16380 81396 16436
rect 80780 16098 80836 16100
rect 80780 16046 80782 16098
rect 80782 16046 80834 16098
rect 80834 16046 80836 16098
rect 80780 16044 80836 16046
rect 81276 15706 81332 15708
rect 81276 15654 81278 15706
rect 81278 15654 81330 15706
rect 81330 15654 81332 15706
rect 81276 15652 81332 15654
rect 81380 15706 81436 15708
rect 81380 15654 81382 15706
rect 81382 15654 81434 15706
rect 81434 15654 81436 15706
rect 81380 15652 81436 15654
rect 81484 15706 81540 15708
rect 81484 15654 81486 15706
rect 81486 15654 81538 15706
rect 81538 15654 81540 15706
rect 81484 15652 81540 15654
rect 81676 15596 81732 15652
rect 80444 14700 80500 14756
rect 80556 14812 80612 14868
rect 80332 14588 80388 14644
rect 81452 14754 81508 14756
rect 81452 14702 81454 14754
rect 81454 14702 81506 14754
rect 81506 14702 81508 14754
rect 81452 14700 81508 14702
rect 81228 14476 81284 14532
rect 80332 14364 80388 14420
rect 81116 14252 81172 14308
rect 81564 14418 81620 14420
rect 81564 14366 81566 14418
rect 81566 14366 81618 14418
rect 81618 14366 81620 14418
rect 81564 14364 81620 14366
rect 81276 14138 81332 14140
rect 81276 14086 81278 14138
rect 81278 14086 81330 14138
rect 81330 14086 81332 14138
rect 81276 14084 81332 14086
rect 81380 14138 81436 14140
rect 81380 14086 81382 14138
rect 81382 14086 81434 14138
rect 81434 14086 81436 14138
rect 81380 14084 81436 14086
rect 81484 14138 81540 14140
rect 81484 14086 81486 14138
rect 81486 14086 81538 14138
rect 81538 14086 81540 14138
rect 81484 14084 81540 14086
rect 80332 13692 80388 13748
rect 79884 13020 79940 13076
rect 80220 12684 80276 12740
rect 80108 12178 80164 12180
rect 80108 12126 80110 12178
rect 80110 12126 80162 12178
rect 80162 12126 80164 12178
rect 80108 12124 80164 12126
rect 79772 11116 79828 11172
rect 79660 10668 79716 10724
rect 79436 9884 79492 9940
rect 79996 9660 80052 9716
rect 79772 9324 79828 9380
rect 79436 8428 79492 8484
rect 80780 12124 80836 12180
rect 81116 13468 81172 13524
rect 81564 13020 81620 13076
rect 81276 12570 81332 12572
rect 81276 12518 81278 12570
rect 81278 12518 81330 12570
rect 81330 12518 81332 12570
rect 81276 12516 81332 12518
rect 81380 12570 81436 12572
rect 81380 12518 81382 12570
rect 81382 12518 81434 12570
rect 81434 12518 81436 12570
rect 81380 12516 81436 12518
rect 81484 12570 81540 12572
rect 81484 12518 81486 12570
rect 81486 12518 81538 12570
rect 81538 12518 81540 12570
rect 81484 12516 81540 12518
rect 81564 12012 81620 12068
rect 82124 17612 82180 17668
rect 82572 19964 82628 20020
rect 82348 18396 82404 18452
rect 83244 17164 83300 17220
rect 82684 16994 82740 16996
rect 82684 16942 82686 16994
rect 82686 16942 82738 16994
rect 82738 16942 82740 16994
rect 82684 16940 82740 16942
rect 82796 16828 82852 16884
rect 82124 16380 82180 16436
rect 82572 15596 82628 15652
rect 81788 14588 81844 14644
rect 81900 14306 81956 14308
rect 81900 14254 81902 14306
rect 81902 14254 81954 14306
rect 81954 14254 81956 14306
rect 81900 14252 81956 14254
rect 81900 13468 81956 13524
rect 81564 11228 81620 11284
rect 80444 11116 80500 11172
rect 80444 10892 80500 10948
rect 81276 11002 81332 11004
rect 81276 10950 81278 11002
rect 81278 10950 81330 11002
rect 81330 10950 81332 11002
rect 81276 10948 81332 10950
rect 81380 11002 81436 11004
rect 81380 10950 81382 11002
rect 81382 10950 81434 11002
rect 81434 10950 81436 11002
rect 81380 10948 81436 10950
rect 81484 11002 81540 11004
rect 81484 10950 81486 11002
rect 81486 10950 81538 11002
rect 81538 10950 81540 11002
rect 81484 10948 81540 10950
rect 81452 10780 81508 10836
rect 81228 10556 81284 10612
rect 81004 10108 81060 10164
rect 80668 9938 80724 9940
rect 80668 9886 80670 9938
rect 80670 9886 80722 9938
rect 80722 9886 80724 9938
rect 80668 9884 80724 9886
rect 80332 9772 80388 9828
rect 80108 9324 80164 9380
rect 79772 7532 79828 7588
rect 79436 7084 79492 7140
rect 80668 7308 80724 7364
rect 80108 6524 80164 6580
rect 79436 6130 79492 6132
rect 79436 6078 79438 6130
rect 79438 6078 79490 6130
rect 79490 6078 79492 6130
rect 79436 6076 79492 6078
rect 79100 4620 79156 4676
rect 77980 3724 78036 3780
rect 79100 4060 79156 4116
rect 78988 3666 79044 3668
rect 78988 3614 78990 3666
rect 78990 3614 79042 3666
rect 79042 3614 79044 3666
rect 78988 3612 79044 3614
rect 79772 4172 79828 4228
rect 80668 5628 80724 5684
rect 80220 4956 80276 5012
rect 80444 4844 80500 4900
rect 79772 2828 79828 2884
rect 81452 10108 81508 10164
rect 81276 9434 81332 9436
rect 81276 9382 81278 9434
rect 81278 9382 81330 9434
rect 81330 9382 81332 9434
rect 81276 9380 81332 9382
rect 81380 9434 81436 9436
rect 81380 9382 81382 9434
rect 81382 9382 81434 9434
rect 81434 9382 81436 9434
rect 81380 9380 81436 9382
rect 81484 9434 81540 9436
rect 81484 9382 81486 9434
rect 81486 9382 81538 9434
rect 81538 9382 81540 9434
rect 81484 9380 81540 9382
rect 81452 8930 81508 8932
rect 81452 8878 81454 8930
rect 81454 8878 81506 8930
rect 81506 8878 81508 8930
rect 81452 8876 81508 8878
rect 81004 8258 81060 8260
rect 81004 8206 81006 8258
rect 81006 8206 81058 8258
rect 81058 8206 81060 8258
rect 81004 8204 81060 8206
rect 81116 8092 81172 8148
rect 81004 6972 81060 7028
rect 81452 8092 81508 8148
rect 81276 7866 81332 7868
rect 81276 7814 81278 7866
rect 81278 7814 81330 7866
rect 81330 7814 81332 7866
rect 81276 7812 81332 7814
rect 81380 7866 81436 7868
rect 81380 7814 81382 7866
rect 81382 7814 81434 7866
rect 81434 7814 81436 7866
rect 81380 7812 81436 7814
rect 81484 7866 81540 7868
rect 81484 7814 81486 7866
rect 81486 7814 81538 7866
rect 81538 7814 81540 7866
rect 81484 7812 81540 7814
rect 81900 10108 81956 10164
rect 82236 10556 82292 10612
rect 84140 22482 84196 22484
rect 84140 22430 84142 22482
rect 84142 22430 84194 22482
rect 84194 22430 84196 22482
rect 84140 22428 84196 22430
rect 85260 22482 85316 22484
rect 85260 22430 85262 22482
rect 85262 22430 85314 22482
rect 85314 22430 85316 22482
rect 85260 22428 85316 22430
rect 84028 19964 84084 20020
rect 84700 22204 84756 22260
rect 83692 18620 83748 18676
rect 83468 18450 83524 18452
rect 83468 18398 83470 18450
rect 83470 18398 83522 18450
rect 83522 18398 83524 18450
rect 83468 18396 83524 18398
rect 83468 17724 83524 17780
rect 83580 16882 83636 16884
rect 83580 16830 83582 16882
rect 83582 16830 83634 16882
rect 83634 16830 83636 16882
rect 83580 16828 83636 16830
rect 83468 16716 83524 16772
rect 83132 15874 83188 15876
rect 83132 15822 83134 15874
rect 83134 15822 83186 15874
rect 83186 15822 83188 15874
rect 83132 15820 83188 15822
rect 83580 15874 83636 15876
rect 83580 15822 83582 15874
rect 83582 15822 83634 15874
rect 83634 15822 83636 15874
rect 83580 15820 83636 15822
rect 83468 15426 83524 15428
rect 83468 15374 83470 15426
rect 83470 15374 83522 15426
rect 83522 15374 83524 15426
rect 83468 15372 83524 15374
rect 82796 15036 82852 15092
rect 82572 14588 82628 14644
rect 82572 14364 82628 14420
rect 83132 14642 83188 14644
rect 83132 14590 83134 14642
rect 83134 14590 83186 14642
rect 83186 14590 83188 14642
rect 83132 14588 83188 14590
rect 83020 14364 83076 14420
rect 83580 14140 83636 14196
rect 83580 13916 83636 13972
rect 82460 10108 82516 10164
rect 82348 9996 82404 10052
rect 82460 9772 82516 9828
rect 82236 8316 82292 8372
rect 81116 6748 81172 6804
rect 81116 6578 81172 6580
rect 81116 6526 81118 6578
rect 81118 6526 81170 6578
rect 81170 6526 81172 6578
rect 81116 6524 81172 6526
rect 81276 6298 81332 6300
rect 81276 6246 81278 6298
rect 81278 6246 81330 6298
rect 81330 6246 81332 6298
rect 81276 6244 81332 6246
rect 81380 6298 81436 6300
rect 81380 6246 81382 6298
rect 81382 6246 81434 6298
rect 81434 6246 81436 6298
rect 81380 6244 81436 6246
rect 81484 6298 81540 6300
rect 81484 6246 81486 6298
rect 81486 6246 81538 6298
rect 81538 6246 81540 6298
rect 81484 6244 81540 6246
rect 81788 6466 81844 6468
rect 81788 6414 81790 6466
rect 81790 6414 81842 6466
rect 81842 6414 81844 6466
rect 81788 6412 81844 6414
rect 81276 4730 81332 4732
rect 81276 4678 81278 4730
rect 81278 4678 81330 4730
rect 81330 4678 81332 4730
rect 81276 4676 81332 4678
rect 81380 4730 81436 4732
rect 81380 4678 81382 4730
rect 81382 4678 81434 4730
rect 81434 4678 81436 4730
rect 81380 4676 81436 4678
rect 81484 4730 81540 4732
rect 81484 4678 81486 4730
rect 81486 4678 81538 4730
rect 81538 4678 81540 4730
rect 81484 4676 81540 4678
rect 81116 4396 81172 4452
rect 81788 3612 81844 3668
rect 81276 3162 81332 3164
rect 81276 3110 81278 3162
rect 81278 3110 81330 3162
rect 81330 3110 81332 3162
rect 81276 3108 81332 3110
rect 81380 3162 81436 3164
rect 81380 3110 81382 3162
rect 81382 3110 81434 3162
rect 81434 3110 81436 3162
rect 81380 3108 81436 3110
rect 81484 3162 81540 3164
rect 81484 3110 81486 3162
rect 81486 3110 81538 3162
rect 81538 3110 81540 3162
rect 81484 3108 81540 3110
rect 80556 2828 80612 2884
rect 80556 924 80612 980
rect 82124 7420 82180 7476
rect 82348 6802 82404 6804
rect 82348 6750 82350 6802
rect 82350 6750 82402 6802
rect 82402 6750 82404 6802
rect 82348 6748 82404 6750
rect 82572 9602 82628 9604
rect 82572 9550 82574 9602
rect 82574 9550 82626 9602
rect 82626 9550 82628 9602
rect 82572 9548 82628 9550
rect 82796 13468 82852 13524
rect 83468 13356 83524 13412
rect 82796 12850 82852 12852
rect 82796 12798 82798 12850
rect 82798 12798 82850 12850
rect 82850 12798 82852 12850
rect 82796 12796 82852 12798
rect 82908 10610 82964 10612
rect 82908 10558 82910 10610
rect 82910 10558 82962 10610
rect 82962 10558 82964 10610
rect 82908 10556 82964 10558
rect 82908 9714 82964 9716
rect 82908 9662 82910 9714
rect 82910 9662 82962 9714
rect 82962 9662 82964 9714
rect 82908 9660 82964 9662
rect 82908 9100 82964 9156
rect 83244 12684 83300 12740
rect 83244 12124 83300 12180
rect 83132 11900 83188 11956
rect 83468 11788 83524 11844
rect 83244 10332 83300 10388
rect 83132 8764 83188 8820
rect 83580 11340 83636 11396
rect 83580 10892 83636 10948
rect 83580 9826 83636 9828
rect 83580 9774 83582 9826
rect 83582 9774 83634 9826
rect 83634 9774 83636 9826
rect 83580 9772 83636 9774
rect 82684 7868 82740 7924
rect 82684 7420 82740 7476
rect 82572 7084 82628 7140
rect 82348 4844 82404 4900
rect 83468 6860 83524 6916
rect 83580 8988 83636 9044
rect 82796 5794 82852 5796
rect 82796 5742 82798 5794
rect 82798 5742 82850 5794
rect 82850 5742 82852 5794
rect 82796 5740 82852 5742
rect 82908 5122 82964 5124
rect 82908 5070 82910 5122
rect 82910 5070 82962 5122
rect 82962 5070 82964 5122
rect 82908 5068 82964 5070
rect 83244 5122 83300 5124
rect 83244 5070 83246 5122
rect 83246 5070 83298 5122
rect 83298 5070 83300 5122
rect 83244 5068 83300 5070
rect 83132 4620 83188 4676
rect 82460 4060 82516 4116
rect 83020 3666 83076 3668
rect 83020 3614 83022 3666
rect 83022 3614 83074 3666
rect 83074 3614 83076 3666
rect 83020 3612 83076 3614
rect 83916 18396 83972 18452
rect 83916 17106 83972 17108
rect 83916 17054 83918 17106
rect 83918 17054 83970 17106
rect 83970 17054 83972 17106
rect 83916 17052 83972 17054
rect 84476 18338 84532 18340
rect 84476 18286 84478 18338
rect 84478 18286 84530 18338
rect 84530 18286 84532 18338
rect 84476 18284 84532 18286
rect 84252 17778 84308 17780
rect 84252 17726 84254 17778
rect 84254 17726 84306 17778
rect 84306 17726 84308 17778
rect 84252 17724 84308 17726
rect 84364 17442 84420 17444
rect 84364 17390 84366 17442
rect 84366 17390 84418 17442
rect 84418 17390 84420 17442
rect 84364 17388 84420 17390
rect 84028 16828 84084 16884
rect 84028 13804 84084 13860
rect 83916 13468 83972 13524
rect 83804 13020 83860 13076
rect 83916 12348 83972 12404
rect 83804 11900 83860 11956
rect 84252 14028 84308 14084
rect 86380 22652 86436 22708
rect 86716 22876 86772 22932
rect 86268 20748 86324 20804
rect 85260 19292 85316 19348
rect 84812 18508 84868 18564
rect 85148 17442 85204 17444
rect 85148 17390 85150 17442
rect 85150 17390 85202 17442
rect 85202 17390 85204 17442
rect 85148 17388 85204 17390
rect 84812 14700 84868 14756
rect 84700 14588 84756 14644
rect 84700 13916 84756 13972
rect 84252 13692 84308 13748
rect 84252 12908 84308 12964
rect 84588 13580 84644 13636
rect 84476 12796 84532 12852
rect 85148 15874 85204 15876
rect 85148 15822 85150 15874
rect 85150 15822 85202 15874
rect 85202 15822 85204 15874
rect 85148 15820 85204 15822
rect 84812 12962 84868 12964
rect 84812 12910 84814 12962
rect 84814 12910 84866 12962
rect 84866 12910 84868 12962
rect 84812 12908 84868 12910
rect 85148 15596 85204 15652
rect 84140 11564 84196 11620
rect 84252 12124 84308 12180
rect 84140 11394 84196 11396
rect 84140 11342 84142 11394
rect 84142 11342 84194 11394
rect 84194 11342 84196 11394
rect 84140 11340 84196 11342
rect 83916 10834 83972 10836
rect 83916 10782 83918 10834
rect 83918 10782 83970 10834
rect 83970 10782 83972 10834
rect 83916 10780 83972 10782
rect 83916 10556 83972 10612
rect 83804 8428 83860 8484
rect 83916 9660 83972 9716
rect 83916 7084 83972 7140
rect 84028 8316 84084 8372
rect 84700 12012 84756 12068
rect 84588 11788 84644 11844
rect 84476 11564 84532 11620
rect 84364 11340 84420 11396
rect 84476 11282 84532 11284
rect 84476 11230 84478 11282
rect 84478 11230 84530 11282
rect 84530 11230 84532 11282
rect 84476 11228 84532 11230
rect 85484 19010 85540 19012
rect 85484 18958 85486 19010
rect 85486 18958 85538 19010
rect 85538 18958 85540 19010
rect 85484 18956 85540 18958
rect 85372 18284 85428 18340
rect 85372 17666 85428 17668
rect 85372 17614 85374 17666
rect 85374 17614 85426 17666
rect 85426 17614 85428 17666
rect 85372 17612 85428 17614
rect 85820 18620 85876 18676
rect 85820 18450 85876 18452
rect 85820 18398 85822 18450
rect 85822 18398 85874 18450
rect 85874 18398 85876 18450
rect 85820 18396 85876 18398
rect 85484 16828 85540 16884
rect 86268 19346 86324 19348
rect 86268 19294 86270 19346
rect 86270 19294 86322 19346
rect 86322 19294 86324 19346
rect 86268 19292 86324 19294
rect 86156 18956 86212 19012
rect 86380 18450 86436 18452
rect 86380 18398 86382 18450
rect 86382 18398 86434 18450
rect 86434 18398 86436 18450
rect 86380 18396 86436 18398
rect 86044 17724 86100 17780
rect 86268 17612 86324 17668
rect 85932 17164 85988 17220
rect 87388 22876 87444 22932
rect 86940 21756 86996 21812
rect 87164 21698 87220 21700
rect 87164 21646 87166 21698
rect 87166 21646 87218 21698
rect 87218 21646 87220 21698
rect 87164 21644 87220 21646
rect 87612 20802 87668 20804
rect 87612 20750 87614 20802
rect 87614 20750 87666 20802
rect 87666 20750 87668 20802
rect 87612 20748 87668 20750
rect 86604 19404 86660 19460
rect 87276 19404 87332 19460
rect 86828 19292 86884 19348
rect 86604 19010 86660 19012
rect 86604 18958 86606 19010
rect 86606 18958 86658 19010
rect 86658 18958 86660 19010
rect 86604 18956 86660 18958
rect 88172 25506 88228 25508
rect 88172 25454 88174 25506
rect 88174 25454 88226 25506
rect 88226 25454 88228 25506
rect 88172 25452 88228 25454
rect 88396 21810 88452 21812
rect 88396 21758 88398 21810
rect 88398 21758 88450 21810
rect 88450 21758 88452 21810
rect 88396 21756 88452 21758
rect 88508 21698 88564 21700
rect 88508 21646 88510 21698
rect 88510 21646 88562 21698
rect 88562 21646 88564 21698
rect 88508 21644 88564 21646
rect 88060 19010 88116 19012
rect 88060 18958 88062 19010
rect 88062 18958 88114 19010
rect 88114 18958 88116 19010
rect 88060 18956 88116 18958
rect 87724 17948 87780 18004
rect 88732 21532 88788 21588
rect 88284 18732 88340 18788
rect 87948 17948 88004 18004
rect 87948 17666 88004 17668
rect 87948 17614 87950 17666
rect 87950 17614 88002 17666
rect 88002 17614 88004 17666
rect 87948 17612 88004 17614
rect 87276 17500 87332 17556
rect 87388 17388 87444 17444
rect 85260 15148 85316 15204
rect 85260 14642 85316 14644
rect 85260 14590 85262 14642
rect 85262 14590 85314 14642
rect 85314 14590 85316 14642
rect 85260 14588 85316 14590
rect 85260 14252 85316 14308
rect 85260 13916 85316 13972
rect 85148 12012 85204 12068
rect 84924 11116 84980 11172
rect 85036 11340 85092 11396
rect 84924 10668 84980 10724
rect 84364 10444 84420 10500
rect 84476 10386 84532 10388
rect 84476 10334 84478 10386
rect 84478 10334 84530 10386
rect 84530 10334 84532 10386
rect 84476 10332 84532 10334
rect 84588 9884 84644 9940
rect 84476 9436 84532 9492
rect 84588 9100 84644 9156
rect 84476 8316 84532 8372
rect 84476 7196 84532 7252
rect 84700 8540 84756 8596
rect 84812 9602 84868 9604
rect 84812 9550 84814 9602
rect 84814 9550 84866 9602
rect 84866 9550 84868 9602
rect 84812 9548 84868 9550
rect 85036 9324 85092 9380
rect 85484 11676 85540 11732
rect 85372 10444 85428 10500
rect 85484 9996 85540 10052
rect 85260 8316 85316 8372
rect 85484 8428 85540 8484
rect 85036 8092 85092 8148
rect 85148 7980 85204 8036
rect 84476 6860 84532 6916
rect 84364 6748 84420 6804
rect 83692 4844 83748 4900
rect 84140 6524 84196 6580
rect 84476 6524 84532 6580
rect 84700 6412 84756 6468
rect 84140 6300 84196 6356
rect 85036 6300 85092 6356
rect 84924 6188 84980 6244
rect 85260 7644 85316 7700
rect 85484 6748 85540 6804
rect 85260 6636 85316 6692
rect 85932 15874 85988 15876
rect 85932 15822 85934 15874
rect 85934 15822 85986 15874
rect 85986 15822 85988 15874
rect 85932 15820 85988 15822
rect 86268 15708 86324 15764
rect 86268 15260 86324 15316
rect 85708 13746 85764 13748
rect 85708 13694 85710 13746
rect 85710 13694 85762 13746
rect 85762 13694 85764 13746
rect 85708 13692 85764 13694
rect 85932 13970 85988 13972
rect 85932 13918 85934 13970
rect 85934 13918 85986 13970
rect 85986 13918 85988 13970
rect 85932 13916 85988 13918
rect 86380 15036 86436 15092
rect 85820 13132 85876 13188
rect 86156 14252 86212 14308
rect 85708 12402 85764 12404
rect 85708 12350 85710 12402
rect 85710 12350 85762 12402
rect 85762 12350 85764 12402
rect 85708 12348 85764 12350
rect 85820 12290 85876 12292
rect 85820 12238 85822 12290
rect 85822 12238 85874 12290
rect 85874 12238 85876 12290
rect 85820 12236 85876 12238
rect 86268 14140 86324 14196
rect 86604 14028 86660 14084
rect 86492 12908 86548 12964
rect 86492 12348 86548 12404
rect 86156 12236 86212 12292
rect 86044 11564 86100 11620
rect 86268 11394 86324 11396
rect 86268 11342 86270 11394
rect 86270 11342 86322 11394
rect 86322 11342 86324 11394
rect 86268 11340 86324 11342
rect 86380 11228 86436 11284
rect 85820 10556 85876 10612
rect 86044 10220 86100 10276
rect 85932 9714 85988 9716
rect 85932 9662 85934 9714
rect 85934 9662 85986 9714
rect 85986 9662 85988 9714
rect 85932 9660 85988 9662
rect 86268 9042 86324 9044
rect 86268 8990 86270 9042
rect 86270 8990 86322 9042
rect 86322 8990 86324 9042
rect 86268 8988 86324 8990
rect 86604 9714 86660 9716
rect 86604 9662 86606 9714
rect 86606 9662 86658 9714
rect 86658 9662 86660 9714
rect 86604 9660 86660 9662
rect 86492 9602 86548 9604
rect 86492 9550 86494 9602
rect 86494 9550 86546 9602
rect 86546 9550 86548 9602
rect 86492 9548 86548 9550
rect 86828 14812 86884 14868
rect 86940 14588 86996 14644
rect 87388 16716 87444 16772
rect 87948 16044 88004 16100
rect 87276 15260 87332 15316
rect 88172 18396 88228 18452
rect 88508 17948 88564 18004
rect 88284 17724 88340 17780
rect 88620 17612 88676 17668
rect 89628 30380 89684 30436
rect 89180 29372 89236 29428
rect 88956 25506 89012 25508
rect 88956 25454 88958 25506
rect 88958 25454 89010 25506
rect 89010 25454 89012 25506
rect 88956 25452 89012 25454
rect 89068 18060 89124 18116
rect 89068 16940 89124 16996
rect 88732 16268 88788 16324
rect 87164 14252 87220 14308
rect 87388 14700 87444 14756
rect 87500 13580 87556 13636
rect 87948 13580 88004 13636
rect 87276 12066 87332 12068
rect 87276 12014 87278 12066
rect 87278 12014 87330 12066
rect 87330 12014 87332 12066
rect 87276 12012 87332 12014
rect 86828 11676 86884 11732
rect 86940 11900 86996 11956
rect 88844 15484 88900 15540
rect 88172 14252 88228 14308
rect 88396 13132 88452 13188
rect 88284 13020 88340 13076
rect 88060 12572 88116 12628
rect 88284 12684 88340 12740
rect 88060 12402 88116 12404
rect 88060 12350 88062 12402
rect 88062 12350 88114 12402
rect 88114 12350 88116 12402
rect 88060 12348 88116 12350
rect 86940 11004 86996 11060
rect 87388 10892 87444 10948
rect 87276 10498 87332 10500
rect 87276 10446 87278 10498
rect 87278 10446 87330 10498
rect 87330 10446 87332 10498
rect 87276 10444 87332 10446
rect 86492 9154 86548 9156
rect 86492 9102 86494 9154
rect 86494 9102 86546 9154
rect 86546 9102 86548 9154
rect 86492 9100 86548 9102
rect 86156 8428 86212 8484
rect 85932 8204 85988 8260
rect 86828 8428 86884 8484
rect 86940 9324 86996 9380
rect 86268 8370 86324 8372
rect 86268 8318 86270 8370
rect 86270 8318 86322 8370
rect 86322 8318 86324 8370
rect 86268 8316 86324 8318
rect 86940 8316 86996 8372
rect 86044 7980 86100 8036
rect 86492 8146 86548 8148
rect 86492 8094 86494 8146
rect 86494 8094 86546 8146
rect 86546 8094 86548 8146
rect 86492 8092 86548 8094
rect 86604 7980 86660 8036
rect 85820 7308 85876 7364
rect 86156 7362 86212 7364
rect 86156 7310 86158 7362
rect 86158 7310 86210 7362
rect 86210 7310 86212 7362
rect 86156 7308 86212 7310
rect 85708 6860 85764 6916
rect 86156 7084 86212 7140
rect 85932 6578 85988 6580
rect 85932 6526 85934 6578
rect 85934 6526 85986 6578
rect 85986 6526 85988 6578
rect 85932 6524 85988 6526
rect 85596 6300 85652 6356
rect 85820 5906 85876 5908
rect 85820 5854 85822 5906
rect 85822 5854 85874 5906
rect 85874 5854 85876 5906
rect 85820 5852 85876 5854
rect 86492 7756 86548 7812
rect 86492 7084 86548 7140
rect 86828 7868 86884 7924
rect 86716 7474 86772 7476
rect 86716 7422 86718 7474
rect 86718 7422 86770 7474
rect 86770 7422 86772 7474
rect 86716 7420 86772 7422
rect 86828 7308 86884 7364
rect 86716 7196 86772 7252
rect 85036 4620 85092 4676
rect 85484 4620 85540 4676
rect 85596 4508 85652 4564
rect 84028 3276 84084 3332
rect 84476 4396 84532 4452
rect 85484 4284 85540 4340
rect 85484 3554 85540 3556
rect 85484 3502 85486 3554
rect 85486 3502 85538 3554
rect 85538 3502 85540 3554
rect 85484 3500 85540 3502
rect 85596 4172 85652 4228
rect 86044 4508 86100 4564
rect 86268 5794 86324 5796
rect 86268 5742 86270 5794
rect 86270 5742 86322 5794
rect 86322 5742 86324 5794
rect 86268 5740 86324 5742
rect 86156 4284 86212 4340
rect 86268 5516 86324 5572
rect 86604 6300 86660 6356
rect 86492 5906 86548 5908
rect 86492 5854 86494 5906
rect 86494 5854 86546 5906
rect 86546 5854 86548 5906
rect 86492 5852 86548 5854
rect 86380 5068 86436 5124
rect 86492 4562 86548 4564
rect 86492 4510 86494 4562
rect 86494 4510 86546 4562
rect 86546 4510 86548 4562
rect 86492 4508 86548 4510
rect 86716 5740 86772 5796
rect 87836 10556 87892 10612
rect 87612 9212 87668 9268
rect 87164 8034 87220 8036
rect 87164 7982 87166 8034
rect 87166 7982 87218 8034
rect 87218 7982 87220 8034
rect 87164 7980 87220 7982
rect 87052 7196 87108 7252
rect 86940 6412 86996 6468
rect 87388 8316 87444 8372
rect 87388 7868 87444 7924
rect 87164 6188 87220 6244
rect 87276 6636 87332 6692
rect 86940 4956 86996 5012
rect 87052 5740 87108 5796
rect 87164 5628 87220 5684
rect 87052 5292 87108 5348
rect 86604 4396 86660 4452
rect 87164 4844 87220 4900
rect 87724 7196 87780 7252
rect 87724 6748 87780 6804
rect 88508 12290 88564 12292
rect 88508 12238 88510 12290
rect 88510 12238 88562 12290
rect 88562 12238 88564 12290
rect 88508 12236 88564 12238
rect 88508 11394 88564 11396
rect 88508 11342 88510 11394
rect 88510 11342 88562 11394
rect 88562 11342 88564 11394
rect 88508 11340 88564 11342
rect 87948 7308 88004 7364
rect 88508 10220 88564 10276
rect 87836 6636 87892 6692
rect 87724 6524 87780 6580
rect 87836 5906 87892 5908
rect 87836 5854 87838 5906
rect 87838 5854 87890 5906
rect 87890 5854 87892 5906
rect 87836 5852 87892 5854
rect 87164 4060 87220 4116
rect 85932 3388 85988 3444
rect 87052 3388 87108 3444
rect 88172 6748 88228 6804
rect 88060 6412 88116 6468
rect 88396 8146 88452 8148
rect 88396 8094 88398 8146
rect 88398 8094 88450 8146
rect 88450 8094 88452 8146
rect 88396 8092 88452 8094
rect 88844 14252 88900 14308
rect 88732 12962 88788 12964
rect 88732 12910 88734 12962
rect 88734 12910 88786 12962
rect 88786 12910 88788 12962
rect 88732 12908 88788 12910
rect 88956 12962 89012 12964
rect 88956 12910 88958 12962
rect 88958 12910 89010 12962
rect 89010 12910 89012 12962
rect 88956 12908 89012 12910
rect 88844 11116 88900 11172
rect 88732 10610 88788 10612
rect 88732 10558 88734 10610
rect 88734 10558 88786 10610
rect 88786 10558 88788 10610
rect 88732 10556 88788 10558
rect 88732 9548 88788 9604
rect 88620 8204 88676 8260
rect 89516 22204 89572 22260
rect 92540 55186 92596 55188
rect 92540 55134 92542 55186
rect 92542 55134 92594 55186
rect 92594 55134 92596 55186
rect 92540 55132 92596 55134
rect 92988 55132 93044 55188
rect 94556 55020 94612 55076
rect 89740 25506 89796 25508
rect 89740 25454 89742 25506
rect 89742 25454 89794 25506
rect 89794 25454 89796 25506
rect 89740 25452 89796 25454
rect 91084 30268 91140 30324
rect 90524 22652 90580 22708
rect 90300 22258 90356 22260
rect 90300 22206 90302 22258
rect 90302 22206 90354 22258
rect 90354 22206 90356 22258
rect 90300 22204 90356 22206
rect 90972 22258 91028 22260
rect 90972 22206 90974 22258
rect 90974 22206 91026 22258
rect 91026 22206 91028 22258
rect 90972 22204 91028 22206
rect 92316 24556 92372 24612
rect 92092 23324 92148 23380
rect 91756 22652 91812 22708
rect 91196 22428 91252 22484
rect 91980 22482 92036 22484
rect 91980 22430 91982 22482
rect 91982 22430 92034 22482
rect 92034 22430 92036 22482
rect 91980 22428 92036 22430
rect 89740 21532 89796 21588
rect 90524 21586 90580 21588
rect 90524 21534 90526 21586
rect 90526 21534 90578 21586
rect 90578 21534 90580 21586
rect 90524 21532 90580 21534
rect 89628 18284 89684 18340
rect 89628 17778 89684 17780
rect 89628 17726 89630 17778
rect 89630 17726 89682 17778
rect 89682 17726 89684 17778
rect 89628 17724 89684 17726
rect 89292 17276 89348 17332
rect 89292 16940 89348 16996
rect 89292 15372 89348 15428
rect 89740 16882 89796 16884
rect 89740 16830 89742 16882
rect 89742 16830 89794 16882
rect 89794 16830 89796 16882
rect 89740 16828 89796 16830
rect 89292 15148 89348 15204
rect 90300 18450 90356 18452
rect 90300 18398 90302 18450
rect 90302 18398 90354 18450
rect 90354 18398 90356 18450
rect 90300 18396 90356 18398
rect 90636 17836 90692 17892
rect 90748 17724 90804 17780
rect 89964 16156 90020 16212
rect 90860 17276 90916 17332
rect 90748 16210 90804 16212
rect 90748 16158 90750 16210
rect 90750 16158 90802 16210
rect 90802 16158 90804 16210
rect 90748 16156 90804 16158
rect 90636 16098 90692 16100
rect 90636 16046 90638 16098
rect 90638 16046 90690 16098
rect 90690 16046 90692 16098
rect 90636 16044 90692 16046
rect 90748 15372 90804 15428
rect 89852 13804 89908 13860
rect 89404 13356 89460 13412
rect 89292 12738 89348 12740
rect 89292 12686 89294 12738
rect 89294 12686 89346 12738
rect 89346 12686 89348 12738
rect 89292 12684 89348 12686
rect 89516 12796 89572 12852
rect 89180 12012 89236 12068
rect 89404 12012 89460 12068
rect 89404 11452 89460 11508
rect 89628 12684 89684 12740
rect 89628 11676 89684 11732
rect 90188 15148 90244 15204
rect 89628 10892 89684 10948
rect 89180 10556 89236 10612
rect 89068 9660 89124 9716
rect 89180 9436 89236 9492
rect 89292 8652 89348 8708
rect 89516 7308 89572 7364
rect 89628 9996 89684 10052
rect 89068 6466 89124 6468
rect 89068 6414 89070 6466
rect 89070 6414 89122 6466
rect 89122 6414 89124 6466
rect 89068 6412 89124 6414
rect 88956 6300 89012 6356
rect 88284 5740 88340 5796
rect 87948 2604 88004 2660
rect 88508 5628 88564 5684
rect 88620 5068 88676 5124
rect 89068 2940 89124 2996
rect 89292 6188 89348 6244
rect 89516 6636 89572 6692
rect 89404 5516 89460 5572
rect 89852 9436 89908 9492
rect 90524 13634 90580 13636
rect 90524 13582 90526 13634
rect 90526 13582 90578 13634
rect 90578 13582 90580 13634
rect 90524 13580 90580 13582
rect 90076 13132 90132 13188
rect 90076 12908 90132 12964
rect 90524 12962 90580 12964
rect 90524 12910 90526 12962
rect 90526 12910 90578 12962
rect 90578 12910 90580 12962
rect 90524 12908 90580 12910
rect 90300 12402 90356 12404
rect 90300 12350 90302 12402
rect 90302 12350 90354 12402
rect 90354 12350 90356 12402
rect 90300 12348 90356 12350
rect 90076 11676 90132 11732
rect 90188 10444 90244 10500
rect 90860 15148 90916 15204
rect 90748 14140 90804 14196
rect 90860 13468 90916 13524
rect 90636 11170 90692 11172
rect 90636 11118 90638 11170
rect 90638 11118 90690 11170
rect 90690 11118 90692 11170
rect 90636 11116 90692 11118
rect 90636 9100 90692 9156
rect 89852 7868 89908 7924
rect 90188 8034 90244 8036
rect 90188 7982 90190 8034
rect 90190 7982 90242 8034
rect 90242 7982 90244 8034
rect 90188 7980 90244 7982
rect 90076 7532 90132 7588
rect 89964 7420 90020 7476
rect 89628 5180 89684 5236
rect 89964 4450 90020 4452
rect 89964 4398 89966 4450
rect 89966 4398 90018 4450
rect 90018 4398 90020 4450
rect 89964 4396 90020 4398
rect 89628 4172 89684 4228
rect 89180 1596 89236 1652
rect 90524 8258 90580 8260
rect 90524 8206 90526 8258
rect 90526 8206 90578 8258
rect 90578 8206 90580 8258
rect 90524 8204 90580 8206
rect 90860 12796 90916 12852
rect 91196 21420 91252 21476
rect 91084 21084 91140 21140
rect 91308 20914 91364 20916
rect 91308 20862 91310 20914
rect 91310 20862 91362 20914
rect 91362 20862 91364 20914
rect 91308 20860 91364 20862
rect 92092 21980 92148 22036
rect 91868 21644 91924 21700
rect 91980 21420 92036 21476
rect 91084 19740 91140 19796
rect 91084 19122 91140 19124
rect 91084 19070 91086 19122
rect 91086 19070 91138 19122
rect 91138 19070 91140 19122
rect 91084 19068 91140 19070
rect 92092 20802 92148 20804
rect 92092 20750 92094 20802
rect 92094 20750 92146 20802
rect 92146 20750 92148 20802
rect 92092 20748 92148 20750
rect 91868 20188 91924 20244
rect 91756 19852 91812 19908
rect 91196 17442 91252 17444
rect 91196 17390 91198 17442
rect 91198 17390 91250 17442
rect 91250 17390 91252 17442
rect 91196 17388 91252 17390
rect 91084 16828 91140 16884
rect 91084 16380 91140 16436
rect 91196 14588 91252 14644
rect 91196 14364 91252 14420
rect 91196 13468 91252 13524
rect 91084 13356 91140 13412
rect 91532 18844 91588 18900
rect 91756 18956 91812 19012
rect 91308 12908 91364 12964
rect 90860 11676 90916 11732
rect 90972 10892 91028 10948
rect 91308 10444 91364 10500
rect 91532 15202 91588 15204
rect 91532 15150 91534 15202
rect 91534 15150 91586 15202
rect 91586 15150 91588 15202
rect 91532 15148 91588 15150
rect 91980 19068 92036 19124
rect 92652 23714 92708 23716
rect 92652 23662 92654 23714
rect 92654 23662 92706 23714
rect 92706 23662 92708 23714
rect 92652 23660 92708 23662
rect 92316 21868 92372 21924
rect 92540 21420 92596 21476
rect 93100 23042 93156 23044
rect 93100 22990 93102 23042
rect 93102 22990 93154 23042
rect 93154 22990 93156 23042
rect 93100 22988 93156 22990
rect 92876 22652 92932 22708
rect 92988 22540 93044 22596
rect 92652 21980 92708 22036
rect 92428 20972 92484 21028
rect 92428 20802 92484 20804
rect 92428 20750 92430 20802
rect 92430 20750 92482 20802
rect 92482 20750 92484 20802
rect 92428 20748 92484 20750
rect 92540 20412 92596 20468
rect 92428 19010 92484 19012
rect 92428 18958 92430 19010
rect 92430 18958 92482 19010
rect 92482 18958 92484 19010
rect 92428 18956 92484 18958
rect 92540 18844 92596 18900
rect 92204 18284 92260 18340
rect 91980 17836 92036 17892
rect 92540 18284 92596 18340
rect 91980 16940 92036 16996
rect 91980 16380 92036 16436
rect 92204 17554 92260 17556
rect 92204 17502 92206 17554
rect 92206 17502 92258 17554
rect 92258 17502 92260 17554
rect 92204 17500 92260 17502
rect 92092 16156 92148 16212
rect 91532 14588 91588 14644
rect 91532 12684 91588 12740
rect 92764 21644 92820 21700
rect 92876 21084 92932 21140
rect 92988 20972 93044 21028
rect 92876 20802 92932 20804
rect 92876 20750 92878 20802
rect 92878 20750 92930 20802
rect 92930 20750 92932 20802
rect 92876 20748 92932 20750
rect 92876 20412 92932 20468
rect 92764 16828 92820 16884
rect 92988 20188 93044 20244
rect 93324 23660 93380 23716
rect 93324 23266 93380 23268
rect 93324 23214 93326 23266
rect 93326 23214 93378 23266
rect 93378 23214 93380 23266
rect 93324 23212 93380 23214
rect 93772 21698 93828 21700
rect 93772 21646 93774 21698
rect 93774 21646 93826 21698
rect 93826 21646 93828 21698
rect 93772 21644 93828 21646
rect 93212 21532 93268 21588
rect 93436 20972 93492 21028
rect 93548 21420 93604 21476
rect 94444 21420 94500 21476
rect 93996 21084 94052 21140
rect 93324 20524 93380 20580
rect 93772 20578 93828 20580
rect 93772 20526 93774 20578
rect 93774 20526 93826 20578
rect 93826 20526 93828 20578
rect 93772 20524 93828 20526
rect 93212 19906 93268 19908
rect 93212 19854 93214 19906
rect 93214 19854 93266 19906
rect 93266 19854 93268 19906
rect 93212 19852 93268 19854
rect 92988 17500 93044 17556
rect 93548 18562 93604 18564
rect 93548 18510 93550 18562
rect 93550 18510 93602 18562
rect 93602 18510 93604 18562
rect 93548 18508 93604 18510
rect 94444 18338 94500 18340
rect 94444 18286 94446 18338
rect 94446 18286 94498 18338
rect 94498 18286 94500 18338
rect 94444 18284 94500 18286
rect 92988 16940 93044 16996
rect 92876 16044 92932 16100
rect 92316 14700 92372 14756
rect 91756 14140 91812 14196
rect 91756 13132 91812 13188
rect 91756 12908 91812 12964
rect 92428 14028 92484 14084
rect 91980 13132 92036 13188
rect 91644 11116 91700 11172
rect 90860 9436 90916 9492
rect 90748 8428 90804 8484
rect 90524 6972 90580 7028
rect 90524 6188 90580 6244
rect 90860 7362 90916 7364
rect 90860 7310 90862 7362
rect 90862 7310 90914 7362
rect 90914 7310 90916 7362
rect 90860 7308 90916 7310
rect 90860 6412 90916 6468
rect 91532 10780 91588 10836
rect 91196 9100 91252 9156
rect 91196 8764 91252 8820
rect 91532 9436 91588 9492
rect 91420 8370 91476 8372
rect 91420 8318 91422 8370
rect 91422 8318 91474 8370
rect 91474 8318 91476 8370
rect 91420 8316 91476 8318
rect 91868 12460 91924 12516
rect 91980 11452 92036 11508
rect 92876 14252 92932 14308
rect 92988 15036 93044 15092
rect 93100 14530 93156 14532
rect 93100 14478 93102 14530
rect 93102 14478 93154 14530
rect 93154 14478 93156 14530
rect 93100 14476 93156 14478
rect 93100 13580 93156 13636
rect 92204 12684 92260 12740
rect 92316 11564 92372 11620
rect 92876 12684 92932 12740
rect 92988 12460 93044 12516
rect 92988 11788 93044 11844
rect 92204 10780 92260 10836
rect 92092 10668 92148 10724
rect 92204 10610 92260 10612
rect 92204 10558 92206 10610
rect 92206 10558 92258 10610
rect 92258 10558 92260 10610
rect 92204 10556 92260 10558
rect 92652 10722 92708 10724
rect 92652 10670 92654 10722
rect 92654 10670 92706 10722
rect 92706 10670 92708 10722
rect 92652 10668 92708 10670
rect 93100 11282 93156 11284
rect 93100 11230 93102 11282
rect 93102 11230 93154 11282
rect 93154 11230 93156 11282
rect 93100 11228 93156 11230
rect 92988 11170 93044 11172
rect 92988 11118 92990 11170
rect 92990 11118 93042 11170
rect 93042 11118 93044 11170
rect 92988 11116 93044 11118
rect 92652 9826 92708 9828
rect 92652 9774 92654 9826
rect 92654 9774 92706 9826
rect 92706 9774 92708 9826
rect 92652 9772 92708 9774
rect 92316 9100 92372 9156
rect 92652 9548 92708 9604
rect 92092 8764 92148 8820
rect 91196 4508 91252 4564
rect 91084 3612 91140 3668
rect 91196 3948 91252 4004
rect 90860 2940 90916 2996
rect 90524 2268 90580 2324
rect 92092 7586 92148 7588
rect 92092 7534 92094 7586
rect 92094 7534 92146 7586
rect 92146 7534 92148 7586
rect 92092 7532 92148 7534
rect 92204 7420 92260 7476
rect 92204 6748 92260 6804
rect 91868 6018 91924 6020
rect 91868 5966 91870 6018
rect 91870 5966 91922 6018
rect 91922 5966 91924 6018
rect 91868 5964 91924 5966
rect 91868 5628 91924 5684
rect 91980 5180 92036 5236
rect 93100 10498 93156 10500
rect 93100 10446 93102 10498
rect 93102 10446 93154 10498
rect 93154 10446 93156 10498
rect 93100 10444 93156 10446
rect 92764 8652 92820 8708
rect 92876 8764 92932 8820
rect 92876 8428 92932 8484
rect 92988 8316 93044 8372
rect 93100 7980 93156 8036
rect 93772 17500 93828 17556
rect 93324 16044 93380 16100
rect 93996 16210 94052 16212
rect 93996 16158 93998 16210
rect 93998 16158 94050 16210
rect 94050 16158 94052 16210
rect 93996 16156 94052 16158
rect 93548 16098 93604 16100
rect 93548 16046 93550 16098
rect 93550 16046 93602 16098
rect 93602 16046 93604 16098
rect 93548 16044 93604 16046
rect 93996 15372 94052 15428
rect 93996 15202 94052 15204
rect 93996 15150 93998 15202
rect 93998 15150 94050 15202
rect 94050 15150 94052 15202
rect 93996 15148 94052 15150
rect 94108 15036 94164 15092
rect 93548 13858 93604 13860
rect 93548 13806 93550 13858
rect 93550 13806 93602 13858
rect 93602 13806 93604 13858
rect 93548 13804 93604 13806
rect 93996 12962 94052 12964
rect 93996 12910 93998 12962
rect 93998 12910 94050 12962
rect 94050 12910 94052 12962
rect 93996 12908 94052 12910
rect 93548 11788 93604 11844
rect 93772 11788 93828 11844
rect 93660 11282 93716 11284
rect 93660 11230 93662 11282
rect 93662 11230 93714 11282
rect 93714 11230 93716 11282
rect 93660 11228 93716 11230
rect 93996 12684 94052 12740
rect 94332 17388 94388 17444
rect 94444 17164 94500 17220
rect 96908 55074 96964 55076
rect 96908 55022 96910 55074
rect 96910 55022 96962 55074
rect 96962 55022 96964 55074
rect 96908 55020 96964 55022
rect 104636 56252 104692 56308
rect 105868 56306 105924 56308
rect 105868 56254 105870 56306
rect 105870 56254 105922 56306
rect 105922 56254 105924 56306
rect 105868 56252 105924 56254
rect 111996 56474 112052 56476
rect 111996 56422 111998 56474
rect 111998 56422 112050 56474
rect 112050 56422 112052 56474
rect 111996 56420 112052 56422
rect 112100 56474 112156 56476
rect 112100 56422 112102 56474
rect 112102 56422 112154 56474
rect 112154 56422 112156 56474
rect 112100 56420 112156 56422
rect 112204 56474 112260 56476
rect 112204 56422 112206 56474
rect 112206 56422 112258 56474
rect 112258 56422 112260 56474
rect 112204 56420 112260 56422
rect 108444 56252 108500 56308
rect 109676 56306 109732 56308
rect 109676 56254 109678 56306
rect 109678 56254 109730 56306
rect 109730 56254 109732 56306
rect 109676 56252 109732 56254
rect 110012 56140 110068 56196
rect 97580 55020 97636 55076
rect 96636 54122 96692 54124
rect 96636 54070 96638 54122
rect 96638 54070 96690 54122
rect 96690 54070 96692 54122
rect 96636 54068 96692 54070
rect 96740 54122 96796 54124
rect 96740 54070 96742 54122
rect 96742 54070 96794 54122
rect 96794 54070 96796 54122
rect 96740 54068 96796 54070
rect 96844 54122 96900 54124
rect 96844 54070 96846 54122
rect 96846 54070 96898 54122
rect 96898 54070 96900 54122
rect 96844 54068 96900 54070
rect 96636 52554 96692 52556
rect 96636 52502 96638 52554
rect 96638 52502 96690 52554
rect 96690 52502 96692 52554
rect 96636 52500 96692 52502
rect 96740 52554 96796 52556
rect 96740 52502 96742 52554
rect 96742 52502 96794 52554
rect 96794 52502 96796 52554
rect 96740 52500 96796 52502
rect 96844 52554 96900 52556
rect 96844 52502 96846 52554
rect 96846 52502 96898 52554
rect 96898 52502 96900 52554
rect 96844 52500 96900 52502
rect 96636 50986 96692 50988
rect 96636 50934 96638 50986
rect 96638 50934 96690 50986
rect 96690 50934 96692 50986
rect 96636 50932 96692 50934
rect 96740 50986 96796 50988
rect 96740 50934 96742 50986
rect 96742 50934 96794 50986
rect 96794 50934 96796 50986
rect 96740 50932 96796 50934
rect 96844 50986 96900 50988
rect 96844 50934 96846 50986
rect 96846 50934 96898 50986
rect 96898 50934 96900 50986
rect 96844 50932 96900 50934
rect 96636 49418 96692 49420
rect 96636 49366 96638 49418
rect 96638 49366 96690 49418
rect 96690 49366 96692 49418
rect 96636 49364 96692 49366
rect 96740 49418 96796 49420
rect 96740 49366 96742 49418
rect 96742 49366 96794 49418
rect 96794 49366 96796 49418
rect 96740 49364 96796 49366
rect 96844 49418 96900 49420
rect 96844 49366 96846 49418
rect 96846 49366 96898 49418
rect 96898 49366 96900 49418
rect 96844 49364 96900 49366
rect 96636 47850 96692 47852
rect 96636 47798 96638 47850
rect 96638 47798 96690 47850
rect 96690 47798 96692 47850
rect 96636 47796 96692 47798
rect 96740 47850 96796 47852
rect 96740 47798 96742 47850
rect 96742 47798 96794 47850
rect 96794 47798 96796 47850
rect 96740 47796 96796 47798
rect 96844 47850 96900 47852
rect 96844 47798 96846 47850
rect 96846 47798 96898 47850
rect 96898 47798 96900 47850
rect 96844 47796 96900 47798
rect 96636 46282 96692 46284
rect 96636 46230 96638 46282
rect 96638 46230 96690 46282
rect 96690 46230 96692 46282
rect 96636 46228 96692 46230
rect 96740 46282 96796 46284
rect 96740 46230 96742 46282
rect 96742 46230 96794 46282
rect 96794 46230 96796 46282
rect 96740 46228 96796 46230
rect 96844 46282 96900 46284
rect 96844 46230 96846 46282
rect 96846 46230 96898 46282
rect 96898 46230 96900 46282
rect 96844 46228 96900 46230
rect 96636 44714 96692 44716
rect 96636 44662 96638 44714
rect 96638 44662 96690 44714
rect 96690 44662 96692 44714
rect 96636 44660 96692 44662
rect 96740 44714 96796 44716
rect 96740 44662 96742 44714
rect 96742 44662 96794 44714
rect 96794 44662 96796 44714
rect 96740 44660 96796 44662
rect 96844 44714 96900 44716
rect 96844 44662 96846 44714
rect 96846 44662 96898 44714
rect 96898 44662 96900 44714
rect 96844 44660 96900 44662
rect 96636 43146 96692 43148
rect 96636 43094 96638 43146
rect 96638 43094 96690 43146
rect 96690 43094 96692 43146
rect 96636 43092 96692 43094
rect 96740 43146 96796 43148
rect 96740 43094 96742 43146
rect 96742 43094 96794 43146
rect 96794 43094 96796 43146
rect 96740 43092 96796 43094
rect 96844 43146 96900 43148
rect 96844 43094 96846 43146
rect 96846 43094 96898 43146
rect 96898 43094 96900 43146
rect 96844 43092 96900 43094
rect 96636 41578 96692 41580
rect 96636 41526 96638 41578
rect 96638 41526 96690 41578
rect 96690 41526 96692 41578
rect 96636 41524 96692 41526
rect 96740 41578 96796 41580
rect 96740 41526 96742 41578
rect 96742 41526 96794 41578
rect 96794 41526 96796 41578
rect 96740 41524 96796 41526
rect 96844 41578 96900 41580
rect 96844 41526 96846 41578
rect 96846 41526 96898 41578
rect 96898 41526 96900 41578
rect 96844 41524 96900 41526
rect 96636 40010 96692 40012
rect 96636 39958 96638 40010
rect 96638 39958 96690 40010
rect 96690 39958 96692 40010
rect 96636 39956 96692 39958
rect 96740 40010 96796 40012
rect 96740 39958 96742 40010
rect 96742 39958 96794 40010
rect 96794 39958 96796 40010
rect 96740 39956 96796 39958
rect 96844 40010 96900 40012
rect 96844 39958 96846 40010
rect 96846 39958 96898 40010
rect 96898 39958 96900 40010
rect 96844 39956 96900 39958
rect 96636 38442 96692 38444
rect 96636 38390 96638 38442
rect 96638 38390 96690 38442
rect 96690 38390 96692 38442
rect 96636 38388 96692 38390
rect 96740 38442 96796 38444
rect 96740 38390 96742 38442
rect 96742 38390 96794 38442
rect 96794 38390 96796 38442
rect 96740 38388 96796 38390
rect 96844 38442 96900 38444
rect 96844 38390 96846 38442
rect 96846 38390 96898 38442
rect 96898 38390 96900 38442
rect 96844 38388 96900 38390
rect 96636 36874 96692 36876
rect 96636 36822 96638 36874
rect 96638 36822 96690 36874
rect 96690 36822 96692 36874
rect 96636 36820 96692 36822
rect 96740 36874 96796 36876
rect 96740 36822 96742 36874
rect 96742 36822 96794 36874
rect 96794 36822 96796 36874
rect 96740 36820 96796 36822
rect 96844 36874 96900 36876
rect 96844 36822 96846 36874
rect 96846 36822 96898 36874
rect 96898 36822 96900 36874
rect 96844 36820 96900 36822
rect 96636 35306 96692 35308
rect 96636 35254 96638 35306
rect 96638 35254 96690 35306
rect 96690 35254 96692 35306
rect 96636 35252 96692 35254
rect 96740 35306 96796 35308
rect 96740 35254 96742 35306
rect 96742 35254 96794 35306
rect 96794 35254 96796 35306
rect 96740 35252 96796 35254
rect 96844 35306 96900 35308
rect 96844 35254 96846 35306
rect 96846 35254 96898 35306
rect 96898 35254 96900 35306
rect 96844 35252 96900 35254
rect 96636 33738 96692 33740
rect 96636 33686 96638 33738
rect 96638 33686 96690 33738
rect 96690 33686 96692 33738
rect 96636 33684 96692 33686
rect 96740 33738 96796 33740
rect 96740 33686 96742 33738
rect 96742 33686 96794 33738
rect 96794 33686 96796 33738
rect 96740 33684 96796 33686
rect 96844 33738 96900 33740
rect 96844 33686 96846 33738
rect 96846 33686 96898 33738
rect 96898 33686 96900 33738
rect 96844 33684 96900 33686
rect 96636 32170 96692 32172
rect 96636 32118 96638 32170
rect 96638 32118 96690 32170
rect 96690 32118 96692 32170
rect 96636 32116 96692 32118
rect 96740 32170 96796 32172
rect 96740 32118 96742 32170
rect 96742 32118 96794 32170
rect 96794 32118 96796 32170
rect 96740 32116 96796 32118
rect 96844 32170 96900 32172
rect 96844 32118 96846 32170
rect 96846 32118 96898 32170
rect 96898 32118 96900 32170
rect 96844 32116 96900 32118
rect 96636 30602 96692 30604
rect 96636 30550 96638 30602
rect 96638 30550 96690 30602
rect 96690 30550 96692 30602
rect 96636 30548 96692 30550
rect 96740 30602 96796 30604
rect 96740 30550 96742 30602
rect 96742 30550 96794 30602
rect 96794 30550 96796 30602
rect 96740 30548 96796 30550
rect 96844 30602 96900 30604
rect 96844 30550 96846 30602
rect 96846 30550 96898 30602
rect 96898 30550 96900 30602
rect 96844 30548 96900 30550
rect 96636 29034 96692 29036
rect 96636 28982 96638 29034
rect 96638 28982 96690 29034
rect 96690 28982 96692 29034
rect 96636 28980 96692 28982
rect 96740 29034 96796 29036
rect 96740 28982 96742 29034
rect 96742 28982 96794 29034
rect 96794 28982 96796 29034
rect 96740 28980 96796 28982
rect 96844 29034 96900 29036
rect 96844 28982 96846 29034
rect 96846 28982 96898 29034
rect 96898 28982 96900 29034
rect 96844 28980 96900 28982
rect 96636 27466 96692 27468
rect 96636 27414 96638 27466
rect 96638 27414 96690 27466
rect 96690 27414 96692 27466
rect 96636 27412 96692 27414
rect 96740 27466 96796 27468
rect 96740 27414 96742 27466
rect 96742 27414 96794 27466
rect 96794 27414 96796 27466
rect 96740 27412 96796 27414
rect 96844 27466 96900 27468
rect 96844 27414 96846 27466
rect 96846 27414 96898 27466
rect 96898 27414 96900 27466
rect 96844 27412 96900 27414
rect 96636 25898 96692 25900
rect 96636 25846 96638 25898
rect 96638 25846 96690 25898
rect 96690 25846 96692 25898
rect 96636 25844 96692 25846
rect 96740 25898 96796 25900
rect 96740 25846 96742 25898
rect 96742 25846 96794 25898
rect 96794 25846 96796 25898
rect 96740 25844 96796 25846
rect 96844 25898 96900 25900
rect 96844 25846 96846 25898
rect 96846 25846 96898 25898
rect 96898 25846 96900 25898
rect 96844 25844 96900 25846
rect 103964 55186 104020 55188
rect 103964 55134 103966 55186
rect 103966 55134 104018 55186
rect 104018 55134 104020 55186
rect 103964 55132 104020 55134
rect 107100 32732 107156 32788
rect 105756 27692 105812 27748
rect 108332 29372 108388 29428
rect 108668 28588 108724 28644
rect 104524 26178 104580 26180
rect 104524 26126 104526 26178
rect 104526 26126 104578 26178
rect 104578 26126 104580 26178
rect 104524 26124 104580 26126
rect 100492 25506 100548 25508
rect 100492 25454 100494 25506
rect 100494 25454 100546 25506
rect 100546 25454 100548 25506
rect 100492 25452 100548 25454
rect 100940 25506 100996 25508
rect 100940 25454 100942 25506
rect 100942 25454 100994 25506
rect 100994 25454 100996 25506
rect 100940 25452 100996 25454
rect 104076 25676 104132 25732
rect 96636 24330 96692 24332
rect 96636 24278 96638 24330
rect 96638 24278 96690 24330
rect 96690 24278 96692 24330
rect 96636 24276 96692 24278
rect 96740 24330 96796 24332
rect 96740 24278 96742 24330
rect 96742 24278 96794 24330
rect 96794 24278 96796 24330
rect 96740 24276 96796 24278
rect 96844 24330 96900 24332
rect 96844 24278 96846 24330
rect 96846 24278 96898 24330
rect 96898 24278 96900 24330
rect 96844 24276 96900 24278
rect 97468 23212 97524 23268
rect 95340 22988 95396 23044
rect 97132 22876 97188 22932
rect 96636 22762 96692 22764
rect 96636 22710 96638 22762
rect 96638 22710 96690 22762
rect 96690 22710 96692 22762
rect 96636 22708 96692 22710
rect 96740 22762 96796 22764
rect 96740 22710 96742 22762
rect 96742 22710 96794 22762
rect 96794 22710 96796 22762
rect 96740 22708 96796 22710
rect 96844 22762 96900 22764
rect 96844 22710 96846 22762
rect 96846 22710 96898 22762
rect 96898 22710 96900 22762
rect 96844 22708 96900 22710
rect 95228 21868 95284 21924
rect 95004 21196 95060 21252
rect 94668 18508 94724 18564
rect 94332 16156 94388 16212
rect 94780 18172 94836 18228
rect 94892 18284 94948 18340
rect 95788 20860 95844 20916
rect 95564 20524 95620 20580
rect 96636 21194 96692 21196
rect 96636 21142 96638 21194
rect 96638 21142 96690 21194
rect 96690 21142 96692 21194
rect 96636 21140 96692 21142
rect 96740 21194 96796 21196
rect 96740 21142 96742 21194
rect 96742 21142 96794 21194
rect 96794 21142 96796 21194
rect 96740 21140 96796 21142
rect 96844 21194 96900 21196
rect 96844 21142 96846 21194
rect 96846 21142 96898 21194
rect 96898 21142 96900 21194
rect 96844 21140 96900 21142
rect 96460 20524 96516 20580
rect 96684 20860 96740 20916
rect 95228 19964 95284 20020
rect 95788 20188 95844 20244
rect 95788 20018 95844 20020
rect 95788 19966 95790 20018
rect 95790 19966 95842 20018
rect 95842 19966 95844 20018
rect 95788 19964 95844 19966
rect 96796 20188 96852 20244
rect 95228 19346 95284 19348
rect 95228 19294 95230 19346
rect 95230 19294 95282 19346
rect 95282 19294 95284 19346
rect 95228 19292 95284 19294
rect 97020 20018 97076 20020
rect 97020 19966 97022 20018
rect 97022 19966 97074 20018
rect 97074 19966 97076 20018
rect 97020 19964 97076 19966
rect 100828 22876 100884 22932
rect 97468 21698 97524 21700
rect 97468 21646 97470 21698
rect 97470 21646 97522 21698
rect 97522 21646 97524 21698
rect 97468 21644 97524 21646
rect 97692 20860 97748 20916
rect 97916 20412 97972 20468
rect 96796 19740 96852 19796
rect 96636 19626 96692 19628
rect 96636 19574 96638 19626
rect 96638 19574 96690 19626
rect 96690 19574 96692 19626
rect 96636 19572 96692 19574
rect 96740 19626 96796 19628
rect 96740 19574 96742 19626
rect 96742 19574 96794 19626
rect 96794 19574 96796 19626
rect 96740 19572 96796 19574
rect 96844 19626 96900 19628
rect 96844 19574 96846 19626
rect 96846 19574 96898 19626
rect 96898 19574 96900 19626
rect 96844 19572 96900 19574
rect 96012 19292 96068 19348
rect 96684 19010 96740 19012
rect 96684 18958 96686 19010
rect 96686 18958 96738 19010
rect 96738 18958 96740 19010
rect 96684 18956 96740 18958
rect 96012 18732 96068 18788
rect 95340 18450 95396 18452
rect 95340 18398 95342 18450
rect 95342 18398 95394 18450
rect 95394 18398 95396 18450
rect 95340 18396 95396 18398
rect 95900 18338 95956 18340
rect 95900 18286 95902 18338
rect 95902 18286 95954 18338
rect 95954 18286 95956 18338
rect 95900 18284 95956 18286
rect 95004 16716 95060 16772
rect 95340 17276 95396 17332
rect 96124 18450 96180 18452
rect 96124 18398 96126 18450
rect 96126 18398 96178 18450
rect 96178 18398 96180 18450
rect 96124 18396 96180 18398
rect 96908 18396 96964 18452
rect 96684 18172 96740 18228
rect 96636 18058 96692 18060
rect 96636 18006 96638 18058
rect 96638 18006 96690 18058
rect 96690 18006 96692 18058
rect 96636 18004 96692 18006
rect 96740 18058 96796 18060
rect 96740 18006 96742 18058
rect 96742 18006 96794 18058
rect 96794 18006 96796 18058
rect 96740 18004 96796 18006
rect 96844 18058 96900 18060
rect 96844 18006 96846 18058
rect 96846 18006 96898 18058
rect 96898 18006 96900 18058
rect 96844 18004 96900 18006
rect 97244 18844 97300 18900
rect 97468 20018 97524 20020
rect 97468 19966 97470 20018
rect 97470 19966 97522 20018
rect 97522 19966 97524 20018
rect 97468 19964 97524 19966
rect 97356 18956 97412 19012
rect 96124 17724 96180 17780
rect 97244 18396 97300 18452
rect 98140 21698 98196 21700
rect 98140 21646 98142 21698
rect 98142 21646 98194 21698
rect 98194 21646 98196 21698
rect 98140 21644 98196 21646
rect 98028 20076 98084 20132
rect 99148 20578 99204 20580
rect 99148 20526 99150 20578
rect 99150 20526 99202 20578
rect 99202 20526 99204 20578
rect 99148 20524 99204 20526
rect 98700 20412 98756 20468
rect 97804 18844 97860 18900
rect 98252 19010 98308 19012
rect 98252 18958 98254 19010
rect 98254 18958 98306 19010
rect 98306 18958 98308 19010
rect 98252 18956 98308 18958
rect 99260 19068 99316 19124
rect 98812 19010 98868 19012
rect 98812 18958 98814 19010
rect 98814 18958 98866 19010
rect 98866 18958 98868 19010
rect 98812 18956 98868 18958
rect 98924 18396 98980 18452
rect 97244 16940 97300 16996
rect 97020 16716 97076 16772
rect 97468 16770 97524 16772
rect 97468 16718 97470 16770
rect 97470 16718 97522 16770
rect 97522 16718 97524 16770
rect 97468 16716 97524 16718
rect 94668 14252 94724 14308
rect 94220 11676 94276 11732
rect 94332 11564 94388 11620
rect 94108 11004 94164 11060
rect 94220 11116 94276 11172
rect 94668 13522 94724 13524
rect 94668 13470 94670 13522
rect 94670 13470 94722 13522
rect 94722 13470 94724 13522
rect 94668 13468 94724 13470
rect 94556 12348 94612 12404
rect 94892 15874 94948 15876
rect 94892 15822 94894 15874
rect 94894 15822 94946 15874
rect 94946 15822 94948 15874
rect 94892 15820 94948 15822
rect 94892 15148 94948 15204
rect 95116 15202 95172 15204
rect 95116 15150 95118 15202
rect 95118 15150 95170 15202
rect 95170 15150 95172 15202
rect 95116 15148 95172 15150
rect 95452 14252 95508 14308
rect 95004 13804 95060 13860
rect 94780 12178 94836 12180
rect 94780 12126 94782 12178
rect 94782 12126 94834 12178
rect 94834 12126 94836 12178
rect 94780 12124 94836 12126
rect 94556 11564 94612 11620
rect 94668 11452 94724 11508
rect 94668 10892 94724 10948
rect 94444 10668 94500 10724
rect 94556 10780 94612 10836
rect 93996 10444 94052 10500
rect 93884 10220 93940 10276
rect 93436 9548 93492 9604
rect 93324 9154 93380 9156
rect 93324 9102 93326 9154
rect 93326 9102 93378 9154
rect 93378 9102 93380 9154
rect 93324 9100 93380 9102
rect 93212 7868 93268 7924
rect 93212 6860 93268 6916
rect 92764 6636 92820 6692
rect 92652 5964 92708 6020
rect 93100 6188 93156 6244
rect 92428 5234 92484 5236
rect 92428 5182 92430 5234
rect 92430 5182 92482 5234
rect 92482 5182 92484 5234
rect 92428 5180 92484 5182
rect 91756 4898 91812 4900
rect 91756 4846 91758 4898
rect 91758 4846 91810 4898
rect 91810 4846 91812 4898
rect 91756 4844 91812 4846
rect 92540 4284 92596 4340
rect 92316 3724 92372 3780
rect 91644 812 91700 868
rect 92764 4060 92820 4116
rect 93436 6412 93492 6468
rect 93660 8204 93716 8260
rect 93324 6076 93380 6132
rect 93548 4226 93604 4228
rect 93548 4174 93550 4226
rect 93550 4174 93602 4226
rect 93602 4174 93604 4226
rect 93548 4172 93604 4174
rect 94220 10498 94276 10500
rect 94220 10446 94222 10498
rect 94222 10446 94274 10498
rect 94274 10446 94276 10498
rect 94220 10444 94276 10446
rect 94332 10610 94388 10612
rect 94332 10558 94334 10610
rect 94334 10558 94386 10610
rect 94386 10558 94388 10610
rect 94332 10556 94388 10558
rect 94108 9548 94164 9604
rect 94108 9042 94164 9044
rect 94108 8990 94110 9042
rect 94110 8990 94162 9042
rect 94162 8990 94164 9042
rect 94108 8988 94164 8990
rect 94332 9436 94388 9492
rect 94556 9996 94612 10052
rect 94556 9548 94612 9604
rect 94108 8316 94164 8372
rect 93996 8204 94052 8260
rect 93996 7532 94052 7588
rect 93884 6636 93940 6692
rect 94220 7196 94276 7252
rect 93884 4396 93940 4452
rect 93884 4060 93940 4116
rect 94220 6130 94276 6132
rect 94220 6078 94222 6130
rect 94222 6078 94274 6130
rect 94274 6078 94276 6130
rect 94220 6076 94276 6078
rect 94220 5852 94276 5908
rect 94108 3948 94164 4004
rect 94108 3500 94164 3556
rect 94108 1484 94164 1540
rect 95228 13634 95284 13636
rect 95228 13582 95230 13634
rect 95230 13582 95282 13634
rect 95282 13582 95284 13634
rect 95228 13580 95284 13582
rect 95228 12066 95284 12068
rect 95228 12014 95230 12066
rect 95230 12014 95282 12066
rect 95282 12014 95284 12066
rect 95228 12012 95284 12014
rect 95340 11676 95396 11732
rect 95228 11506 95284 11508
rect 95228 11454 95230 11506
rect 95230 11454 95282 11506
rect 95282 11454 95284 11506
rect 95228 11452 95284 11454
rect 95116 9996 95172 10052
rect 95340 10780 95396 10836
rect 95228 9826 95284 9828
rect 95228 9774 95230 9826
rect 95230 9774 95282 9826
rect 95282 9774 95284 9826
rect 95228 9772 95284 9774
rect 95228 9548 95284 9604
rect 94556 8764 94612 8820
rect 94892 9100 94948 9156
rect 94556 7756 94612 7812
rect 94668 8092 94724 8148
rect 94780 8034 94836 8036
rect 94780 7982 94782 8034
rect 94782 7982 94834 8034
rect 94834 7982 94836 8034
rect 94780 7980 94836 7982
rect 95228 8876 95284 8932
rect 94556 7532 94612 7588
rect 94556 6300 94612 6356
rect 94668 6636 94724 6692
rect 94556 4450 94612 4452
rect 94556 4398 94558 4450
rect 94558 4398 94610 4450
rect 94610 4398 94612 4450
rect 94556 4396 94612 4398
rect 95004 7474 95060 7476
rect 95004 7422 95006 7474
rect 95006 7422 95058 7474
rect 95058 7422 95060 7474
rect 95004 7420 95060 7422
rect 94892 7308 94948 7364
rect 94892 6466 94948 6468
rect 94892 6414 94894 6466
rect 94894 6414 94946 6466
rect 94946 6414 94948 6466
rect 94892 6412 94948 6414
rect 95228 6412 95284 6468
rect 95228 6130 95284 6132
rect 95228 6078 95230 6130
rect 95230 6078 95282 6130
rect 95282 6078 95284 6130
rect 95228 6076 95284 6078
rect 95116 6018 95172 6020
rect 95116 5966 95118 6018
rect 95118 5966 95170 6018
rect 95170 5966 95172 6018
rect 95116 5964 95172 5966
rect 95004 5852 95060 5908
rect 95004 5068 95060 5124
rect 95564 12236 95620 12292
rect 96636 16490 96692 16492
rect 96636 16438 96638 16490
rect 96638 16438 96690 16490
rect 96690 16438 96692 16490
rect 96636 16436 96692 16438
rect 96740 16490 96796 16492
rect 96740 16438 96742 16490
rect 96742 16438 96794 16490
rect 96794 16438 96796 16490
rect 96740 16436 96796 16438
rect 96844 16490 96900 16492
rect 96844 16438 96846 16490
rect 96846 16438 96898 16490
rect 96898 16438 96900 16490
rect 96844 16436 96900 16438
rect 97244 16492 97300 16548
rect 96012 15596 96068 15652
rect 95788 12124 95844 12180
rect 95900 15202 95956 15204
rect 95900 15150 95902 15202
rect 95902 15150 95954 15202
rect 95954 15150 95956 15202
rect 95900 15148 95956 15150
rect 96636 14922 96692 14924
rect 96636 14870 96638 14922
rect 96638 14870 96690 14922
rect 96690 14870 96692 14922
rect 96636 14868 96692 14870
rect 96740 14922 96796 14924
rect 96740 14870 96742 14922
rect 96742 14870 96794 14922
rect 96794 14870 96796 14922
rect 96740 14868 96796 14870
rect 96844 14922 96900 14924
rect 96844 14870 96846 14922
rect 96846 14870 96898 14922
rect 96898 14870 96900 14922
rect 96844 14868 96900 14870
rect 97132 14588 97188 14644
rect 96124 13916 96180 13972
rect 96012 13746 96068 13748
rect 96012 13694 96014 13746
rect 96014 13694 96066 13746
rect 96066 13694 96068 13746
rect 96012 13692 96068 13694
rect 96348 13356 96404 13412
rect 96348 12962 96404 12964
rect 96348 12910 96350 12962
rect 96350 12910 96402 12962
rect 96402 12910 96404 12962
rect 96348 12908 96404 12910
rect 96124 11900 96180 11956
rect 96636 13354 96692 13356
rect 96636 13302 96638 13354
rect 96638 13302 96690 13354
rect 96690 13302 96692 13354
rect 96636 13300 96692 13302
rect 96740 13354 96796 13356
rect 96740 13302 96742 13354
rect 96742 13302 96794 13354
rect 96794 13302 96796 13354
rect 96740 13300 96796 13302
rect 96844 13354 96900 13356
rect 96844 13302 96846 13354
rect 96846 13302 96898 13354
rect 96898 13302 96900 13354
rect 96844 13300 96900 13302
rect 96636 11786 96692 11788
rect 96636 11734 96638 11786
rect 96638 11734 96690 11786
rect 96690 11734 96692 11786
rect 96636 11732 96692 11734
rect 96740 11786 96796 11788
rect 96740 11734 96742 11786
rect 96742 11734 96794 11786
rect 96794 11734 96796 11786
rect 96740 11732 96796 11734
rect 96844 11786 96900 11788
rect 96844 11734 96846 11786
rect 96846 11734 96898 11786
rect 96898 11734 96900 11786
rect 96844 11732 96900 11734
rect 95788 11452 95844 11508
rect 95564 9996 95620 10052
rect 96012 9436 96068 9492
rect 95900 9100 95956 9156
rect 95900 8818 95956 8820
rect 95900 8766 95902 8818
rect 95902 8766 95954 8818
rect 95954 8766 95956 8818
rect 95900 8764 95956 8766
rect 95676 8428 95732 8484
rect 95676 8204 95732 8260
rect 95788 7980 95844 8036
rect 95452 7532 95508 7588
rect 95788 7644 95844 7700
rect 96348 11170 96404 11172
rect 96348 11118 96350 11170
rect 96350 11118 96402 11170
rect 96402 11118 96404 11170
rect 96348 11116 96404 11118
rect 96796 10780 96852 10836
rect 97580 16156 97636 16212
rect 97468 14306 97524 14308
rect 97468 14254 97470 14306
rect 97470 14254 97522 14306
rect 97522 14254 97524 14306
rect 97468 14252 97524 14254
rect 98700 17442 98756 17444
rect 98700 17390 98702 17442
rect 98702 17390 98754 17442
rect 98754 17390 98756 17442
rect 98700 17388 98756 17390
rect 98252 17276 98308 17332
rect 97916 17164 97972 17220
rect 98252 16994 98308 16996
rect 98252 16942 98254 16994
rect 98254 16942 98306 16994
rect 98306 16942 98308 16994
rect 98252 16940 98308 16942
rect 97916 15932 97972 15988
rect 97804 14476 97860 14532
rect 98252 14700 98308 14756
rect 97804 13746 97860 13748
rect 97804 13694 97806 13746
rect 97806 13694 97858 13746
rect 97858 13694 97860 13746
rect 97804 13692 97860 13694
rect 97356 13186 97412 13188
rect 97356 13134 97358 13186
rect 97358 13134 97410 13186
rect 97410 13134 97412 13186
rect 97356 13132 97412 13134
rect 97804 12908 97860 12964
rect 96908 10444 96964 10500
rect 97020 11116 97076 11172
rect 96636 10218 96692 10220
rect 96636 10166 96638 10218
rect 96638 10166 96690 10218
rect 96690 10166 96692 10218
rect 96636 10164 96692 10166
rect 96740 10218 96796 10220
rect 96740 10166 96742 10218
rect 96742 10166 96794 10218
rect 96794 10166 96796 10218
rect 96740 10164 96796 10166
rect 96844 10218 96900 10220
rect 96844 10166 96846 10218
rect 96846 10166 96898 10218
rect 96898 10166 96900 10218
rect 96844 10164 96900 10166
rect 96124 8316 96180 8372
rect 96236 9772 96292 9828
rect 96460 9996 96516 10052
rect 97020 9996 97076 10052
rect 96684 9436 96740 9492
rect 96348 9154 96404 9156
rect 96348 9102 96350 9154
rect 96350 9102 96402 9154
rect 96402 9102 96404 9154
rect 96348 9100 96404 9102
rect 96572 8764 96628 8820
rect 96636 8650 96692 8652
rect 96636 8598 96638 8650
rect 96638 8598 96690 8650
rect 96690 8598 96692 8650
rect 96636 8596 96692 8598
rect 96740 8650 96796 8652
rect 96740 8598 96742 8650
rect 96742 8598 96794 8650
rect 96794 8598 96796 8650
rect 96740 8596 96796 8598
rect 96844 8650 96900 8652
rect 96844 8598 96846 8650
rect 96846 8598 96898 8650
rect 96898 8598 96900 8650
rect 96844 8596 96900 8598
rect 96572 7196 96628 7252
rect 97020 7756 97076 7812
rect 96636 7082 96692 7084
rect 96636 7030 96638 7082
rect 96638 7030 96690 7082
rect 96690 7030 96692 7082
rect 96636 7028 96692 7030
rect 96740 7082 96796 7084
rect 96740 7030 96742 7082
rect 96742 7030 96794 7082
rect 96794 7030 96796 7082
rect 96740 7028 96796 7030
rect 96844 7082 96900 7084
rect 96844 7030 96846 7082
rect 96846 7030 96898 7082
rect 96898 7030 96900 7082
rect 96844 7028 96900 7030
rect 95564 5852 95620 5908
rect 95564 5122 95620 5124
rect 95564 5070 95566 5122
rect 95566 5070 95618 5122
rect 95618 5070 95620 5122
rect 95564 5068 95620 5070
rect 96236 6300 96292 6356
rect 96012 4956 96068 5012
rect 95340 4732 95396 4788
rect 96636 5514 96692 5516
rect 96636 5462 96638 5514
rect 96638 5462 96690 5514
rect 96690 5462 96692 5514
rect 96636 5460 96692 5462
rect 96740 5514 96796 5516
rect 96740 5462 96742 5514
rect 96742 5462 96794 5514
rect 96794 5462 96796 5514
rect 96740 5460 96796 5462
rect 96844 5514 96900 5516
rect 96844 5462 96846 5514
rect 96846 5462 96898 5514
rect 96898 5462 96900 5514
rect 96844 5460 96900 5462
rect 96124 4732 96180 4788
rect 96236 4844 96292 4900
rect 96236 4284 96292 4340
rect 96012 4114 96068 4116
rect 96012 4062 96014 4114
rect 96014 4062 96066 4114
rect 96066 4062 96068 4114
rect 96012 4060 96068 4062
rect 96636 3946 96692 3948
rect 96636 3894 96638 3946
rect 96638 3894 96690 3946
rect 96690 3894 96692 3946
rect 96636 3892 96692 3894
rect 96740 3946 96796 3948
rect 96740 3894 96742 3946
rect 96742 3894 96794 3946
rect 96794 3894 96796 3946
rect 96740 3892 96796 3894
rect 96844 3946 96900 3948
rect 96844 3894 96846 3946
rect 96846 3894 96898 3946
rect 96898 3894 96900 3946
rect 96844 3892 96900 3894
rect 97020 3836 97076 3892
rect 96908 3612 96964 3668
rect 94780 1372 94836 1428
rect 96572 3388 96628 3444
rect 94444 1260 94500 1316
rect 97244 10444 97300 10500
rect 97244 9660 97300 9716
rect 97356 9548 97412 9604
rect 97804 11788 97860 11844
rect 97916 11676 97972 11732
rect 97916 11452 97972 11508
rect 97580 9660 97636 9716
rect 97692 9324 97748 9380
rect 97804 10332 97860 10388
rect 97580 9212 97636 9268
rect 97468 8428 97524 8484
rect 97244 6412 97300 6468
rect 97916 9548 97972 9604
rect 97916 8316 97972 8372
rect 97916 7756 97972 7812
rect 98252 13692 98308 13748
rect 99708 18732 99764 18788
rect 99484 18284 99540 18340
rect 98588 16492 98644 16548
rect 98140 12236 98196 12292
rect 98812 16210 98868 16212
rect 98812 16158 98814 16210
rect 98814 16158 98866 16210
rect 98866 16158 98868 16210
rect 98812 16156 98868 16158
rect 98812 15090 98868 15092
rect 98812 15038 98814 15090
rect 98814 15038 98866 15090
rect 98866 15038 98868 15090
rect 98812 15036 98868 15038
rect 98364 11676 98420 11732
rect 98476 11564 98532 11620
rect 98252 11004 98308 11060
rect 98252 10220 98308 10276
rect 98252 9212 98308 9268
rect 98140 8876 98196 8932
rect 97916 6076 97972 6132
rect 97804 5516 97860 5572
rect 97244 5404 97300 5460
rect 98924 14476 98980 14532
rect 98812 13522 98868 13524
rect 98812 13470 98814 13522
rect 98814 13470 98866 13522
rect 98866 13470 98868 13522
rect 98812 13468 98868 13470
rect 98812 13244 98868 13300
rect 98812 12124 98868 12180
rect 98812 11954 98868 11956
rect 98812 11902 98814 11954
rect 98814 11902 98866 11954
rect 98866 11902 98868 11954
rect 98812 11900 98868 11902
rect 99708 18284 99764 18340
rect 101276 20524 101332 20580
rect 100828 20076 100884 20132
rect 103964 21474 104020 21476
rect 103964 21422 103966 21474
rect 103966 21422 104018 21474
rect 104018 21422 104020 21474
rect 103964 21420 104020 21422
rect 103292 20578 103348 20580
rect 103292 20526 103294 20578
rect 103294 20526 103346 20578
rect 103346 20526 103348 20578
rect 103292 20524 103348 20526
rect 103068 20188 103124 20244
rect 99932 19122 99988 19124
rect 99932 19070 99934 19122
rect 99934 19070 99986 19122
rect 99986 19070 99988 19122
rect 99932 19068 99988 19070
rect 104188 20188 104244 20244
rect 104972 26124 105028 26180
rect 105532 26124 105588 26180
rect 105980 26124 106036 26180
rect 106092 25506 106148 25508
rect 106092 25454 106094 25506
rect 106094 25454 106146 25506
rect 106146 25454 106148 25506
rect 106092 25452 106148 25454
rect 106540 25506 106596 25508
rect 106540 25454 106542 25506
rect 106542 25454 106594 25506
rect 106594 25454 106596 25506
rect 106540 25452 106596 25454
rect 105420 21420 105476 21476
rect 104076 19068 104132 19124
rect 99820 18396 99876 18452
rect 100044 18284 100100 18340
rect 99820 17106 99876 17108
rect 99820 17054 99822 17106
rect 99822 17054 99874 17106
rect 99874 17054 99876 17106
rect 99820 17052 99876 17054
rect 100044 17052 100100 17108
rect 100044 16716 100100 16772
rect 100828 18956 100884 19012
rect 100380 18396 100436 18452
rect 101948 18450 102004 18452
rect 101948 18398 101950 18450
rect 101950 18398 102002 18450
rect 102002 18398 102004 18450
rect 101948 18396 102004 18398
rect 101724 18284 101780 18340
rect 101724 17388 101780 17444
rect 99260 14476 99316 14532
rect 100380 16882 100436 16884
rect 100380 16830 100382 16882
rect 100382 16830 100434 16882
rect 100434 16830 100436 16882
rect 100380 16828 100436 16830
rect 99148 11564 99204 11620
rect 99372 13692 99428 13748
rect 100492 16716 100548 16772
rect 100380 15596 100436 15652
rect 100156 14700 100212 14756
rect 100044 14588 100100 14644
rect 99932 14476 99988 14532
rect 99596 13244 99652 13300
rect 99708 12908 99764 12964
rect 99820 11170 99876 11172
rect 99820 11118 99822 11170
rect 99822 11118 99874 11170
rect 99874 11118 99876 11170
rect 99820 11116 99876 11118
rect 99036 10556 99092 10612
rect 99148 9996 99204 10052
rect 99036 9714 99092 9716
rect 99036 9662 99038 9714
rect 99038 9662 99090 9714
rect 99090 9662 99092 9714
rect 99036 9660 99092 9662
rect 99148 9324 99204 9380
rect 99036 8988 99092 9044
rect 98364 8316 98420 8372
rect 98476 8764 98532 8820
rect 98364 8146 98420 8148
rect 98364 8094 98366 8146
rect 98366 8094 98418 8146
rect 98418 8094 98420 8146
rect 98364 8092 98420 8094
rect 98252 5068 98308 5124
rect 97244 4732 97300 4788
rect 98700 8652 98756 8708
rect 99148 8258 99204 8260
rect 99148 8206 99150 8258
rect 99150 8206 99202 8258
rect 99202 8206 99204 8258
rect 99148 8204 99204 8206
rect 98700 5346 98756 5348
rect 98700 5294 98702 5346
rect 98702 5294 98754 5346
rect 98754 5294 98756 5346
rect 98700 5292 98756 5294
rect 98924 5122 98980 5124
rect 98924 5070 98926 5122
rect 98926 5070 98978 5122
rect 98978 5070 98980 5122
rect 98924 5068 98980 5070
rect 99036 5010 99092 5012
rect 99036 4958 99038 5010
rect 99038 4958 99090 5010
rect 99090 4958 99092 5010
rect 99036 4956 99092 4958
rect 99036 4450 99092 4452
rect 99036 4398 99038 4450
rect 99038 4398 99090 4450
rect 99090 4398 99092 4450
rect 99036 4396 99092 4398
rect 97132 2492 97188 2548
rect 99036 3388 99092 3444
rect 99820 10780 99876 10836
rect 99820 10444 99876 10500
rect 99708 9324 99764 9380
rect 99708 6860 99764 6916
rect 101388 17164 101444 17220
rect 100828 16882 100884 16884
rect 100828 16830 100830 16882
rect 100830 16830 100882 16882
rect 100882 16830 100884 16882
rect 100828 16828 100884 16830
rect 101052 16716 101108 16772
rect 100828 15596 100884 15652
rect 100492 15484 100548 15540
rect 100044 14028 100100 14084
rect 100268 13746 100324 13748
rect 100268 13694 100270 13746
rect 100270 13694 100322 13746
rect 100322 13694 100324 13746
rect 100268 13692 100324 13694
rect 100156 12908 100212 12964
rect 100268 12850 100324 12852
rect 100268 12798 100270 12850
rect 100270 12798 100322 12850
rect 100322 12798 100324 12850
rect 100268 12796 100324 12798
rect 100044 11900 100100 11956
rect 100156 12012 100212 12068
rect 100828 12962 100884 12964
rect 100828 12910 100830 12962
rect 100830 12910 100882 12962
rect 100882 12910 100884 12962
rect 100828 12908 100884 12910
rect 101052 15932 101108 15988
rect 101500 16268 101556 16324
rect 101724 17052 101780 17108
rect 102508 18450 102564 18452
rect 102508 18398 102510 18450
rect 102510 18398 102562 18450
rect 102562 18398 102564 18450
rect 102508 18396 102564 18398
rect 105196 20018 105252 20020
rect 105196 19966 105198 20018
rect 105198 19966 105250 20018
rect 105250 19966 105252 20018
rect 105196 19964 105252 19966
rect 104972 19292 105028 19348
rect 106988 25394 107044 25396
rect 106988 25342 106990 25394
rect 106990 25342 107042 25394
rect 107042 25342 107044 25394
rect 106988 25340 107044 25342
rect 107324 25340 107380 25396
rect 105756 20188 105812 20244
rect 104972 19122 105028 19124
rect 104972 19070 104974 19122
rect 104974 19070 105026 19122
rect 105026 19070 105028 19122
rect 104972 19068 105028 19070
rect 104636 18396 104692 18452
rect 105868 20130 105924 20132
rect 105868 20078 105870 20130
rect 105870 20078 105922 20130
rect 105922 20078 105924 20130
rect 105868 20076 105924 20078
rect 105980 20018 106036 20020
rect 105980 19966 105982 20018
rect 105982 19966 106034 20018
rect 106034 19966 106036 20018
rect 105980 19964 106036 19966
rect 106428 20018 106484 20020
rect 106428 19966 106430 20018
rect 106430 19966 106482 20018
rect 106482 19966 106484 20018
rect 106428 19964 106484 19966
rect 105868 19292 105924 19348
rect 106652 20076 106708 20132
rect 106428 19292 106484 19348
rect 106092 19068 106148 19124
rect 106204 18396 106260 18452
rect 101948 17164 102004 17220
rect 102508 17612 102564 17668
rect 102508 17106 102564 17108
rect 102508 17054 102510 17106
rect 102510 17054 102562 17106
rect 102562 17054 102564 17106
rect 102508 17052 102564 17054
rect 104860 17388 104916 17444
rect 105420 17106 105476 17108
rect 105420 17054 105422 17106
rect 105422 17054 105474 17106
rect 105474 17054 105476 17106
rect 105420 17052 105476 17054
rect 105308 16994 105364 16996
rect 105308 16942 105310 16994
rect 105310 16942 105362 16994
rect 105362 16942 105364 16994
rect 105308 16940 105364 16942
rect 101724 15538 101780 15540
rect 101724 15486 101726 15538
rect 101726 15486 101778 15538
rect 101778 15486 101780 15538
rect 101724 15484 101780 15486
rect 103964 16828 104020 16884
rect 102508 15932 102564 15988
rect 101612 15426 101668 15428
rect 101612 15374 101614 15426
rect 101614 15374 101666 15426
rect 101666 15374 101668 15426
rect 101612 15372 101668 15374
rect 102284 15314 102340 15316
rect 102284 15262 102286 15314
rect 102286 15262 102338 15314
rect 102338 15262 102340 15314
rect 102284 15260 102340 15262
rect 101500 14700 101556 14756
rect 101388 14588 101444 14644
rect 102956 16156 103012 16212
rect 102956 14812 103012 14868
rect 103516 15036 103572 15092
rect 103628 14588 103684 14644
rect 101388 13804 101444 13860
rect 101276 12796 101332 12852
rect 100940 11564 100996 11620
rect 101276 12124 101332 12180
rect 100604 11506 100660 11508
rect 100604 11454 100606 11506
rect 100606 11454 100658 11506
rect 100658 11454 100660 11506
rect 100604 11452 100660 11454
rect 100380 10332 100436 10388
rect 100380 9212 100436 9268
rect 100268 8316 100324 8372
rect 100156 7980 100212 8036
rect 100380 8092 100436 8148
rect 100156 7532 100212 7588
rect 100044 5180 100100 5236
rect 99372 3164 99428 3220
rect 100268 7644 100324 7700
rect 100268 6802 100324 6804
rect 100268 6750 100270 6802
rect 100270 6750 100322 6802
rect 100322 6750 100324 6802
rect 100268 6748 100324 6750
rect 101164 10780 101220 10836
rect 100716 9884 100772 9940
rect 100828 8818 100884 8820
rect 100828 8766 100830 8818
rect 100830 8766 100882 8818
rect 100882 8766 100884 8818
rect 100828 8764 100884 8766
rect 100604 7980 100660 8036
rect 100716 8316 100772 8372
rect 101164 10108 101220 10164
rect 101276 10556 101332 10612
rect 102732 13746 102788 13748
rect 102732 13694 102734 13746
rect 102734 13694 102786 13746
rect 102786 13694 102788 13746
rect 102732 13692 102788 13694
rect 102508 13244 102564 13300
rect 101836 11452 101892 11508
rect 101388 7644 101444 7700
rect 101612 10556 101668 10612
rect 101500 9548 101556 9604
rect 101052 7532 101108 7588
rect 101500 7420 101556 7476
rect 101836 9938 101892 9940
rect 101836 9886 101838 9938
rect 101838 9886 101890 9938
rect 101890 9886 101892 9938
rect 101836 9884 101892 9886
rect 101724 8258 101780 8260
rect 101724 8206 101726 8258
rect 101726 8206 101778 8258
rect 101778 8206 101780 8258
rect 101724 8204 101780 8206
rect 101612 7980 101668 8036
rect 100940 6524 100996 6580
rect 100492 6412 100548 6468
rect 100156 4620 100212 4676
rect 100492 5516 100548 5572
rect 101612 5516 101668 5572
rect 101724 5292 101780 5348
rect 100716 4732 100772 4788
rect 101948 8316 102004 8372
rect 102060 6748 102116 6804
rect 102508 12348 102564 12404
rect 102844 12908 102900 12964
rect 103180 13356 103236 13412
rect 103292 14476 103348 14532
rect 103292 13132 103348 13188
rect 103516 13356 103572 13412
rect 102620 12236 102676 12292
rect 102732 11732 102788 11788
rect 102508 11116 102564 11172
rect 102396 10556 102452 10612
rect 102620 10444 102676 10500
rect 102956 11788 103012 11844
rect 102956 11340 103012 11396
rect 102844 11228 102900 11284
rect 102844 10892 102900 10948
rect 102844 10444 102900 10500
rect 102844 10108 102900 10164
rect 103628 12572 103684 12628
rect 103628 12348 103684 12404
rect 103628 11788 103684 11844
rect 103404 11228 103460 11284
rect 103068 10108 103124 10164
rect 103292 10892 103348 10948
rect 102844 9884 102900 9940
rect 103068 9826 103124 9828
rect 103068 9774 103070 9826
rect 103070 9774 103122 9826
rect 103122 9774 103124 9826
rect 103068 9772 103124 9774
rect 103068 9324 103124 9380
rect 102844 9154 102900 9156
rect 102844 9102 102846 9154
rect 102846 9102 102898 9154
rect 102898 9102 102900 9154
rect 102844 9100 102900 9102
rect 102396 8930 102452 8932
rect 102396 8878 102398 8930
rect 102398 8878 102450 8930
rect 102450 8878 102452 8930
rect 102396 8876 102452 8878
rect 102508 8652 102564 8708
rect 102844 8764 102900 8820
rect 102508 7474 102564 7476
rect 102508 7422 102510 7474
rect 102510 7422 102562 7474
rect 102562 7422 102564 7474
rect 102508 7420 102564 7422
rect 102508 6972 102564 7028
rect 102396 6690 102452 6692
rect 102396 6638 102398 6690
rect 102398 6638 102450 6690
rect 102450 6638 102452 6690
rect 102396 6636 102452 6638
rect 102732 6748 102788 6804
rect 102956 8204 103012 8260
rect 102956 7420 103012 7476
rect 103068 7644 103124 7700
rect 102844 6188 102900 6244
rect 102844 5516 102900 5572
rect 103628 10610 103684 10612
rect 103628 10558 103630 10610
rect 103630 10558 103682 10610
rect 103682 10558 103684 10610
rect 103628 10556 103684 10558
rect 103516 10444 103572 10500
rect 103292 9996 103348 10052
rect 104860 16828 104916 16884
rect 104188 16268 104244 16324
rect 103964 16044 104020 16100
rect 105644 16882 105700 16884
rect 105644 16830 105646 16882
rect 105646 16830 105698 16882
rect 105698 16830 105700 16882
rect 105644 16828 105700 16830
rect 106204 17666 106260 17668
rect 106204 17614 106206 17666
rect 106206 17614 106258 17666
rect 106258 17614 106260 17666
rect 106204 17612 106260 17614
rect 106428 17612 106484 17668
rect 107212 20018 107268 20020
rect 107212 19966 107214 20018
rect 107214 19966 107266 20018
rect 107266 19966 107268 20018
rect 107212 19964 107268 19966
rect 106988 18450 107044 18452
rect 106988 18398 106990 18450
rect 106990 18398 107042 18450
rect 107042 18398 107044 18450
rect 106988 18396 107044 18398
rect 106764 17724 106820 17780
rect 105756 16604 105812 16660
rect 104300 15372 104356 15428
rect 103964 14812 104020 14868
rect 103964 14364 104020 14420
rect 104748 15260 104804 15316
rect 104636 13858 104692 13860
rect 104636 13806 104638 13858
rect 104638 13806 104690 13858
rect 104690 13806 104692 13858
rect 104636 13804 104692 13806
rect 103964 13468 104020 13524
rect 104524 13580 104580 13636
rect 103964 12178 104020 12180
rect 103964 12126 103966 12178
rect 103966 12126 104018 12178
rect 104018 12126 104020 12178
rect 103964 12124 104020 12126
rect 103852 11116 103908 11172
rect 103964 11788 104020 11844
rect 103852 10780 103908 10836
rect 103852 10220 103908 10276
rect 104076 11340 104132 11396
rect 105644 16156 105700 16212
rect 105756 15874 105812 15876
rect 105756 15822 105758 15874
rect 105758 15822 105810 15874
rect 105810 15822 105812 15874
rect 105756 15820 105812 15822
rect 106316 15874 106372 15876
rect 106316 15822 106318 15874
rect 106318 15822 106370 15874
rect 106370 15822 106372 15874
rect 106316 15820 106372 15822
rect 106764 17554 106820 17556
rect 106764 17502 106766 17554
rect 106766 17502 106818 17554
rect 106818 17502 106820 17554
rect 106764 17500 106820 17502
rect 106540 15708 106596 15764
rect 105644 15148 105700 15204
rect 106428 15484 106484 15540
rect 105532 14700 105588 14756
rect 106092 14700 106148 14756
rect 106876 17276 106932 17332
rect 106652 15314 106708 15316
rect 106652 15262 106654 15314
rect 106654 15262 106706 15314
rect 106706 15262 106708 15314
rect 106652 15260 106708 15262
rect 106652 14306 106708 14308
rect 106652 14254 106654 14306
rect 106654 14254 106706 14306
rect 106706 14254 106708 14306
rect 106652 14252 106708 14254
rect 106652 13858 106708 13860
rect 106652 13806 106654 13858
rect 106654 13806 106706 13858
rect 106706 13806 106708 13858
rect 106652 13804 106708 13806
rect 104860 12572 104916 12628
rect 104188 9996 104244 10052
rect 104300 11116 104356 11172
rect 103964 8316 104020 8372
rect 104524 10556 104580 10612
rect 104524 10332 104580 10388
rect 105308 13132 105364 13188
rect 105308 11900 105364 11956
rect 105196 11564 105252 11620
rect 105084 11452 105140 11508
rect 105420 11452 105476 11508
rect 103964 7644 104020 7700
rect 104300 7980 104356 8036
rect 103404 6578 103460 6580
rect 103404 6526 103406 6578
rect 103406 6526 103458 6578
rect 103458 6526 103460 6578
rect 103404 6524 103460 6526
rect 103516 6412 103572 6468
rect 102172 4956 102228 5012
rect 103740 5794 103796 5796
rect 103740 5742 103742 5794
rect 103742 5742 103794 5794
rect 103794 5742 103796 5794
rect 103740 5740 103796 5742
rect 103740 5010 103796 5012
rect 103740 4958 103742 5010
rect 103742 4958 103794 5010
rect 103794 4958 103796 5010
rect 103740 4956 103796 4958
rect 103628 4844 103684 4900
rect 101948 4732 102004 4788
rect 103740 4732 103796 4788
rect 100604 3388 100660 3444
rect 102956 4226 103012 4228
rect 102956 4174 102958 4226
rect 102958 4174 103010 4226
rect 103010 4174 103012 4226
rect 102956 4172 103012 4174
rect 103292 3948 103348 4004
rect 104188 6524 104244 6580
rect 104188 4732 104244 4788
rect 104636 8540 104692 8596
rect 105308 9602 105364 9604
rect 105308 9550 105310 9602
rect 105310 9550 105362 9602
rect 105362 9550 105364 9602
rect 105308 9548 105364 9550
rect 105644 13522 105700 13524
rect 105644 13470 105646 13522
rect 105646 13470 105698 13522
rect 105698 13470 105700 13522
rect 105644 13468 105700 13470
rect 105644 12124 105700 12180
rect 106204 13580 106260 13636
rect 105980 12402 106036 12404
rect 105980 12350 105982 12402
rect 105982 12350 106034 12402
rect 106034 12350 106036 12402
rect 105980 12348 106036 12350
rect 105532 11004 105588 11060
rect 105196 8764 105252 8820
rect 104860 8204 104916 8260
rect 105196 8316 105252 8372
rect 106540 12908 106596 12964
rect 106428 12684 106484 12740
rect 106316 11564 106372 11620
rect 106092 10668 106148 10724
rect 106204 11282 106260 11284
rect 106204 11230 106206 11282
rect 106206 11230 106258 11282
rect 106258 11230 106260 11282
rect 106204 11228 106260 11230
rect 106428 11676 106484 11732
rect 106316 10780 106372 10836
rect 106204 10556 106260 10612
rect 105868 9826 105924 9828
rect 105868 9774 105870 9826
rect 105870 9774 105922 9826
rect 105922 9774 105924 9826
rect 105868 9772 105924 9774
rect 105756 9154 105812 9156
rect 105756 9102 105758 9154
rect 105758 9102 105810 9154
rect 105810 9102 105812 9154
rect 105756 9100 105812 9102
rect 105980 8988 106036 9044
rect 105644 8540 105700 8596
rect 106092 10108 106148 10164
rect 105084 7532 105140 7588
rect 104860 6972 104916 7028
rect 104860 6802 104916 6804
rect 104860 6750 104862 6802
rect 104862 6750 104914 6802
rect 104914 6750 104916 6802
rect 104860 6748 104916 6750
rect 106540 9884 106596 9940
rect 106988 15874 107044 15876
rect 106988 15822 106990 15874
rect 106990 15822 107042 15874
rect 107042 15822 107044 15874
rect 106988 15820 107044 15822
rect 106988 15372 107044 15428
rect 107660 25506 107716 25508
rect 107660 25454 107662 25506
rect 107662 25454 107714 25506
rect 107714 25454 107716 25506
rect 107660 25452 107716 25454
rect 116060 56252 116116 56308
rect 117292 56306 117348 56308
rect 117292 56254 117294 56306
rect 117294 56254 117346 56306
rect 117346 56254 117348 56306
rect 117292 56252 117348 56254
rect 119868 56252 119924 56308
rect 121100 56306 121156 56308
rect 121100 56254 121102 56306
rect 121102 56254 121154 56306
rect 121154 56254 121156 56306
rect 121100 56252 121156 56254
rect 112476 56194 112532 56196
rect 112476 56142 112478 56194
rect 112478 56142 112530 56194
rect 112530 56142 112532 56194
rect 112476 56140 112532 56142
rect 115052 56140 115108 56196
rect 111996 54906 112052 54908
rect 111996 54854 111998 54906
rect 111998 54854 112050 54906
rect 112050 54854 112052 54906
rect 111996 54852 112052 54854
rect 112100 54906 112156 54908
rect 112100 54854 112102 54906
rect 112102 54854 112154 54906
rect 112154 54854 112156 54906
rect 112100 54852 112156 54854
rect 112204 54906 112260 54908
rect 112204 54854 112206 54906
rect 112206 54854 112258 54906
rect 112258 54854 112260 54906
rect 112204 54852 112260 54854
rect 111996 53338 112052 53340
rect 111996 53286 111998 53338
rect 111998 53286 112050 53338
rect 112050 53286 112052 53338
rect 111996 53284 112052 53286
rect 112100 53338 112156 53340
rect 112100 53286 112102 53338
rect 112102 53286 112154 53338
rect 112154 53286 112156 53338
rect 112100 53284 112156 53286
rect 112204 53338 112260 53340
rect 112204 53286 112206 53338
rect 112206 53286 112258 53338
rect 112258 53286 112260 53338
rect 112204 53284 112260 53286
rect 111996 51770 112052 51772
rect 111996 51718 111998 51770
rect 111998 51718 112050 51770
rect 112050 51718 112052 51770
rect 111996 51716 112052 51718
rect 112100 51770 112156 51772
rect 112100 51718 112102 51770
rect 112102 51718 112154 51770
rect 112154 51718 112156 51770
rect 112100 51716 112156 51718
rect 112204 51770 112260 51772
rect 112204 51718 112206 51770
rect 112206 51718 112258 51770
rect 112258 51718 112260 51770
rect 112204 51716 112260 51718
rect 111996 50202 112052 50204
rect 111996 50150 111998 50202
rect 111998 50150 112050 50202
rect 112050 50150 112052 50202
rect 111996 50148 112052 50150
rect 112100 50202 112156 50204
rect 112100 50150 112102 50202
rect 112102 50150 112154 50202
rect 112154 50150 112156 50202
rect 112100 50148 112156 50150
rect 112204 50202 112260 50204
rect 112204 50150 112206 50202
rect 112206 50150 112258 50202
rect 112258 50150 112260 50202
rect 112204 50148 112260 50150
rect 111996 48634 112052 48636
rect 111996 48582 111998 48634
rect 111998 48582 112050 48634
rect 112050 48582 112052 48634
rect 111996 48580 112052 48582
rect 112100 48634 112156 48636
rect 112100 48582 112102 48634
rect 112102 48582 112154 48634
rect 112154 48582 112156 48634
rect 112100 48580 112156 48582
rect 112204 48634 112260 48636
rect 112204 48582 112206 48634
rect 112206 48582 112258 48634
rect 112258 48582 112260 48634
rect 112204 48580 112260 48582
rect 111996 47066 112052 47068
rect 111996 47014 111998 47066
rect 111998 47014 112050 47066
rect 112050 47014 112052 47066
rect 111996 47012 112052 47014
rect 112100 47066 112156 47068
rect 112100 47014 112102 47066
rect 112102 47014 112154 47066
rect 112154 47014 112156 47066
rect 112100 47012 112156 47014
rect 112204 47066 112260 47068
rect 112204 47014 112206 47066
rect 112206 47014 112258 47066
rect 112258 47014 112260 47066
rect 112204 47012 112260 47014
rect 111996 45498 112052 45500
rect 111996 45446 111998 45498
rect 111998 45446 112050 45498
rect 112050 45446 112052 45498
rect 111996 45444 112052 45446
rect 112100 45498 112156 45500
rect 112100 45446 112102 45498
rect 112102 45446 112154 45498
rect 112154 45446 112156 45498
rect 112100 45444 112156 45446
rect 112204 45498 112260 45500
rect 112204 45446 112206 45498
rect 112206 45446 112258 45498
rect 112258 45446 112260 45498
rect 112204 45444 112260 45446
rect 111996 43930 112052 43932
rect 111996 43878 111998 43930
rect 111998 43878 112050 43930
rect 112050 43878 112052 43930
rect 111996 43876 112052 43878
rect 112100 43930 112156 43932
rect 112100 43878 112102 43930
rect 112102 43878 112154 43930
rect 112154 43878 112156 43930
rect 112100 43876 112156 43878
rect 112204 43930 112260 43932
rect 112204 43878 112206 43930
rect 112206 43878 112258 43930
rect 112258 43878 112260 43930
rect 112204 43876 112260 43878
rect 111996 42362 112052 42364
rect 111996 42310 111998 42362
rect 111998 42310 112050 42362
rect 112050 42310 112052 42362
rect 111996 42308 112052 42310
rect 112100 42362 112156 42364
rect 112100 42310 112102 42362
rect 112102 42310 112154 42362
rect 112154 42310 112156 42362
rect 112100 42308 112156 42310
rect 112204 42362 112260 42364
rect 112204 42310 112206 42362
rect 112206 42310 112258 42362
rect 112258 42310 112260 42362
rect 112204 42308 112260 42310
rect 111996 40794 112052 40796
rect 111996 40742 111998 40794
rect 111998 40742 112050 40794
rect 112050 40742 112052 40794
rect 111996 40740 112052 40742
rect 112100 40794 112156 40796
rect 112100 40742 112102 40794
rect 112102 40742 112154 40794
rect 112154 40742 112156 40794
rect 112100 40740 112156 40742
rect 112204 40794 112260 40796
rect 112204 40742 112206 40794
rect 112206 40742 112258 40794
rect 112258 40742 112260 40794
rect 112204 40740 112260 40742
rect 111996 39226 112052 39228
rect 111996 39174 111998 39226
rect 111998 39174 112050 39226
rect 112050 39174 112052 39226
rect 111996 39172 112052 39174
rect 112100 39226 112156 39228
rect 112100 39174 112102 39226
rect 112102 39174 112154 39226
rect 112154 39174 112156 39226
rect 112100 39172 112156 39174
rect 112204 39226 112260 39228
rect 112204 39174 112206 39226
rect 112206 39174 112258 39226
rect 112258 39174 112260 39226
rect 112204 39172 112260 39174
rect 111996 37658 112052 37660
rect 111996 37606 111998 37658
rect 111998 37606 112050 37658
rect 112050 37606 112052 37658
rect 111996 37604 112052 37606
rect 112100 37658 112156 37660
rect 112100 37606 112102 37658
rect 112102 37606 112154 37658
rect 112154 37606 112156 37658
rect 112100 37604 112156 37606
rect 112204 37658 112260 37660
rect 112204 37606 112206 37658
rect 112206 37606 112258 37658
rect 112258 37606 112260 37658
rect 112204 37604 112260 37606
rect 111996 36090 112052 36092
rect 111996 36038 111998 36090
rect 111998 36038 112050 36090
rect 112050 36038 112052 36090
rect 111996 36036 112052 36038
rect 112100 36090 112156 36092
rect 112100 36038 112102 36090
rect 112102 36038 112154 36090
rect 112154 36038 112156 36090
rect 112100 36036 112156 36038
rect 112204 36090 112260 36092
rect 112204 36038 112206 36090
rect 112206 36038 112258 36090
rect 112258 36038 112260 36090
rect 112204 36036 112260 36038
rect 111996 34522 112052 34524
rect 111996 34470 111998 34522
rect 111998 34470 112050 34522
rect 112050 34470 112052 34522
rect 111996 34468 112052 34470
rect 112100 34522 112156 34524
rect 112100 34470 112102 34522
rect 112102 34470 112154 34522
rect 112154 34470 112156 34522
rect 112100 34468 112156 34470
rect 112204 34522 112260 34524
rect 112204 34470 112206 34522
rect 112206 34470 112258 34522
rect 112258 34470 112260 34522
rect 112204 34468 112260 34470
rect 111996 32954 112052 32956
rect 111996 32902 111998 32954
rect 111998 32902 112050 32954
rect 112050 32902 112052 32954
rect 111996 32900 112052 32902
rect 112100 32954 112156 32956
rect 112100 32902 112102 32954
rect 112102 32902 112154 32954
rect 112154 32902 112156 32954
rect 112100 32900 112156 32902
rect 112204 32954 112260 32956
rect 112204 32902 112206 32954
rect 112206 32902 112258 32954
rect 112258 32902 112260 32954
rect 112204 32900 112260 32902
rect 111996 31386 112052 31388
rect 111996 31334 111998 31386
rect 111998 31334 112050 31386
rect 112050 31334 112052 31386
rect 111996 31332 112052 31334
rect 112100 31386 112156 31388
rect 112100 31334 112102 31386
rect 112102 31334 112154 31386
rect 112154 31334 112156 31386
rect 112100 31332 112156 31334
rect 112204 31386 112260 31388
rect 112204 31334 112206 31386
rect 112206 31334 112258 31386
rect 112258 31334 112260 31386
rect 112204 31332 112260 31334
rect 111996 29818 112052 29820
rect 111996 29766 111998 29818
rect 111998 29766 112050 29818
rect 112050 29766 112052 29818
rect 111996 29764 112052 29766
rect 112100 29818 112156 29820
rect 112100 29766 112102 29818
rect 112102 29766 112154 29818
rect 112154 29766 112156 29818
rect 112100 29764 112156 29766
rect 112204 29818 112260 29820
rect 112204 29766 112206 29818
rect 112206 29766 112258 29818
rect 112258 29766 112260 29818
rect 112204 29764 112260 29766
rect 127484 56252 127540 56308
rect 128716 56306 128772 56308
rect 128716 56254 128718 56306
rect 128718 56254 128770 56306
rect 128770 56254 128772 56306
rect 128716 56252 128772 56254
rect 131292 56252 131348 56308
rect 132524 56306 132580 56308
rect 132524 56254 132526 56306
rect 132526 56254 132578 56306
rect 132578 56254 132580 56306
rect 132524 56252 132580 56254
rect 123900 56194 123956 56196
rect 123900 56142 123902 56194
rect 123902 56142 123954 56194
rect 123954 56142 123956 56194
rect 123900 56140 123956 56142
rect 125132 55916 125188 55972
rect 115724 55298 115780 55300
rect 115724 55246 115726 55298
rect 115726 55246 115778 55298
rect 115778 55246 115780 55298
rect 115724 55244 115780 55246
rect 115836 54348 115892 54404
rect 116620 54402 116676 54404
rect 116620 54350 116622 54402
rect 116622 54350 116674 54402
rect 116674 54350 116676 54402
rect 116620 54348 116676 54350
rect 115052 28588 115108 28644
rect 111996 28250 112052 28252
rect 111996 28198 111998 28250
rect 111998 28198 112050 28250
rect 112050 28198 112052 28250
rect 111996 28196 112052 28198
rect 112100 28250 112156 28252
rect 112100 28198 112102 28250
rect 112102 28198 112154 28250
rect 112154 28198 112156 28250
rect 112100 28196 112156 28198
rect 112204 28250 112260 28252
rect 112204 28198 112206 28250
rect 112206 28198 112258 28250
rect 112258 28198 112260 28250
rect 112204 28196 112260 28198
rect 111996 26682 112052 26684
rect 111996 26630 111998 26682
rect 111998 26630 112050 26682
rect 112050 26630 112052 26682
rect 111996 26628 112052 26630
rect 112100 26682 112156 26684
rect 112100 26630 112102 26682
rect 112102 26630 112154 26682
rect 112154 26630 112156 26682
rect 112100 26628 112156 26630
rect 112204 26682 112260 26684
rect 112204 26630 112206 26682
rect 112206 26630 112258 26682
rect 112258 26630 112260 26682
rect 112204 26628 112260 26630
rect 110012 25340 110068 25396
rect 107772 20130 107828 20132
rect 107772 20078 107774 20130
rect 107774 20078 107826 20130
rect 107826 20078 107828 20130
rect 107772 20076 107828 20078
rect 111996 25114 112052 25116
rect 111996 25062 111998 25114
rect 111998 25062 112050 25114
rect 112050 25062 112052 25114
rect 111996 25060 112052 25062
rect 112100 25114 112156 25116
rect 112100 25062 112102 25114
rect 112102 25062 112154 25114
rect 112154 25062 112156 25114
rect 112100 25060 112156 25062
rect 112204 25114 112260 25116
rect 112204 25062 112206 25114
rect 112206 25062 112258 25114
rect 112258 25062 112260 25114
rect 112204 25060 112260 25062
rect 111996 23546 112052 23548
rect 111996 23494 111998 23546
rect 111998 23494 112050 23546
rect 112050 23494 112052 23546
rect 111996 23492 112052 23494
rect 112100 23546 112156 23548
rect 112100 23494 112102 23546
rect 112102 23494 112154 23546
rect 112154 23494 112156 23546
rect 112100 23492 112156 23494
rect 112204 23546 112260 23548
rect 112204 23494 112206 23546
rect 112206 23494 112258 23546
rect 112258 23494 112260 23546
rect 112204 23492 112260 23494
rect 108892 22876 108948 22932
rect 107996 20578 108052 20580
rect 107996 20526 107998 20578
rect 107998 20526 108050 20578
rect 108050 20526 108052 20578
rect 107996 20524 108052 20526
rect 108556 20130 108612 20132
rect 108556 20078 108558 20130
rect 108558 20078 108610 20130
rect 108610 20078 108612 20130
rect 108556 20076 108612 20078
rect 107884 19794 107940 19796
rect 107884 19742 107886 19794
rect 107886 19742 107938 19794
rect 107938 19742 107940 19794
rect 107884 19740 107940 19742
rect 107884 19122 107940 19124
rect 107884 19070 107886 19122
rect 107886 19070 107938 19122
rect 107938 19070 107940 19122
rect 107884 19068 107940 19070
rect 107548 17724 107604 17780
rect 107996 17612 108052 17668
rect 107660 17554 107716 17556
rect 107660 17502 107662 17554
rect 107662 17502 107714 17554
rect 107714 17502 107716 17554
rect 107660 17500 107716 17502
rect 107772 16716 107828 16772
rect 108220 20018 108276 20020
rect 108220 19966 108222 20018
rect 108222 19966 108274 20018
rect 108274 19966 108276 20018
rect 108220 19964 108276 19966
rect 108780 19852 108836 19908
rect 111996 21978 112052 21980
rect 111996 21926 111998 21978
rect 111998 21926 112050 21978
rect 112050 21926 112052 21978
rect 111996 21924 112052 21926
rect 112100 21978 112156 21980
rect 112100 21926 112102 21978
rect 112102 21926 112154 21978
rect 112154 21926 112156 21978
rect 112100 21924 112156 21926
rect 112204 21978 112260 21980
rect 112204 21926 112206 21978
rect 112206 21926 112258 21978
rect 112258 21926 112260 21978
rect 112204 21924 112260 21926
rect 110796 21532 110852 21588
rect 109788 20018 109844 20020
rect 109788 19966 109790 20018
rect 109790 19966 109842 20018
rect 109842 19966 109844 20018
rect 109788 19964 109844 19966
rect 110012 20018 110068 20020
rect 110012 19966 110014 20018
rect 110014 19966 110066 20018
rect 110066 19966 110068 20018
rect 110012 19964 110068 19966
rect 109788 19628 109844 19684
rect 109452 19234 109508 19236
rect 109452 19182 109454 19234
rect 109454 19182 109506 19234
rect 109506 19182 109508 19234
rect 109452 19180 109508 19182
rect 110236 19852 110292 19908
rect 111692 20524 111748 20580
rect 111996 20410 112052 20412
rect 111996 20358 111998 20410
rect 111998 20358 112050 20410
rect 112050 20358 112052 20410
rect 111996 20356 112052 20358
rect 112100 20410 112156 20412
rect 112100 20358 112102 20410
rect 112102 20358 112154 20410
rect 112154 20358 112156 20410
rect 112100 20356 112156 20358
rect 112204 20410 112260 20412
rect 112204 20358 112206 20410
rect 112206 20358 112258 20410
rect 112258 20358 112260 20410
rect 112204 20356 112260 20358
rect 112476 20076 112532 20132
rect 113372 20130 113428 20132
rect 113372 20078 113374 20130
rect 113374 20078 113426 20130
rect 113426 20078 113428 20130
rect 113372 20076 113428 20078
rect 111356 19964 111412 20020
rect 110908 19906 110964 19908
rect 110908 19854 110910 19906
rect 110910 19854 110962 19906
rect 110962 19854 110964 19906
rect 110908 19852 110964 19854
rect 110796 19740 110852 19796
rect 112364 20018 112420 20020
rect 112364 19966 112366 20018
rect 112366 19966 112418 20018
rect 112418 19966 112420 20018
rect 112364 19964 112420 19966
rect 111916 19852 111972 19908
rect 111356 19292 111412 19348
rect 112476 19906 112532 19908
rect 112476 19854 112478 19906
rect 112478 19854 112530 19906
rect 112530 19854 112532 19906
rect 112476 19852 112532 19854
rect 112924 19852 112980 19908
rect 112588 19628 112644 19684
rect 109116 18338 109172 18340
rect 109116 18286 109118 18338
rect 109118 18286 109170 18338
rect 109170 18286 109172 18338
rect 109116 18284 109172 18286
rect 109340 18172 109396 18228
rect 109228 17612 109284 17668
rect 108892 16828 108948 16884
rect 108780 16716 108836 16772
rect 107772 15708 107828 15764
rect 107436 15484 107492 15540
rect 107100 15202 107156 15204
rect 107100 15150 107102 15202
rect 107102 15150 107154 15202
rect 107154 15150 107156 15202
rect 107100 15148 107156 15150
rect 107660 15148 107716 15204
rect 109564 17388 109620 17444
rect 109788 18284 109844 18340
rect 110236 19180 110292 19236
rect 112364 19180 112420 19236
rect 113148 19180 113204 19236
rect 111996 18842 112052 18844
rect 111996 18790 111998 18842
rect 111998 18790 112050 18842
rect 112050 18790 112052 18842
rect 111996 18788 112052 18790
rect 112100 18842 112156 18844
rect 112100 18790 112102 18842
rect 112102 18790 112154 18842
rect 112154 18790 112156 18842
rect 112100 18788 112156 18790
rect 112204 18842 112260 18844
rect 112204 18790 112206 18842
rect 112206 18790 112258 18842
rect 112258 18790 112260 18842
rect 112204 18788 112260 18790
rect 111020 18396 111076 18452
rect 111692 18450 111748 18452
rect 111692 18398 111694 18450
rect 111694 18398 111746 18450
rect 111746 18398 111748 18450
rect 111692 18396 111748 18398
rect 112140 18450 112196 18452
rect 112140 18398 112142 18450
rect 112142 18398 112194 18450
rect 112194 18398 112196 18450
rect 112140 18396 112196 18398
rect 111916 18338 111972 18340
rect 111916 18286 111918 18338
rect 111918 18286 111970 18338
rect 111970 18286 111972 18338
rect 111916 18284 111972 18286
rect 112140 18172 112196 18228
rect 112812 18284 112868 18340
rect 111020 17836 111076 17892
rect 112252 17442 112308 17444
rect 112252 17390 112254 17442
rect 112254 17390 112306 17442
rect 112306 17390 112308 17442
rect 112252 17388 112308 17390
rect 111996 17274 112052 17276
rect 111996 17222 111998 17274
rect 111998 17222 112050 17274
rect 112050 17222 112052 17274
rect 111996 17220 112052 17222
rect 112100 17274 112156 17276
rect 112100 17222 112102 17274
rect 112102 17222 112154 17274
rect 112154 17222 112156 17274
rect 112100 17220 112156 17222
rect 112204 17274 112260 17276
rect 112204 17222 112206 17274
rect 112206 17222 112258 17274
rect 112258 17222 112260 17274
rect 112204 17220 112260 17222
rect 111916 16882 111972 16884
rect 111916 16830 111918 16882
rect 111918 16830 111970 16882
rect 111970 16830 111972 16882
rect 111916 16828 111972 16830
rect 107884 15484 107940 15540
rect 107212 14364 107268 14420
rect 108108 14252 108164 14308
rect 107548 13580 107604 13636
rect 108780 15538 108836 15540
rect 108780 15486 108782 15538
rect 108782 15486 108834 15538
rect 108834 15486 108836 15538
rect 108780 15484 108836 15486
rect 110236 16716 110292 16772
rect 112588 17052 112644 17108
rect 108892 15426 108948 15428
rect 108892 15374 108894 15426
rect 108894 15374 108946 15426
rect 108946 15374 108948 15426
rect 108892 15372 108948 15374
rect 109788 15202 109844 15204
rect 109788 15150 109790 15202
rect 109790 15150 109842 15202
rect 109842 15150 109844 15202
rect 109788 15148 109844 15150
rect 109004 14588 109060 14644
rect 108444 14364 108500 14420
rect 108332 14028 108388 14084
rect 109004 13580 109060 13636
rect 107660 13020 107716 13076
rect 108108 13468 108164 13524
rect 106988 12684 107044 12740
rect 107660 12738 107716 12740
rect 107660 12686 107662 12738
rect 107662 12686 107714 12738
rect 107714 12686 107716 12738
rect 107660 12684 107716 12686
rect 107884 12738 107940 12740
rect 107884 12686 107886 12738
rect 107886 12686 107938 12738
rect 107938 12686 107940 12738
rect 107884 12684 107940 12686
rect 108668 13244 108724 13300
rect 108220 13074 108276 13076
rect 108220 13022 108222 13074
rect 108222 13022 108274 13074
rect 108274 13022 108276 13074
rect 108220 13020 108276 13022
rect 108892 13132 108948 13188
rect 107324 12178 107380 12180
rect 107324 12126 107326 12178
rect 107326 12126 107378 12178
rect 107378 12126 107380 12178
rect 107324 12124 107380 12126
rect 106652 10668 106708 10724
rect 106204 9212 106260 9268
rect 106428 8764 106484 8820
rect 106204 8370 106260 8372
rect 106204 8318 106206 8370
rect 106206 8318 106258 8370
rect 106258 8318 106260 8370
rect 106204 8316 106260 8318
rect 105532 7474 105588 7476
rect 105532 7422 105534 7474
rect 105534 7422 105586 7474
rect 105586 7422 105588 7474
rect 105532 7420 105588 7422
rect 105756 6860 105812 6916
rect 106204 6972 106260 7028
rect 105420 6636 105476 6692
rect 104748 5516 104804 5572
rect 104860 5964 104916 6020
rect 104524 5068 104580 5124
rect 103964 3724 104020 3780
rect 103964 3554 104020 3556
rect 103964 3502 103966 3554
rect 103966 3502 104018 3554
rect 104018 3502 104020 3554
rect 103964 3500 104020 3502
rect 104636 3948 104692 4004
rect 105644 4620 105700 4676
rect 105868 4562 105924 4564
rect 105868 4510 105870 4562
rect 105870 4510 105922 4562
rect 105922 4510 105924 4562
rect 105868 4508 105924 4510
rect 104412 2828 104468 2884
rect 106540 6860 106596 6916
rect 106652 6412 106708 6468
rect 107100 9996 107156 10052
rect 106988 7980 107044 8036
rect 107996 12290 108052 12292
rect 107996 12238 107998 12290
rect 107998 12238 108050 12290
rect 108050 12238 108052 12290
rect 107996 12236 108052 12238
rect 107548 11282 107604 11284
rect 107548 11230 107550 11282
rect 107550 11230 107602 11282
rect 107602 11230 107604 11282
rect 107548 11228 107604 11230
rect 107436 9212 107492 9268
rect 107212 6524 107268 6580
rect 107436 8428 107492 8484
rect 107436 6412 107492 6468
rect 108108 11900 108164 11956
rect 107996 10108 108052 10164
rect 107884 9100 107940 9156
rect 107996 9826 108052 9828
rect 107996 9774 107998 9826
rect 107998 9774 108050 9826
rect 108050 9774 108052 9826
rect 107996 9772 108052 9774
rect 107884 8428 107940 8484
rect 107660 8316 107716 8372
rect 107660 8034 107716 8036
rect 107660 7982 107662 8034
rect 107662 7982 107714 8034
rect 107714 7982 107716 8034
rect 107660 7980 107716 7982
rect 107884 8034 107940 8036
rect 107884 7982 107886 8034
rect 107886 7982 107938 8034
rect 107938 7982 107940 8034
rect 107884 7980 107940 7982
rect 106876 6076 106932 6132
rect 106764 5010 106820 5012
rect 106764 4958 106766 5010
rect 106766 4958 106818 5010
rect 106818 4958 106820 5010
rect 106764 4956 106820 4958
rect 107324 4844 107380 4900
rect 105644 2716 105700 2772
rect 105980 4060 106036 4116
rect 107212 4114 107268 4116
rect 107212 4062 107214 4114
rect 107214 4062 107266 4114
rect 107266 4062 107268 4114
rect 107212 4060 107268 4062
rect 106876 3442 106932 3444
rect 106876 3390 106878 3442
rect 106878 3390 106930 3442
rect 106930 3390 106932 3442
rect 106876 3388 106932 3390
rect 107436 4732 107492 4788
rect 107884 6018 107940 6020
rect 107884 5966 107886 6018
rect 107886 5966 107938 6018
rect 107938 5966 107940 6018
rect 107884 5964 107940 5966
rect 107660 5010 107716 5012
rect 107660 4958 107662 5010
rect 107662 4958 107714 5010
rect 107714 4958 107716 5010
rect 107660 4956 107716 4958
rect 107548 4172 107604 4228
rect 108668 12348 108724 12404
rect 108556 12290 108612 12292
rect 108556 12238 108558 12290
rect 108558 12238 108610 12290
rect 108610 12238 108612 12290
rect 108556 12236 108612 12238
rect 108444 11900 108500 11956
rect 108556 12012 108612 12068
rect 108668 11788 108724 11844
rect 108332 10108 108388 10164
rect 108780 11282 108836 11284
rect 108780 11230 108782 11282
rect 108782 11230 108834 11282
rect 108834 11230 108836 11282
rect 108780 11228 108836 11230
rect 108780 10556 108836 10612
rect 112476 15874 112532 15876
rect 112476 15822 112478 15874
rect 112478 15822 112530 15874
rect 112530 15822 112532 15874
rect 112476 15820 112532 15822
rect 111996 15706 112052 15708
rect 111996 15654 111998 15706
rect 111998 15654 112050 15706
rect 112050 15654 112052 15706
rect 111996 15652 112052 15654
rect 112100 15706 112156 15708
rect 112100 15654 112102 15706
rect 112102 15654 112154 15706
rect 112154 15654 112156 15706
rect 112100 15652 112156 15654
rect 112204 15706 112260 15708
rect 112204 15654 112206 15706
rect 112206 15654 112258 15706
rect 112258 15654 112260 15706
rect 112204 15652 112260 15654
rect 113484 19740 113540 19796
rect 114940 19852 114996 19908
rect 114044 19346 114100 19348
rect 114044 19294 114046 19346
rect 114046 19294 114098 19346
rect 114098 19294 114100 19346
rect 114044 19292 114100 19294
rect 114156 19010 114212 19012
rect 114156 18958 114158 19010
rect 114158 18958 114210 19010
rect 114210 18958 114212 19010
rect 114156 18956 114212 18958
rect 113260 18396 113316 18452
rect 117964 18284 118020 18340
rect 115052 18226 115108 18228
rect 115052 18174 115054 18226
rect 115054 18174 115106 18226
rect 115106 18174 115108 18226
rect 115052 18172 115108 18174
rect 112924 17052 112980 17108
rect 115276 17106 115332 17108
rect 115276 17054 115278 17106
rect 115278 17054 115330 17106
rect 115330 17054 115332 17106
rect 115276 17052 115332 17054
rect 114940 15820 114996 15876
rect 112588 14924 112644 14980
rect 110572 14642 110628 14644
rect 110572 14590 110574 14642
rect 110574 14590 110626 14642
rect 110626 14590 110628 14642
rect 110572 14588 110628 14590
rect 110460 14252 110516 14308
rect 110348 13468 110404 13524
rect 109116 13132 109172 13188
rect 110348 13020 110404 13076
rect 109564 12962 109620 12964
rect 109564 12910 109566 12962
rect 109566 12910 109618 12962
rect 109618 12910 109620 12962
rect 109564 12908 109620 12910
rect 110012 12962 110068 12964
rect 110012 12910 110014 12962
rect 110014 12910 110066 12962
rect 110066 12910 110068 12962
rect 110012 12908 110068 12910
rect 109676 12684 109732 12740
rect 109340 12402 109396 12404
rect 109340 12350 109342 12402
rect 109342 12350 109394 12402
rect 109394 12350 109396 12402
rect 109340 12348 109396 12350
rect 109452 11452 109508 11508
rect 109116 9996 109172 10052
rect 109228 9938 109284 9940
rect 109228 9886 109230 9938
rect 109230 9886 109282 9938
rect 109282 9886 109284 9938
rect 109228 9884 109284 9886
rect 108780 8540 108836 8596
rect 109004 9042 109060 9044
rect 109004 8990 109006 9042
rect 109006 8990 109058 9042
rect 109058 8990 109060 9042
rect 109004 8988 109060 8990
rect 108556 8316 108612 8372
rect 108892 7980 108948 8036
rect 108444 7756 108500 7812
rect 108444 7084 108500 7140
rect 108780 6130 108836 6132
rect 108780 6078 108782 6130
rect 108782 6078 108834 6130
rect 108834 6078 108836 6130
rect 108780 6076 108836 6078
rect 108108 4284 108164 4340
rect 108556 5292 108612 5348
rect 108332 3836 108388 3892
rect 107548 3276 107604 3332
rect 109004 7084 109060 7140
rect 109228 6412 109284 6468
rect 109452 10722 109508 10724
rect 109452 10670 109454 10722
rect 109454 10670 109506 10722
rect 109506 10670 109508 10722
rect 109452 10668 109508 10670
rect 109900 12066 109956 12068
rect 109900 12014 109902 12066
rect 109902 12014 109954 12066
rect 109954 12014 109956 12066
rect 109900 12012 109956 12014
rect 111468 14252 111524 14308
rect 111996 14138 112052 14140
rect 111996 14086 111998 14138
rect 111998 14086 112050 14138
rect 112050 14086 112052 14138
rect 111996 14084 112052 14086
rect 112100 14138 112156 14140
rect 112100 14086 112102 14138
rect 112102 14086 112154 14138
rect 112154 14086 112156 14138
rect 112100 14084 112156 14086
rect 112204 14138 112260 14140
rect 112204 14086 112206 14138
rect 112206 14086 112258 14138
rect 112258 14086 112260 14138
rect 112204 14084 112260 14086
rect 111132 13468 111188 13524
rect 110012 11788 110068 11844
rect 109900 11676 109956 11732
rect 109676 9548 109732 9604
rect 109676 8428 109732 8484
rect 109564 7420 109620 7476
rect 110012 10722 110068 10724
rect 110012 10670 110014 10722
rect 110014 10670 110066 10722
rect 110066 10670 110068 10722
rect 110012 10668 110068 10670
rect 109900 10556 109956 10612
rect 110348 10332 110404 10388
rect 110124 9548 110180 9604
rect 110236 9996 110292 10052
rect 109900 8764 109956 8820
rect 109564 5516 109620 5572
rect 110236 7362 110292 7364
rect 110236 7310 110238 7362
rect 110238 7310 110290 7362
rect 110290 7310 110292 7362
rect 110236 7308 110292 7310
rect 110236 6748 110292 6804
rect 110348 6690 110404 6692
rect 110348 6638 110350 6690
rect 110350 6638 110402 6690
rect 110402 6638 110404 6690
rect 110348 6636 110404 6638
rect 110124 5234 110180 5236
rect 110124 5182 110126 5234
rect 110126 5182 110178 5234
rect 110178 5182 110180 5234
rect 110124 5180 110180 5182
rect 110012 4732 110068 4788
rect 110124 4620 110180 4676
rect 109228 3500 109284 3556
rect 109676 3836 109732 3892
rect 106876 2828 106932 2884
rect 110124 3724 110180 3780
rect 110908 12572 110964 12628
rect 110796 12460 110852 12516
rect 110572 10892 110628 10948
rect 110572 10556 110628 10612
rect 111020 11452 111076 11508
rect 110908 10834 110964 10836
rect 110908 10782 110910 10834
rect 110910 10782 110962 10834
rect 110962 10782 110964 10834
rect 110908 10780 110964 10782
rect 110796 10332 110852 10388
rect 110572 8652 110628 8708
rect 110684 8876 110740 8932
rect 110684 8540 110740 8596
rect 110684 8258 110740 8260
rect 110684 8206 110686 8258
rect 110686 8206 110738 8258
rect 110738 8206 110740 8258
rect 110684 8204 110740 8206
rect 110572 7420 110628 7476
rect 111244 12738 111300 12740
rect 111244 12686 111246 12738
rect 111246 12686 111298 12738
rect 111298 12686 111300 12738
rect 111244 12684 111300 12686
rect 111692 12850 111748 12852
rect 111692 12798 111694 12850
rect 111694 12798 111746 12850
rect 111746 12798 111748 12850
rect 111692 12796 111748 12798
rect 111580 11676 111636 11732
rect 111468 9884 111524 9940
rect 111580 10610 111636 10612
rect 111580 10558 111582 10610
rect 111582 10558 111634 10610
rect 111634 10558 111636 10610
rect 111580 10556 111636 10558
rect 111244 9772 111300 9828
rect 111356 9100 111412 9156
rect 112140 12962 112196 12964
rect 112140 12910 112142 12962
rect 112142 12910 112194 12962
rect 112194 12910 112196 12962
rect 112140 12908 112196 12910
rect 112700 12850 112756 12852
rect 112700 12798 112702 12850
rect 112702 12798 112754 12850
rect 112754 12798 112756 12850
rect 112700 12796 112756 12798
rect 111996 12570 112052 12572
rect 111996 12518 111998 12570
rect 111998 12518 112050 12570
rect 112050 12518 112052 12570
rect 111996 12516 112052 12518
rect 112100 12570 112156 12572
rect 112100 12518 112102 12570
rect 112102 12518 112154 12570
rect 112154 12518 112156 12570
rect 112100 12516 112156 12518
rect 112204 12570 112260 12572
rect 112204 12518 112206 12570
rect 112206 12518 112258 12570
rect 112258 12518 112260 12570
rect 112204 12516 112260 12518
rect 112700 12348 112756 12404
rect 112140 11394 112196 11396
rect 112140 11342 112142 11394
rect 112142 11342 112194 11394
rect 112194 11342 112196 11394
rect 112140 11340 112196 11342
rect 111916 11228 111972 11284
rect 111996 11002 112052 11004
rect 111996 10950 111998 11002
rect 111998 10950 112050 11002
rect 112050 10950 112052 11002
rect 111996 10948 112052 10950
rect 112100 11002 112156 11004
rect 112100 10950 112102 11002
rect 112102 10950 112154 11002
rect 112154 10950 112156 11002
rect 112100 10948 112156 10950
rect 112204 11002 112260 11004
rect 112204 10950 112206 11002
rect 112206 10950 112258 11002
rect 112258 10950 112260 11002
rect 112204 10948 112260 10950
rect 112140 10220 112196 10276
rect 111804 10108 111860 10164
rect 112924 12066 112980 12068
rect 112924 12014 112926 12066
rect 112926 12014 112978 12066
rect 112978 12014 112980 12066
rect 112924 12012 112980 12014
rect 112476 11900 112532 11956
rect 112028 9996 112084 10052
rect 112812 11452 112868 11508
rect 111996 9434 112052 9436
rect 111996 9382 111998 9434
rect 111998 9382 112050 9434
rect 112050 9382 112052 9434
rect 111996 9380 112052 9382
rect 112100 9434 112156 9436
rect 112100 9382 112102 9434
rect 112102 9382 112154 9434
rect 112154 9382 112156 9434
rect 112100 9380 112156 9382
rect 112204 9434 112260 9436
rect 112204 9382 112206 9434
rect 112206 9382 112258 9434
rect 112258 9382 112260 9434
rect 112204 9380 112260 9382
rect 111692 9212 111748 9268
rect 111132 8428 111188 8484
rect 111020 7980 111076 8036
rect 110908 7868 110964 7924
rect 111356 8540 111412 8596
rect 111356 8092 111412 8148
rect 112476 9548 112532 9604
rect 112476 9212 112532 9268
rect 112364 8988 112420 9044
rect 112476 8652 112532 8708
rect 112140 8204 112196 8260
rect 112364 8428 112420 8484
rect 112700 9212 112756 9268
rect 113036 11170 113092 11172
rect 113036 11118 113038 11170
rect 113038 11118 113090 11170
rect 113090 11118 113092 11170
rect 113036 11116 113092 11118
rect 113820 12684 113876 12740
rect 113148 10108 113204 10164
rect 113148 9436 113204 9492
rect 112924 9324 112980 9380
rect 113036 8988 113092 9044
rect 113372 9548 113428 9604
rect 113708 9884 113764 9940
rect 113932 9714 113988 9716
rect 113932 9662 113934 9714
rect 113934 9662 113986 9714
rect 113986 9662 113988 9714
rect 113932 9660 113988 9662
rect 113820 9436 113876 9492
rect 113484 9042 113540 9044
rect 113484 8990 113486 9042
rect 113486 8990 113538 9042
rect 113538 8990 113540 9042
rect 113484 8988 113540 8990
rect 111996 7866 112052 7868
rect 111996 7814 111998 7866
rect 111998 7814 112050 7866
rect 112050 7814 112052 7866
rect 111996 7812 112052 7814
rect 112100 7866 112156 7868
rect 112100 7814 112102 7866
rect 112102 7814 112154 7866
rect 112154 7814 112156 7866
rect 112100 7812 112156 7814
rect 112204 7866 112260 7868
rect 112204 7814 112206 7866
rect 112206 7814 112258 7866
rect 112258 7814 112260 7866
rect 112204 7812 112260 7814
rect 110684 6018 110740 6020
rect 110684 5966 110686 6018
rect 110686 5966 110738 6018
rect 110738 5966 110740 6018
rect 110684 5964 110740 5966
rect 111356 6018 111412 6020
rect 111356 5966 111358 6018
rect 111358 5966 111410 6018
rect 111410 5966 111412 6018
rect 111356 5964 111412 5966
rect 111244 5516 111300 5572
rect 111580 5852 111636 5908
rect 110908 4508 110964 4564
rect 111356 5180 111412 5236
rect 111356 4508 111412 4564
rect 110572 4338 110628 4340
rect 110572 4286 110574 4338
rect 110574 4286 110626 4338
rect 110626 4286 110628 4338
rect 110572 4284 110628 4286
rect 110460 3612 110516 3668
rect 109676 3164 109732 3220
rect 112028 6972 112084 7028
rect 112364 6578 112420 6580
rect 112364 6526 112366 6578
rect 112366 6526 112418 6578
rect 112418 6526 112420 6578
rect 112364 6524 112420 6526
rect 111996 6298 112052 6300
rect 111996 6246 111998 6298
rect 111998 6246 112050 6298
rect 112050 6246 112052 6298
rect 111996 6244 112052 6246
rect 112100 6298 112156 6300
rect 112100 6246 112102 6298
rect 112102 6246 112154 6298
rect 112154 6246 112156 6298
rect 112100 6244 112156 6246
rect 112204 6298 112260 6300
rect 112204 6246 112206 6298
rect 112206 6246 112258 6298
rect 112258 6246 112260 6298
rect 112204 6244 112260 6246
rect 112364 6300 112420 6356
rect 111804 5292 111860 5348
rect 112364 5180 112420 5236
rect 111916 5122 111972 5124
rect 111916 5070 111918 5122
rect 111918 5070 111970 5122
rect 111970 5070 111972 5122
rect 111916 5068 111972 5070
rect 111804 4898 111860 4900
rect 111804 4846 111806 4898
rect 111806 4846 111858 4898
rect 111858 4846 111860 4898
rect 111804 4844 111860 4846
rect 111996 4730 112052 4732
rect 111996 4678 111998 4730
rect 111998 4678 112050 4730
rect 112050 4678 112052 4730
rect 111996 4676 112052 4678
rect 112100 4730 112156 4732
rect 112100 4678 112102 4730
rect 112102 4678 112154 4730
rect 112154 4678 112156 4730
rect 112100 4676 112156 4678
rect 112204 4730 112260 4732
rect 112204 4678 112206 4730
rect 112206 4678 112258 4730
rect 112258 4678 112260 4730
rect 112204 4676 112260 4678
rect 111692 4172 111748 4228
rect 112252 4226 112308 4228
rect 112252 4174 112254 4226
rect 112254 4174 112306 4226
rect 112306 4174 112308 4226
rect 112252 4172 112308 4174
rect 112924 6524 112980 6580
rect 112588 4844 112644 4900
rect 112700 5964 112756 6020
rect 111996 3162 112052 3164
rect 111996 3110 111998 3162
rect 111998 3110 112050 3162
rect 112050 3110 112052 3162
rect 111996 3108 112052 3110
rect 112100 3162 112156 3164
rect 112100 3110 112102 3162
rect 112102 3110 112154 3162
rect 112154 3110 112156 3162
rect 112100 3108 112156 3110
rect 112204 3162 112260 3164
rect 112204 3110 112206 3162
rect 112206 3110 112258 3162
rect 112258 3110 112260 3162
rect 112204 3108 112260 3110
rect 111468 2940 111524 2996
rect 112924 5852 112980 5908
rect 113484 8370 113540 8372
rect 113484 8318 113486 8370
rect 113486 8318 113538 8370
rect 113538 8318 113540 8370
rect 113484 8316 113540 8318
rect 113932 9042 113988 9044
rect 113932 8990 113934 9042
rect 113934 8990 113986 9042
rect 113986 8990 113988 9042
rect 113932 8988 113988 8990
rect 113820 7980 113876 8036
rect 114156 9884 114212 9940
rect 114156 9154 114212 9156
rect 114156 9102 114158 9154
rect 114158 9102 114210 9154
rect 114210 9102 114212 9154
rect 114156 9100 114212 9102
rect 114380 10444 114436 10500
rect 114828 10332 114884 10388
rect 114492 9826 114548 9828
rect 114492 9774 114494 9826
rect 114494 9774 114546 9826
rect 114546 9774 114548 9826
rect 114492 9772 114548 9774
rect 114268 8258 114324 8260
rect 114268 8206 114270 8258
rect 114270 8206 114322 8258
rect 114322 8206 114324 8258
rect 114268 8204 114324 8206
rect 114044 7756 114100 7812
rect 114604 8316 114660 8372
rect 114604 7868 114660 7924
rect 114828 7980 114884 8036
rect 114716 7420 114772 7476
rect 115500 10498 115556 10500
rect 115500 10446 115502 10498
rect 115502 10446 115554 10498
rect 115554 10446 115556 10498
rect 115500 10444 115556 10446
rect 115612 9826 115668 9828
rect 115612 9774 115614 9826
rect 115614 9774 115666 9826
rect 115666 9774 115668 9826
rect 115612 9772 115668 9774
rect 115500 9602 115556 9604
rect 115500 9550 115502 9602
rect 115502 9550 115554 9602
rect 115554 9550 115556 9602
rect 115500 9548 115556 9550
rect 115388 9266 115444 9268
rect 115388 9214 115390 9266
rect 115390 9214 115442 9266
rect 115442 9214 115444 9266
rect 115388 9212 115444 9214
rect 115276 9100 115332 9156
rect 115500 8428 115556 8484
rect 115276 8204 115332 8260
rect 115612 8092 115668 8148
rect 115724 7532 115780 7588
rect 115052 7084 115108 7140
rect 115612 7308 115668 7364
rect 113708 6524 113764 6580
rect 114268 6748 114324 6804
rect 113484 6300 113540 6356
rect 114716 6578 114772 6580
rect 114716 6526 114718 6578
rect 114718 6526 114770 6578
rect 114770 6526 114772 6578
rect 114716 6524 114772 6526
rect 115500 6578 115556 6580
rect 115500 6526 115502 6578
rect 115502 6526 115554 6578
rect 115554 6526 115556 6578
rect 115500 6524 115556 6526
rect 114268 6076 114324 6132
rect 114380 6412 114436 6468
rect 115164 6076 115220 6132
rect 113260 4844 113316 4900
rect 113036 4508 113092 4564
rect 113260 4284 113316 4340
rect 112924 3666 112980 3668
rect 112924 3614 112926 3666
rect 112926 3614 112978 3666
rect 112978 3614 112980 3666
rect 112924 3612 112980 3614
rect 113820 4508 113876 4564
rect 113372 3052 113428 3108
rect 115164 4226 115220 4228
rect 115164 4174 115166 4226
rect 115166 4174 115218 4226
rect 115218 4174 115220 4226
rect 115164 4172 115220 4174
rect 115388 4338 115444 4340
rect 115388 4286 115390 4338
rect 115390 4286 115442 4338
rect 115442 4286 115444 4338
rect 115388 4284 115444 4286
rect 113932 2716 113988 2772
rect 114044 3388 114100 3444
rect 114604 3330 114660 3332
rect 114604 3278 114606 3330
rect 114606 3278 114658 3330
rect 114658 3278 114660 3330
rect 114604 3276 114660 3278
rect 115500 2940 115556 2996
rect 116060 11564 116116 11620
rect 115948 10498 116004 10500
rect 115948 10446 115950 10498
rect 115950 10446 116002 10498
rect 116002 10446 116004 10498
rect 115948 10444 116004 10446
rect 117292 10668 117348 10724
rect 115948 9660 116004 9716
rect 116396 9548 116452 9604
rect 116172 9154 116228 9156
rect 116172 9102 116174 9154
rect 116174 9102 116226 9154
rect 116226 9102 116228 9154
rect 116172 9100 116228 9102
rect 116284 8764 116340 8820
rect 116396 7586 116452 7588
rect 116396 7534 116398 7586
rect 116398 7534 116450 7586
rect 116450 7534 116452 7586
rect 116396 7532 116452 7534
rect 116284 6860 116340 6916
rect 115948 4844 116004 4900
rect 116732 8204 116788 8260
rect 116396 5516 116452 5572
rect 116844 5964 116900 6020
rect 117180 8764 117236 8820
rect 117292 8034 117348 8036
rect 117292 7982 117294 8034
rect 117294 7982 117346 8034
rect 117346 7982 117348 8034
rect 117292 7980 117348 7982
rect 117628 8930 117684 8932
rect 117628 8878 117630 8930
rect 117630 8878 117682 8930
rect 117682 8878 117684 8930
rect 117628 8876 117684 8878
rect 118412 14924 118468 14980
rect 118300 10780 118356 10836
rect 117516 8316 117572 8372
rect 117404 7362 117460 7364
rect 117404 7310 117406 7362
rect 117406 7310 117458 7362
rect 117458 7310 117460 7362
rect 117404 7308 117460 7310
rect 117292 6466 117348 6468
rect 117292 6414 117294 6466
rect 117294 6414 117346 6466
rect 117346 6414 117348 6466
rect 117292 6412 117348 6414
rect 117740 7308 117796 7364
rect 117852 6748 117908 6804
rect 117964 6972 118020 7028
rect 117628 6076 117684 6132
rect 117852 5906 117908 5908
rect 117852 5854 117854 5906
rect 117854 5854 117906 5906
rect 117906 5854 117908 5906
rect 117852 5852 117908 5854
rect 117068 5740 117124 5796
rect 117628 5628 117684 5684
rect 117852 5516 117908 5572
rect 116956 4844 117012 4900
rect 116620 3948 116676 4004
rect 116732 4620 116788 4676
rect 115052 2604 115108 2660
rect 117852 4898 117908 4900
rect 117852 4846 117854 4898
rect 117854 4846 117906 4898
rect 117906 4846 117908 4898
rect 117852 4844 117908 4846
rect 118300 8258 118356 8260
rect 118300 8206 118302 8258
rect 118302 8206 118354 8258
rect 118354 8206 118356 8258
rect 118300 8204 118356 8206
rect 118188 7362 118244 7364
rect 118188 7310 118190 7362
rect 118190 7310 118242 7362
rect 118242 7310 118244 7362
rect 118188 7308 118244 7310
rect 127356 55690 127412 55692
rect 127356 55638 127358 55690
rect 127358 55638 127410 55690
rect 127410 55638 127412 55690
rect 127356 55636 127412 55638
rect 127460 55690 127516 55692
rect 127460 55638 127462 55690
rect 127462 55638 127514 55690
rect 127514 55638 127516 55690
rect 127460 55636 127516 55638
rect 127564 55690 127620 55692
rect 127564 55638 127566 55690
rect 127566 55638 127618 55690
rect 127618 55638 127620 55690
rect 127564 55636 127620 55638
rect 126812 55186 126868 55188
rect 126812 55134 126814 55186
rect 126814 55134 126866 55186
rect 126866 55134 126868 55186
rect 126812 55132 126868 55134
rect 127260 55132 127316 55188
rect 126812 54348 126868 54404
rect 142716 57036 142772 57092
rect 144508 57036 144564 57092
rect 142716 56474 142772 56476
rect 142716 56422 142718 56474
rect 142718 56422 142770 56474
rect 142770 56422 142772 56474
rect 142716 56420 142772 56422
rect 142820 56474 142876 56476
rect 142820 56422 142822 56474
rect 142822 56422 142874 56474
rect 142874 56422 142876 56474
rect 142820 56420 142876 56422
rect 142924 56474 142980 56476
rect 142924 56422 142926 56474
rect 142926 56422 142978 56474
rect 142978 56422 142980 56474
rect 142924 56420 142980 56422
rect 138908 56252 138964 56308
rect 140140 56306 140196 56308
rect 140140 56254 140142 56306
rect 140142 56254 140194 56306
rect 140194 56254 140196 56306
rect 140140 56252 140196 56254
rect 135772 55970 135828 55972
rect 135772 55918 135774 55970
rect 135774 55918 135826 55970
rect 135826 55918 135828 55970
rect 135772 55916 135828 55918
rect 136892 55916 136948 55972
rect 127356 54122 127412 54124
rect 127356 54070 127358 54122
rect 127358 54070 127410 54122
rect 127410 54070 127412 54122
rect 127356 54068 127412 54070
rect 127460 54122 127516 54124
rect 127460 54070 127462 54122
rect 127462 54070 127514 54122
rect 127514 54070 127516 54122
rect 127460 54068 127516 54070
rect 127564 54122 127620 54124
rect 127564 54070 127566 54122
rect 127566 54070 127618 54122
rect 127618 54070 127620 54122
rect 127564 54068 127620 54070
rect 127356 52554 127412 52556
rect 127356 52502 127358 52554
rect 127358 52502 127410 52554
rect 127410 52502 127412 52554
rect 127356 52500 127412 52502
rect 127460 52554 127516 52556
rect 127460 52502 127462 52554
rect 127462 52502 127514 52554
rect 127514 52502 127516 52554
rect 127460 52500 127516 52502
rect 127564 52554 127620 52556
rect 127564 52502 127566 52554
rect 127566 52502 127618 52554
rect 127618 52502 127620 52554
rect 127564 52500 127620 52502
rect 127356 50986 127412 50988
rect 127356 50934 127358 50986
rect 127358 50934 127410 50986
rect 127410 50934 127412 50986
rect 127356 50932 127412 50934
rect 127460 50986 127516 50988
rect 127460 50934 127462 50986
rect 127462 50934 127514 50986
rect 127514 50934 127516 50986
rect 127460 50932 127516 50934
rect 127564 50986 127620 50988
rect 127564 50934 127566 50986
rect 127566 50934 127618 50986
rect 127618 50934 127620 50986
rect 127564 50932 127620 50934
rect 127356 49418 127412 49420
rect 127356 49366 127358 49418
rect 127358 49366 127410 49418
rect 127410 49366 127412 49418
rect 127356 49364 127412 49366
rect 127460 49418 127516 49420
rect 127460 49366 127462 49418
rect 127462 49366 127514 49418
rect 127514 49366 127516 49418
rect 127460 49364 127516 49366
rect 127564 49418 127620 49420
rect 127564 49366 127566 49418
rect 127566 49366 127618 49418
rect 127618 49366 127620 49418
rect 127564 49364 127620 49366
rect 127356 47850 127412 47852
rect 127356 47798 127358 47850
rect 127358 47798 127410 47850
rect 127410 47798 127412 47850
rect 127356 47796 127412 47798
rect 127460 47850 127516 47852
rect 127460 47798 127462 47850
rect 127462 47798 127514 47850
rect 127514 47798 127516 47850
rect 127460 47796 127516 47798
rect 127564 47850 127620 47852
rect 127564 47798 127566 47850
rect 127566 47798 127618 47850
rect 127618 47798 127620 47850
rect 127564 47796 127620 47798
rect 127356 46282 127412 46284
rect 127356 46230 127358 46282
rect 127358 46230 127410 46282
rect 127410 46230 127412 46282
rect 127356 46228 127412 46230
rect 127460 46282 127516 46284
rect 127460 46230 127462 46282
rect 127462 46230 127514 46282
rect 127514 46230 127516 46282
rect 127460 46228 127516 46230
rect 127564 46282 127620 46284
rect 127564 46230 127566 46282
rect 127566 46230 127618 46282
rect 127618 46230 127620 46282
rect 127564 46228 127620 46230
rect 127356 44714 127412 44716
rect 127356 44662 127358 44714
rect 127358 44662 127410 44714
rect 127410 44662 127412 44714
rect 127356 44660 127412 44662
rect 127460 44714 127516 44716
rect 127460 44662 127462 44714
rect 127462 44662 127514 44714
rect 127514 44662 127516 44714
rect 127460 44660 127516 44662
rect 127564 44714 127620 44716
rect 127564 44662 127566 44714
rect 127566 44662 127618 44714
rect 127618 44662 127620 44714
rect 127564 44660 127620 44662
rect 127356 43146 127412 43148
rect 127356 43094 127358 43146
rect 127358 43094 127410 43146
rect 127410 43094 127412 43146
rect 127356 43092 127412 43094
rect 127460 43146 127516 43148
rect 127460 43094 127462 43146
rect 127462 43094 127514 43146
rect 127514 43094 127516 43146
rect 127460 43092 127516 43094
rect 127564 43146 127620 43148
rect 127564 43094 127566 43146
rect 127566 43094 127618 43146
rect 127618 43094 127620 43146
rect 127564 43092 127620 43094
rect 127356 41578 127412 41580
rect 127356 41526 127358 41578
rect 127358 41526 127410 41578
rect 127410 41526 127412 41578
rect 127356 41524 127412 41526
rect 127460 41578 127516 41580
rect 127460 41526 127462 41578
rect 127462 41526 127514 41578
rect 127514 41526 127516 41578
rect 127460 41524 127516 41526
rect 127564 41578 127620 41580
rect 127564 41526 127566 41578
rect 127566 41526 127618 41578
rect 127618 41526 127620 41578
rect 127564 41524 127620 41526
rect 127356 40010 127412 40012
rect 127356 39958 127358 40010
rect 127358 39958 127410 40010
rect 127410 39958 127412 40010
rect 127356 39956 127412 39958
rect 127460 40010 127516 40012
rect 127460 39958 127462 40010
rect 127462 39958 127514 40010
rect 127514 39958 127516 40010
rect 127460 39956 127516 39958
rect 127564 40010 127620 40012
rect 127564 39958 127566 40010
rect 127566 39958 127618 40010
rect 127618 39958 127620 40010
rect 127564 39956 127620 39958
rect 127356 38442 127412 38444
rect 127356 38390 127358 38442
rect 127358 38390 127410 38442
rect 127410 38390 127412 38442
rect 127356 38388 127412 38390
rect 127460 38442 127516 38444
rect 127460 38390 127462 38442
rect 127462 38390 127514 38442
rect 127514 38390 127516 38442
rect 127460 38388 127516 38390
rect 127564 38442 127620 38444
rect 127564 38390 127566 38442
rect 127566 38390 127618 38442
rect 127618 38390 127620 38442
rect 127564 38388 127620 38390
rect 127356 36874 127412 36876
rect 127356 36822 127358 36874
rect 127358 36822 127410 36874
rect 127410 36822 127412 36874
rect 127356 36820 127412 36822
rect 127460 36874 127516 36876
rect 127460 36822 127462 36874
rect 127462 36822 127514 36874
rect 127514 36822 127516 36874
rect 127460 36820 127516 36822
rect 127564 36874 127620 36876
rect 127564 36822 127566 36874
rect 127566 36822 127618 36874
rect 127618 36822 127620 36874
rect 127564 36820 127620 36822
rect 127356 35306 127412 35308
rect 127356 35254 127358 35306
rect 127358 35254 127410 35306
rect 127410 35254 127412 35306
rect 127356 35252 127412 35254
rect 127460 35306 127516 35308
rect 127460 35254 127462 35306
rect 127462 35254 127514 35306
rect 127514 35254 127516 35306
rect 127460 35252 127516 35254
rect 127564 35306 127620 35308
rect 127564 35254 127566 35306
rect 127566 35254 127618 35306
rect 127618 35254 127620 35306
rect 127564 35252 127620 35254
rect 127356 33738 127412 33740
rect 127356 33686 127358 33738
rect 127358 33686 127410 33738
rect 127410 33686 127412 33738
rect 127356 33684 127412 33686
rect 127460 33738 127516 33740
rect 127460 33686 127462 33738
rect 127462 33686 127514 33738
rect 127514 33686 127516 33738
rect 127460 33684 127516 33686
rect 127564 33738 127620 33740
rect 127564 33686 127566 33738
rect 127566 33686 127618 33738
rect 127618 33686 127620 33738
rect 127564 33684 127620 33686
rect 125132 32732 125188 32788
rect 127356 32170 127412 32172
rect 127356 32118 127358 32170
rect 127358 32118 127410 32170
rect 127410 32118 127412 32170
rect 127356 32116 127412 32118
rect 127460 32170 127516 32172
rect 127460 32118 127462 32170
rect 127462 32118 127514 32170
rect 127514 32118 127516 32170
rect 127460 32116 127516 32118
rect 127564 32170 127620 32172
rect 127564 32118 127566 32170
rect 127566 32118 127618 32170
rect 127618 32118 127620 32170
rect 127564 32116 127620 32118
rect 127356 30602 127412 30604
rect 127356 30550 127358 30602
rect 127358 30550 127410 30602
rect 127410 30550 127412 30602
rect 127356 30548 127412 30550
rect 127460 30602 127516 30604
rect 127460 30550 127462 30602
rect 127462 30550 127514 30602
rect 127514 30550 127516 30602
rect 127460 30548 127516 30550
rect 127564 30602 127620 30604
rect 127564 30550 127566 30602
rect 127566 30550 127618 30602
rect 127618 30550 127620 30602
rect 127564 30548 127620 30550
rect 127356 29034 127412 29036
rect 127356 28982 127358 29034
rect 127358 28982 127410 29034
rect 127410 28982 127412 29034
rect 127356 28980 127412 28982
rect 127460 29034 127516 29036
rect 127460 28982 127462 29034
rect 127462 28982 127514 29034
rect 127514 28982 127516 29034
rect 127460 28980 127516 28982
rect 127564 29034 127620 29036
rect 127564 28982 127566 29034
rect 127566 28982 127618 29034
rect 127618 28982 127620 29034
rect 127564 28980 127620 28982
rect 127356 27466 127412 27468
rect 127356 27414 127358 27466
rect 127358 27414 127410 27466
rect 127410 27414 127412 27466
rect 127356 27412 127412 27414
rect 127460 27466 127516 27468
rect 127460 27414 127462 27466
rect 127462 27414 127514 27466
rect 127514 27414 127516 27466
rect 127460 27412 127516 27414
rect 127564 27466 127620 27468
rect 127564 27414 127566 27466
rect 127566 27414 127618 27466
rect 127618 27414 127620 27466
rect 127564 27412 127620 27414
rect 127356 25898 127412 25900
rect 127356 25846 127358 25898
rect 127358 25846 127410 25898
rect 127410 25846 127412 25898
rect 127356 25844 127412 25846
rect 127460 25898 127516 25900
rect 127460 25846 127462 25898
rect 127462 25846 127514 25898
rect 127514 25846 127516 25898
rect 127460 25844 127516 25846
rect 127564 25898 127620 25900
rect 127564 25846 127566 25898
rect 127566 25846 127618 25898
rect 127618 25846 127620 25898
rect 127564 25844 127620 25846
rect 127356 24330 127412 24332
rect 127356 24278 127358 24330
rect 127358 24278 127410 24330
rect 127410 24278 127412 24330
rect 127356 24276 127412 24278
rect 127460 24330 127516 24332
rect 127460 24278 127462 24330
rect 127462 24278 127514 24330
rect 127514 24278 127516 24330
rect 127460 24276 127516 24278
rect 127564 24330 127620 24332
rect 127564 24278 127566 24330
rect 127566 24278 127618 24330
rect 127618 24278 127620 24330
rect 127564 24276 127620 24278
rect 127356 22762 127412 22764
rect 127356 22710 127358 22762
rect 127358 22710 127410 22762
rect 127410 22710 127412 22762
rect 127356 22708 127412 22710
rect 127460 22762 127516 22764
rect 127460 22710 127462 22762
rect 127462 22710 127514 22762
rect 127514 22710 127516 22762
rect 127460 22708 127516 22710
rect 127564 22762 127620 22764
rect 127564 22710 127566 22762
rect 127566 22710 127618 22762
rect 127618 22710 127620 22762
rect 127564 22708 127620 22710
rect 127356 21194 127412 21196
rect 127356 21142 127358 21194
rect 127358 21142 127410 21194
rect 127410 21142 127412 21194
rect 127356 21140 127412 21142
rect 127460 21194 127516 21196
rect 127460 21142 127462 21194
rect 127462 21142 127514 21194
rect 127514 21142 127516 21194
rect 127460 21140 127516 21142
rect 127564 21194 127620 21196
rect 127564 21142 127566 21194
rect 127566 21142 127618 21194
rect 127618 21142 127620 21194
rect 127564 21140 127620 21142
rect 127356 19626 127412 19628
rect 127356 19574 127358 19626
rect 127358 19574 127410 19626
rect 127410 19574 127412 19626
rect 127356 19572 127412 19574
rect 127460 19626 127516 19628
rect 127460 19574 127462 19626
rect 127462 19574 127514 19626
rect 127514 19574 127516 19626
rect 127460 19572 127516 19574
rect 127564 19626 127620 19628
rect 127564 19574 127566 19626
rect 127566 19574 127618 19626
rect 127618 19574 127620 19626
rect 127564 19572 127620 19574
rect 119756 14476 119812 14532
rect 120092 18172 120148 18228
rect 119532 13916 119588 13972
rect 118748 8258 118804 8260
rect 118748 8206 118750 8258
rect 118750 8206 118802 8258
rect 118802 8206 118804 8258
rect 118748 8204 118804 8206
rect 118748 7698 118804 7700
rect 118748 7646 118750 7698
rect 118750 7646 118802 7698
rect 118802 7646 118804 7698
rect 118748 7644 118804 7646
rect 118636 6412 118692 6468
rect 118636 5682 118692 5684
rect 118636 5630 118638 5682
rect 118638 5630 118690 5682
rect 118690 5630 118692 5682
rect 118636 5628 118692 5630
rect 118524 5516 118580 5572
rect 119084 5964 119140 6020
rect 118748 4620 118804 4676
rect 118412 4114 118468 4116
rect 118412 4062 118414 4114
rect 118414 4062 118466 4114
rect 118466 4062 118468 4114
rect 118412 4060 118468 4062
rect 118076 3612 118132 3668
rect 117628 3442 117684 3444
rect 117628 3390 117630 3442
rect 117630 3390 117682 3442
rect 117682 3390 117684 3442
rect 117628 3388 117684 3390
rect 119420 5794 119476 5796
rect 119420 5742 119422 5794
rect 119422 5742 119474 5794
rect 119474 5742 119476 5794
rect 119420 5740 119476 5742
rect 119308 5068 119364 5124
rect 119420 3948 119476 4004
rect 118860 3442 118916 3444
rect 118860 3390 118862 3442
rect 118862 3390 118914 3442
rect 118914 3390 118916 3442
rect 118860 3388 118916 3390
rect 119868 7698 119924 7700
rect 119868 7646 119870 7698
rect 119870 7646 119922 7698
rect 119922 7646 119924 7698
rect 119868 7644 119924 7646
rect 119644 5906 119700 5908
rect 119644 5854 119646 5906
rect 119646 5854 119698 5906
rect 119698 5854 119700 5906
rect 119644 5852 119700 5854
rect 127356 18058 127412 18060
rect 127356 18006 127358 18058
rect 127358 18006 127410 18058
rect 127410 18006 127412 18058
rect 127356 18004 127412 18006
rect 127460 18058 127516 18060
rect 127460 18006 127462 18058
rect 127462 18006 127514 18058
rect 127514 18006 127516 18058
rect 127460 18004 127516 18006
rect 127564 18058 127620 18060
rect 127564 18006 127566 18058
rect 127566 18006 127618 18058
rect 127618 18006 127620 18058
rect 127564 18004 127620 18006
rect 127356 16490 127412 16492
rect 127356 16438 127358 16490
rect 127358 16438 127410 16490
rect 127410 16438 127412 16490
rect 127356 16436 127412 16438
rect 127460 16490 127516 16492
rect 127460 16438 127462 16490
rect 127462 16438 127514 16490
rect 127514 16438 127516 16490
rect 127460 16436 127516 16438
rect 127564 16490 127620 16492
rect 127564 16438 127566 16490
rect 127566 16438 127618 16490
rect 127618 16438 127620 16490
rect 127564 16436 127620 16438
rect 127356 14922 127412 14924
rect 127356 14870 127358 14922
rect 127358 14870 127410 14922
rect 127410 14870 127412 14922
rect 127356 14868 127412 14870
rect 127460 14922 127516 14924
rect 127460 14870 127462 14922
rect 127462 14870 127514 14922
rect 127514 14870 127516 14922
rect 127460 14868 127516 14870
rect 127564 14922 127620 14924
rect 127564 14870 127566 14922
rect 127566 14870 127618 14922
rect 127618 14870 127620 14922
rect 127564 14868 127620 14870
rect 138348 55186 138404 55188
rect 138348 55134 138350 55186
rect 138350 55134 138402 55186
rect 138402 55134 138404 55186
rect 138348 55132 138404 55134
rect 139020 55132 139076 55188
rect 150332 56252 150388 56308
rect 151564 56306 151620 56308
rect 151564 56254 151566 56306
rect 151566 56254 151618 56306
rect 151618 56254 151620 56306
rect 151564 56252 151620 56254
rect 154140 56252 154196 56308
rect 155372 56306 155428 56308
rect 155372 56254 155374 56306
rect 155374 56254 155426 56306
rect 155426 56254 155428 56306
rect 155372 56252 155428 56254
rect 147196 55970 147252 55972
rect 147196 55918 147198 55970
rect 147198 55918 147250 55970
rect 147250 55918 147252 55970
rect 147196 55916 147252 55918
rect 136892 27692 136948 27748
rect 149772 55356 149828 55412
rect 158076 55690 158132 55692
rect 158076 55638 158078 55690
rect 158078 55638 158130 55690
rect 158130 55638 158132 55690
rect 158076 55636 158132 55638
rect 158180 55690 158236 55692
rect 158180 55638 158182 55690
rect 158182 55638 158234 55690
rect 158234 55638 158236 55690
rect 158180 55636 158236 55638
rect 158284 55690 158340 55692
rect 158284 55638 158286 55690
rect 158286 55638 158338 55690
rect 158338 55638 158340 55690
rect 158284 55636 158340 55638
rect 150780 55356 150836 55412
rect 142716 54906 142772 54908
rect 142716 54854 142718 54906
rect 142718 54854 142770 54906
rect 142770 54854 142772 54906
rect 142716 54852 142772 54854
rect 142820 54906 142876 54908
rect 142820 54854 142822 54906
rect 142822 54854 142874 54906
rect 142874 54854 142876 54906
rect 142820 54852 142876 54854
rect 142924 54906 142980 54908
rect 142924 54854 142926 54906
rect 142926 54854 142978 54906
rect 142978 54854 142980 54906
rect 142924 54852 142980 54854
rect 142716 53338 142772 53340
rect 142716 53286 142718 53338
rect 142718 53286 142770 53338
rect 142770 53286 142772 53338
rect 142716 53284 142772 53286
rect 142820 53338 142876 53340
rect 142820 53286 142822 53338
rect 142822 53286 142874 53338
rect 142874 53286 142876 53338
rect 142820 53284 142876 53286
rect 142924 53338 142980 53340
rect 142924 53286 142926 53338
rect 142926 53286 142978 53338
rect 142978 53286 142980 53338
rect 142924 53284 142980 53286
rect 142716 51770 142772 51772
rect 142716 51718 142718 51770
rect 142718 51718 142770 51770
rect 142770 51718 142772 51770
rect 142716 51716 142772 51718
rect 142820 51770 142876 51772
rect 142820 51718 142822 51770
rect 142822 51718 142874 51770
rect 142874 51718 142876 51770
rect 142820 51716 142876 51718
rect 142924 51770 142980 51772
rect 142924 51718 142926 51770
rect 142926 51718 142978 51770
rect 142978 51718 142980 51770
rect 142924 51716 142980 51718
rect 142716 50202 142772 50204
rect 142716 50150 142718 50202
rect 142718 50150 142770 50202
rect 142770 50150 142772 50202
rect 142716 50148 142772 50150
rect 142820 50202 142876 50204
rect 142820 50150 142822 50202
rect 142822 50150 142874 50202
rect 142874 50150 142876 50202
rect 142820 50148 142876 50150
rect 142924 50202 142980 50204
rect 142924 50150 142926 50202
rect 142926 50150 142978 50202
rect 142978 50150 142980 50202
rect 142924 50148 142980 50150
rect 142716 48634 142772 48636
rect 142716 48582 142718 48634
rect 142718 48582 142770 48634
rect 142770 48582 142772 48634
rect 142716 48580 142772 48582
rect 142820 48634 142876 48636
rect 142820 48582 142822 48634
rect 142822 48582 142874 48634
rect 142874 48582 142876 48634
rect 142820 48580 142876 48582
rect 142924 48634 142980 48636
rect 142924 48582 142926 48634
rect 142926 48582 142978 48634
rect 142978 48582 142980 48634
rect 142924 48580 142980 48582
rect 142716 47066 142772 47068
rect 142716 47014 142718 47066
rect 142718 47014 142770 47066
rect 142770 47014 142772 47066
rect 142716 47012 142772 47014
rect 142820 47066 142876 47068
rect 142820 47014 142822 47066
rect 142822 47014 142874 47066
rect 142874 47014 142876 47066
rect 142820 47012 142876 47014
rect 142924 47066 142980 47068
rect 142924 47014 142926 47066
rect 142926 47014 142978 47066
rect 142978 47014 142980 47066
rect 142924 47012 142980 47014
rect 142716 45498 142772 45500
rect 142716 45446 142718 45498
rect 142718 45446 142770 45498
rect 142770 45446 142772 45498
rect 142716 45444 142772 45446
rect 142820 45498 142876 45500
rect 142820 45446 142822 45498
rect 142822 45446 142874 45498
rect 142874 45446 142876 45498
rect 142820 45444 142876 45446
rect 142924 45498 142980 45500
rect 142924 45446 142926 45498
rect 142926 45446 142978 45498
rect 142978 45446 142980 45498
rect 142924 45444 142980 45446
rect 142716 43930 142772 43932
rect 142716 43878 142718 43930
rect 142718 43878 142770 43930
rect 142770 43878 142772 43930
rect 142716 43876 142772 43878
rect 142820 43930 142876 43932
rect 142820 43878 142822 43930
rect 142822 43878 142874 43930
rect 142874 43878 142876 43930
rect 142820 43876 142876 43878
rect 142924 43930 142980 43932
rect 142924 43878 142926 43930
rect 142926 43878 142978 43930
rect 142978 43878 142980 43930
rect 142924 43876 142980 43878
rect 142716 42362 142772 42364
rect 142716 42310 142718 42362
rect 142718 42310 142770 42362
rect 142770 42310 142772 42362
rect 142716 42308 142772 42310
rect 142820 42362 142876 42364
rect 142820 42310 142822 42362
rect 142822 42310 142874 42362
rect 142874 42310 142876 42362
rect 142820 42308 142876 42310
rect 142924 42362 142980 42364
rect 142924 42310 142926 42362
rect 142926 42310 142978 42362
rect 142978 42310 142980 42362
rect 142924 42308 142980 42310
rect 142716 40794 142772 40796
rect 142716 40742 142718 40794
rect 142718 40742 142770 40794
rect 142770 40742 142772 40794
rect 142716 40740 142772 40742
rect 142820 40794 142876 40796
rect 142820 40742 142822 40794
rect 142822 40742 142874 40794
rect 142874 40742 142876 40794
rect 142820 40740 142876 40742
rect 142924 40794 142980 40796
rect 142924 40742 142926 40794
rect 142926 40742 142978 40794
rect 142978 40742 142980 40794
rect 142924 40740 142980 40742
rect 142716 39226 142772 39228
rect 142716 39174 142718 39226
rect 142718 39174 142770 39226
rect 142770 39174 142772 39226
rect 142716 39172 142772 39174
rect 142820 39226 142876 39228
rect 142820 39174 142822 39226
rect 142822 39174 142874 39226
rect 142874 39174 142876 39226
rect 142820 39172 142876 39174
rect 142924 39226 142980 39228
rect 142924 39174 142926 39226
rect 142926 39174 142978 39226
rect 142978 39174 142980 39226
rect 142924 39172 142980 39174
rect 142716 37658 142772 37660
rect 142716 37606 142718 37658
rect 142718 37606 142770 37658
rect 142770 37606 142772 37658
rect 142716 37604 142772 37606
rect 142820 37658 142876 37660
rect 142820 37606 142822 37658
rect 142822 37606 142874 37658
rect 142874 37606 142876 37658
rect 142820 37604 142876 37606
rect 142924 37658 142980 37660
rect 142924 37606 142926 37658
rect 142926 37606 142978 37658
rect 142978 37606 142980 37658
rect 142924 37604 142980 37606
rect 142716 36090 142772 36092
rect 142716 36038 142718 36090
rect 142718 36038 142770 36090
rect 142770 36038 142772 36090
rect 142716 36036 142772 36038
rect 142820 36090 142876 36092
rect 142820 36038 142822 36090
rect 142822 36038 142874 36090
rect 142874 36038 142876 36090
rect 142820 36036 142876 36038
rect 142924 36090 142980 36092
rect 142924 36038 142926 36090
rect 142926 36038 142978 36090
rect 142978 36038 142980 36090
rect 142924 36036 142980 36038
rect 142716 34522 142772 34524
rect 142716 34470 142718 34522
rect 142718 34470 142770 34522
rect 142770 34470 142772 34522
rect 142716 34468 142772 34470
rect 142820 34522 142876 34524
rect 142820 34470 142822 34522
rect 142822 34470 142874 34522
rect 142874 34470 142876 34522
rect 142820 34468 142876 34470
rect 142924 34522 142980 34524
rect 142924 34470 142926 34522
rect 142926 34470 142978 34522
rect 142978 34470 142980 34522
rect 142924 34468 142980 34470
rect 142716 32954 142772 32956
rect 142716 32902 142718 32954
rect 142718 32902 142770 32954
rect 142770 32902 142772 32954
rect 142716 32900 142772 32902
rect 142820 32954 142876 32956
rect 142820 32902 142822 32954
rect 142822 32902 142874 32954
rect 142874 32902 142876 32954
rect 142820 32900 142876 32902
rect 142924 32954 142980 32956
rect 142924 32902 142926 32954
rect 142926 32902 142978 32954
rect 142978 32902 142980 32954
rect 142924 32900 142980 32902
rect 142716 31386 142772 31388
rect 142716 31334 142718 31386
rect 142718 31334 142770 31386
rect 142770 31334 142772 31386
rect 142716 31332 142772 31334
rect 142820 31386 142876 31388
rect 142820 31334 142822 31386
rect 142822 31334 142874 31386
rect 142874 31334 142876 31386
rect 142820 31332 142876 31334
rect 142924 31386 142980 31388
rect 142924 31334 142926 31386
rect 142926 31334 142978 31386
rect 142978 31334 142980 31386
rect 142924 31332 142980 31334
rect 142716 29818 142772 29820
rect 142716 29766 142718 29818
rect 142718 29766 142770 29818
rect 142770 29766 142772 29818
rect 142716 29764 142772 29766
rect 142820 29818 142876 29820
rect 142820 29766 142822 29818
rect 142822 29766 142874 29818
rect 142874 29766 142876 29818
rect 142820 29764 142876 29766
rect 142924 29818 142980 29820
rect 142924 29766 142926 29818
rect 142926 29766 142978 29818
rect 142978 29766 142980 29818
rect 142924 29764 142980 29766
rect 142716 28250 142772 28252
rect 142716 28198 142718 28250
rect 142718 28198 142770 28250
rect 142770 28198 142772 28250
rect 142716 28196 142772 28198
rect 142820 28250 142876 28252
rect 142820 28198 142822 28250
rect 142822 28198 142874 28250
rect 142874 28198 142876 28250
rect 142820 28196 142876 28198
rect 142924 28250 142980 28252
rect 142924 28198 142926 28250
rect 142926 28198 142978 28250
rect 142978 28198 142980 28250
rect 142924 28196 142980 28198
rect 142716 26682 142772 26684
rect 142716 26630 142718 26682
rect 142718 26630 142770 26682
rect 142770 26630 142772 26682
rect 142716 26628 142772 26630
rect 142820 26682 142876 26684
rect 142820 26630 142822 26682
rect 142822 26630 142874 26682
rect 142874 26630 142876 26682
rect 142820 26628 142876 26630
rect 142924 26682 142980 26684
rect 142924 26630 142926 26682
rect 142926 26630 142978 26682
rect 142978 26630 142980 26682
rect 142924 26628 142980 26630
rect 142716 25114 142772 25116
rect 142716 25062 142718 25114
rect 142718 25062 142770 25114
rect 142770 25062 142772 25114
rect 142716 25060 142772 25062
rect 142820 25114 142876 25116
rect 142820 25062 142822 25114
rect 142822 25062 142874 25114
rect 142874 25062 142876 25114
rect 142820 25060 142876 25062
rect 142924 25114 142980 25116
rect 142924 25062 142926 25114
rect 142926 25062 142978 25114
rect 142978 25062 142980 25114
rect 142924 25060 142980 25062
rect 142716 23546 142772 23548
rect 142716 23494 142718 23546
rect 142718 23494 142770 23546
rect 142770 23494 142772 23546
rect 142716 23492 142772 23494
rect 142820 23546 142876 23548
rect 142820 23494 142822 23546
rect 142822 23494 142874 23546
rect 142874 23494 142876 23546
rect 142820 23492 142876 23494
rect 142924 23546 142980 23548
rect 142924 23494 142926 23546
rect 142926 23494 142978 23546
rect 142978 23494 142980 23546
rect 142924 23492 142980 23494
rect 142716 21978 142772 21980
rect 142716 21926 142718 21978
rect 142718 21926 142770 21978
rect 142770 21926 142772 21978
rect 142716 21924 142772 21926
rect 142820 21978 142876 21980
rect 142820 21926 142822 21978
rect 142822 21926 142874 21978
rect 142874 21926 142876 21978
rect 142820 21924 142876 21926
rect 142924 21978 142980 21980
rect 142924 21926 142926 21978
rect 142926 21926 142978 21978
rect 142978 21926 142980 21978
rect 142924 21924 142980 21926
rect 142716 20410 142772 20412
rect 142716 20358 142718 20410
rect 142718 20358 142770 20410
rect 142770 20358 142772 20410
rect 142716 20356 142772 20358
rect 142820 20410 142876 20412
rect 142820 20358 142822 20410
rect 142822 20358 142874 20410
rect 142874 20358 142876 20410
rect 142820 20356 142876 20358
rect 142924 20410 142980 20412
rect 142924 20358 142926 20410
rect 142926 20358 142978 20410
rect 142978 20358 142980 20410
rect 142924 20356 142980 20358
rect 142716 18842 142772 18844
rect 142716 18790 142718 18842
rect 142718 18790 142770 18842
rect 142770 18790 142772 18842
rect 142716 18788 142772 18790
rect 142820 18842 142876 18844
rect 142820 18790 142822 18842
rect 142822 18790 142874 18842
rect 142874 18790 142876 18842
rect 142820 18788 142876 18790
rect 142924 18842 142980 18844
rect 142924 18790 142926 18842
rect 142926 18790 142978 18842
rect 142978 18790 142980 18842
rect 142924 18788 142980 18790
rect 142716 17274 142772 17276
rect 142716 17222 142718 17274
rect 142718 17222 142770 17274
rect 142770 17222 142772 17274
rect 142716 17220 142772 17222
rect 142820 17274 142876 17276
rect 142820 17222 142822 17274
rect 142822 17222 142874 17274
rect 142874 17222 142876 17274
rect 142820 17220 142876 17222
rect 142924 17274 142980 17276
rect 142924 17222 142926 17274
rect 142926 17222 142978 17274
rect 142978 17222 142980 17274
rect 142924 17220 142980 17222
rect 142604 16156 142660 16212
rect 158076 54122 158132 54124
rect 158076 54070 158078 54122
rect 158078 54070 158130 54122
rect 158130 54070 158132 54122
rect 158076 54068 158132 54070
rect 158180 54122 158236 54124
rect 158180 54070 158182 54122
rect 158182 54070 158234 54122
rect 158234 54070 158236 54122
rect 158180 54068 158236 54070
rect 158284 54122 158340 54124
rect 158284 54070 158286 54122
rect 158286 54070 158338 54122
rect 158338 54070 158340 54122
rect 158284 54068 158340 54070
rect 158076 52554 158132 52556
rect 158076 52502 158078 52554
rect 158078 52502 158130 52554
rect 158130 52502 158132 52554
rect 158076 52500 158132 52502
rect 158180 52554 158236 52556
rect 158180 52502 158182 52554
rect 158182 52502 158234 52554
rect 158234 52502 158236 52554
rect 158180 52500 158236 52502
rect 158284 52554 158340 52556
rect 158284 52502 158286 52554
rect 158286 52502 158338 52554
rect 158338 52502 158340 52554
rect 158284 52500 158340 52502
rect 158076 50986 158132 50988
rect 158076 50934 158078 50986
rect 158078 50934 158130 50986
rect 158130 50934 158132 50986
rect 158076 50932 158132 50934
rect 158180 50986 158236 50988
rect 158180 50934 158182 50986
rect 158182 50934 158234 50986
rect 158234 50934 158236 50986
rect 158180 50932 158236 50934
rect 158284 50986 158340 50988
rect 158284 50934 158286 50986
rect 158286 50934 158338 50986
rect 158338 50934 158340 50986
rect 158284 50932 158340 50934
rect 158076 49418 158132 49420
rect 158076 49366 158078 49418
rect 158078 49366 158130 49418
rect 158130 49366 158132 49418
rect 158076 49364 158132 49366
rect 158180 49418 158236 49420
rect 158180 49366 158182 49418
rect 158182 49366 158234 49418
rect 158234 49366 158236 49418
rect 158180 49364 158236 49366
rect 158284 49418 158340 49420
rect 158284 49366 158286 49418
rect 158286 49366 158338 49418
rect 158338 49366 158340 49418
rect 158284 49364 158340 49366
rect 158076 47850 158132 47852
rect 158076 47798 158078 47850
rect 158078 47798 158130 47850
rect 158130 47798 158132 47850
rect 158076 47796 158132 47798
rect 158180 47850 158236 47852
rect 158180 47798 158182 47850
rect 158182 47798 158234 47850
rect 158234 47798 158236 47850
rect 158180 47796 158236 47798
rect 158284 47850 158340 47852
rect 158284 47798 158286 47850
rect 158286 47798 158338 47850
rect 158338 47798 158340 47850
rect 158284 47796 158340 47798
rect 158076 46282 158132 46284
rect 158076 46230 158078 46282
rect 158078 46230 158130 46282
rect 158130 46230 158132 46282
rect 158076 46228 158132 46230
rect 158180 46282 158236 46284
rect 158180 46230 158182 46282
rect 158182 46230 158234 46282
rect 158234 46230 158236 46282
rect 158180 46228 158236 46230
rect 158284 46282 158340 46284
rect 158284 46230 158286 46282
rect 158286 46230 158338 46282
rect 158338 46230 158340 46282
rect 158284 46228 158340 46230
rect 158076 44714 158132 44716
rect 158076 44662 158078 44714
rect 158078 44662 158130 44714
rect 158130 44662 158132 44714
rect 158076 44660 158132 44662
rect 158180 44714 158236 44716
rect 158180 44662 158182 44714
rect 158182 44662 158234 44714
rect 158234 44662 158236 44714
rect 158180 44660 158236 44662
rect 158284 44714 158340 44716
rect 158284 44662 158286 44714
rect 158286 44662 158338 44714
rect 158338 44662 158340 44714
rect 158284 44660 158340 44662
rect 158076 43146 158132 43148
rect 158076 43094 158078 43146
rect 158078 43094 158130 43146
rect 158130 43094 158132 43146
rect 158076 43092 158132 43094
rect 158180 43146 158236 43148
rect 158180 43094 158182 43146
rect 158182 43094 158234 43146
rect 158234 43094 158236 43146
rect 158180 43092 158236 43094
rect 158284 43146 158340 43148
rect 158284 43094 158286 43146
rect 158286 43094 158338 43146
rect 158338 43094 158340 43146
rect 158284 43092 158340 43094
rect 158076 41578 158132 41580
rect 158076 41526 158078 41578
rect 158078 41526 158130 41578
rect 158130 41526 158132 41578
rect 158076 41524 158132 41526
rect 158180 41578 158236 41580
rect 158180 41526 158182 41578
rect 158182 41526 158234 41578
rect 158234 41526 158236 41578
rect 158180 41524 158236 41526
rect 158284 41578 158340 41580
rect 158284 41526 158286 41578
rect 158286 41526 158338 41578
rect 158338 41526 158340 41578
rect 158284 41524 158340 41526
rect 158076 40010 158132 40012
rect 158076 39958 158078 40010
rect 158078 39958 158130 40010
rect 158130 39958 158132 40010
rect 158076 39956 158132 39958
rect 158180 40010 158236 40012
rect 158180 39958 158182 40010
rect 158182 39958 158234 40010
rect 158234 39958 158236 40010
rect 158180 39956 158236 39958
rect 158284 40010 158340 40012
rect 158284 39958 158286 40010
rect 158286 39958 158338 40010
rect 158338 39958 158340 40010
rect 158284 39956 158340 39958
rect 158076 38442 158132 38444
rect 158076 38390 158078 38442
rect 158078 38390 158130 38442
rect 158130 38390 158132 38442
rect 158076 38388 158132 38390
rect 158180 38442 158236 38444
rect 158180 38390 158182 38442
rect 158182 38390 158234 38442
rect 158234 38390 158236 38442
rect 158180 38388 158236 38390
rect 158284 38442 158340 38444
rect 158284 38390 158286 38442
rect 158286 38390 158338 38442
rect 158338 38390 158340 38442
rect 158284 38388 158340 38390
rect 158076 36874 158132 36876
rect 158076 36822 158078 36874
rect 158078 36822 158130 36874
rect 158130 36822 158132 36874
rect 158076 36820 158132 36822
rect 158180 36874 158236 36876
rect 158180 36822 158182 36874
rect 158182 36822 158234 36874
rect 158234 36822 158236 36874
rect 158180 36820 158236 36822
rect 158284 36874 158340 36876
rect 158284 36822 158286 36874
rect 158286 36822 158338 36874
rect 158338 36822 158340 36874
rect 158284 36820 158340 36822
rect 158076 35306 158132 35308
rect 158076 35254 158078 35306
rect 158078 35254 158130 35306
rect 158130 35254 158132 35306
rect 158076 35252 158132 35254
rect 158180 35306 158236 35308
rect 158180 35254 158182 35306
rect 158182 35254 158234 35306
rect 158234 35254 158236 35306
rect 158180 35252 158236 35254
rect 158284 35306 158340 35308
rect 158284 35254 158286 35306
rect 158286 35254 158338 35306
rect 158338 35254 158340 35306
rect 158284 35252 158340 35254
rect 158076 33738 158132 33740
rect 158076 33686 158078 33738
rect 158078 33686 158130 33738
rect 158130 33686 158132 33738
rect 158076 33684 158132 33686
rect 158180 33738 158236 33740
rect 158180 33686 158182 33738
rect 158182 33686 158234 33738
rect 158234 33686 158236 33738
rect 158180 33684 158236 33686
rect 158284 33738 158340 33740
rect 158284 33686 158286 33738
rect 158286 33686 158338 33738
rect 158338 33686 158340 33738
rect 158284 33684 158340 33686
rect 158076 32170 158132 32172
rect 158076 32118 158078 32170
rect 158078 32118 158130 32170
rect 158130 32118 158132 32170
rect 158076 32116 158132 32118
rect 158180 32170 158236 32172
rect 158180 32118 158182 32170
rect 158182 32118 158234 32170
rect 158234 32118 158236 32170
rect 158180 32116 158236 32118
rect 158284 32170 158340 32172
rect 158284 32118 158286 32170
rect 158286 32118 158338 32170
rect 158338 32118 158340 32170
rect 158284 32116 158340 32118
rect 158076 30602 158132 30604
rect 158076 30550 158078 30602
rect 158078 30550 158130 30602
rect 158130 30550 158132 30602
rect 158076 30548 158132 30550
rect 158180 30602 158236 30604
rect 158180 30550 158182 30602
rect 158182 30550 158234 30602
rect 158234 30550 158236 30602
rect 158180 30548 158236 30550
rect 158284 30602 158340 30604
rect 158284 30550 158286 30602
rect 158286 30550 158338 30602
rect 158338 30550 158340 30602
rect 158284 30548 158340 30550
rect 158076 29034 158132 29036
rect 158076 28982 158078 29034
rect 158078 28982 158130 29034
rect 158130 28982 158132 29034
rect 158076 28980 158132 28982
rect 158180 29034 158236 29036
rect 158180 28982 158182 29034
rect 158182 28982 158234 29034
rect 158234 28982 158236 29034
rect 158180 28980 158236 28982
rect 158284 29034 158340 29036
rect 158284 28982 158286 29034
rect 158286 28982 158338 29034
rect 158338 28982 158340 29034
rect 158284 28980 158340 28982
rect 158076 27466 158132 27468
rect 158076 27414 158078 27466
rect 158078 27414 158130 27466
rect 158130 27414 158132 27466
rect 158076 27412 158132 27414
rect 158180 27466 158236 27468
rect 158180 27414 158182 27466
rect 158182 27414 158234 27466
rect 158234 27414 158236 27466
rect 158180 27412 158236 27414
rect 158284 27466 158340 27468
rect 158284 27414 158286 27466
rect 158286 27414 158338 27466
rect 158338 27414 158340 27466
rect 158284 27412 158340 27414
rect 158076 25898 158132 25900
rect 158076 25846 158078 25898
rect 158078 25846 158130 25898
rect 158130 25846 158132 25898
rect 158076 25844 158132 25846
rect 158180 25898 158236 25900
rect 158180 25846 158182 25898
rect 158182 25846 158234 25898
rect 158234 25846 158236 25898
rect 158180 25844 158236 25846
rect 158284 25898 158340 25900
rect 158284 25846 158286 25898
rect 158286 25846 158338 25898
rect 158338 25846 158340 25898
rect 158284 25844 158340 25846
rect 158076 24330 158132 24332
rect 158076 24278 158078 24330
rect 158078 24278 158130 24330
rect 158130 24278 158132 24330
rect 158076 24276 158132 24278
rect 158180 24330 158236 24332
rect 158180 24278 158182 24330
rect 158182 24278 158234 24330
rect 158234 24278 158236 24330
rect 158180 24276 158236 24278
rect 158284 24330 158340 24332
rect 158284 24278 158286 24330
rect 158286 24278 158338 24330
rect 158338 24278 158340 24330
rect 158284 24276 158340 24278
rect 158076 22762 158132 22764
rect 158076 22710 158078 22762
rect 158078 22710 158130 22762
rect 158130 22710 158132 22762
rect 158076 22708 158132 22710
rect 158180 22762 158236 22764
rect 158180 22710 158182 22762
rect 158182 22710 158234 22762
rect 158234 22710 158236 22762
rect 158180 22708 158236 22710
rect 158284 22762 158340 22764
rect 158284 22710 158286 22762
rect 158286 22710 158338 22762
rect 158338 22710 158340 22762
rect 158284 22708 158340 22710
rect 158076 21194 158132 21196
rect 158076 21142 158078 21194
rect 158078 21142 158130 21194
rect 158130 21142 158132 21194
rect 158076 21140 158132 21142
rect 158180 21194 158236 21196
rect 158180 21142 158182 21194
rect 158182 21142 158234 21194
rect 158234 21142 158236 21194
rect 158180 21140 158236 21142
rect 158284 21194 158340 21196
rect 158284 21142 158286 21194
rect 158286 21142 158338 21194
rect 158338 21142 158340 21194
rect 158284 21140 158340 21142
rect 158076 19626 158132 19628
rect 158076 19574 158078 19626
rect 158078 19574 158130 19626
rect 158130 19574 158132 19626
rect 158076 19572 158132 19574
rect 158180 19626 158236 19628
rect 158180 19574 158182 19626
rect 158182 19574 158234 19626
rect 158234 19574 158236 19626
rect 158180 19572 158236 19574
rect 158284 19626 158340 19628
rect 158284 19574 158286 19626
rect 158286 19574 158338 19626
rect 158338 19574 158340 19626
rect 158284 19572 158340 19574
rect 158076 18058 158132 18060
rect 158076 18006 158078 18058
rect 158078 18006 158130 18058
rect 158130 18006 158132 18058
rect 158076 18004 158132 18006
rect 158180 18058 158236 18060
rect 158180 18006 158182 18058
rect 158182 18006 158234 18058
rect 158234 18006 158236 18058
rect 158180 18004 158236 18006
rect 158284 18058 158340 18060
rect 158284 18006 158286 18058
rect 158286 18006 158338 18058
rect 158338 18006 158340 18058
rect 158284 18004 158340 18006
rect 158076 16490 158132 16492
rect 158076 16438 158078 16490
rect 158078 16438 158130 16490
rect 158130 16438 158132 16490
rect 158076 16436 158132 16438
rect 158180 16490 158236 16492
rect 158180 16438 158182 16490
rect 158182 16438 158234 16490
rect 158234 16438 158236 16490
rect 158180 16436 158236 16438
rect 158284 16490 158340 16492
rect 158284 16438 158286 16490
rect 158286 16438 158338 16490
rect 158338 16438 158340 16490
rect 158284 16436 158340 16438
rect 154028 16044 154084 16100
rect 142716 15706 142772 15708
rect 142716 15654 142718 15706
rect 142718 15654 142770 15706
rect 142770 15654 142772 15706
rect 142716 15652 142772 15654
rect 142820 15706 142876 15708
rect 142820 15654 142822 15706
rect 142822 15654 142874 15706
rect 142874 15654 142876 15706
rect 142820 15652 142876 15654
rect 142924 15706 142980 15708
rect 142924 15654 142926 15706
rect 142926 15654 142978 15706
rect 142978 15654 142980 15706
rect 142924 15652 142980 15654
rect 158076 14922 158132 14924
rect 158076 14870 158078 14922
rect 158078 14870 158130 14922
rect 158130 14870 158132 14922
rect 158076 14868 158132 14870
rect 158180 14922 158236 14924
rect 158180 14870 158182 14922
rect 158182 14870 158234 14922
rect 158234 14870 158236 14922
rect 158180 14868 158236 14870
rect 158284 14922 158340 14924
rect 158284 14870 158286 14922
rect 158286 14870 158338 14922
rect 158338 14870 158340 14922
rect 158284 14868 158340 14870
rect 131180 14364 131236 14420
rect 142716 14138 142772 14140
rect 142716 14086 142718 14138
rect 142718 14086 142770 14138
rect 142770 14086 142772 14138
rect 142716 14084 142772 14086
rect 142820 14138 142876 14140
rect 142820 14086 142822 14138
rect 142822 14086 142874 14138
rect 142874 14086 142876 14138
rect 142820 14084 142876 14086
rect 142924 14138 142980 14140
rect 142924 14086 142926 14138
rect 142926 14086 142978 14138
rect 142978 14086 142980 14138
rect 142924 14084 142980 14086
rect 127356 13354 127412 13356
rect 127356 13302 127358 13354
rect 127358 13302 127410 13354
rect 127410 13302 127412 13354
rect 127356 13300 127412 13302
rect 127460 13354 127516 13356
rect 127460 13302 127462 13354
rect 127462 13302 127514 13354
rect 127514 13302 127516 13354
rect 127460 13300 127516 13302
rect 127564 13354 127620 13356
rect 127564 13302 127566 13354
rect 127566 13302 127618 13354
rect 127618 13302 127620 13354
rect 127564 13300 127620 13302
rect 158076 13354 158132 13356
rect 158076 13302 158078 13354
rect 158078 13302 158130 13354
rect 158130 13302 158132 13354
rect 158076 13300 158132 13302
rect 158180 13354 158236 13356
rect 158180 13302 158182 13354
rect 158182 13302 158234 13354
rect 158234 13302 158236 13354
rect 158180 13300 158236 13302
rect 158284 13354 158340 13356
rect 158284 13302 158286 13354
rect 158286 13302 158338 13354
rect 158338 13302 158340 13354
rect 158284 13300 158340 13302
rect 121772 12796 121828 12852
rect 142716 12570 142772 12572
rect 142716 12518 142718 12570
rect 142718 12518 142770 12570
rect 142770 12518 142772 12570
rect 142716 12516 142772 12518
rect 142820 12570 142876 12572
rect 142820 12518 142822 12570
rect 142822 12518 142874 12570
rect 142874 12518 142876 12570
rect 142820 12516 142876 12518
rect 142924 12570 142980 12572
rect 142924 12518 142926 12570
rect 142926 12518 142978 12570
rect 142978 12518 142980 12570
rect 142924 12516 142980 12518
rect 145516 12012 145572 12068
rect 122668 11900 122724 11956
rect 127356 11786 127412 11788
rect 127356 11734 127358 11786
rect 127358 11734 127410 11786
rect 127410 11734 127412 11786
rect 127356 11732 127412 11734
rect 127460 11786 127516 11788
rect 127460 11734 127462 11786
rect 127462 11734 127514 11786
rect 127514 11734 127516 11786
rect 127460 11732 127516 11734
rect 127564 11786 127620 11788
rect 127564 11734 127566 11786
rect 127566 11734 127618 11786
rect 127618 11734 127620 11786
rect 127564 11732 127620 11734
rect 142716 11002 142772 11004
rect 142716 10950 142718 11002
rect 142718 10950 142770 11002
rect 142770 10950 142772 11002
rect 142716 10948 142772 10950
rect 142820 11002 142876 11004
rect 142820 10950 142822 11002
rect 142822 10950 142874 11002
rect 142874 10950 142876 11002
rect 142820 10948 142876 10950
rect 142924 11002 142980 11004
rect 142924 10950 142926 11002
rect 142926 10950 142978 11002
rect 142978 10950 142980 11002
rect 142924 10948 142980 10950
rect 127356 10218 127412 10220
rect 127356 10166 127358 10218
rect 127358 10166 127410 10218
rect 127410 10166 127412 10218
rect 127356 10164 127412 10166
rect 127460 10218 127516 10220
rect 127460 10166 127462 10218
rect 127462 10166 127514 10218
rect 127514 10166 127516 10218
rect 127460 10164 127516 10166
rect 127564 10218 127620 10220
rect 127564 10166 127566 10218
rect 127566 10166 127618 10218
rect 127618 10166 127620 10218
rect 127564 10164 127620 10166
rect 142716 9434 142772 9436
rect 142716 9382 142718 9434
rect 142718 9382 142770 9434
rect 142770 9382 142772 9434
rect 142716 9380 142772 9382
rect 142820 9434 142876 9436
rect 142820 9382 142822 9434
rect 142822 9382 142874 9434
rect 142874 9382 142876 9434
rect 142820 9380 142876 9382
rect 142924 9434 142980 9436
rect 142924 9382 142926 9434
rect 142926 9382 142978 9434
rect 142978 9382 142980 9434
rect 142924 9380 142980 9382
rect 122668 9212 122724 9268
rect 137900 9212 137956 9268
rect 121772 8316 121828 8372
rect 126476 9100 126532 9156
rect 121324 7756 121380 7812
rect 120316 7586 120372 7588
rect 120316 7534 120318 7586
rect 120318 7534 120370 7586
rect 120370 7534 120372 7586
rect 120316 7532 120372 7534
rect 120316 5404 120372 5460
rect 119756 4060 119812 4116
rect 120764 4226 120820 4228
rect 120764 4174 120766 4226
rect 120766 4174 120818 4226
rect 120818 4174 120820 4226
rect 120764 4172 120820 4174
rect 120652 3500 120708 3556
rect 119532 3388 119588 3444
rect 120764 3388 120820 3444
rect 121212 4396 121268 4452
rect 122668 7420 122724 7476
rect 121660 5516 121716 5572
rect 122556 4620 122612 4676
rect 122108 3948 122164 4004
rect 122332 3836 122388 3892
rect 121884 3724 121940 3780
rect 120988 3666 121044 3668
rect 120988 3614 120990 3666
rect 120990 3614 121042 3666
rect 121042 3614 121044 3666
rect 120988 3612 121044 3614
rect 122108 3612 122164 3668
rect 120876 2828 120932 2884
rect 122556 3388 122612 3444
rect 122892 5404 122948 5460
rect 122780 4450 122836 4452
rect 122780 4398 122782 4450
rect 122782 4398 122834 4450
rect 122834 4398 122836 4450
rect 122780 4396 122836 4398
rect 122892 4172 122948 4228
rect 124796 4956 124852 5012
rect 124572 4396 124628 4452
rect 124572 3666 124628 3668
rect 124572 3614 124574 3666
rect 124574 3614 124626 3666
rect 124626 3614 124628 3666
rect 124572 3612 124628 3614
rect 123564 3554 123620 3556
rect 123564 3502 123566 3554
rect 123566 3502 123618 3554
rect 123618 3502 123620 3554
rect 123564 3500 123620 3502
rect 125580 4956 125636 5012
rect 125244 4620 125300 4676
rect 126140 4508 126196 4564
rect 126140 3612 126196 3668
rect 127356 8650 127412 8652
rect 127356 8598 127358 8650
rect 127358 8598 127410 8650
rect 127410 8598 127412 8650
rect 127356 8596 127412 8598
rect 127460 8650 127516 8652
rect 127460 8598 127462 8650
rect 127462 8598 127514 8650
rect 127514 8598 127516 8650
rect 127460 8596 127516 8598
rect 127564 8650 127620 8652
rect 127564 8598 127566 8650
rect 127566 8598 127618 8650
rect 127618 8598 127620 8650
rect 127564 8596 127620 8598
rect 128828 8316 128884 8372
rect 127356 7082 127412 7084
rect 127356 7030 127358 7082
rect 127358 7030 127410 7082
rect 127410 7030 127412 7082
rect 127356 7028 127412 7030
rect 127460 7082 127516 7084
rect 127460 7030 127462 7082
rect 127462 7030 127514 7082
rect 127514 7030 127516 7082
rect 127460 7028 127516 7030
rect 127564 7082 127620 7084
rect 127564 7030 127566 7082
rect 127566 7030 127618 7082
rect 127618 7030 127620 7082
rect 127564 7028 127620 7030
rect 127148 5628 127204 5684
rect 127356 5514 127412 5516
rect 127356 5462 127358 5514
rect 127358 5462 127410 5514
rect 127410 5462 127412 5514
rect 127356 5460 127412 5462
rect 127460 5514 127516 5516
rect 127460 5462 127462 5514
rect 127462 5462 127514 5514
rect 127514 5462 127516 5514
rect 127460 5460 127516 5462
rect 127564 5514 127620 5516
rect 127564 5462 127566 5514
rect 127566 5462 127618 5514
rect 127618 5462 127620 5514
rect 127564 5460 127620 5462
rect 128044 5010 128100 5012
rect 128044 4958 128046 5010
rect 128046 4958 128098 5010
rect 128098 4958 128100 5010
rect 128044 4956 128100 4958
rect 134092 6412 134148 6468
rect 127260 4450 127316 4452
rect 127260 4398 127262 4450
rect 127262 4398 127314 4450
rect 127314 4398 127316 4450
rect 127260 4396 127316 4398
rect 127932 4396 127988 4452
rect 127356 3946 127412 3948
rect 127356 3894 127358 3946
rect 127358 3894 127410 3946
rect 127410 3894 127412 3946
rect 127356 3892 127412 3894
rect 127460 3946 127516 3948
rect 127460 3894 127462 3946
rect 127462 3894 127514 3946
rect 127514 3894 127516 3946
rect 127460 3892 127516 3894
rect 127564 3946 127620 3948
rect 127564 3894 127566 3946
rect 127566 3894 127618 3946
rect 127618 3894 127620 3946
rect 127564 3892 127620 3894
rect 131180 4732 131236 4788
rect 129948 4450 130004 4452
rect 129948 4398 129950 4450
rect 129950 4398 130002 4450
rect 130002 4398 130004 4450
rect 129948 4396 130004 4398
rect 129164 4172 129220 4228
rect 130732 4226 130788 4228
rect 130732 4174 130734 4226
rect 130734 4174 130786 4226
rect 130786 4174 130788 4226
rect 130732 4172 130788 4174
rect 128380 3666 128436 3668
rect 128380 3614 128382 3666
rect 128382 3614 128434 3666
rect 128434 3614 128436 3666
rect 128380 3612 128436 3614
rect 128828 3500 128884 3556
rect 130396 3554 130452 3556
rect 130396 3502 130398 3554
rect 130398 3502 130450 3554
rect 130450 3502 130452 3554
rect 130396 3500 130452 3502
rect 131516 4284 131572 4340
rect 130172 3388 130228 3444
rect 132524 4562 132580 4564
rect 132524 4510 132526 4562
rect 132526 4510 132578 4562
rect 132578 4510 132580 4562
rect 132524 4508 132580 4510
rect 132300 4284 132356 4340
rect 132748 4338 132804 4340
rect 132748 4286 132750 4338
rect 132750 4286 132802 4338
rect 132802 4286 132804 4338
rect 132748 4284 132804 4286
rect 131740 3500 131796 3556
rect 132748 3442 132804 3444
rect 132748 3390 132750 3442
rect 132750 3390 132802 3442
rect 132802 3390 132804 3442
rect 132748 3388 132804 3390
rect 136220 5292 136276 5348
rect 134204 3612 134260 3668
rect 135772 5068 135828 5124
rect 137340 5180 137396 5236
rect 136892 4396 136948 4452
rect 134988 2940 135044 2996
rect 136108 3666 136164 3668
rect 136108 3614 136110 3666
rect 136110 3614 136162 3666
rect 136162 3614 136164 3666
rect 136108 3612 136164 3614
rect 137676 4396 137732 4452
rect 142716 7866 142772 7868
rect 142716 7814 142718 7866
rect 142718 7814 142770 7866
rect 142770 7814 142772 7866
rect 142716 7812 142772 7814
rect 142820 7866 142876 7868
rect 142820 7814 142822 7866
rect 142822 7814 142874 7866
rect 142874 7814 142876 7866
rect 142820 7812 142876 7814
rect 142924 7866 142980 7868
rect 142924 7814 142926 7866
rect 142926 7814 142978 7866
rect 142978 7814 142980 7866
rect 142924 7812 142980 7814
rect 141036 7644 141092 7700
rect 138908 5404 138964 5460
rect 138236 5122 138292 5124
rect 138236 5070 138238 5122
rect 138238 5070 138290 5122
rect 138290 5070 138292 5122
rect 138236 5068 138292 5070
rect 138348 4898 138404 4900
rect 138348 4846 138350 4898
rect 138350 4846 138402 4898
rect 138402 4846 138404 4898
rect 138348 4844 138404 4846
rect 140140 5234 140196 5236
rect 140140 5182 140142 5234
rect 140142 5182 140194 5234
rect 140194 5182 140196 5234
rect 140140 5180 140196 5182
rect 139020 4284 139076 4340
rect 138348 3612 138404 3668
rect 140924 3724 140980 3780
rect 139804 3666 139860 3668
rect 139804 3614 139806 3666
rect 139806 3614 139858 3666
rect 139858 3614 139860 3666
rect 139804 3612 139860 3614
rect 139244 3554 139300 3556
rect 139244 3502 139246 3554
rect 139246 3502 139298 3554
rect 139298 3502 139300 3554
rect 139244 3500 139300 3502
rect 139580 3500 139636 3556
rect 142716 6298 142772 6300
rect 142716 6246 142718 6298
rect 142718 6246 142770 6298
rect 142770 6246 142772 6298
rect 142716 6244 142772 6246
rect 142820 6298 142876 6300
rect 142820 6246 142822 6298
rect 142822 6246 142874 6298
rect 142874 6246 142876 6298
rect 142820 6244 142876 6246
rect 142924 6298 142980 6300
rect 142924 6246 142926 6298
rect 142926 6246 142978 6298
rect 142978 6246 142980 6298
rect 142924 6244 142980 6246
rect 142940 5404 142996 5460
rect 142044 5292 142100 5348
rect 141708 5068 141764 5124
rect 141484 4844 141540 4900
rect 141932 4338 141988 4340
rect 141932 4286 141934 4338
rect 141934 4286 141986 4338
rect 141986 4286 141988 4338
rect 141932 4284 141988 4286
rect 142156 5180 142212 5236
rect 142940 5234 142996 5236
rect 142940 5182 142942 5234
rect 142942 5182 142994 5234
rect 142994 5182 142996 5234
rect 142940 5180 142996 5182
rect 142716 4844 142772 4900
rect 142716 4730 142772 4732
rect 142716 4678 142718 4730
rect 142718 4678 142770 4730
rect 142770 4678 142772 4730
rect 142716 4676 142772 4678
rect 142820 4730 142876 4732
rect 142820 4678 142822 4730
rect 142822 4678 142874 4730
rect 142874 4678 142876 4730
rect 142820 4676 142876 4678
rect 142924 4730 142980 4732
rect 142924 4678 142926 4730
rect 142926 4678 142978 4730
rect 142978 4678 142980 4730
rect 142924 4676 142980 4678
rect 143052 4338 143108 4340
rect 143052 4286 143054 4338
rect 143054 4286 143106 4338
rect 143106 4286 143108 4338
rect 143052 4284 143108 4286
rect 142492 3724 142548 3780
rect 142604 4172 142660 4228
rect 142268 3612 142324 3668
rect 141036 3388 141092 3444
rect 141708 3442 141764 3444
rect 141708 3390 141710 3442
rect 141710 3390 141762 3442
rect 141762 3390 141764 3442
rect 141708 3388 141764 3390
rect 143612 4226 143668 4228
rect 143612 4174 143614 4226
rect 143614 4174 143666 4226
rect 143666 4174 143668 4226
rect 143612 4172 143668 4174
rect 143612 3666 143668 3668
rect 143612 3614 143614 3666
rect 143614 3614 143666 3666
rect 143666 3614 143668 3666
rect 143612 3612 143668 3614
rect 143052 3500 143108 3556
rect 143948 4844 144004 4900
rect 144732 5068 144788 5124
rect 144284 4284 144340 4340
rect 144956 4172 145012 4228
rect 142380 3052 142436 3108
rect 142716 3162 142772 3164
rect 142716 3110 142718 3162
rect 142718 3110 142770 3162
rect 142770 3110 142772 3162
rect 142716 3108 142772 3110
rect 142820 3162 142876 3164
rect 142820 3110 142822 3162
rect 142822 3110 142874 3162
rect 142874 3110 142876 3162
rect 142820 3108 142876 3110
rect 142924 3162 142980 3164
rect 142924 3110 142926 3162
rect 142926 3110 142978 3162
rect 142978 3110 142980 3162
rect 142924 3108 142980 3110
rect 158076 11786 158132 11788
rect 158076 11734 158078 11786
rect 158078 11734 158130 11786
rect 158130 11734 158132 11786
rect 158076 11732 158132 11734
rect 158180 11786 158236 11788
rect 158180 11734 158182 11786
rect 158182 11734 158234 11786
rect 158234 11734 158236 11786
rect 158180 11732 158236 11734
rect 158284 11786 158340 11788
rect 158284 11734 158286 11786
rect 158286 11734 158338 11786
rect 158338 11734 158340 11786
rect 158284 11732 158340 11734
rect 158076 10218 158132 10220
rect 158076 10166 158078 10218
rect 158078 10166 158130 10218
rect 158130 10166 158132 10218
rect 158076 10164 158132 10166
rect 158180 10218 158236 10220
rect 158180 10166 158182 10218
rect 158182 10166 158234 10218
rect 158234 10166 158236 10218
rect 158180 10164 158236 10166
rect 158284 10218 158340 10220
rect 158284 10166 158286 10218
rect 158286 10166 158338 10218
rect 158338 10166 158340 10218
rect 158284 10164 158340 10166
rect 158076 8650 158132 8652
rect 158076 8598 158078 8650
rect 158078 8598 158130 8650
rect 158130 8598 158132 8650
rect 158076 8596 158132 8598
rect 158180 8650 158236 8652
rect 158180 8598 158182 8650
rect 158182 8598 158234 8650
rect 158234 8598 158236 8650
rect 158180 8596 158236 8598
rect 158284 8650 158340 8652
rect 158284 8598 158286 8650
rect 158286 8598 158338 8650
rect 158338 8598 158340 8650
rect 158284 8596 158340 8598
rect 158076 7082 158132 7084
rect 158076 7030 158078 7082
rect 158078 7030 158130 7082
rect 158130 7030 158132 7082
rect 158076 7028 158132 7030
rect 158180 7082 158236 7084
rect 158180 7030 158182 7082
rect 158182 7030 158234 7082
rect 158234 7030 158236 7082
rect 158180 7028 158236 7030
rect 158284 7082 158340 7084
rect 158284 7030 158286 7082
rect 158286 7030 158338 7082
rect 158338 7030 158340 7082
rect 158284 7028 158340 7030
rect 158076 5514 158132 5516
rect 158076 5462 158078 5514
rect 158078 5462 158130 5514
rect 158130 5462 158132 5514
rect 158076 5460 158132 5462
rect 158180 5514 158236 5516
rect 158180 5462 158182 5514
rect 158182 5462 158234 5514
rect 158234 5462 158236 5514
rect 158180 5460 158236 5462
rect 158284 5514 158340 5516
rect 158284 5462 158286 5514
rect 158286 5462 158338 5514
rect 158338 5462 158340 5514
rect 158284 5460 158340 5462
rect 147868 5292 147924 5348
rect 147644 5122 147700 5124
rect 147644 5070 147646 5122
rect 147646 5070 147698 5122
rect 147698 5070 147700 5122
rect 147644 5068 147700 5070
rect 147532 4226 147588 4228
rect 147532 4174 147534 4226
rect 147534 4174 147586 4226
rect 147586 4174 147588 4226
rect 147532 4172 147588 4174
rect 145852 3554 145908 3556
rect 145852 3502 145854 3554
rect 145854 3502 145906 3554
rect 145906 3502 145908 3554
rect 145852 3500 145908 3502
rect 145964 2716 146020 2772
rect 146300 3388 146356 3444
rect 147532 3388 147588 3444
rect 148092 5122 148148 5124
rect 148092 5070 148094 5122
rect 148094 5070 148146 5122
rect 148146 5070 148148 5122
rect 148092 5068 148148 5070
rect 148876 4172 148932 4228
rect 147756 3500 147812 3556
rect 149772 4956 149828 5012
rect 158076 3946 158132 3948
rect 158076 3894 158078 3946
rect 158078 3894 158130 3946
rect 158130 3894 158132 3946
rect 158076 3892 158132 3894
rect 158180 3946 158236 3948
rect 158180 3894 158182 3946
rect 158182 3894 158234 3946
rect 158234 3894 158236 3946
rect 158180 3892 158236 3894
rect 158284 3946 158340 3948
rect 158284 3894 158286 3946
rect 158286 3894 158338 3946
rect 158338 3894 158340 3946
rect 158284 3892 158340 3894
rect 149772 3500 149828 3556
rect 150332 3612 150388 3668
rect 149660 1596 149716 1652
rect 151564 3666 151620 3668
rect 151564 3614 151566 3666
rect 151566 3614 151618 3666
rect 151618 3614 151620 3666
rect 151564 3612 151620 3614
rect 150556 3554 150612 3556
rect 150556 3502 150558 3554
rect 150558 3502 150610 3554
rect 150610 3502 150612 3554
rect 150556 3500 150612 3502
<< metal3 >>
rect 142706 57036 142716 57092
rect 142772 57036 144508 57092
rect 144564 57036 144574 57092
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 81266 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81550 56476
rect 111986 56420 111996 56476
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 112260 56420 112270 56476
rect 142706 56420 142716 56476
rect 142772 56420 142820 56476
rect 142876 56420 142924 56476
rect 142980 56420 142990 56476
rect 28466 56252 28476 56308
rect 28532 56252 29708 56308
rect 29764 56252 29774 56308
rect 51314 56252 51324 56308
rect 51380 56252 52556 56308
rect 52612 56252 52622 56308
rect 62738 56252 62748 56308
rect 62804 56252 63980 56308
rect 64036 56252 64046 56308
rect 70354 56252 70364 56308
rect 70420 56252 71596 56308
rect 71652 56252 71662 56308
rect 81778 56252 81788 56308
rect 81844 56252 83020 56308
rect 83076 56252 83086 56308
rect 93202 56252 93212 56308
rect 93268 56252 94444 56308
rect 94500 56252 94510 56308
rect 97010 56252 97020 56308
rect 97076 56252 98252 56308
rect 98308 56252 98318 56308
rect 104626 56252 104636 56308
rect 104692 56252 105868 56308
rect 105924 56252 105934 56308
rect 108434 56252 108444 56308
rect 108500 56252 109676 56308
rect 109732 56252 109742 56308
rect 116050 56252 116060 56308
rect 116116 56252 117292 56308
rect 117348 56252 117358 56308
rect 119858 56252 119868 56308
rect 119924 56252 121100 56308
rect 121156 56252 121166 56308
rect 127474 56252 127484 56308
rect 127540 56252 128716 56308
rect 128772 56252 128782 56308
rect 131282 56252 131292 56308
rect 131348 56252 132524 56308
rect 132580 56252 132590 56308
rect 138898 56252 138908 56308
rect 138964 56252 140140 56308
rect 140196 56252 140206 56308
rect 150322 56252 150332 56308
rect 150388 56252 151564 56308
rect 151620 56252 151630 56308
rect 154130 56252 154140 56308
rect 154196 56252 155372 56308
rect 155428 56252 155438 56308
rect 6178 56140 6188 56196
rect 6244 56140 9212 56196
rect 9268 56140 9278 56196
rect 67106 56140 67116 56196
rect 67172 56140 68012 56196
rect 68068 56140 68078 56196
rect 110002 56140 110012 56196
rect 110068 56140 112476 56196
rect 112532 56140 112542 56196
rect 115042 56140 115052 56196
rect 115108 56140 123900 56196
rect 123956 56140 123966 56196
rect 50082 56028 50092 56084
rect 50148 56028 51548 56084
rect 51604 56028 51614 56084
rect 61282 56028 61292 56084
rect 61348 56028 62972 56084
rect 63028 56028 63038 56084
rect 19842 55916 19852 55972
rect 19908 55916 20972 55972
rect 21028 55916 27916 55972
rect 27972 55916 27982 55972
rect 42690 55916 42700 55972
rect 42756 55916 43820 55972
rect 43876 55916 43886 55972
rect 125122 55916 125132 55972
rect 125188 55916 135772 55972
rect 135828 55916 135838 55972
rect 136882 55916 136892 55972
rect 136948 55916 147196 55972
rect 147252 55916 147262 55972
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 96626 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96910 55692
rect 127346 55636 127356 55692
rect 127412 55636 127460 55692
rect 127516 55636 127564 55692
rect 127620 55636 127630 55692
rect 158066 55636 158076 55692
rect 158132 55636 158180 55692
rect 158236 55636 158284 55692
rect 158340 55636 158350 55692
rect 149492 55356 149772 55412
rect 149828 55356 150780 55412
rect 150836 55356 150846 55412
rect 60946 55244 60956 55300
rect 61012 55244 61740 55300
rect 61796 55244 62188 55300
rect 62244 55244 62254 55300
rect 62962 55244 62972 55300
rect 63028 55244 69804 55300
rect 69860 55244 71036 55300
rect 71092 55244 115724 55300
rect 115780 55244 115790 55300
rect 149492 55188 149548 55356
rect 70130 55132 70140 55188
rect 70196 55132 70700 55188
rect 70756 55132 71484 55188
rect 71540 55132 81116 55188
rect 81172 55132 81564 55188
rect 81620 55132 92540 55188
rect 92596 55132 92988 55188
rect 93044 55132 103964 55188
rect 104020 55132 104030 55188
rect 126802 55132 126812 55188
rect 126868 55132 127260 55188
rect 127316 55132 138348 55188
rect 138404 55132 139020 55188
rect 139076 55132 149548 55188
rect 28466 55020 28476 55076
rect 28532 55020 29372 55076
rect 29428 55020 29438 55076
rect 43698 55020 43708 55076
rect 43764 55020 49644 55076
rect 49700 55020 49710 55076
rect 50978 55020 50988 55076
rect 51044 55020 59948 55076
rect 60004 55020 60508 55076
rect 60564 55020 60574 55076
rect 94546 55020 94556 55076
rect 94612 55020 96908 55076
rect 96964 55020 97580 55076
rect 97636 55020 97646 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 81266 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81550 54908
rect 111986 54852 111996 54908
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 112260 54852 112270 54908
rect 142706 54852 142716 54908
rect 142772 54852 142820 54908
rect 142876 54852 142924 54908
rect 142980 54852 142990 54908
rect 115826 54348 115836 54404
rect 115892 54348 116620 54404
rect 116676 54348 126812 54404
rect 126868 54348 126878 54404
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 96626 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96910 54124
rect 127346 54068 127356 54124
rect 127412 54068 127460 54124
rect 127516 54068 127564 54124
rect 127620 54068 127630 54124
rect 158066 54068 158076 54124
rect 158132 54068 158180 54124
rect 158236 54068 158284 54124
rect 158340 54068 158350 54124
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 81266 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81550 53340
rect 111986 53284 111996 53340
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 112260 53284 112270 53340
rect 142706 53284 142716 53340
rect 142772 53284 142820 53340
rect 142876 53284 142924 53340
rect 142980 53284 142990 53340
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 96626 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96910 52556
rect 127346 52500 127356 52556
rect 127412 52500 127460 52556
rect 127516 52500 127564 52556
rect 127620 52500 127630 52556
rect 158066 52500 158076 52556
rect 158132 52500 158180 52556
rect 158236 52500 158284 52556
rect 158340 52500 158350 52556
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 81266 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81550 51772
rect 111986 51716 111996 51772
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 112260 51716 112270 51772
rect 142706 51716 142716 51772
rect 142772 51716 142820 51772
rect 142876 51716 142924 51772
rect 142980 51716 142990 51772
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 96626 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96910 50988
rect 127346 50932 127356 50988
rect 127412 50932 127460 50988
rect 127516 50932 127564 50988
rect 127620 50932 127630 50988
rect 158066 50932 158076 50988
rect 158132 50932 158180 50988
rect 158236 50932 158284 50988
rect 158340 50932 158350 50988
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 81266 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81550 50204
rect 111986 50148 111996 50204
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 112260 50148 112270 50204
rect 142706 50148 142716 50204
rect 142772 50148 142820 50204
rect 142876 50148 142924 50204
rect 142980 50148 142990 50204
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 96626 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96910 49420
rect 127346 49364 127356 49420
rect 127412 49364 127460 49420
rect 127516 49364 127564 49420
rect 127620 49364 127630 49420
rect 158066 49364 158076 49420
rect 158132 49364 158180 49420
rect 158236 49364 158284 49420
rect 158340 49364 158350 49420
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 81266 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81550 48636
rect 111986 48580 111996 48636
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 112260 48580 112270 48636
rect 142706 48580 142716 48636
rect 142772 48580 142820 48636
rect 142876 48580 142924 48636
rect 142980 48580 142990 48636
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 96626 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96910 47852
rect 127346 47796 127356 47852
rect 127412 47796 127460 47852
rect 127516 47796 127564 47852
rect 127620 47796 127630 47852
rect 158066 47796 158076 47852
rect 158132 47796 158180 47852
rect 158236 47796 158284 47852
rect 158340 47796 158350 47852
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 81266 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81550 47068
rect 111986 47012 111996 47068
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 112260 47012 112270 47068
rect 142706 47012 142716 47068
rect 142772 47012 142820 47068
rect 142876 47012 142924 47068
rect 142980 47012 142990 47068
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 96626 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96910 46284
rect 127346 46228 127356 46284
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127620 46228 127630 46284
rect 158066 46228 158076 46284
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158340 46228 158350 46284
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 81266 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81550 45500
rect 111986 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112270 45500
rect 142706 45444 142716 45500
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142980 45444 142990 45500
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 96626 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96910 44716
rect 127346 44660 127356 44716
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127620 44660 127630 44716
rect 158066 44660 158076 44716
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158340 44660 158350 44716
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 81266 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81550 43932
rect 111986 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112270 43932
rect 142706 43876 142716 43932
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142980 43876 142990 43932
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 96626 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96910 43148
rect 127346 43092 127356 43148
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127620 43092 127630 43148
rect 158066 43092 158076 43148
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158340 43092 158350 43148
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 81266 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81550 42364
rect 111986 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112270 42364
rect 142706 42308 142716 42364
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142980 42308 142990 42364
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 96626 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96910 41580
rect 127346 41524 127356 41580
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127620 41524 127630 41580
rect 158066 41524 158076 41580
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158340 41524 158350 41580
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 81266 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81550 40796
rect 111986 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112270 40796
rect 142706 40740 142716 40796
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142980 40740 142990 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 96626 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96910 40012
rect 127346 39956 127356 40012
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127620 39956 127630 40012
rect 158066 39956 158076 40012
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158340 39956 158350 40012
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 81266 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81550 39228
rect 111986 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112270 39228
rect 142706 39172 142716 39228
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142980 39172 142990 39228
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 96626 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96910 38444
rect 127346 38388 127356 38444
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127620 38388 127630 38444
rect 158066 38388 158076 38444
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158340 38388 158350 38444
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 81266 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81550 37660
rect 111986 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112270 37660
rect 142706 37604 142716 37660
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142980 37604 142990 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 96626 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96910 36876
rect 127346 36820 127356 36876
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127620 36820 127630 36876
rect 158066 36820 158076 36876
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158340 36820 158350 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 81266 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81550 36092
rect 111986 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112270 36092
rect 142706 36036 142716 36092
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142980 36036 142990 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 96626 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96910 35308
rect 127346 35252 127356 35308
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127620 35252 127630 35308
rect 158066 35252 158076 35308
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158340 35252 158350 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 81266 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81550 34524
rect 111986 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112270 34524
rect 142706 34468 142716 34524
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142980 34468 142990 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 96626 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96910 33740
rect 127346 33684 127356 33740
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127620 33684 127630 33740
rect 158066 33684 158076 33740
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158340 33684 158350 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 81266 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81550 32956
rect 111986 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112270 32956
rect 142706 32900 142716 32956
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142980 32900 142990 32956
rect 107090 32732 107100 32788
rect 107156 32732 125132 32788
rect 125188 32732 125198 32788
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 96626 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96910 32172
rect 127346 32116 127356 32172
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127620 32116 127630 32172
rect 158066 32116 158076 32172
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158340 32116 158350 32172
rect 46834 31948 46844 32004
rect 46900 31948 60956 32004
rect 61012 31948 61022 32004
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 81266 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81550 31388
rect 111986 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112270 31388
rect 142706 31332 142716 31388
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142980 31332 142990 31388
rect 48290 30940 48300 30996
rect 48356 30940 74620 30996
rect 74676 30940 74686 30996
rect 37874 30828 37884 30884
rect 37940 30828 74060 30884
rect 74116 30828 74126 30884
rect 49746 30716 49756 30772
rect 49812 30716 69468 30772
rect 69524 30716 69534 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 96626 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96910 30604
rect 127346 30548 127356 30604
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127620 30548 127630 30604
rect 158066 30548 158076 30604
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158340 30548 158350 30604
rect 68002 30492 68012 30548
rect 68068 30492 73388 30548
rect 73444 30492 73454 30548
rect 51986 30380 51996 30436
rect 52052 30380 89628 30436
rect 89684 30380 89694 30436
rect 32834 30268 32844 30324
rect 32900 30268 91084 30324
rect 91140 30268 91150 30324
rect 54786 30156 54796 30212
rect 54852 30156 55916 30212
rect 55972 30156 55982 30212
rect 49298 29932 49308 29988
rect 49364 29932 51100 29988
rect 51156 29932 52780 29988
rect 52836 29932 54124 29988
rect 54180 29932 55468 29988
rect 55524 29932 55534 29988
rect 62066 29820 62076 29876
rect 62132 29820 62972 29876
rect 63028 29820 63038 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 81266 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81550 29820
rect 111986 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112270 29820
rect 142706 29764 142716 29820
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142980 29764 142990 29820
rect 52098 29484 52108 29540
rect 52164 29484 54572 29540
rect 54628 29484 55020 29540
rect 55076 29484 55086 29540
rect 45154 29372 45164 29428
rect 45220 29372 46172 29428
rect 46228 29372 46238 29428
rect 77186 29372 77196 29428
rect 77252 29372 83244 29428
rect 83300 29372 83310 29428
rect 89170 29372 89180 29428
rect 89236 29372 108332 29428
rect 108388 29372 108398 29428
rect 46050 29260 46060 29316
rect 46116 29260 47292 29316
rect 47348 29260 49084 29316
rect 49140 29260 49150 29316
rect 50978 29260 50988 29316
rect 51044 29260 51772 29316
rect 51828 29260 51838 29316
rect 53890 29260 53900 29316
rect 53956 29260 55244 29316
rect 55300 29260 56588 29316
rect 56644 29260 56654 29316
rect 53788 29148 56812 29204
rect 56868 29148 56878 29204
rect 53788 29092 53844 29148
rect 36866 29036 36876 29092
rect 36932 29036 49420 29092
rect 49476 29036 49486 29092
rect 50530 29036 50540 29092
rect 50596 29036 53788 29092
rect 53844 29036 53854 29092
rect 54908 29036 55804 29092
rect 55860 29036 55870 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 54908 28980 54964 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 96626 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96910 29036
rect 127346 28980 127356 29036
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127620 28980 127630 29036
rect 158066 28980 158076 29036
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158340 28980 158350 29036
rect 49298 28924 49308 28980
rect 49364 28924 54908 28980
rect 54964 28924 54974 28980
rect 55122 28924 55132 28980
rect 55188 28924 56476 28980
rect 56532 28924 59388 28980
rect 59444 28924 59454 28980
rect 43362 28812 43372 28868
rect 43428 28812 68236 28868
rect 68292 28812 68302 28868
rect 53004 28700 53900 28756
rect 53956 28700 53966 28756
rect 55682 28700 55692 28756
rect 55748 28700 57820 28756
rect 57876 28700 58492 28756
rect 58548 28700 59388 28756
rect 59444 28700 59454 28756
rect 62132 28700 88060 28756
rect 88116 28700 88126 28756
rect 53004 28644 53060 28700
rect 62132 28644 62188 28700
rect 49410 28588 49420 28644
rect 49476 28588 53004 28644
rect 53060 28588 53070 28644
rect 53442 28588 53452 28644
rect 53508 28588 54348 28644
rect 54404 28588 54414 28644
rect 55906 28588 55916 28644
rect 55972 28588 56924 28644
rect 56980 28588 56990 28644
rect 57148 28588 62188 28644
rect 108658 28588 108668 28644
rect 108724 28588 115052 28644
rect 115108 28588 115118 28644
rect 57148 28532 57204 28588
rect 48514 28476 48524 28532
rect 48580 28476 49644 28532
rect 49700 28476 49710 28532
rect 49858 28476 49868 28532
rect 49924 28476 50988 28532
rect 51044 28476 51054 28532
rect 55346 28476 55356 28532
rect 55412 28476 57204 28532
rect 46722 28364 46732 28420
rect 46788 28364 49980 28420
rect 50036 28364 50046 28420
rect 57026 28364 57036 28420
rect 57092 28364 57820 28420
rect 57876 28364 57886 28420
rect 58034 28364 58044 28420
rect 58100 28364 59052 28420
rect 59108 28364 59118 28420
rect 67666 28364 67676 28420
rect 67732 28364 69356 28420
rect 69412 28364 72716 28420
rect 72772 28364 72782 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 81266 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81550 28252
rect 111986 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112270 28252
rect 142706 28196 142716 28252
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142980 28196 142990 28252
rect 63196 28140 66108 28196
rect 66164 28140 66174 28196
rect 63196 28084 63252 28140
rect 32610 28028 32620 28084
rect 32676 28028 33404 28084
rect 33460 28028 33470 28084
rect 50306 28028 50316 28084
rect 50372 28028 50540 28084
rect 50596 28028 50606 28084
rect 51090 28028 51100 28084
rect 51156 28028 51436 28084
rect 51492 28028 51502 28084
rect 55356 28028 56364 28084
rect 56420 28028 63196 28084
rect 63252 28028 63262 28084
rect 63634 28028 63644 28084
rect 63700 28028 64764 28084
rect 64820 28028 64830 28084
rect 65650 28028 65660 28084
rect 65716 28028 71372 28084
rect 71428 28028 71438 28084
rect 55356 27972 55412 28028
rect 30930 27916 30940 27972
rect 30996 27916 31612 27972
rect 31668 27916 34188 27972
rect 34244 27916 35756 27972
rect 35812 27916 35822 27972
rect 46050 27916 46060 27972
rect 46116 27916 55412 27972
rect 55570 27916 55580 27972
rect 55636 27916 57148 27972
rect 57204 27916 57214 27972
rect 63746 27916 63756 27972
rect 63812 27916 65324 27972
rect 65380 27916 65996 27972
rect 66052 27916 66062 27972
rect 31714 27804 31724 27860
rect 31780 27804 33180 27860
rect 33236 27804 35868 27860
rect 35924 27804 35934 27860
rect 49634 27804 49644 27860
rect 49700 27804 50316 27860
rect 50372 27804 53228 27860
rect 53284 27804 53294 27860
rect 54338 27804 54348 27860
rect 54404 27804 55132 27860
rect 55188 27804 55198 27860
rect 58818 27804 58828 27860
rect 58884 27804 59836 27860
rect 59892 27804 60620 27860
rect 60676 27804 61068 27860
rect 61124 27804 61134 27860
rect 65090 27804 65100 27860
rect 65156 27804 65884 27860
rect 65940 27804 65950 27860
rect 66210 27804 66220 27860
rect 66276 27804 67228 27860
rect 70354 27804 70364 27860
rect 70420 27804 77308 27860
rect 77364 27804 77374 27860
rect 26898 27692 26908 27748
rect 26964 27692 29820 27748
rect 29876 27692 30156 27748
rect 30212 27692 30222 27748
rect 45042 27692 45052 27748
rect 45108 27692 46172 27748
rect 46228 27692 46238 27748
rect 51314 27692 51324 27748
rect 51380 27692 51772 27748
rect 51828 27692 51838 27748
rect 67172 27636 67228 27804
rect 74274 27692 74284 27748
rect 74340 27692 75852 27748
rect 75908 27692 75918 27748
rect 105746 27692 105756 27748
rect 105812 27692 136892 27748
rect 136948 27692 136958 27748
rect 29698 27580 29708 27636
rect 29764 27580 30716 27636
rect 30772 27580 30782 27636
rect 44818 27580 44828 27636
rect 44884 27580 45724 27636
rect 45780 27580 45790 27636
rect 45938 27580 45948 27636
rect 46004 27580 48860 27636
rect 48916 27580 48926 27636
rect 50082 27580 50092 27636
rect 50148 27580 50764 27636
rect 50820 27580 50830 27636
rect 50978 27580 50988 27636
rect 51044 27580 52108 27636
rect 52164 27580 52174 27636
rect 52658 27580 52668 27636
rect 52724 27580 57820 27636
rect 57876 27580 63308 27636
rect 63364 27580 63374 27636
rect 67172 27580 70700 27636
rect 70756 27580 73948 27636
rect 74004 27580 77196 27636
rect 77252 27580 77644 27636
rect 77700 27580 77710 27636
rect 48626 27468 48636 27524
rect 48692 27468 51100 27524
rect 51156 27468 51548 27524
rect 51604 27468 60844 27524
rect 60900 27468 62748 27524
rect 62804 27468 62814 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 96626 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96910 27468
rect 127346 27412 127356 27468
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127620 27412 127630 27468
rect 158066 27412 158076 27468
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158340 27412 158350 27468
rect 45042 27356 45052 27412
rect 45108 27356 59388 27412
rect 59444 27356 60508 27412
rect 60564 27356 60574 27412
rect 70130 27356 70140 27412
rect 70196 27356 71148 27412
rect 71204 27356 75292 27412
rect 75348 27356 75358 27412
rect 49718 27244 49756 27300
rect 49812 27244 49822 27300
rect 50418 27244 50428 27300
rect 50484 27244 50988 27300
rect 51044 27244 51054 27300
rect 51202 27244 51212 27300
rect 51268 27244 51772 27300
rect 51828 27244 51838 27300
rect 51958 27244 51996 27300
rect 52052 27244 52062 27300
rect 61170 27244 61180 27300
rect 61236 27244 67228 27300
rect 71586 27244 71596 27300
rect 71652 27244 72380 27300
rect 72436 27244 73612 27300
rect 73668 27244 73678 27300
rect 67172 27188 67228 27244
rect 45714 27132 45724 27188
rect 45780 27132 46732 27188
rect 46788 27132 46798 27188
rect 59042 27132 59052 27188
rect 59108 27132 61628 27188
rect 61684 27132 61694 27188
rect 63634 27132 63644 27188
rect 63700 27132 66444 27188
rect 66500 27132 66510 27188
rect 67172 27132 69580 27188
rect 69636 27132 74172 27188
rect 74228 27132 74732 27188
rect 74788 27132 74798 27188
rect 75170 27132 75180 27188
rect 75236 27132 78540 27188
rect 78596 27132 78606 27188
rect 31378 27020 31388 27076
rect 31444 27020 31724 27076
rect 31780 27020 31790 27076
rect 46162 27020 46172 27076
rect 46228 27020 49252 27076
rect 49410 27020 49420 27076
rect 49476 27020 51436 27076
rect 51492 27020 51502 27076
rect 53330 27020 53340 27076
rect 53396 27020 55020 27076
rect 55076 27020 57708 27076
rect 57764 27020 58044 27076
rect 58100 27020 58110 27076
rect 63186 27020 63196 27076
rect 63252 27020 63980 27076
rect 64036 27020 64046 27076
rect 64754 27020 64764 27076
rect 64820 27020 68460 27076
rect 68516 27020 70364 27076
rect 70420 27020 70430 27076
rect 71698 27020 71708 27076
rect 71764 27020 73276 27076
rect 73332 27020 76188 27076
rect 76244 27020 76254 27076
rect 77298 27020 77308 27076
rect 77364 27020 78876 27076
rect 78932 27020 78942 27076
rect 49196 26964 49252 27020
rect 35606 26908 35644 26964
rect 35700 26908 39900 26964
rect 39956 26908 39966 26964
rect 40114 26908 40124 26964
rect 40180 26908 40796 26964
rect 40852 26908 40862 26964
rect 45826 26908 45836 26964
rect 45892 26908 47964 26964
rect 48020 26908 48748 26964
rect 48804 26908 48814 26964
rect 49196 26908 50204 26964
rect 50260 26908 50270 26964
rect 59490 26908 59500 26964
rect 59556 26908 61852 26964
rect 61908 26908 61918 26964
rect 67890 26908 67900 26964
rect 67956 26908 69804 26964
rect 69860 26908 69870 26964
rect 71250 26908 71260 26964
rect 71316 26908 73724 26964
rect 73780 26908 73790 26964
rect 73938 26908 73948 26964
rect 74004 26908 74956 26964
rect 75012 26908 75022 26964
rect 24434 26796 24444 26852
rect 24500 26796 25788 26852
rect 25844 26796 26348 26852
rect 26404 26796 47852 26852
rect 47908 26796 47918 26852
rect 50642 26796 50652 26852
rect 50708 26796 51436 26852
rect 51492 26796 51502 26852
rect 53666 26796 53676 26852
rect 53732 26796 54124 26852
rect 54180 26796 54190 26852
rect 61282 26796 61292 26852
rect 61348 26796 61964 26852
rect 62020 26796 62030 26852
rect 64194 26796 64204 26852
rect 64260 26796 67788 26852
rect 67844 26796 70252 26852
rect 70308 26796 72828 26852
rect 72884 26796 72894 26852
rect 74050 26796 74060 26852
rect 74116 26796 75068 26852
rect 75124 26796 75134 26852
rect 38546 26684 38556 26740
rect 38612 26684 40572 26740
rect 40628 26684 40638 26740
rect 50978 26684 50988 26740
rect 51044 26684 51884 26740
rect 51940 26684 51950 26740
rect 60498 26684 60508 26740
rect 60564 26684 62636 26740
rect 62692 26684 64428 26740
rect 64484 26684 65436 26740
rect 65492 26684 65502 26740
rect 67442 26684 67452 26740
rect 67508 26684 69188 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 69132 26628 69188 26684
rect 81266 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81550 26684
rect 111986 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112270 26684
rect 142706 26628 142716 26684
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142980 26628 142990 26684
rect 25330 26572 25340 26628
rect 25396 26572 26684 26628
rect 26740 26572 27020 26628
rect 27076 26572 28364 26628
rect 28420 26572 28430 26628
rect 31826 26572 31836 26628
rect 31892 26572 38332 26628
rect 38388 26572 38398 26628
rect 38612 26572 45388 26628
rect 45444 26572 45454 26628
rect 49718 26572 49756 26628
rect 49812 26572 49822 26628
rect 53890 26572 53900 26628
rect 53956 26572 54572 26628
rect 54628 26572 54638 26628
rect 56914 26572 56924 26628
rect 56980 26572 58156 26628
rect 58212 26572 58222 26628
rect 63634 26572 63644 26628
rect 63700 26572 67564 26628
rect 67620 26572 68796 26628
rect 68852 26572 68862 26628
rect 69122 26572 69132 26628
rect 69188 26572 70476 26628
rect 70532 26572 70542 26628
rect 38612 26516 38668 26572
rect 26002 26460 26012 26516
rect 26068 26460 27132 26516
rect 27188 26460 38668 26516
rect 39890 26460 39900 26516
rect 39956 26460 41916 26516
rect 41972 26460 41982 26516
rect 48850 26460 48860 26516
rect 48916 26460 50316 26516
rect 50372 26460 50764 26516
rect 50820 26460 50830 26516
rect 63746 26460 63756 26516
rect 63812 26460 67004 26516
rect 67060 26460 69748 26516
rect 71698 26460 71708 26516
rect 71764 26460 72156 26516
rect 72212 26460 86660 26516
rect 69692 26404 69748 26460
rect 34626 26348 34636 26404
rect 34692 26348 36540 26404
rect 36596 26348 36606 26404
rect 38322 26348 38332 26404
rect 38388 26348 38668 26404
rect 39442 26348 39452 26404
rect 39508 26348 40236 26404
rect 40292 26348 42028 26404
rect 42084 26348 42588 26404
rect 42644 26348 43260 26404
rect 43316 26348 43326 26404
rect 49410 26348 49420 26404
rect 49476 26348 49644 26404
rect 49700 26348 50652 26404
rect 50708 26348 50718 26404
rect 53106 26348 53116 26404
rect 53172 26348 53900 26404
rect 53956 26348 54460 26404
rect 54516 26348 55916 26404
rect 55972 26348 55982 26404
rect 58706 26348 58716 26404
rect 58772 26348 68348 26404
rect 68404 26348 69468 26404
rect 69524 26348 69534 26404
rect 69692 26348 73948 26404
rect 74004 26348 74014 26404
rect 38612 26292 38668 26348
rect 24770 26236 24780 26292
rect 24836 26236 25564 26292
rect 25620 26236 25630 26292
rect 30258 26236 30268 26292
rect 30324 26236 30940 26292
rect 30996 26236 31006 26292
rect 35522 26236 35532 26292
rect 35588 26236 37436 26292
rect 37492 26236 37502 26292
rect 37986 26236 37996 26292
rect 38052 26236 38444 26292
rect 38500 26236 38510 26292
rect 38612 26236 39788 26292
rect 39844 26236 39854 26292
rect 40012 26236 41468 26292
rect 41524 26236 41534 26292
rect 42802 26236 42812 26292
rect 42868 26236 43596 26292
rect 43652 26236 44268 26292
rect 44324 26236 44604 26292
rect 44660 26236 44670 26292
rect 48066 26236 48076 26292
rect 48132 26236 48860 26292
rect 48916 26236 50876 26292
rect 50932 26236 50942 26292
rect 55682 26236 55692 26292
rect 55748 26236 56140 26292
rect 56196 26236 57148 26292
rect 57204 26236 58044 26292
rect 58100 26236 58110 26292
rect 61170 26236 61180 26292
rect 61236 26236 61246 26292
rect 61954 26236 61964 26292
rect 62020 26236 63196 26292
rect 63252 26236 63262 26292
rect 72818 26236 72828 26292
rect 72884 26236 73836 26292
rect 73892 26236 73902 26292
rect 74386 26236 74396 26292
rect 74452 26236 75516 26292
rect 75572 26236 75582 26292
rect 40012 26180 40068 26236
rect 61180 26180 61236 26236
rect 86604 26180 86660 26460
rect 35746 26124 35756 26180
rect 35812 26124 36652 26180
rect 36708 26124 36718 26180
rect 37762 26124 37772 26180
rect 37828 26124 39004 26180
rect 39060 26124 39676 26180
rect 39732 26124 40068 26180
rect 41346 26124 41356 26180
rect 41412 26124 44716 26180
rect 44772 26124 44782 26180
rect 49074 26124 49084 26180
rect 49140 26124 49868 26180
rect 49924 26124 49934 26180
rect 50372 26124 61236 26180
rect 71698 26124 71708 26180
rect 71764 26124 76860 26180
rect 76916 26124 77756 26180
rect 77812 26124 86156 26180
rect 86212 26124 86222 26180
rect 86594 26124 86604 26180
rect 86660 26124 104524 26180
rect 104580 26124 104972 26180
rect 105028 26124 105532 26180
rect 105588 26124 105980 26180
rect 106036 26124 106046 26180
rect 50372 26068 50428 26124
rect 86156 26068 86212 26124
rect 30482 26012 30492 26068
rect 30548 26012 31836 26068
rect 31892 26012 34748 26068
rect 34804 26012 35812 26068
rect 36754 26012 36764 26068
rect 36820 26012 37548 26068
rect 37604 26012 37614 26068
rect 48626 26012 48636 26068
rect 48692 26012 48972 26068
rect 49028 26012 50428 26068
rect 50866 26012 50876 26068
rect 50932 26012 51212 26068
rect 51268 26012 51278 26068
rect 52098 26012 52108 26068
rect 52164 26012 52892 26068
rect 52948 26012 52958 26068
rect 59602 26012 59612 26068
rect 59668 26012 60956 26068
rect 61012 26012 61516 26068
rect 61572 26012 61582 26068
rect 86156 26012 86940 26068
rect 86996 26012 87006 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 35756 25844 35812 26012
rect 45154 25900 45164 25956
rect 45220 25900 46508 25956
rect 46564 25900 61180 25956
rect 61236 25900 61246 25956
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 96626 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96910 25900
rect 127346 25844 127356 25900
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127620 25844 127630 25900
rect 158066 25844 158076 25900
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158340 25844 158350 25900
rect 35746 25788 35756 25844
rect 35812 25788 35822 25844
rect 48178 25788 48188 25844
rect 48244 25788 62188 25844
rect 62244 25788 62254 25844
rect 35186 25676 35196 25732
rect 35252 25676 36316 25732
rect 36372 25676 36382 25732
rect 44034 25676 44044 25732
rect 44100 25676 44828 25732
rect 44884 25676 47292 25732
rect 47348 25676 47358 25732
rect 48066 25676 48076 25732
rect 48132 25676 49644 25732
rect 49700 25676 51660 25732
rect 51716 25676 51726 25732
rect 74834 25676 74844 25732
rect 74900 25676 104076 25732
rect 104132 25676 104142 25732
rect 45266 25564 45276 25620
rect 45332 25564 48972 25620
rect 49028 25564 49038 25620
rect 50754 25564 50764 25620
rect 50820 25564 52780 25620
rect 52836 25564 52846 25620
rect 53004 25564 54012 25620
rect 54068 25564 54078 25620
rect 70466 25564 70476 25620
rect 70532 25564 71596 25620
rect 71652 25564 71662 25620
rect 53004 25508 53060 25564
rect 23426 25452 23436 25508
rect 23492 25452 24556 25508
rect 24612 25452 24622 25508
rect 31938 25452 31948 25508
rect 32004 25452 34860 25508
rect 34916 25452 34926 25508
rect 38770 25452 38780 25508
rect 38836 25452 39564 25508
rect 39620 25452 39630 25508
rect 40338 25452 40348 25508
rect 40404 25452 41244 25508
rect 41300 25452 41310 25508
rect 45378 25452 45388 25508
rect 45444 25452 50092 25508
rect 50148 25452 50158 25508
rect 50530 25452 50540 25508
rect 50596 25452 51100 25508
rect 51156 25452 53004 25508
rect 53060 25452 53070 25508
rect 53330 25452 53340 25508
rect 53396 25452 56812 25508
rect 56868 25452 56878 25508
rect 59490 25452 59500 25508
rect 59556 25452 60508 25508
rect 60564 25452 60574 25508
rect 64978 25452 64988 25508
rect 65044 25452 70700 25508
rect 70756 25452 72044 25508
rect 72100 25452 72110 25508
rect 88162 25452 88172 25508
rect 88228 25452 88956 25508
rect 89012 25452 89740 25508
rect 89796 25452 100492 25508
rect 100548 25452 100940 25508
rect 100996 25452 106092 25508
rect 106148 25452 106540 25508
rect 106596 25452 107660 25508
rect 107716 25452 107726 25508
rect 53340 25396 53396 25452
rect 33954 25340 33964 25396
rect 34020 25340 37996 25396
rect 38052 25340 38062 25396
rect 38882 25340 38892 25396
rect 38948 25340 40460 25396
rect 40516 25340 42084 25396
rect 43138 25340 43148 25396
rect 43204 25340 43820 25396
rect 43876 25340 43886 25396
rect 44594 25340 44604 25396
rect 44660 25340 50316 25396
rect 50372 25340 50382 25396
rect 52098 25340 52108 25396
rect 52164 25340 53396 25396
rect 54450 25340 54460 25396
rect 54516 25340 58156 25396
rect 58212 25340 58222 25396
rect 69906 25340 69916 25396
rect 69972 25340 72716 25396
rect 72772 25340 72782 25396
rect 106978 25340 106988 25396
rect 107044 25340 107324 25396
rect 107380 25340 110012 25396
rect 110068 25340 110078 25396
rect 42028 25284 42084 25340
rect 23426 25228 23436 25284
rect 23492 25228 33628 25284
rect 33684 25228 33694 25284
rect 36082 25228 36092 25284
rect 36148 25228 36988 25284
rect 37044 25228 38220 25284
rect 38276 25228 38286 25284
rect 40114 25228 40124 25284
rect 40180 25228 41020 25284
rect 41076 25228 41086 25284
rect 42028 25228 43708 25284
rect 43764 25228 45164 25284
rect 45220 25228 45230 25284
rect 46610 25228 46620 25284
rect 46676 25228 47740 25284
rect 47796 25228 54236 25284
rect 54292 25228 60732 25284
rect 60788 25228 61628 25284
rect 61684 25228 61694 25284
rect 68898 25228 68908 25284
rect 68964 25228 69468 25284
rect 69524 25228 69534 25284
rect 70018 25228 70028 25284
rect 70084 25228 70588 25284
rect 70644 25228 70654 25284
rect 79650 25228 79660 25284
rect 79716 25228 80668 25284
rect 80724 25228 80734 25284
rect 56018 25116 56028 25172
rect 56084 25116 57148 25172
rect 57204 25116 57214 25172
rect 59154 25116 59164 25172
rect 59220 25116 66724 25172
rect 68002 25116 68012 25172
rect 68068 25116 68684 25172
rect 68740 25116 69244 25172
rect 69300 25116 69580 25172
rect 69636 25116 70364 25172
rect 70420 25116 70430 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 59164 25060 59220 25116
rect 38612 25004 39452 25060
rect 39508 25004 39518 25060
rect 51286 25004 51324 25060
rect 51380 25004 59220 25060
rect 28354 24892 28364 24948
rect 28420 24892 31388 24948
rect 31444 24892 38444 24948
rect 38500 24892 38510 24948
rect 38612 24836 38668 25004
rect 66668 24948 66724 25116
rect 81266 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81550 25116
rect 111986 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112270 25116
rect 142706 25060 142716 25116
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142980 25060 142990 25116
rect 69346 25004 69356 25060
rect 69412 25004 72492 25060
rect 72548 25004 72558 25060
rect 74162 25004 74172 25060
rect 74228 25004 76524 25060
rect 76580 25004 80780 25060
rect 80836 25004 80846 25060
rect 45042 24892 45052 24948
rect 45108 24892 46396 24948
rect 46452 24892 46462 24948
rect 48626 24892 48636 24948
rect 48692 24892 50764 24948
rect 50820 24892 51548 24948
rect 51604 24892 51614 24948
rect 55794 24892 55804 24948
rect 55860 24892 58492 24948
rect 58548 24892 59500 24948
rect 59556 24892 59566 24948
rect 60274 24892 60284 24948
rect 60340 24892 62860 24948
rect 62916 24892 64316 24948
rect 64372 24892 65436 24948
rect 65492 24892 65502 24948
rect 66658 24892 66668 24948
rect 66724 24892 66734 24948
rect 68898 24892 68908 24948
rect 68964 24892 71260 24948
rect 71316 24892 72604 24948
rect 72660 24892 72670 24948
rect 74386 24892 74396 24948
rect 74452 24892 74732 24948
rect 74788 24892 75628 24948
rect 75684 24892 75694 24948
rect 78418 24892 78428 24948
rect 78484 24892 79100 24948
rect 79156 24892 80444 24948
rect 80500 24892 80510 24948
rect 31266 24780 31276 24836
rect 31332 24780 31836 24836
rect 31892 24780 31902 24836
rect 35298 24780 35308 24836
rect 35364 24780 35644 24836
rect 35700 24780 35756 24836
rect 35812 24780 35822 24836
rect 36978 24780 36988 24836
rect 37044 24780 38668 24836
rect 45490 24780 45500 24836
rect 45556 24780 46508 24836
rect 46564 24780 55916 24836
rect 55972 24780 55982 24836
rect 57026 24780 57036 24836
rect 57092 24780 58268 24836
rect 58324 24780 58334 24836
rect 64754 24780 64764 24836
rect 64820 24780 71148 24836
rect 71204 24780 71708 24836
rect 71764 24780 71774 24836
rect 74162 24780 74172 24836
rect 74228 24780 74844 24836
rect 74900 24780 74910 24836
rect 81106 24780 81116 24836
rect 81172 24780 81900 24836
rect 81956 24780 81966 24836
rect 32610 24668 32620 24724
rect 32676 24668 34748 24724
rect 34804 24668 34814 24724
rect 36194 24668 36204 24724
rect 36260 24668 37100 24724
rect 37156 24668 40236 24724
rect 40292 24668 40302 24724
rect 41122 24668 41132 24724
rect 41188 24668 50428 24724
rect 50484 24668 50494 24724
rect 50988 24668 51324 24724
rect 51380 24668 51390 24724
rect 55346 24668 55356 24724
rect 55412 24668 56924 24724
rect 56980 24668 57708 24724
rect 57764 24668 58828 24724
rect 58884 24668 58894 24724
rect 67778 24668 67788 24724
rect 67844 24668 68348 24724
rect 68404 24668 68908 24724
rect 68964 24668 70364 24724
rect 70420 24668 70430 24724
rect 73378 24668 73388 24724
rect 73444 24668 74732 24724
rect 74788 24668 74798 24724
rect 76850 24668 76860 24724
rect 76916 24668 78204 24724
rect 78260 24668 78270 24724
rect 82786 24668 82796 24724
rect 82852 24668 83804 24724
rect 83860 24668 83870 24724
rect 50988 24612 51044 24668
rect 26898 24556 26908 24612
rect 26964 24556 27244 24612
rect 27300 24556 30492 24612
rect 30548 24556 30558 24612
rect 32050 24556 32060 24612
rect 32116 24556 36988 24612
rect 37044 24556 37054 24612
rect 49186 24556 49196 24612
rect 49252 24556 49868 24612
rect 49924 24556 51044 24612
rect 51202 24556 51212 24612
rect 51268 24556 51660 24612
rect 51716 24556 51726 24612
rect 65762 24556 65772 24612
rect 65828 24556 69468 24612
rect 69524 24556 69534 24612
rect 75282 24556 75292 24612
rect 75348 24556 92316 24612
rect 92372 24556 92382 24612
rect 36306 24444 36316 24500
rect 36372 24444 37436 24500
rect 37492 24444 37502 24500
rect 38546 24444 38556 24500
rect 38612 24444 52388 24500
rect 52546 24444 52556 24500
rect 52612 24444 53564 24500
rect 53620 24444 53630 24500
rect 66658 24444 66668 24500
rect 66724 24444 71372 24500
rect 71428 24444 71438 24500
rect 52332 24388 52388 24444
rect 44818 24332 44828 24388
rect 44884 24332 52276 24388
rect 52332 24332 55356 24388
rect 55412 24332 55422 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 52220 24276 52276 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 96626 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96910 24332
rect 127346 24276 127356 24332
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127620 24276 127630 24332
rect 158066 24276 158076 24332
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158340 24276 158350 24332
rect 50978 24220 50988 24276
rect 51044 24220 51828 24276
rect 52220 24220 53900 24276
rect 53956 24220 53966 24276
rect 54114 24220 54124 24276
rect 54180 24220 64428 24276
rect 64484 24220 64494 24276
rect 51772 24164 51828 24220
rect 45388 24108 46732 24164
rect 46788 24108 46798 24164
rect 47170 24108 47180 24164
rect 47236 24108 47908 24164
rect 49410 24108 49420 24164
rect 49476 24108 50204 24164
rect 50260 24108 50270 24164
rect 50418 24108 50428 24164
rect 50484 24108 51548 24164
rect 51604 24108 51614 24164
rect 51772 24108 52780 24164
rect 52836 24108 60956 24164
rect 61012 24108 62188 24164
rect 45388 24052 45444 24108
rect 47852 24052 47908 24108
rect 34962 23996 34972 24052
rect 35028 23996 43820 24052
rect 43876 23996 43886 24052
rect 45378 23996 45388 24052
rect 45444 23996 45454 24052
rect 46050 23996 46060 24052
rect 46116 23996 47628 24052
rect 47684 23996 47694 24052
rect 47852 23996 53676 24052
rect 53732 23996 53742 24052
rect 53890 23996 53900 24052
rect 53956 23996 54684 24052
rect 54740 23996 57708 24052
rect 57764 23996 58604 24052
rect 58660 23996 58670 24052
rect 37538 23884 37548 23940
rect 37604 23884 39564 23940
rect 39620 23884 39630 23940
rect 44482 23884 44492 23940
rect 44548 23884 46564 23940
rect 46722 23884 46732 23940
rect 46788 23884 47292 23940
rect 47348 23884 47358 23940
rect 50754 23884 50764 23940
rect 50820 23884 51772 23940
rect 51828 23884 57148 23940
rect 57204 23884 57214 23940
rect 46508 23828 46564 23884
rect 62132 23828 62188 24108
rect 67778 23996 67788 24052
rect 67844 23996 69020 24052
rect 69076 23996 69244 24052
rect 69300 23996 69310 24052
rect 73042 23996 73052 24052
rect 73108 23996 74172 24052
rect 74228 23996 74238 24052
rect 75618 23884 75628 23940
rect 75684 23884 76076 23940
rect 76132 23884 84588 23940
rect 84644 23884 84654 23940
rect 27794 23772 27804 23828
rect 27860 23772 32172 23828
rect 32228 23772 32238 23828
rect 40002 23772 40012 23828
rect 40068 23772 40460 23828
rect 40516 23772 42252 23828
rect 42308 23772 42318 23828
rect 42578 23772 42588 23828
rect 42644 23772 44604 23828
rect 44660 23772 44670 23828
rect 45154 23772 45164 23828
rect 45220 23772 46284 23828
rect 46340 23772 46350 23828
rect 46508 23772 58380 23828
rect 58436 23772 58446 23828
rect 60050 23772 60060 23828
rect 60116 23772 60956 23828
rect 61012 23772 61022 23828
rect 62132 23772 68012 23828
rect 68068 23772 68078 23828
rect 68786 23772 68796 23828
rect 68852 23772 69356 23828
rect 69412 23772 69422 23828
rect 75068 23772 86828 23828
rect 86884 23772 86894 23828
rect 75068 23716 75124 23772
rect 30482 23660 30492 23716
rect 30548 23660 31164 23716
rect 31220 23660 33068 23716
rect 33124 23660 34412 23716
rect 34468 23660 34478 23716
rect 39442 23660 39452 23716
rect 39508 23660 46396 23716
rect 46452 23660 46462 23716
rect 51202 23660 51212 23716
rect 51268 23660 51324 23716
rect 51380 23660 51390 23716
rect 51958 23660 51996 23716
rect 52052 23660 52062 23716
rect 52322 23660 52332 23716
rect 52388 23660 55188 23716
rect 55346 23660 55356 23716
rect 55412 23660 55692 23716
rect 55748 23660 55758 23716
rect 75058 23660 75068 23716
rect 75124 23660 75134 23716
rect 80658 23660 80668 23716
rect 80724 23660 83356 23716
rect 83412 23660 84364 23716
rect 84420 23660 84430 23716
rect 84578 23660 84588 23716
rect 84644 23660 92652 23716
rect 92708 23660 93324 23716
rect 93380 23660 93390 23716
rect 55132 23604 55188 23660
rect 37426 23548 37436 23604
rect 37492 23548 38556 23604
rect 38612 23548 42812 23604
rect 42868 23548 43204 23604
rect 43362 23548 43372 23604
rect 43428 23548 45388 23604
rect 45444 23548 45454 23604
rect 46274 23548 46284 23604
rect 46340 23548 48636 23604
rect 48692 23548 48702 23604
rect 51090 23548 51100 23604
rect 51156 23548 51212 23604
rect 51268 23548 51278 23604
rect 51398 23548 51436 23604
rect 51492 23548 51502 23604
rect 51762 23548 51772 23604
rect 51828 23548 52892 23604
rect 52948 23548 52958 23604
rect 55122 23548 55132 23604
rect 55188 23548 56476 23604
rect 56532 23548 56542 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 43148 23492 43204 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 81266 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81550 23548
rect 111986 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112270 23548
rect 142706 23492 142716 23548
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142980 23492 142990 23548
rect 35634 23436 35644 23492
rect 35700 23436 38332 23492
rect 38388 23436 40796 23492
rect 40852 23436 41916 23492
rect 41972 23436 41982 23492
rect 43148 23436 43708 23492
rect 43764 23436 43774 23492
rect 45042 23436 45052 23492
rect 45108 23436 47180 23492
rect 47236 23436 47246 23492
rect 51538 23436 51548 23492
rect 51604 23436 52220 23492
rect 52276 23436 52286 23492
rect 52770 23436 52780 23492
rect 52836 23436 53676 23492
rect 53732 23436 68572 23492
rect 68628 23436 68638 23492
rect 24658 23324 24668 23380
rect 24724 23324 25340 23380
rect 25396 23324 41132 23380
rect 41188 23324 42028 23380
rect 42084 23324 42094 23380
rect 42364 23324 51660 23380
rect 51716 23324 51726 23380
rect 52630 23324 52668 23380
rect 52724 23324 52734 23380
rect 53666 23324 53676 23380
rect 53732 23324 55692 23380
rect 55748 23324 58268 23380
rect 58324 23324 58334 23380
rect 61394 23324 61404 23380
rect 61460 23324 92092 23380
rect 92148 23324 92158 23380
rect 42364 23268 42420 23324
rect 34066 23212 34076 23268
rect 34132 23212 36428 23268
rect 36484 23212 36494 23268
rect 41010 23212 41020 23268
rect 41076 23212 42140 23268
rect 42196 23212 42206 23268
rect 42354 23212 42364 23268
rect 42420 23212 42430 23268
rect 46946 23212 46956 23268
rect 47012 23212 47852 23268
rect 47908 23212 47918 23268
rect 50306 23212 50316 23268
rect 50372 23212 50596 23268
rect 50540 23156 50596 23212
rect 51100 23212 53900 23268
rect 53956 23212 54684 23268
rect 54740 23212 54750 23268
rect 55234 23212 55244 23268
rect 55300 23212 55804 23268
rect 55860 23212 55870 23268
rect 56028 23212 57820 23268
rect 57876 23212 59948 23268
rect 60004 23212 62188 23268
rect 78306 23212 78316 23268
rect 78372 23212 78988 23268
rect 79044 23212 79054 23268
rect 80210 23212 80220 23268
rect 80276 23212 81564 23268
rect 81620 23212 81630 23268
rect 93314 23212 93324 23268
rect 93380 23212 97468 23268
rect 97524 23212 97534 23268
rect 27234 23100 27244 23156
rect 27300 23100 27804 23156
rect 27860 23100 27870 23156
rect 33506 23100 33516 23156
rect 33572 23100 34188 23156
rect 34244 23100 45276 23156
rect 45332 23100 45342 23156
rect 47618 23100 47628 23156
rect 47684 23100 50428 23156
rect 50540 23100 50876 23156
rect 50932 23100 50942 23156
rect 50372 23044 50428 23100
rect 51100 23044 51156 23212
rect 56028 23156 56084 23212
rect 62132 23156 62188 23212
rect 52546 23100 52556 23156
rect 52612 23100 52892 23156
rect 52948 23100 52958 23156
rect 53330 23100 53340 23156
rect 53396 23100 54012 23156
rect 54068 23100 54078 23156
rect 55010 23100 55020 23156
rect 55076 23100 56084 23156
rect 56914 23100 56924 23156
rect 56980 23100 57932 23156
rect 57988 23100 57998 23156
rect 59826 23100 59836 23156
rect 59892 23100 60284 23156
rect 60340 23100 60350 23156
rect 62132 23100 72268 23156
rect 72324 23100 72334 23156
rect 72482 23100 72492 23156
rect 72548 23100 75628 23156
rect 75684 23100 75694 23156
rect 76514 23100 76524 23156
rect 76580 23100 77532 23156
rect 77588 23100 78428 23156
rect 78484 23100 78494 23156
rect 82226 23100 82236 23156
rect 82292 23100 83580 23156
rect 83636 23100 83646 23156
rect 22530 22988 22540 23044
rect 22596 22988 23324 23044
rect 23380 22988 23390 23044
rect 40786 22988 40796 23044
rect 40852 22988 41804 23044
rect 41860 22988 41870 23044
rect 48178 22988 48188 23044
rect 48244 22988 49532 23044
rect 49588 22988 49598 23044
rect 50372 22988 51156 23044
rect 51314 22988 51324 23044
rect 51380 22988 51884 23044
rect 51940 22988 51950 23044
rect 52098 22988 52108 23044
rect 52164 22988 52174 23044
rect 52322 22988 52332 23044
rect 52388 22988 53116 23044
rect 53172 22988 53182 23044
rect 59154 22988 59164 23044
rect 59220 22988 60396 23044
rect 60452 22988 60462 23044
rect 61058 22988 61068 23044
rect 61124 22988 63084 23044
rect 63140 22988 63150 23044
rect 73042 22988 73052 23044
rect 73108 22988 76188 23044
rect 76244 22988 76254 23044
rect 80882 22988 80892 23044
rect 80948 22988 82684 23044
rect 82740 22988 82750 23044
rect 83346 22988 83356 23044
rect 83412 22988 84476 23044
rect 84532 22988 86156 23044
rect 86212 22988 86222 23044
rect 93090 22988 93100 23044
rect 93156 22988 95340 23044
rect 95396 22988 95406 23044
rect 52108 22932 52164 22988
rect 23762 22876 23772 22932
rect 23828 22876 25340 22932
rect 25396 22876 25406 22932
rect 41906 22876 41916 22932
rect 41972 22876 43484 22932
rect 43540 22876 43550 22932
rect 49074 22876 49084 22932
rect 49140 22876 50652 22932
rect 50708 22876 50718 22932
rect 50866 22876 50876 22932
rect 50932 22876 52164 22932
rect 52434 22876 52444 22932
rect 52500 22876 53564 22932
rect 53620 22876 54348 22932
rect 54404 22876 54414 22932
rect 75142 22876 75180 22932
rect 75236 22876 75246 22932
rect 81666 22876 81676 22932
rect 81732 22876 82124 22932
rect 82180 22876 82190 22932
rect 82450 22876 82460 22932
rect 82516 22876 84028 22932
rect 84084 22876 84094 22932
rect 85652 22876 86716 22932
rect 86772 22876 87388 22932
rect 87444 22876 97132 22932
rect 97188 22876 100828 22932
rect 100884 22876 108892 22932
rect 108948 22876 108958 22932
rect 85652 22820 85708 22876
rect 36978 22764 36988 22820
rect 37044 22764 37996 22820
rect 38052 22764 47404 22820
rect 47460 22764 48076 22820
rect 48132 22764 48142 22820
rect 49522 22764 49532 22820
rect 49588 22764 50540 22820
rect 50596 22764 58940 22820
rect 58996 22764 59006 22820
rect 63858 22764 63868 22820
rect 63924 22764 64764 22820
rect 64820 22764 65324 22820
rect 65380 22764 65390 22820
rect 78866 22764 78876 22820
rect 78932 22764 79548 22820
rect 79604 22764 85708 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 96626 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96910 22764
rect 127346 22708 127356 22764
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127620 22708 127630 22764
rect 158066 22708 158076 22764
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158340 22708 158350 22764
rect 41458 22652 41468 22708
rect 41524 22652 42588 22708
rect 42644 22652 42654 22708
rect 43698 22652 43708 22708
rect 43764 22652 53788 22708
rect 53844 22652 55804 22708
rect 55860 22652 55870 22708
rect 57026 22652 57036 22708
rect 57092 22652 59052 22708
rect 59108 22652 59118 22708
rect 74610 22652 74620 22708
rect 74676 22652 75740 22708
rect 75796 22652 75806 22708
rect 86370 22652 86380 22708
rect 86436 22652 90524 22708
rect 90580 22652 91756 22708
rect 91812 22652 92876 22708
rect 92932 22652 92942 22708
rect 29362 22540 29372 22596
rect 29428 22540 31500 22596
rect 31556 22540 31566 22596
rect 42690 22540 42700 22596
rect 42756 22540 47180 22596
rect 47236 22540 47246 22596
rect 50082 22540 50092 22596
rect 50148 22540 51324 22596
rect 51380 22540 51390 22596
rect 52210 22540 52220 22596
rect 52276 22540 55020 22596
rect 55076 22540 55086 22596
rect 65426 22540 65436 22596
rect 65492 22540 92988 22596
rect 93044 22540 93054 22596
rect 23660 22428 27020 22484
rect 27076 22428 28140 22484
rect 28196 22428 28206 22484
rect 31826 22428 31836 22484
rect 31892 22428 32732 22484
rect 32788 22428 32798 22484
rect 36418 22428 36428 22484
rect 36484 22428 38668 22484
rect 39778 22428 39788 22484
rect 39844 22428 40348 22484
rect 40404 22428 41916 22484
rect 41972 22428 47068 22484
rect 47124 22428 47134 22484
rect 49858 22428 49868 22484
rect 49924 22428 49934 22484
rect 51510 22428 51548 22484
rect 51604 22428 51614 22484
rect 55458 22428 55468 22484
rect 55524 22428 57036 22484
rect 57092 22428 59836 22484
rect 59892 22428 59902 22484
rect 75618 22428 75628 22484
rect 75684 22428 76412 22484
rect 76468 22428 76478 22484
rect 83458 22428 83468 22484
rect 83524 22428 84140 22484
rect 84196 22428 85260 22484
rect 85316 22428 85326 22484
rect 91186 22428 91196 22484
rect 91252 22428 91980 22484
rect 92036 22428 92046 22484
rect 23660 22260 23716 22428
rect 38612 22372 38668 22428
rect 49868 22372 49924 22428
rect 25442 22316 25452 22372
rect 25508 22316 26684 22372
rect 26740 22316 29372 22372
rect 29428 22316 33740 22372
rect 33796 22316 33806 22372
rect 38612 22316 49924 22372
rect 50978 22316 50988 22372
rect 51044 22316 52668 22372
rect 52724 22316 52734 22372
rect 63522 22316 63532 22372
rect 63588 22316 79156 22372
rect 79314 22316 79324 22372
rect 79380 22316 89572 22372
rect 79100 22260 79156 22316
rect 89516 22260 89572 22316
rect 23650 22204 23660 22260
rect 23716 22204 23726 22260
rect 23874 22204 23884 22260
rect 23940 22204 24780 22260
rect 24836 22204 24846 22260
rect 28018 22204 28028 22260
rect 28084 22204 29036 22260
rect 29092 22204 29102 22260
rect 37202 22204 37212 22260
rect 37268 22204 39116 22260
rect 39172 22204 39182 22260
rect 43362 22204 43372 22260
rect 43428 22204 50204 22260
rect 50260 22204 50270 22260
rect 58370 22204 58380 22260
rect 58436 22204 59836 22260
rect 59892 22204 59902 22260
rect 73826 22204 73836 22260
rect 73892 22204 76300 22260
rect 76356 22204 76366 22260
rect 79100 22204 84700 22260
rect 84756 22204 84766 22260
rect 89506 22204 89516 22260
rect 89572 22204 90300 22260
rect 90356 22204 90972 22260
rect 91028 22204 91038 22260
rect 28130 22092 28140 22148
rect 28196 22092 29148 22148
rect 29204 22092 29214 22148
rect 45378 22092 45388 22148
rect 45444 22092 46844 22148
rect 46900 22092 50092 22148
rect 50148 22092 50158 22148
rect 50372 22092 51548 22148
rect 51604 22092 52332 22148
rect 52388 22092 52398 22148
rect 57138 22092 57148 22148
rect 57204 22092 58604 22148
rect 58660 22092 58670 22148
rect 59378 22092 59388 22148
rect 59444 22092 60956 22148
rect 61012 22092 63868 22148
rect 63924 22092 63934 22148
rect 74498 22092 74508 22148
rect 74564 22092 77868 22148
rect 77924 22092 77934 22148
rect 27682 21980 27692 22036
rect 27748 21980 27758 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 26226 21868 26236 21924
rect 26292 21868 26852 21924
rect 26796 21812 26852 21868
rect 27692 21812 27748 21980
rect 50372 21812 50428 22092
rect 51650 21980 51660 22036
rect 51716 21980 52108 22036
rect 52164 21980 52174 22036
rect 92082 21980 92092 22036
rect 92148 21980 92652 22036
rect 92708 21980 92718 22036
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 81266 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81550 21980
rect 111986 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112270 21980
rect 142706 21924 142716 21980
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142980 21924 142990 21980
rect 55794 21868 55804 21924
rect 55860 21868 56588 21924
rect 56644 21868 56654 21924
rect 59042 21868 59052 21924
rect 59108 21868 60060 21924
rect 60116 21868 60126 21924
rect 81666 21868 81676 21924
rect 81732 21868 82684 21924
rect 82740 21868 82750 21924
rect 92306 21868 92316 21924
rect 92372 21868 95228 21924
rect 95284 21868 95294 21924
rect 21074 21756 21084 21812
rect 21140 21756 21868 21812
rect 21924 21756 21934 21812
rect 26796 21756 27748 21812
rect 29810 21756 29820 21812
rect 29876 21756 50204 21812
rect 50260 21756 50428 21812
rect 51958 21756 51996 21812
rect 52052 21756 52062 21812
rect 52658 21756 52668 21812
rect 52724 21756 52892 21812
rect 52948 21756 53676 21812
rect 53732 21756 53742 21812
rect 57362 21756 57372 21812
rect 57428 21756 58828 21812
rect 58884 21756 58894 21812
rect 60834 21756 60844 21812
rect 60900 21756 63644 21812
rect 63700 21756 63710 21812
rect 76402 21756 76412 21812
rect 76468 21756 80220 21812
rect 80276 21756 80286 21812
rect 80434 21756 80444 21812
rect 80500 21756 81452 21812
rect 81508 21756 82012 21812
rect 82068 21756 82078 21812
rect 86930 21756 86940 21812
rect 86996 21756 88396 21812
rect 88452 21756 88462 21812
rect 23986 21644 23996 21700
rect 24052 21644 26012 21700
rect 26068 21644 26078 21700
rect 30706 21644 30716 21700
rect 30772 21644 31612 21700
rect 31668 21644 31678 21700
rect 33394 21644 33404 21700
rect 33460 21644 34412 21700
rect 34468 21644 34478 21700
rect 45602 21644 45612 21700
rect 45668 21644 46620 21700
rect 46676 21644 46686 21700
rect 46834 21644 46844 21700
rect 46900 21644 48748 21700
rect 48804 21644 48814 21700
rect 51090 21644 51100 21700
rect 51156 21644 52668 21700
rect 52724 21644 52734 21700
rect 55346 21644 55356 21700
rect 55412 21644 69132 21700
rect 69188 21644 69198 21700
rect 74722 21644 74732 21700
rect 74788 21644 74956 21700
rect 75012 21644 75022 21700
rect 87154 21644 87164 21700
rect 87220 21644 88508 21700
rect 88564 21644 91868 21700
rect 91924 21644 92764 21700
rect 92820 21644 93772 21700
rect 93828 21644 93838 21700
rect 97458 21644 97468 21700
rect 97524 21644 98140 21700
rect 98196 21644 110852 21700
rect 110796 21588 110852 21644
rect 25890 21532 25900 21588
rect 25956 21532 26684 21588
rect 26740 21532 26908 21588
rect 34626 21532 34636 21588
rect 34692 21532 35644 21588
rect 35700 21532 35710 21588
rect 42018 21532 42028 21588
rect 42084 21532 51212 21588
rect 51268 21532 51278 21588
rect 51762 21532 51772 21588
rect 51828 21532 52556 21588
rect 52612 21532 52622 21588
rect 59490 21532 59500 21588
rect 59556 21532 60956 21588
rect 61012 21532 61022 21588
rect 74162 21532 74172 21588
rect 74228 21532 75404 21588
rect 75460 21532 77420 21588
rect 77476 21532 77486 21588
rect 88722 21532 88732 21588
rect 88788 21532 89740 21588
rect 89796 21532 90524 21588
rect 90580 21532 93212 21588
rect 93268 21532 93278 21588
rect 110786 21532 110796 21588
rect 110852 21532 110862 21588
rect 26852 21476 26908 21532
rect 51772 21476 51828 21532
rect 21858 21420 21868 21476
rect 21924 21420 23324 21476
rect 23380 21420 23390 21476
rect 26852 21420 30044 21476
rect 30100 21420 33628 21476
rect 33684 21420 34412 21476
rect 34468 21420 35532 21476
rect 35588 21420 36652 21476
rect 36708 21420 36718 21476
rect 38612 21420 41468 21476
rect 41524 21420 41534 21476
rect 47058 21420 47068 21476
rect 47124 21420 48188 21476
rect 48244 21420 48860 21476
rect 48916 21420 48926 21476
rect 51314 21420 51324 21476
rect 51380 21420 51828 21476
rect 72818 21420 72828 21476
rect 72884 21420 73948 21476
rect 74004 21420 74014 21476
rect 78530 21420 78540 21476
rect 78596 21420 79548 21476
rect 79604 21420 79614 21476
rect 91186 21420 91196 21476
rect 91252 21420 91980 21476
rect 92036 21420 92046 21476
rect 92530 21420 92540 21476
rect 92596 21420 93548 21476
rect 93604 21420 94444 21476
rect 94500 21420 103964 21476
rect 104020 21420 105420 21476
rect 105476 21420 105486 21476
rect 38612 21364 38668 21420
rect 23986 21308 23996 21364
rect 24052 21308 24444 21364
rect 24500 21308 38668 21364
rect 51548 21308 54908 21364
rect 54964 21308 54974 21364
rect 60610 21308 60620 21364
rect 60676 21308 89628 21364
rect 89684 21308 89694 21364
rect 51548 21252 51604 21308
rect 23874 21196 23884 21252
rect 23940 21196 24220 21252
rect 24276 21196 24286 21252
rect 43922 21196 43932 21252
rect 43988 21196 47068 21252
rect 48738 21196 48748 21252
rect 48804 21196 51604 21252
rect 51762 21196 51772 21252
rect 51828 21196 52332 21252
rect 52388 21196 57372 21252
rect 57428 21196 57438 21252
rect 70466 21196 70476 21252
rect 70532 21196 73948 21252
rect 74004 21196 74014 21252
rect 75506 21196 75516 21252
rect 75572 21196 95004 21252
rect 95060 21196 95070 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 47012 21028 47068 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 96626 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96910 21196
rect 127346 21140 127356 21196
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127620 21140 127630 21196
rect 158066 21140 158076 21196
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158340 21140 158350 21196
rect 47394 21084 47404 21140
rect 47460 21084 53676 21140
rect 53732 21084 53742 21140
rect 55122 21084 55132 21140
rect 55188 21084 56028 21140
rect 56084 21084 64092 21140
rect 64148 21084 64158 21140
rect 91074 21084 91084 21140
rect 91140 21084 92876 21140
rect 92932 21084 93996 21140
rect 94052 21084 94062 21140
rect 23650 20972 23660 21028
rect 23716 20972 25004 21028
rect 25060 20972 27132 21028
rect 27188 20972 27580 21028
rect 27636 20972 27646 21028
rect 47012 20972 50036 21028
rect 50194 20972 50204 21028
rect 50260 20972 63308 21028
rect 63364 20972 63374 21028
rect 68002 20972 68012 21028
rect 68068 20972 92428 21028
rect 92484 20972 92494 21028
rect 92978 20972 92988 21028
rect 93044 20972 93436 21028
rect 93492 20972 93502 21028
rect 49980 20916 50036 20972
rect 21970 20860 21980 20916
rect 22036 20860 24556 20916
rect 24612 20860 25900 20916
rect 25956 20860 25966 20916
rect 41682 20860 41692 20916
rect 41748 20860 45612 20916
rect 45668 20860 45678 20916
rect 45826 20860 45836 20916
rect 45892 20860 47740 20916
rect 47796 20860 47806 20916
rect 49980 20860 51660 20916
rect 51716 20860 51726 20916
rect 52098 20860 52108 20916
rect 52164 20860 52556 20916
rect 52612 20860 52622 20916
rect 57474 20860 57484 20916
rect 57540 20860 58268 20916
rect 58324 20860 59052 20916
rect 59108 20860 59118 20916
rect 59938 20860 59948 20916
rect 60004 20860 60508 20916
rect 60564 20860 60574 20916
rect 64418 20860 64428 20916
rect 64484 20860 66556 20916
rect 66612 20860 66622 20916
rect 77746 20860 77756 20916
rect 77812 20860 79324 20916
rect 79380 20860 79390 20916
rect 85652 20860 91308 20916
rect 91364 20860 95788 20916
rect 95844 20860 95854 20916
rect 96674 20860 96684 20916
rect 96740 20860 97692 20916
rect 97748 20860 97758 20916
rect 51660 20804 51716 20860
rect 28578 20748 28588 20804
rect 28644 20748 29372 20804
rect 29428 20748 30044 20804
rect 30100 20748 30110 20804
rect 44258 20748 44268 20804
rect 44324 20748 45948 20804
rect 46004 20748 46014 20804
rect 46722 20748 46732 20804
rect 46788 20748 51324 20804
rect 51380 20748 51390 20804
rect 51660 20748 52164 20804
rect 53330 20748 53340 20804
rect 53396 20748 54348 20804
rect 54404 20748 54796 20804
rect 54852 20748 54862 20804
rect 59378 20748 59388 20804
rect 59444 20748 59724 20804
rect 59780 20748 60620 20804
rect 60676 20748 60686 20804
rect 60946 20748 60956 20804
rect 61012 20748 64652 20804
rect 64708 20748 65212 20804
rect 65268 20748 65278 20804
rect 77074 20748 77084 20804
rect 77140 20748 78764 20804
rect 78820 20748 81116 20804
rect 81172 20748 81564 20804
rect 81620 20748 81630 20804
rect 52108 20692 52164 20748
rect 85652 20692 85708 20860
rect 92092 20804 92148 20860
rect 86258 20748 86268 20804
rect 86324 20748 87612 20804
rect 87668 20748 87678 20804
rect 92082 20748 92092 20804
rect 92148 20748 92158 20804
rect 92418 20748 92428 20804
rect 92484 20748 92876 20804
rect 92932 20748 92942 20804
rect 37538 20636 37548 20692
rect 37604 20636 38444 20692
rect 38500 20636 38510 20692
rect 44034 20636 44044 20692
rect 44100 20636 45388 20692
rect 45444 20636 46844 20692
rect 46900 20636 48188 20692
rect 48244 20636 48254 20692
rect 50372 20636 51660 20692
rect 51716 20636 51726 20692
rect 52098 20636 52108 20692
rect 52164 20636 54684 20692
rect 54740 20636 55916 20692
rect 55972 20636 55982 20692
rect 75394 20636 75404 20692
rect 75460 20636 85708 20692
rect 50372 20580 50428 20636
rect 47058 20524 47068 20580
rect 47124 20524 50428 20580
rect 50754 20524 50764 20580
rect 50820 20524 52724 20580
rect 52882 20524 52892 20580
rect 52948 20524 57484 20580
rect 57540 20524 57550 20580
rect 58818 20524 58828 20580
rect 58884 20524 59388 20580
rect 59444 20524 59454 20580
rect 74162 20524 74172 20580
rect 74228 20524 74732 20580
rect 74788 20524 75180 20580
rect 75236 20524 75246 20580
rect 78082 20524 78092 20580
rect 78148 20524 78540 20580
rect 78596 20524 78606 20580
rect 80546 20524 80556 20580
rect 80612 20524 81564 20580
rect 81620 20524 81630 20580
rect 93314 20524 93324 20580
rect 93380 20524 93772 20580
rect 93828 20524 95564 20580
rect 95620 20524 96460 20580
rect 96516 20524 99148 20580
rect 99204 20524 101276 20580
rect 101332 20524 103292 20580
rect 103348 20524 107996 20580
rect 108052 20524 111692 20580
rect 111748 20524 111758 20580
rect 52668 20468 52724 20524
rect 52668 20412 52780 20468
rect 52836 20412 52846 20468
rect 59042 20412 59052 20468
rect 59108 20412 59724 20468
rect 59780 20412 59790 20468
rect 64082 20412 64092 20468
rect 64148 20412 66332 20468
rect 66388 20412 66398 20468
rect 77858 20412 77868 20468
rect 77924 20412 78316 20468
rect 78372 20412 78382 20468
rect 92530 20412 92540 20468
rect 92596 20412 92876 20468
rect 92932 20412 92942 20468
rect 97906 20412 97916 20468
rect 97972 20412 98700 20468
rect 98756 20412 98766 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 81266 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81550 20412
rect 111986 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112270 20412
rect 142706 20356 142716 20412
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142980 20356 142990 20412
rect 23874 20300 23884 20356
rect 23940 20300 24668 20356
rect 24724 20300 24734 20356
rect 27906 20300 27916 20356
rect 27972 20300 29148 20356
rect 29204 20300 29214 20356
rect 34850 20300 34860 20356
rect 34916 20300 50428 20356
rect 50372 20244 50428 20300
rect 51996 20300 64484 20356
rect 74386 20300 74396 20356
rect 74452 20300 74620 20356
rect 74676 20300 74686 20356
rect 51996 20244 52052 20300
rect 64428 20244 64484 20300
rect 21970 20188 21980 20244
rect 22036 20188 23324 20244
rect 23380 20188 23390 20244
rect 23986 20188 23996 20244
rect 24052 20188 40012 20244
rect 40068 20188 40078 20244
rect 45602 20188 45612 20244
rect 45668 20188 47292 20244
rect 47348 20188 47358 20244
rect 50372 20188 52052 20244
rect 53330 20188 53340 20244
rect 53396 20188 53564 20244
rect 53620 20188 54124 20244
rect 54180 20188 60732 20244
rect 60788 20188 62524 20244
rect 62580 20188 62590 20244
rect 64428 20188 68908 20244
rect 68964 20188 68974 20244
rect 72930 20188 72940 20244
rect 72996 20188 74844 20244
rect 74900 20188 74910 20244
rect 91858 20188 91868 20244
rect 91924 20188 92988 20244
rect 93044 20188 93054 20244
rect 95778 20188 95788 20244
rect 95844 20188 96796 20244
rect 96852 20188 96862 20244
rect 103058 20188 103068 20244
rect 103124 20188 104188 20244
rect 104244 20188 105756 20244
rect 105812 20188 105822 20244
rect 24322 20076 24332 20132
rect 24388 20076 26460 20132
rect 26516 20076 26526 20132
rect 31714 20076 31724 20132
rect 31780 20076 32284 20132
rect 32340 20076 34188 20132
rect 34244 20076 38108 20132
rect 38164 20076 38174 20132
rect 38434 20076 38444 20132
rect 38500 20076 39004 20132
rect 39060 20076 39070 20132
rect 47954 20076 47964 20132
rect 48020 20076 50204 20132
rect 50260 20076 50270 20132
rect 52994 20076 53004 20132
rect 53060 20076 53070 20132
rect 60050 20076 60060 20132
rect 60116 20076 60956 20132
rect 61012 20076 61022 20132
rect 65314 20076 65324 20132
rect 65380 20076 66892 20132
rect 66948 20076 66958 20132
rect 74582 20076 74620 20132
rect 74676 20076 74686 20132
rect 77186 20076 77196 20132
rect 77252 20076 77756 20132
rect 77812 20076 78652 20132
rect 78708 20076 78718 20132
rect 81778 20076 81788 20132
rect 81844 20076 82236 20132
rect 82292 20076 82302 20132
rect 98018 20076 98028 20132
rect 98084 20076 100828 20132
rect 100884 20076 100894 20132
rect 105858 20076 105868 20132
rect 105924 20076 106652 20132
rect 106708 20076 107772 20132
rect 107828 20076 107838 20132
rect 108546 20076 108556 20132
rect 108612 20076 109228 20132
rect 112466 20076 112476 20132
rect 112532 20076 113372 20132
rect 113428 20076 113438 20132
rect 53004 20020 53060 20076
rect 109172 20020 109228 20076
rect 26226 19964 26236 20020
rect 26292 19964 26302 20020
rect 30258 19964 30268 20020
rect 30324 19964 30940 20020
rect 30996 19964 31006 20020
rect 33394 19964 33404 20020
rect 33460 19964 33852 20020
rect 33908 19964 33918 20020
rect 36082 19964 36092 20020
rect 36148 19964 50428 20020
rect 50866 19964 50876 20020
rect 50932 19964 51884 20020
rect 51940 19964 51950 20020
rect 52210 19964 52220 20020
rect 52276 19964 53060 20020
rect 59154 19964 59164 20020
rect 59220 19964 60172 20020
rect 60228 19964 60238 20020
rect 76514 19964 76524 20020
rect 76580 19964 77644 20020
rect 77700 19964 77710 20020
rect 78764 19964 80892 20020
rect 80948 19964 82572 20020
rect 82628 19964 82638 20020
rect 84018 19964 84028 20020
rect 84084 19964 87948 20020
rect 88004 19964 88014 20020
rect 95218 19964 95228 20020
rect 95284 19964 95788 20020
rect 95844 19964 95854 20020
rect 97010 19964 97020 20020
rect 97076 19964 97468 20020
rect 97524 19964 97534 20020
rect 105186 19964 105196 20020
rect 105252 19964 105980 20020
rect 106036 19964 106046 20020
rect 106418 19964 106428 20020
rect 106484 19964 107212 20020
rect 107268 19964 108220 20020
rect 108276 19964 108286 20020
rect 109172 19964 109788 20020
rect 109844 19964 109854 20020
rect 110002 19964 110012 20020
rect 110068 19964 111356 20020
rect 111412 19964 111422 20020
rect 112354 19964 112364 20020
rect 112420 19964 114268 20020
rect 19842 19852 19852 19908
rect 19908 19852 22764 19908
rect 22820 19852 22830 19908
rect 26236 19796 26292 19964
rect 50372 19908 50428 19964
rect 78764 19908 78820 19964
rect 114212 19908 114268 19964
rect 28578 19852 28588 19908
rect 28644 19852 31164 19908
rect 31220 19852 31230 19908
rect 31602 19852 31612 19908
rect 31668 19852 32396 19908
rect 32452 19852 33628 19908
rect 33684 19852 33694 19908
rect 35858 19852 35868 19908
rect 35924 19852 37100 19908
rect 37156 19852 37166 19908
rect 37986 19852 37996 19908
rect 38052 19852 39004 19908
rect 39060 19852 49084 19908
rect 49140 19852 49150 19908
rect 50372 19852 51996 19908
rect 52052 19852 53900 19908
rect 53956 19852 53966 19908
rect 64988 19852 67004 19908
rect 67060 19852 67070 19908
rect 69906 19852 69916 19908
rect 69972 19852 76748 19908
rect 76804 19852 78820 19908
rect 78876 19852 91756 19908
rect 91812 19852 93212 19908
rect 93268 19852 93278 19908
rect 97412 19852 108780 19908
rect 108836 19852 108846 19908
rect 110226 19852 110236 19908
rect 110292 19852 110908 19908
rect 110964 19852 111916 19908
rect 111972 19852 111982 19908
rect 112466 19852 112476 19908
rect 112532 19852 112924 19908
rect 112980 19852 112990 19908
rect 114212 19852 114940 19908
rect 114996 19852 115006 19908
rect 64988 19796 65044 19852
rect 26236 19740 31948 19796
rect 32004 19740 32172 19796
rect 32228 19740 32238 19796
rect 34066 19740 34076 19796
rect 34132 19740 38668 19796
rect 51426 19740 51436 19796
rect 51492 19740 51772 19796
rect 51828 19740 59836 19796
rect 59892 19740 59902 19796
rect 63858 19740 63868 19796
rect 63924 19740 64988 19796
rect 65044 19740 65054 19796
rect 65548 19740 66220 19796
rect 66276 19740 67676 19796
rect 67732 19740 67742 19796
rect 74162 19740 74172 19796
rect 74228 19740 75852 19796
rect 75908 19740 75918 19796
rect 38612 19684 38668 19740
rect 65548 19684 65604 19740
rect 38612 19628 46284 19684
rect 46340 19628 46350 19684
rect 49186 19628 49196 19684
rect 49252 19628 50204 19684
rect 50260 19628 52892 19684
rect 52948 19628 52958 19684
rect 53106 19628 53116 19684
rect 53172 19628 53564 19684
rect 53620 19628 53630 19684
rect 65426 19628 65436 19684
rect 65492 19628 65604 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 52892 19572 52948 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 78876 19572 78932 19852
rect 97412 19796 97468 19852
rect 81554 19740 81564 19796
rect 81620 19740 82012 19796
rect 82068 19740 91084 19796
rect 91140 19740 91150 19796
rect 96786 19740 96796 19796
rect 96852 19740 97468 19796
rect 107874 19740 107884 19796
rect 107940 19740 110124 19796
rect 110180 19740 110190 19796
rect 110786 19740 110796 19796
rect 110852 19740 113484 19796
rect 113540 19740 113550 19796
rect 81218 19628 81228 19684
rect 81284 19628 81676 19684
rect 81732 19628 82236 19684
rect 82292 19628 82302 19684
rect 86156 19628 94892 19684
rect 94948 19628 94958 19684
rect 109778 19628 109788 19684
rect 109844 19628 112588 19684
rect 112644 19628 112654 19684
rect 40226 19516 40236 19572
rect 40292 19516 41020 19572
rect 41076 19516 42028 19572
rect 42084 19516 43260 19572
rect 43316 19516 43326 19572
rect 44706 19516 44716 19572
rect 44772 19516 52444 19572
rect 52500 19516 52510 19572
rect 52892 19516 58268 19572
rect 58324 19516 58334 19572
rect 59042 19516 59052 19572
rect 59108 19516 59388 19572
rect 59444 19516 62188 19572
rect 68226 19516 68236 19572
rect 68292 19516 78932 19572
rect 62132 19460 62188 19516
rect 86156 19460 86212 19628
rect 96626 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96910 19628
rect 127346 19572 127356 19628
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127620 19572 127630 19628
rect 158066 19572 158076 19628
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158340 19572 158350 19628
rect 27010 19404 27020 19460
rect 27076 19404 28476 19460
rect 28532 19404 39116 19460
rect 39172 19404 42140 19460
rect 42196 19404 42206 19460
rect 50372 19404 53172 19460
rect 53330 19404 53340 19460
rect 53396 19404 55132 19460
rect 55188 19404 55198 19460
rect 57260 19404 59276 19460
rect 59332 19404 59342 19460
rect 62132 19404 67844 19460
rect 71250 19404 71260 19460
rect 71316 19404 86212 19460
rect 86594 19404 86604 19460
rect 86660 19404 87276 19460
rect 87332 19404 87342 19460
rect 33618 19292 33628 19348
rect 33684 19292 34356 19348
rect 37314 19292 37324 19348
rect 37380 19292 38220 19348
rect 38276 19292 38286 19348
rect 42354 19292 42364 19348
rect 42420 19292 43372 19348
rect 43428 19292 43438 19348
rect 34300 19236 34356 19292
rect 50372 19236 50428 19404
rect 53116 19348 53172 19404
rect 57260 19348 57316 19404
rect 51314 19292 51324 19348
rect 51380 19292 52220 19348
rect 52276 19292 52286 19348
rect 53116 19292 57316 19348
rect 57474 19292 57484 19348
rect 57540 19292 66780 19348
rect 66836 19292 66846 19348
rect 67788 19236 67844 19404
rect 68002 19292 68012 19348
rect 68068 19292 85260 19348
rect 85316 19292 86268 19348
rect 86324 19292 86828 19348
rect 86884 19292 86894 19348
rect 95218 19292 95228 19348
rect 95284 19292 96012 19348
rect 96068 19292 96078 19348
rect 104962 19292 104972 19348
rect 105028 19292 105868 19348
rect 105924 19292 106428 19348
rect 106484 19292 106494 19348
rect 111346 19292 111356 19348
rect 111412 19292 114044 19348
rect 114100 19292 114110 19348
rect 23426 19180 23436 19236
rect 23492 19180 23884 19236
rect 23940 19180 24332 19236
rect 24388 19180 24398 19236
rect 31826 19180 31836 19236
rect 31892 19180 33852 19236
rect 33908 19180 33918 19236
rect 34290 19180 34300 19236
rect 34356 19180 37548 19236
rect 37604 19180 37996 19236
rect 38052 19180 38062 19236
rect 39890 19180 39900 19236
rect 39956 19180 43708 19236
rect 43764 19180 43774 19236
rect 46050 19180 46060 19236
rect 46116 19180 48972 19236
rect 49028 19180 49038 19236
rect 49186 19180 49196 19236
rect 49252 19180 50428 19236
rect 51986 19180 51996 19236
rect 52052 19180 55972 19236
rect 56578 19180 56588 19236
rect 56644 19180 62412 19236
rect 62468 19180 62478 19236
rect 64194 19180 64204 19236
rect 64260 19180 64652 19236
rect 64708 19180 64718 19236
rect 66994 19180 67004 19236
rect 67060 19180 67564 19236
rect 67620 19180 67630 19236
rect 67788 19180 68292 19236
rect 68562 19180 68572 19236
rect 68628 19180 71372 19236
rect 71428 19180 72044 19236
rect 72100 19180 72110 19236
rect 73892 19180 109452 19236
rect 109508 19180 110236 19236
rect 110292 19180 110302 19236
rect 112354 19180 112364 19236
rect 112420 19180 113148 19236
rect 113204 19180 113214 19236
rect 55916 19124 55972 19180
rect 25330 19068 25340 19124
rect 25396 19068 27804 19124
rect 27860 19068 28812 19124
rect 28868 19068 30268 19124
rect 30324 19068 30334 19124
rect 41570 19068 41580 19124
rect 41636 19068 42812 19124
rect 42868 19068 43148 19124
rect 43204 19068 43214 19124
rect 49074 19068 49084 19124
rect 49140 19068 53564 19124
rect 53620 19068 54012 19124
rect 54068 19068 54078 19124
rect 55346 19068 55356 19124
rect 55412 19068 55692 19124
rect 55748 19068 55758 19124
rect 55916 19068 58268 19124
rect 58324 19068 58334 19124
rect 60722 19068 60732 19124
rect 60788 19068 62300 19124
rect 62356 19068 62366 19124
rect 64530 19068 64540 19124
rect 64596 19068 65772 19124
rect 65828 19068 66556 19124
rect 66612 19068 66622 19124
rect 68236 19012 68292 19180
rect 73892 19124 73948 19180
rect 73714 19068 73724 19124
rect 73780 19068 73948 19124
rect 74386 19068 74396 19124
rect 74452 19068 75292 19124
rect 75348 19068 75358 19124
rect 91074 19068 91084 19124
rect 91140 19068 91980 19124
rect 92036 19068 92046 19124
rect 99250 19068 99260 19124
rect 99316 19068 99932 19124
rect 99988 19068 99998 19124
rect 104066 19068 104076 19124
rect 104132 19068 104972 19124
rect 105028 19068 106092 19124
rect 106148 19068 107884 19124
rect 107940 19068 107950 19124
rect 31042 18956 31052 19012
rect 31108 18956 32956 19012
rect 33012 18956 33022 19012
rect 38612 18956 45388 19012
rect 45444 18956 46284 19012
rect 46340 18956 46350 19012
rect 49522 18956 49532 19012
rect 49588 18956 49980 19012
rect 50036 18956 50046 19012
rect 50306 18956 50316 19012
rect 50372 18956 51436 19012
rect 51492 18956 51502 19012
rect 53106 18956 53116 19012
rect 53172 18956 56028 19012
rect 56084 18956 56094 19012
rect 60162 18956 60172 19012
rect 60228 18956 61292 19012
rect 61348 18956 61358 19012
rect 68002 18956 68012 19012
rect 68068 18956 68078 19012
rect 68236 18956 73948 19012
rect 74834 18956 74844 19012
rect 74900 18956 75068 19012
rect 75124 18956 76188 19012
rect 76244 18956 76254 19012
rect 85446 18956 85484 19012
rect 85540 18956 85550 19012
rect 86146 18956 86156 19012
rect 86212 18956 86604 19012
rect 86660 18956 88060 19012
rect 88116 18956 88126 19012
rect 91746 18956 91756 19012
rect 91812 18956 92428 19012
rect 92484 18956 92494 19012
rect 96674 18956 96684 19012
rect 96740 18956 97356 19012
rect 97412 18956 98252 19012
rect 98308 18956 98318 19012
rect 98802 18956 98812 19012
rect 98868 18956 100828 19012
rect 100884 18956 100894 19012
rect 114146 18956 114156 19012
rect 114212 18956 116004 19012
rect 38612 18900 38668 18956
rect 68012 18900 68068 18956
rect 29250 18844 29260 18900
rect 29316 18844 38668 18900
rect 58146 18844 58156 18900
rect 58212 18844 68068 18900
rect 68226 18844 68236 18900
rect 68292 18844 68302 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 68236 18788 68292 18844
rect 44706 18732 44716 18788
rect 44772 18732 44782 18788
rect 46834 18732 46844 18788
rect 46900 18732 48412 18788
rect 48468 18732 50428 18788
rect 60610 18732 60620 18788
rect 60676 18732 68292 18788
rect 22866 18620 22876 18676
rect 22932 18620 24444 18676
rect 24500 18620 24780 18676
rect 24836 18620 26516 18676
rect 32050 18620 32060 18676
rect 32116 18620 33180 18676
rect 33236 18620 33246 18676
rect 42578 18620 42588 18676
rect 42644 18620 43372 18676
rect 43428 18620 43438 18676
rect 26460 18564 26516 18620
rect 44716 18564 44772 18732
rect 50372 18676 50428 18732
rect 48178 18620 48188 18676
rect 48244 18620 49756 18676
rect 49812 18620 49822 18676
rect 50372 18620 58380 18676
rect 58436 18620 58446 18676
rect 63410 18620 63420 18676
rect 63476 18620 64764 18676
rect 64820 18620 65100 18676
rect 65156 18620 65166 18676
rect 73892 18564 73948 18956
rect 88060 18900 88116 18956
rect 88060 18844 91532 18900
rect 91588 18844 91598 18900
rect 92530 18844 92540 18900
rect 92596 18844 97244 18900
rect 97300 18844 97804 18900
rect 97860 18844 97870 18900
rect 81266 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81550 18844
rect 111986 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112270 18844
rect 88274 18732 88284 18788
rect 88340 18732 88732 18788
rect 88788 18732 88798 18788
rect 96002 18732 96012 18788
rect 96068 18732 99708 18788
rect 99764 18732 99774 18788
rect 83682 18620 83692 18676
rect 83748 18620 85820 18676
rect 85876 18620 85886 18676
rect 19170 18508 19180 18564
rect 19236 18508 21532 18564
rect 21588 18508 22428 18564
rect 22484 18508 25340 18564
rect 25396 18508 25406 18564
rect 26450 18508 26460 18564
rect 26516 18508 26526 18564
rect 31378 18508 31388 18564
rect 31444 18508 35532 18564
rect 35588 18508 35598 18564
rect 38612 18508 44772 18564
rect 58594 18508 58604 18564
rect 58660 18508 59724 18564
rect 59780 18508 59790 18564
rect 61170 18508 61180 18564
rect 61236 18508 64204 18564
rect 64260 18508 66444 18564
rect 66500 18508 66510 18564
rect 67330 18508 67340 18564
rect 67396 18508 71932 18564
rect 71988 18508 71998 18564
rect 73892 18508 84812 18564
rect 84868 18508 84878 18564
rect 93538 18508 93548 18564
rect 93604 18508 94668 18564
rect 94724 18508 94734 18564
rect 26460 18452 26516 18508
rect 26460 18396 26908 18452
rect 28690 18396 28700 18452
rect 28756 18396 29596 18452
rect 29652 18396 30268 18452
rect 30324 18396 30334 18452
rect 30482 18396 30492 18452
rect 30548 18396 34748 18452
rect 34804 18396 34814 18452
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 26852 17892 26908 18396
rect 38612 18340 38668 18508
rect 41010 18396 41020 18452
rect 41076 18396 41804 18452
rect 41860 18396 44268 18452
rect 44324 18396 44334 18452
rect 46498 18396 46508 18452
rect 46564 18396 47740 18452
rect 47796 18396 47806 18452
rect 48066 18396 48076 18452
rect 48132 18396 48860 18452
rect 48916 18396 50092 18452
rect 50148 18396 50158 18452
rect 50978 18396 50988 18452
rect 51044 18396 52668 18452
rect 52724 18396 52734 18452
rect 55906 18396 55916 18452
rect 55972 18396 59500 18452
rect 59556 18396 61068 18452
rect 61124 18396 61134 18452
rect 66546 18396 66556 18452
rect 66612 18396 66622 18452
rect 69458 18396 69468 18452
rect 69524 18396 70700 18452
rect 70756 18396 73724 18452
rect 73780 18396 73790 18452
rect 75730 18396 75740 18452
rect 75796 18396 78988 18452
rect 79044 18396 79054 18452
rect 82338 18396 82348 18452
rect 82404 18396 83468 18452
rect 83524 18396 83534 18452
rect 83906 18396 83916 18452
rect 83972 18396 85820 18452
rect 85876 18396 86380 18452
rect 86436 18396 86446 18452
rect 88162 18396 88172 18452
rect 88228 18396 90300 18452
rect 90356 18396 90366 18452
rect 90962 18396 90972 18452
rect 91028 18396 95340 18452
rect 95396 18396 96124 18452
rect 96180 18396 96190 18452
rect 96898 18396 96908 18452
rect 96964 18396 97244 18452
rect 97300 18396 97310 18452
rect 98914 18396 98924 18452
rect 98980 18396 99820 18452
rect 99876 18396 99886 18452
rect 100370 18396 100380 18452
rect 100436 18396 101948 18452
rect 102004 18396 102014 18452
rect 102498 18396 102508 18452
rect 102564 18396 104636 18452
rect 104692 18396 104702 18452
rect 106194 18396 106204 18452
rect 106260 18396 106988 18452
rect 107044 18396 107054 18452
rect 111010 18396 111020 18452
rect 111076 18396 111692 18452
rect 111748 18396 111758 18452
rect 112130 18396 112140 18452
rect 112196 18396 113260 18452
rect 113316 18396 113326 18452
rect 31826 18284 31836 18340
rect 31892 18284 33740 18340
rect 33796 18284 38668 18340
rect 41906 18284 41916 18340
rect 41972 18284 43148 18340
rect 43204 18284 43214 18340
rect 47506 18284 47516 18340
rect 47572 18284 49420 18340
rect 49476 18284 49486 18340
rect 51762 18284 51772 18340
rect 51828 18284 53004 18340
rect 53060 18284 53070 18340
rect 56802 18284 56812 18340
rect 56868 18284 57820 18340
rect 57876 18284 57886 18340
rect 58482 18284 58492 18340
rect 58548 18284 60732 18340
rect 60788 18284 60798 18340
rect 61954 18284 61964 18340
rect 62020 18284 63084 18340
rect 63140 18284 63150 18340
rect 49420 18228 49476 18284
rect 66556 18228 66612 18396
rect 102508 18340 102564 18396
rect 115948 18340 116004 18956
rect 142706 18788 142716 18844
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142980 18788 142990 18844
rect 69794 18284 69804 18340
rect 69860 18284 72268 18340
rect 72324 18284 72334 18340
rect 73892 18284 76860 18340
rect 76916 18284 76926 18340
rect 84466 18284 84476 18340
rect 84532 18284 85372 18340
rect 85428 18284 89628 18340
rect 89684 18284 89694 18340
rect 92194 18284 92204 18340
rect 92260 18284 92540 18340
rect 92596 18284 92606 18340
rect 94406 18284 94444 18340
rect 94500 18284 94510 18340
rect 94882 18284 94892 18340
rect 94948 18284 95900 18340
rect 95956 18284 95966 18340
rect 96684 18284 99484 18340
rect 99540 18284 99550 18340
rect 99698 18284 99708 18340
rect 99764 18284 100044 18340
rect 100100 18284 100110 18340
rect 101714 18284 101724 18340
rect 101780 18284 102564 18340
rect 109106 18284 109116 18340
rect 109172 18284 109788 18340
rect 109844 18284 109854 18340
rect 111906 18284 111916 18340
rect 111972 18284 112812 18340
rect 112868 18284 112878 18340
rect 115948 18284 117964 18340
rect 118020 18284 118030 18340
rect 73892 18228 73948 18284
rect 96684 18228 96740 18284
rect 101724 18228 101780 18284
rect 33506 18172 33516 18228
rect 33572 18172 36204 18228
rect 36260 18172 36270 18228
rect 49420 18172 51660 18228
rect 51716 18172 51726 18228
rect 51884 18172 52892 18228
rect 52948 18172 52958 18228
rect 56578 18172 56588 18228
rect 56644 18172 57372 18228
rect 57428 18172 57438 18228
rect 59714 18172 59724 18228
rect 59780 18172 60620 18228
rect 60676 18172 66612 18228
rect 73266 18172 73276 18228
rect 73332 18172 73948 18228
rect 74946 18172 74956 18228
rect 75012 18172 75180 18228
rect 75236 18172 75246 18228
rect 76626 18172 76636 18228
rect 76692 18172 79548 18228
rect 79604 18172 82012 18228
rect 82068 18172 94780 18228
rect 94836 18172 96684 18228
rect 96740 18172 96750 18228
rect 97020 18172 101780 18228
rect 109330 18172 109340 18228
rect 109396 18172 112140 18228
rect 112196 18172 112206 18228
rect 115042 18172 115052 18228
rect 115108 18172 120092 18228
rect 120148 18172 120158 18228
rect 51884 18116 51940 18172
rect 48290 18060 48300 18116
rect 48356 18060 49308 18116
rect 49364 18060 50428 18116
rect 51538 18060 51548 18116
rect 51604 18060 51940 18116
rect 52770 18060 52780 18116
rect 52836 18060 53340 18116
rect 53396 18060 57260 18116
rect 57316 18060 57326 18116
rect 61058 18060 61068 18116
rect 61124 18060 65548 18116
rect 65604 18060 65614 18116
rect 72930 18060 72940 18116
rect 72996 18060 77196 18116
rect 77252 18060 77262 18116
rect 77410 18060 77420 18116
rect 77476 18060 89068 18116
rect 89124 18060 89134 18116
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 50372 18004 50428 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 96626 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96910 18060
rect 32610 17948 32620 18004
rect 32676 17948 33628 18004
rect 33684 17948 33694 18004
rect 36194 17948 36204 18004
rect 36260 17948 48412 18004
rect 48468 17948 48478 18004
rect 50372 17948 51212 18004
rect 51268 17948 56252 18004
rect 56308 17948 56318 18004
rect 64306 17948 64316 18004
rect 64372 17948 65772 18004
rect 65828 17948 65838 18004
rect 72258 17948 72268 18004
rect 72324 17948 79212 18004
rect 79268 17948 79278 18004
rect 85652 17948 87724 18004
rect 87780 17948 87948 18004
rect 88004 17948 88508 18004
rect 88564 17948 88574 18004
rect 85652 17892 85708 17948
rect 97020 17892 97076 18172
rect 127346 18004 127356 18060
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127620 18004 127630 18060
rect 158066 18004 158076 18060
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158340 18004 158350 18060
rect 23314 17836 23324 17892
rect 23380 17836 23772 17892
rect 23828 17836 23838 17892
rect 26852 17836 27356 17892
rect 27412 17836 45724 17892
rect 45780 17836 54684 17892
rect 54740 17836 54750 17892
rect 54908 17836 85708 17892
rect 88284 17836 90636 17892
rect 90692 17836 90702 17892
rect 91970 17836 91980 17892
rect 92036 17836 97076 17892
rect 97412 17836 111020 17892
rect 111076 17836 111086 17892
rect 54908 17780 54964 17836
rect 88284 17780 88340 17836
rect 97412 17780 97468 17836
rect 23538 17724 23548 17780
rect 23604 17724 24556 17780
rect 24612 17724 24622 17780
rect 35634 17724 35644 17780
rect 35700 17724 42364 17780
rect 42420 17724 42430 17780
rect 50372 17724 51548 17780
rect 51604 17724 51614 17780
rect 54002 17724 54012 17780
rect 54068 17724 54964 17780
rect 55234 17724 55244 17780
rect 55300 17724 56140 17780
rect 56196 17724 56206 17780
rect 62850 17724 62860 17780
rect 62916 17724 69692 17780
rect 69748 17724 69758 17780
rect 77186 17724 77196 17780
rect 77252 17724 77262 17780
rect 83458 17724 83468 17780
rect 83524 17724 84252 17780
rect 84308 17724 84318 17780
rect 86034 17724 86044 17780
rect 86100 17724 88284 17780
rect 88340 17724 88350 17780
rect 89618 17724 89628 17780
rect 89684 17724 90748 17780
rect 90804 17724 90814 17780
rect 96114 17724 96124 17780
rect 96180 17724 97468 17780
rect 106754 17724 106764 17780
rect 106820 17724 107548 17780
rect 107604 17724 107614 17780
rect 22754 17612 22764 17668
rect 22820 17612 24108 17668
rect 24164 17612 28700 17668
rect 28756 17612 28766 17668
rect 33170 17612 33180 17668
rect 33236 17612 34524 17668
rect 34580 17612 34590 17668
rect 39442 17612 39452 17668
rect 39508 17612 41580 17668
rect 41636 17612 41646 17668
rect 45826 17612 45836 17668
rect 45892 17612 46284 17668
rect 46340 17612 47292 17668
rect 47348 17612 48860 17668
rect 48916 17612 49532 17668
rect 49588 17612 49598 17668
rect 50372 17556 50428 17724
rect 52882 17612 52892 17668
rect 52948 17612 55580 17668
rect 55636 17612 56700 17668
rect 56756 17612 56766 17668
rect 63858 17612 63868 17668
rect 63924 17612 65100 17668
rect 65156 17612 65660 17668
rect 65716 17612 65726 17668
rect 68898 17612 68908 17668
rect 68964 17612 69356 17668
rect 69412 17612 70476 17668
rect 70532 17612 70924 17668
rect 70980 17612 71820 17668
rect 71876 17612 71886 17668
rect 77196 17556 77252 17724
rect 79762 17612 79772 17668
rect 79828 17612 79996 17668
rect 80052 17612 80444 17668
rect 80500 17612 80510 17668
rect 80770 17612 80780 17668
rect 80836 17612 82124 17668
rect 82180 17612 82190 17668
rect 85362 17612 85372 17668
rect 85428 17612 86268 17668
rect 86324 17612 86334 17668
rect 87910 17612 87948 17668
rect 88004 17612 88620 17668
rect 88676 17612 88686 17668
rect 102498 17612 102508 17668
rect 102564 17612 106204 17668
rect 106260 17612 106270 17668
rect 106418 17612 106428 17668
rect 106484 17612 107996 17668
rect 108052 17612 109228 17668
rect 109284 17612 109294 17668
rect 38994 17500 39004 17556
rect 39060 17500 39564 17556
rect 39620 17500 40236 17556
rect 40292 17500 41020 17556
rect 41076 17500 41086 17556
rect 49858 17500 49868 17556
rect 49924 17500 50428 17556
rect 50978 17500 50988 17556
rect 51044 17500 51660 17556
rect 51716 17500 51726 17556
rect 52434 17500 52444 17556
rect 52500 17500 56812 17556
rect 56868 17500 58940 17556
rect 58996 17500 59500 17556
rect 59556 17500 62188 17556
rect 65762 17500 65772 17556
rect 65828 17500 68684 17556
rect 68740 17500 68750 17556
rect 77196 17500 87276 17556
rect 87332 17500 92204 17556
rect 92260 17500 92988 17556
rect 93044 17500 93772 17556
rect 93828 17500 93838 17556
rect 106754 17500 106764 17556
rect 106820 17500 107660 17556
rect 107716 17500 107726 17556
rect 62132 17444 62188 17500
rect 27794 17388 27804 17444
rect 27860 17388 30828 17444
rect 30884 17388 30894 17444
rect 34850 17388 34860 17444
rect 34916 17388 34926 17444
rect 38210 17388 38220 17444
rect 38276 17388 39228 17444
rect 39284 17388 39294 17444
rect 50082 17388 50092 17444
rect 50148 17388 57148 17444
rect 57204 17388 57214 17444
rect 62132 17388 62580 17444
rect 67778 17388 67788 17444
rect 67844 17388 69580 17444
rect 69636 17388 72492 17444
rect 72548 17388 72558 17444
rect 73714 17388 73724 17444
rect 73780 17388 74284 17444
rect 74340 17388 74350 17444
rect 84326 17388 84364 17444
rect 84420 17388 84430 17444
rect 85110 17388 85148 17444
rect 85204 17388 85214 17444
rect 87378 17388 87388 17444
rect 87444 17388 91196 17444
rect 91252 17388 94332 17444
rect 94388 17388 98700 17444
rect 98756 17388 101724 17444
rect 101780 17388 104860 17444
rect 104916 17388 104926 17444
rect 109554 17388 109564 17444
rect 109620 17388 112252 17444
rect 112308 17388 112318 17444
rect 34860 17332 34916 17388
rect 34860 17276 39004 17332
rect 39060 17276 39070 17332
rect 51090 17276 51100 17332
rect 51156 17276 52332 17332
rect 52388 17276 57596 17332
rect 57652 17276 59948 17332
rect 60004 17276 60396 17332
rect 60452 17276 62188 17332
rect 62244 17276 62254 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 22642 17164 22652 17220
rect 22708 17164 45724 17220
rect 45780 17164 45790 17220
rect 46162 17164 46172 17220
rect 46228 17164 46956 17220
rect 47012 17164 47404 17220
rect 47460 17164 50428 17220
rect 51314 17164 51324 17220
rect 51380 17164 51884 17220
rect 51940 17164 51950 17220
rect 57250 17164 57260 17220
rect 57316 17164 61964 17220
rect 62020 17164 62030 17220
rect 50372 17108 50428 17164
rect 62524 17108 62580 17388
rect 74162 17276 74172 17332
rect 74228 17276 77420 17332
rect 77476 17276 77486 17332
rect 89254 17276 89292 17332
rect 89348 17276 89358 17332
rect 90850 17276 90860 17332
rect 90916 17276 95340 17332
rect 95396 17276 95406 17332
rect 98242 17276 98252 17332
rect 98308 17276 106876 17332
rect 106932 17276 106942 17332
rect 81266 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81550 17276
rect 111986 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112270 17276
rect 142706 17220 142716 17276
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142980 17220 142990 17276
rect 62738 17164 62748 17220
rect 62804 17164 81172 17220
rect 81890 17164 81900 17220
rect 81956 17164 83244 17220
rect 83300 17164 85932 17220
rect 85988 17164 91140 17220
rect 94434 17164 94444 17220
rect 94500 17164 97916 17220
rect 97972 17164 97982 17220
rect 101378 17164 101388 17220
rect 101444 17164 101948 17220
rect 102004 17164 102014 17220
rect 81116 17108 81172 17164
rect 91084 17108 91140 17164
rect 9202 17052 9212 17108
rect 9268 17052 19628 17108
rect 19684 17052 20188 17108
rect 20244 17052 20254 17108
rect 31154 17052 31164 17108
rect 31220 17052 37772 17108
rect 37828 17052 37838 17108
rect 48402 17052 48412 17108
rect 48468 17052 49868 17108
rect 49924 17052 50204 17108
rect 50260 17052 50270 17108
rect 50372 17052 52556 17108
rect 52612 17052 52622 17108
rect 56690 17052 56700 17108
rect 56756 17052 58716 17108
rect 58772 17052 58782 17108
rect 62524 17052 63756 17108
rect 63812 17052 64540 17108
rect 64596 17052 68460 17108
rect 68516 17052 68526 17108
rect 75506 17052 75516 17108
rect 75572 17052 75740 17108
rect 75796 17052 75806 17108
rect 79202 17052 79212 17108
rect 79268 17052 80108 17108
rect 80164 17052 80174 17108
rect 81116 17052 83916 17108
rect 83972 17052 83982 17108
rect 91084 17052 99652 17108
rect 99810 17052 99820 17108
rect 99876 17052 100044 17108
rect 100100 17052 100110 17108
rect 101714 17052 101724 17108
rect 101780 17052 102508 17108
rect 102564 17052 102574 17108
rect 105410 17052 105420 17108
rect 105476 17052 112588 17108
rect 112644 17052 112654 17108
rect 112914 17052 112924 17108
rect 112980 17052 115276 17108
rect 115332 17052 115342 17108
rect 75516 16996 75572 17052
rect 99596 16996 99652 17052
rect 101724 16996 101780 17052
rect 21634 16940 21644 16996
rect 21700 16940 45948 16996
rect 46004 16940 46508 16996
rect 46564 16940 46574 16996
rect 47618 16940 47628 16996
rect 47684 16940 48524 16996
rect 48580 16940 48590 16996
rect 50306 16940 50316 16996
rect 50372 16940 50876 16996
rect 50932 16940 50942 16996
rect 53890 16940 53900 16996
rect 53956 16940 55020 16996
rect 55076 16940 68908 16996
rect 68964 16940 68974 16996
rect 71586 16940 71596 16996
rect 71652 16940 72492 16996
rect 72548 16940 75572 16996
rect 79986 16940 79996 16996
rect 80052 16940 80892 16996
rect 80948 16940 80958 16996
rect 81106 16940 81116 16996
rect 81172 16940 82684 16996
rect 82740 16940 82750 16996
rect 89058 16940 89068 16996
rect 89124 16940 89292 16996
rect 89348 16940 89358 16996
rect 91970 16940 91980 16996
rect 92036 16940 92988 16996
rect 93044 16940 93054 16996
rect 97234 16940 97244 16996
rect 97300 16940 98252 16996
rect 98308 16940 98318 16996
rect 99596 16940 101780 16996
rect 103964 16940 105308 16996
rect 105364 16940 105374 16996
rect 68908 16884 68964 16940
rect 92988 16884 93044 16940
rect 103964 16884 104020 16940
rect 29922 16828 29932 16884
rect 29988 16828 30716 16884
rect 30772 16828 31500 16884
rect 31556 16828 31566 16884
rect 31826 16828 31836 16884
rect 31892 16828 32396 16884
rect 32452 16828 33740 16884
rect 33796 16828 33806 16884
rect 35970 16828 35980 16884
rect 36036 16828 36876 16884
rect 36932 16828 36942 16884
rect 37202 16828 37212 16884
rect 37268 16828 38668 16884
rect 38724 16828 38734 16884
rect 46050 16828 46060 16884
rect 46116 16828 47852 16884
rect 47908 16828 47918 16884
rect 48066 16828 48076 16884
rect 48132 16828 49532 16884
rect 49588 16828 49598 16884
rect 50194 16828 50204 16884
rect 50260 16828 51100 16884
rect 51156 16828 51166 16884
rect 55682 16828 55692 16884
rect 55748 16828 56588 16884
rect 56644 16828 57036 16884
rect 57092 16828 58828 16884
rect 58884 16828 58894 16884
rect 59154 16828 59164 16884
rect 59220 16828 60732 16884
rect 60788 16828 60798 16884
rect 60946 16828 60956 16884
rect 61012 16828 61404 16884
rect 61460 16828 62076 16884
rect 62132 16828 62142 16884
rect 62402 16828 62412 16884
rect 62468 16828 63420 16884
rect 63476 16828 63486 16884
rect 64530 16828 64540 16884
rect 64596 16828 65548 16884
rect 65604 16828 65614 16884
rect 68908 16828 76636 16884
rect 76692 16828 76702 16884
rect 76850 16828 76860 16884
rect 76916 16828 77644 16884
rect 77700 16828 77710 16884
rect 82786 16828 82796 16884
rect 82852 16828 83580 16884
rect 83636 16828 84028 16884
rect 84084 16828 84094 16884
rect 85446 16828 85484 16884
rect 85540 16828 85550 16884
rect 89730 16828 89740 16884
rect 89796 16828 91084 16884
rect 91140 16828 91150 16884
rect 92418 16828 92428 16884
rect 92484 16828 92764 16884
rect 92820 16828 92830 16884
rect 92988 16828 100380 16884
rect 100436 16828 100446 16884
rect 100818 16828 100828 16884
rect 100884 16828 103964 16884
rect 104020 16828 104030 16884
rect 104850 16828 104860 16884
rect 104916 16828 105644 16884
rect 105700 16828 108892 16884
rect 108948 16828 111916 16884
rect 111972 16828 111982 16884
rect 19282 16716 19292 16772
rect 19348 16716 20300 16772
rect 20356 16716 20366 16772
rect 22754 16716 22764 16772
rect 22820 16716 24892 16772
rect 24948 16716 24958 16772
rect 30370 16716 30380 16772
rect 30436 16716 31052 16772
rect 31108 16716 31118 16772
rect 32162 16716 32172 16772
rect 32228 16716 34636 16772
rect 34692 16716 34702 16772
rect 47282 16716 47292 16772
rect 47348 16716 48860 16772
rect 48916 16716 48926 16772
rect 62850 16716 62860 16772
rect 62916 16716 67340 16772
rect 67396 16716 67406 16772
rect 73602 16716 73612 16772
rect 73668 16716 76300 16772
rect 76356 16716 76366 16772
rect 83458 16716 83468 16772
rect 83524 16716 87388 16772
rect 87444 16716 87454 16772
rect 94966 16716 95004 16772
rect 95060 16716 95070 16772
rect 97010 16716 97020 16772
rect 97076 16716 97468 16772
rect 97524 16716 97534 16772
rect 100034 16716 100044 16772
rect 100100 16716 100492 16772
rect 100548 16716 101052 16772
rect 101108 16716 101118 16772
rect 107762 16716 107772 16772
rect 107828 16716 108780 16772
rect 108836 16716 110236 16772
rect 110292 16716 110302 16772
rect 32172 16660 32228 16716
rect 27122 16604 27132 16660
rect 27188 16604 27916 16660
rect 27972 16604 32228 16660
rect 38210 16604 38220 16660
rect 38276 16604 72044 16660
rect 72100 16604 73276 16660
rect 73332 16604 73342 16660
rect 77186 16604 77196 16660
rect 77252 16604 105756 16660
rect 105812 16604 105822 16660
rect 48290 16492 48300 16548
rect 48356 16492 49868 16548
rect 49924 16492 49934 16548
rect 52882 16492 52892 16548
rect 52948 16492 53676 16548
rect 53732 16492 53742 16548
rect 76178 16492 76188 16548
rect 76244 16492 77420 16548
rect 77476 16492 77486 16548
rect 97234 16492 97244 16548
rect 97300 16492 98588 16548
rect 98644 16492 98654 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 96626 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96910 16492
rect 127346 16436 127356 16492
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127620 16436 127630 16492
rect 158066 16436 158076 16492
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158340 16436 158350 16492
rect 43250 16380 43260 16436
rect 43316 16380 55916 16436
rect 55972 16380 56588 16436
rect 56644 16380 56654 16436
rect 73892 16380 81340 16436
rect 81396 16380 82124 16436
rect 82180 16380 82190 16436
rect 85652 16380 91084 16436
rect 91140 16380 91980 16436
rect 92036 16380 92046 16436
rect 73892 16324 73948 16380
rect 85652 16324 85708 16380
rect 33394 16268 33404 16324
rect 33460 16268 34972 16324
rect 35028 16268 35038 16324
rect 38322 16268 38332 16324
rect 38388 16268 41356 16324
rect 41412 16268 42140 16324
rect 42196 16268 42812 16324
rect 42868 16268 42878 16324
rect 49634 16268 49644 16324
rect 49700 16268 56028 16324
rect 56084 16268 56094 16324
rect 61058 16268 61068 16324
rect 61124 16268 62076 16324
rect 62132 16268 62142 16324
rect 63074 16268 63084 16324
rect 63140 16268 73948 16324
rect 75282 16268 75292 16324
rect 75348 16268 76412 16324
rect 76468 16268 77308 16324
rect 77364 16268 77374 16324
rect 77634 16268 77644 16324
rect 77700 16268 78428 16324
rect 78484 16268 85708 16324
rect 88722 16268 88732 16324
rect 88788 16268 100212 16324
rect 101490 16268 101500 16324
rect 101556 16268 104188 16324
rect 104244 16268 104254 16324
rect 100156 16212 100212 16268
rect 20738 16156 20748 16212
rect 20804 16156 22876 16212
rect 22932 16156 22942 16212
rect 28802 16156 28812 16212
rect 28868 16156 36428 16212
rect 36484 16156 36988 16212
rect 37044 16156 37054 16212
rect 40898 16156 40908 16212
rect 40964 16156 41692 16212
rect 41748 16156 41758 16212
rect 46498 16156 46508 16212
rect 46564 16156 60620 16212
rect 60676 16156 60686 16212
rect 62132 16156 76804 16212
rect 77970 16156 77980 16212
rect 78036 16156 85708 16212
rect 89954 16156 89964 16212
rect 90020 16156 90748 16212
rect 90804 16156 90814 16212
rect 92082 16156 92092 16212
rect 92148 16156 93996 16212
rect 94052 16156 94332 16212
rect 94388 16156 94398 16212
rect 97570 16156 97580 16212
rect 97636 16156 98812 16212
rect 98868 16156 98878 16212
rect 100156 16156 102956 16212
rect 103012 16156 103022 16212
rect 105634 16156 105644 16212
rect 105700 16156 142604 16212
rect 142660 16156 142670 16212
rect 62132 16100 62188 16156
rect 17938 16044 17948 16100
rect 18004 16044 20412 16100
rect 20468 16044 21644 16100
rect 21700 16044 21710 16100
rect 24882 16044 24892 16100
rect 24948 16044 29820 16100
rect 29876 16044 30492 16100
rect 30548 16044 30558 16100
rect 31042 16044 31052 16100
rect 31108 16044 31836 16100
rect 31892 16044 32508 16100
rect 32564 16044 32574 16100
rect 40562 16044 40572 16100
rect 40628 16044 41804 16100
rect 41860 16044 41870 16100
rect 48626 16044 48636 16100
rect 48692 16044 49756 16100
rect 49812 16044 49822 16100
rect 52770 16044 52780 16100
rect 52836 16044 57484 16100
rect 57540 16044 59276 16100
rect 59332 16044 62188 16100
rect 9202 15932 9212 15988
rect 9268 15932 66444 15988
rect 66500 15932 66510 15988
rect 68338 15932 68348 15988
rect 68404 15932 69132 15988
rect 69188 15932 69198 15988
rect 73042 15932 73052 15988
rect 73108 15932 74172 15988
rect 74228 15932 74956 15988
rect 75012 15932 75022 15988
rect 75618 15932 75628 15988
rect 75684 15932 76412 15988
rect 76468 15932 76478 15988
rect 76748 15876 76804 16156
rect 85652 16100 85708 16156
rect 79538 16044 79548 16100
rect 79604 16044 79884 16100
rect 79940 16044 80780 16100
rect 80836 16044 80846 16100
rect 85652 16044 87948 16100
rect 88004 16044 90636 16100
rect 90692 16044 90702 16100
rect 92866 16044 92876 16100
rect 92932 16044 93324 16100
rect 93380 16044 93548 16100
rect 93604 16044 93614 16100
rect 103954 16044 103964 16100
rect 104020 16044 154028 16100
rect 154084 16044 154094 16100
rect 80098 15932 80108 15988
rect 80164 15932 85708 15988
rect 97906 15932 97916 15988
rect 97972 15932 101052 15988
rect 101108 15932 102508 15988
rect 102564 15932 102574 15988
rect 85652 15876 85708 15932
rect 29586 15820 29596 15876
rect 29652 15820 31052 15876
rect 31108 15820 31118 15876
rect 34402 15820 34412 15876
rect 34468 15820 35644 15876
rect 35700 15820 35710 15876
rect 36082 15820 36092 15876
rect 36148 15820 36988 15876
rect 37044 15820 37054 15876
rect 40338 15820 40348 15876
rect 40404 15820 43820 15876
rect 43876 15820 47180 15876
rect 47236 15820 47246 15876
rect 47394 15820 47404 15876
rect 47460 15820 48188 15876
rect 48244 15820 48254 15876
rect 49186 15820 49196 15876
rect 49252 15820 52500 15876
rect 52658 15820 52668 15876
rect 52724 15820 54124 15876
rect 54180 15820 54190 15876
rect 75170 15820 75180 15876
rect 75236 15820 75852 15876
rect 75908 15820 75918 15876
rect 76290 15820 76300 15876
rect 76356 15820 76366 15876
rect 76738 15820 76748 15876
rect 76804 15820 76814 15876
rect 76962 15820 76972 15876
rect 77028 15820 77420 15876
rect 77476 15820 77980 15876
rect 78036 15820 78046 15876
rect 83094 15820 83132 15876
rect 83188 15820 83198 15876
rect 83542 15820 83580 15876
rect 83636 15820 83646 15876
rect 84466 15820 84476 15876
rect 84532 15820 85148 15876
rect 85204 15820 85214 15876
rect 85652 15820 85932 15876
rect 85988 15820 85998 15876
rect 94854 15820 94892 15876
rect 94948 15820 94958 15876
rect 105718 15820 105756 15876
rect 105812 15820 105822 15876
rect 106306 15820 106316 15876
rect 106372 15820 106988 15876
rect 107044 15820 107054 15876
rect 112466 15820 112476 15876
rect 112532 15820 114940 15876
rect 114996 15820 115006 15876
rect 52444 15764 52500 15820
rect 76300 15764 76356 15820
rect 30370 15708 30380 15764
rect 30436 15708 30446 15764
rect 37650 15708 37660 15764
rect 37716 15708 38332 15764
rect 38388 15708 38398 15764
rect 38612 15708 40796 15764
rect 40852 15708 40862 15764
rect 41682 15708 41692 15764
rect 41748 15708 41758 15764
rect 48066 15708 48076 15764
rect 48132 15708 48972 15764
rect 49028 15708 49038 15764
rect 52444 15708 56252 15764
rect 56308 15708 60508 15764
rect 60564 15708 61404 15764
rect 61460 15708 61470 15764
rect 70578 15708 70588 15764
rect 70644 15708 72940 15764
rect 72996 15708 73836 15764
rect 73892 15708 76356 15764
rect 76626 15708 76636 15764
rect 76692 15708 79772 15764
rect 79828 15708 79838 15764
rect 86258 15708 86268 15764
rect 86324 15708 97468 15764
rect 106530 15708 106540 15764
rect 106596 15708 107772 15764
rect 107828 15708 107838 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 30380 15652 30436 15708
rect 38612 15652 38668 15708
rect 30380 15596 38668 15652
rect 41692 15540 41748 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 81266 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81550 15708
rect 97412 15652 97468 15708
rect 111986 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112270 15708
rect 142706 15652 142716 15708
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142980 15652 142990 15708
rect 70130 15596 70140 15652
rect 70196 15596 70812 15652
rect 70868 15596 70878 15652
rect 81666 15596 81676 15652
rect 81732 15596 82572 15652
rect 82628 15596 82638 15652
rect 85138 15596 85148 15652
rect 85204 15596 96012 15652
rect 96068 15596 96078 15652
rect 97412 15596 100380 15652
rect 100436 15596 100828 15652
rect 100884 15596 106484 15652
rect 106428 15540 106484 15596
rect 18610 15484 18620 15540
rect 18676 15484 20748 15540
rect 20804 15484 20814 15540
rect 20962 15484 20972 15540
rect 21028 15484 22764 15540
rect 22820 15484 22830 15540
rect 23314 15484 23324 15540
rect 23380 15484 25788 15540
rect 25844 15484 25854 15540
rect 26114 15484 26124 15540
rect 26180 15484 31836 15540
rect 31892 15484 34860 15540
rect 34916 15484 35532 15540
rect 35588 15484 35868 15540
rect 35924 15484 35934 15540
rect 38322 15484 38332 15540
rect 38388 15484 41748 15540
rect 44258 15484 44268 15540
rect 44324 15484 45276 15540
rect 45332 15484 48300 15540
rect 48356 15484 48366 15540
rect 48850 15484 48860 15540
rect 48916 15484 49420 15540
rect 49476 15484 49486 15540
rect 49970 15484 49980 15540
rect 50036 15484 50764 15540
rect 50820 15484 50830 15540
rect 54114 15484 54124 15540
rect 54180 15484 55132 15540
rect 55188 15484 59388 15540
rect 59444 15484 59454 15540
rect 69682 15484 69692 15540
rect 69748 15484 71260 15540
rect 71316 15484 71326 15540
rect 71474 15484 71484 15540
rect 71540 15484 72380 15540
rect 72436 15484 72446 15540
rect 78530 15484 78540 15540
rect 78596 15484 79548 15540
rect 79604 15484 80108 15540
rect 80164 15484 80174 15540
rect 88834 15484 88844 15540
rect 88900 15484 90804 15540
rect 100482 15484 100492 15540
rect 100548 15484 101724 15540
rect 101780 15484 101790 15540
rect 106418 15484 106428 15540
rect 106484 15484 107436 15540
rect 107492 15484 107502 15540
rect 107874 15484 107884 15540
rect 107940 15484 108780 15540
rect 108836 15484 108846 15540
rect 90748 15428 90804 15484
rect 22194 15372 22204 15428
rect 22260 15372 25228 15428
rect 25284 15372 25294 15428
rect 33954 15372 33964 15428
rect 34020 15372 36316 15428
rect 36372 15372 36382 15428
rect 41346 15372 41356 15428
rect 41412 15372 50876 15428
rect 50932 15372 51772 15428
rect 51828 15372 52668 15428
rect 52724 15372 52734 15428
rect 57138 15372 57148 15428
rect 57204 15372 62188 15428
rect 62244 15372 63644 15428
rect 63700 15372 63710 15428
rect 68236 15372 72492 15428
rect 72548 15372 73052 15428
rect 73108 15372 73118 15428
rect 74274 15372 74284 15428
rect 74340 15372 78932 15428
rect 79090 15372 79100 15428
rect 79156 15372 83468 15428
rect 83524 15372 83534 15428
rect 85820 15372 89292 15428
rect 89348 15372 89358 15428
rect 90738 15372 90748 15428
rect 90804 15372 93996 15428
rect 94052 15372 94062 15428
rect 101602 15372 101612 15428
rect 101668 15372 104300 15428
rect 104356 15372 104366 15428
rect 106978 15372 106988 15428
rect 107044 15372 108892 15428
rect 108948 15372 108958 15428
rect 68236 15316 68292 15372
rect 78876 15316 78932 15372
rect 19618 15260 19628 15316
rect 19684 15260 20636 15316
rect 20692 15260 22428 15316
rect 22484 15260 22494 15316
rect 24546 15260 24556 15316
rect 24612 15260 25340 15316
rect 25396 15260 26684 15316
rect 26740 15260 29036 15316
rect 29092 15260 29102 15316
rect 35634 15260 35644 15316
rect 35700 15260 36204 15316
rect 36260 15260 37996 15316
rect 38052 15260 38062 15316
rect 61618 15260 61628 15316
rect 61684 15260 63196 15316
rect 63252 15260 63262 15316
rect 63746 15260 63756 15316
rect 63812 15260 68292 15316
rect 68450 15260 68460 15316
rect 68516 15260 70700 15316
rect 70756 15260 70766 15316
rect 70914 15260 70924 15316
rect 70980 15260 74956 15316
rect 75012 15260 75022 15316
rect 78876 15260 85316 15316
rect 85260 15204 85316 15260
rect 85820 15204 85876 15372
rect 86258 15260 86268 15316
rect 86324 15260 87276 15316
rect 87332 15260 87342 15316
rect 102274 15260 102284 15316
rect 102340 15260 104748 15316
rect 104804 15260 106652 15316
rect 106708 15260 106718 15316
rect 38994 15148 39004 15204
rect 39060 15148 39340 15204
rect 39396 15148 39406 15204
rect 52882 15148 52892 15204
rect 52948 15148 54236 15204
rect 54292 15148 54302 15204
rect 63074 15148 63084 15204
rect 63140 15148 68012 15204
rect 68068 15148 68078 15204
rect 69122 15148 69132 15204
rect 69188 15148 74620 15204
rect 74676 15148 74686 15204
rect 77186 15148 77196 15204
rect 77252 15148 77980 15204
rect 78036 15148 78046 15204
rect 85250 15148 85260 15204
rect 85316 15148 85876 15204
rect 89068 15148 89292 15204
rect 89348 15148 89358 15204
rect 90178 15148 90188 15204
rect 90244 15148 90860 15204
rect 90916 15148 91532 15204
rect 91588 15148 91598 15204
rect 93986 15148 93996 15204
rect 94052 15148 94892 15204
rect 94948 15148 94958 15204
rect 95106 15148 95116 15204
rect 95172 15148 95900 15204
rect 95956 15148 95966 15204
rect 103292 15148 105644 15204
rect 105700 15148 105710 15204
rect 105868 15148 107100 15204
rect 107156 15148 107660 15204
rect 107716 15148 109788 15204
rect 109844 15148 109854 15204
rect 89068 15092 89124 15148
rect 103292 15092 103348 15148
rect 105868 15092 105924 15148
rect 28466 15036 28476 15092
rect 28532 15036 31948 15092
rect 32004 15036 32014 15092
rect 34290 15036 34300 15092
rect 34356 15036 51660 15092
rect 51716 15036 51726 15092
rect 52210 15036 52220 15092
rect 52276 15036 53116 15092
rect 53172 15036 53182 15092
rect 54124 15036 58436 15092
rect 58706 15036 58716 15092
rect 58772 15036 63308 15092
rect 63364 15036 63374 15092
rect 66658 15036 66668 15092
rect 66724 15036 67340 15092
rect 67396 15036 74564 15092
rect 74722 15036 74732 15092
rect 74788 15036 82796 15092
rect 82852 15036 82862 15092
rect 83010 15036 83020 15092
rect 83076 15036 86380 15092
rect 86436 15036 86446 15092
rect 89068 15036 92988 15092
rect 93044 15036 93054 15092
rect 94098 15036 94108 15092
rect 94164 15036 94444 15092
rect 94500 15036 94510 15092
rect 98802 15036 98812 15092
rect 98868 15036 103348 15092
rect 103506 15036 103516 15092
rect 103572 15036 105924 15092
rect 54124 14980 54180 15036
rect 58380 14980 58436 15036
rect 46386 14924 46396 14980
rect 46452 14924 54180 14980
rect 54236 14924 58156 14980
rect 58212 14924 58222 14980
rect 58380 14924 62076 14980
rect 62132 14924 62860 14980
rect 62916 14924 62926 14980
rect 66322 14924 66332 14980
rect 66388 14924 74284 14980
rect 74340 14924 74350 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 47170 14812 47180 14868
rect 47236 14812 54012 14868
rect 54068 14812 54078 14868
rect 54236 14756 54292 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 74508 14868 74564 15036
rect 78642 14924 78652 14980
rect 78708 14924 85708 14980
rect 112578 14924 112588 14980
rect 112644 14924 118412 14980
rect 118468 14924 118478 14980
rect 85652 14868 85708 14924
rect 96626 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96910 14924
rect 127346 14868 127356 14924
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127620 14868 127630 14924
rect 158066 14868 158076 14924
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158340 14868 158350 14924
rect 42130 14700 42140 14756
rect 42196 14700 45388 14756
rect 45444 14700 45454 14756
rect 49186 14700 49196 14756
rect 49252 14700 54292 14756
rect 58772 14812 62748 14868
rect 62804 14812 62814 14868
rect 64530 14812 64540 14868
rect 64596 14812 65324 14868
rect 65380 14812 65390 14868
rect 74508 14812 80556 14868
rect 80612 14812 80622 14868
rect 85652 14812 86828 14868
rect 86884 14812 86894 14868
rect 102946 14812 102956 14868
rect 103012 14812 103964 14868
rect 104020 14812 104030 14868
rect 42354 14588 42364 14644
rect 42420 14588 52780 14644
rect 52836 14588 52846 14644
rect 58772 14532 58828 14812
rect 60610 14700 60620 14756
rect 60676 14700 67788 14756
rect 67844 14700 67854 14756
rect 68012 14700 70028 14756
rect 70084 14700 74116 14756
rect 80434 14700 80444 14756
rect 80500 14700 81452 14756
rect 81508 14700 81518 14756
rect 84802 14700 84812 14756
rect 84868 14700 85708 14756
rect 87378 14700 87388 14756
rect 87444 14700 92316 14756
rect 92372 14700 92382 14756
rect 97412 14700 98252 14756
rect 98308 14700 100156 14756
rect 100212 14700 100222 14756
rect 101490 14700 101500 14756
rect 101556 14700 105532 14756
rect 105588 14700 106092 14756
rect 106148 14700 106158 14756
rect 68012 14644 68068 14700
rect 63746 14588 63756 14644
rect 63812 14588 68068 14644
rect 69010 14588 69020 14644
rect 69076 14588 72380 14644
rect 72436 14588 72446 14644
rect 37090 14476 37100 14532
rect 37156 14476 37324 14532
rect 37380 14476 44940 14532
rect 44996 14476 45006 14532
rect 49746 14476 49756 14532
rect 49812 14476 58828 14532
rect 60722 14476 60732 14532
rect 60788 14476 60798 14532
rect 61366 14476 61404 14532
rect 61460 14476 61470 14532
rect 61618 14476 61628 14532
rect 61684 14476 62188 14532
rect 62244 14476 62524 14532
rect 62580 14476 62590 14532
rect 63634 14476 63644 14532
rect 63700 14476 72492 14532
rect 72548 14476 72558 14532
rect 60732 14420 60788 14476
rect 74060 14420 74116 14700
rect 85652 14644 85708 14700
rect 97412 14644 97468 14700
rect 75282 14588 75292 14644
rect 75348 14588 80332 14644
rect 80388 14588 80398 14644
rect 81778 14588 81788 14644
rect 81844 14588 82572 14644
rect 82628 14588 83132 14644
rect 83188 14588 84700 14644
rect 84756 14588 85260 14644
rect 85316 14588 85326 14644
rect 85652 14588 86940 14644
rect 86996 14588 87006 14644
rect 91186 14588 91196 14644
rect 91252 14588 91532 14644
rect 91588 14588 91598 14644
rect 97122 14588 97132 14644
rect 97188 14588 97468 14644
rect 100034 14588 100044 14644
rect 100100 14588 101388 14644
rect 101444 14588 103628 14644
rect 103684 14588 103694 14644
rect 108994 14588 109004 14644
rect 109060 14588 110572 14644
rect 110628 14588 110638 14644
rect 74274 14476 74284 14532
rect 74340 14476 80388 14532
rect 81218 14476 81228 14532
rect 81284 14476 93100 14532
rect 93156 14476 93166 14532
rect 97794 14476 97804 14532
rect 97860 14476 98924 14532
rect 98980 14476 98990 14532
rect 99250 14476 99260 14532
rect 99316 14476 99932 14532
rect 99988 14476 99998 14532
rect 103282 14476 103292 14532
rect 103348 14476 119756 14532
rect 119812 14476 119822 14532
rect 80332 14420 80388 14476
rect 29138 14364 29148 14420
rect 29204 14364 30156 14420
rect 30212 14364 30222 14420
rect 35746 14364 35756 14420
rect 35812 14364 38444 14420
rect 38500 14364 38668 14420
rect 50306 14364 50316 14420
rect 50372 14364 60788 14420
rect 65314 14364 65324 14420
rect 65380 14364 66444 14420
rect 66500 14364 66510 14420
rect 74060 14364 74900 14420
rect 80322 14364 80332 14420
rect 80388 14364 80398 14420
rect 81554 14364 81564 14420
rect 81620 14364 82572 14420
rect 82628 14364 83020 14420
rect 83076 14364 83086 14420
rect 86940 14364 91196 14420
rect 91252 14364 97468 14420
rect 103954 14364 103964 14420
rect 104020 14364 107212 14420
rect 107268 14364 108444 14420
rect 108500 14364 108510 14420
rect 108892 14364 131180 14420
rect 131236 14364 131246 14420
rect 38612 14308 38668 14364
rect 74844 14308 74900 14364
rect 17154 14252 17164 14308
rect 17220 14252 20412 14308
rect 20468 14252 22652 14308
rect 22708 14252 25676 14308
rect 25732 14252 26684 14308
rect 26740 14252 29708 14308
rect 29764 14252 31052 14308
rect 31108 14252 32508 14308
rect 32564 14252 33516 14308
rect 33572 14252 34412 14308
rect 34468 14252 37100 14308
rect 37156 14252 37436 14308
rect 37492 14252 37502 14308
rect 38612 14252 39564 14308
rect 39620 14252 39630 14308
rect 54562 14252 54572 14308
rect 54628 14252 62188 14308
rect 62132 14196 62188 14252
rect 64540 14252 68908 14308
rect 68964 14252 68974 14308
rect 73266 14252 73276 14308
rect 73332 14252 74284 14308
rect 74340 14252 74350 14308
rect 74834 14252 74844 14308
rect 74900 14252 75628 14308
rect 75684 14252 75694 14308
rect 81106 14252 81116 14308
rect 81172 14252 81900 14308
rect 81956 14252 81966 14308
rect 85250 14252 85260 14308
rect 85316 14252 86156 14308
rect 86212 14252 86222 14308
rect 64540 14196 64596 14252
rect 86940 14196 86996 14364
rect 87154 14252 87164 14308
rect 87220 14252 88172 14308
rect 88228 14252 88844 14308
rect 88900 14252 92876 14308
rect 92932 14252 92942 14308
rect 94658 14252 94668 14308
rect 94724 14252 95452 14308
rect 95508 14252 95518 14308
rect 25218 14140 25228 14196
rect 25284 14140 25788 14196
rect 25844 14140 39676 14196
rect 39732 14140 39742 14196
rect 62132 14140 64596 14196
rect 64754 14140 64764 14196
rect 64820 14140 66668 14196
rect 66724 14140 79100 14196
rect 79156 14140 79166 14196
rect 83570 14140 83580 14196
rect 83636 14140 83692 14196
rect 83748 14140 83758 14196
rect 83906 14140 83916 14196
rect 83972 14140 86268 14196
rect 86324 14140 86996 14196
rect 90738 14140 90748 14196
rect 90804 14140 91756 14196
rect 91812 14140 91822 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 81266 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81550 14140
rect 24994 14028 25004 14084
rect 25060 14028 30492 14084
rect 30548 14028 30558 14084
rect 30940 14028 39452 14084
rect 39508 14028 39518 14084
rect 39890 14028 39900 14084
rect 39956 14028 40124 14084
rect 40180 14028 42588 14084
rect 42644 14028 44492 14084
rect 44548 14028 44558 14084
rect 61058 14028 61068 14084
rect 61124 14028 62076 14084
rect 62132 14028 62142 14084
rect 62850 14028 62860 14084
rect 62916 14028 65772 14084
rect 65828 14028 66780 14084
rect 66836 14028 66846 14084
rect 84242 14028 84252 14084
rect 84308 14028 85708 14084
rect 86594 14028 86604 14084
rect 86660 14028 92428 14084
rect 92484 14028 92494 14084
rect 20066 13916 20076 13972
rect 20132 13916 30492 13972
rect 30548 13916 30558 13972
rect 30940 13860 30996 14028
rect 35298 13916 35308 13972
rect 35364 13916 35868 13972
rect 35924 13916 38220 13972
rect 38276 13916 38286 13972
rect 39554 13916 39564 13972
rect 39620 13916 42140 13972
rect 42196 13916 42206 13972
rect 46386 13916 46396 13972
rect 46452 13916 49532 13972
rect 49588 13916 50204 13972
rect 50260 13916 50270 13972
rect 61954 13916 61964 13972
rect 62020 13916 63756 13972
rect 63812 13916 63822 13972
rect 65538 13916 65548 13972
rect 65604 13916 66220 13972
rect 66276 13916 68684 13972
rect 68740 13916 69804 13972
rect 69860 13916 69870 13972
rect 71250 13916 71260 13972
rect 71316 13916 71820 13972
rect 71876 13916 77868 13972
rect 77924 13916 77934 13972
rect 78418 13916 78428 13972
rect 78484 13916 83020 13972
rect 83076 13916 83086 13972
rect 83542 13916 83580 13972
rect 83636 13916 83646 13972
rect 84690 13916 84700 13972
rect 84756 13916 85260 13972
rect 85316 13916 85326 13972
rect 26852 13804 30996 13860
rect 31154 13804 31164 13860
rect 31220 13804 31500 13860
rect 31556 13804 52108 13860
rect 52164 13804 52174 13860
rect 52444 13804 53116 13860
rect 53172 13804 62524 13860
rect 62580 13804 62590 13860
rect 65650 13804 65660 13860
rect 65716 13804 66332 13860
rect 66388 13804 66398 13860
rect 72930 13804 72940 13860
rect 72996 13804 74732 13860
rect 74788 13804 74798 13860
rect 75506 13804 75516 13860
rect 75572 13804 84028 13860
rect 84084 13804 84980 13860
rect 26852 13524 26908 13804
rect 52444 13748 52500 13804
rect 30370 13692 30380 13748
rect 30436 13692 31388 13748
rect 31444 13692 34636 13748
rect 34692 13692 36652 13748
rect 36708 13692 36718 13748
rect 37090 13692 37100 13748
rect 37156 13692 38108 13748
rect 38164 13692 38174 13748
rect 41010 13692 41020 13748
rect 41076 13692 41692 13748
rect 41748 13692 41758 13748
rect 50306 13692 50316 13748
rect 50372 13692 52500 13748
rect 52658 13692 52668 13748
rect 52724 13692 55132 13748
rect 55188 13692 55198 13748
rect 56802 13692 56812 13748
rect 56868 13692 57596 13748
rect 57652 13692 57662 13748
rect 61628 13692 64428 13748
rect 64484 13692 64494 13748
rect 69570 13692 69580 13748
rect 69636 13692 71036 13748
rect 71092 13692 71102 13748
rect 75394 13692 75404 13748
rect 75460 13692 76412 13748
rect 76468 13692 76478 13748
rect 80322 13692 80332 13748
rect 80388 13692 84252 13748
rect 84308 13692 84318 13748
rect 27346 13580 27356 13636
rect 27412 13580 30268 13636
rect 30324 13580 30334 13636
rect 30482 13580 30492 13636
rect 30548 13580 33516 13636
rect 33572 13580 34300 13636
rect 34356 13580 34366 13636
rect 36754 13580 36764 13636
rect 36820 13580 37548 13636
rect 37604 13580 37614 13636
rect 40338 13580 40348 13636
rect 40404 13580 48188 13636
rect 48244 13580 48254 13636
rect 55234 13580 55244 13636
rect 55300 13580 56700 13636
rect 56756 13580 56766 13636
rect 57138 13580 57148 13636
rect 57204 13580 58044 13636
rect 58100 13580 58110 13636
rect 61628 13524 61684 13692
rect 84924 13636 84980 13804
rect 85652 13692 85708 14028
rect 97412 13972 97468 14364
rect 97524 14252 97544 14308
rect 106642 14252 106652 14308
rect 106708 14252 108108 14308
rect 108164 14252 108174 14308
rect 108892 14196 108948 14364
rect 100044 14140 108948 14196
rect 109172 14252 110460 14308
rect 110516 14252 111468 14308
rect 111524 14252 111534 14308
rect 100044 14084 100100 14140
rect 109172 14084 109228 14252
rect 111986 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112270 14140
rect 142706 14084 142716 14140
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142980 14084 142990 14140
rect 100034 14028 100044 14084
rect 100100 14028 100110 14084
rect 108322 14028 108332 14084
rect 108388 14028 109228 14084
rect 85922 13916 85932 13972
rect 85988 13916 96124 13972
rect 96180 13916 96190 13972
rect 97412 13916 119532 13972
rect 119588 13916 119598 13972
rect 89842 13804 89852 13860
rect 89908 13804 93548 13860
rect 93604 13804 93614 13860
rect 94966 13804 95004 13860
rect 95060 13804 95070 13860
rect 101378 13804 101388 13860
rect 101444 13804 104636 13860
rect 104692 13804 106652 13860
rect 106708 13804 106718 13860
rect 85764 13692 85774 13748
rect 87724 13692 96012 13748
rect 96068 13692 96078 13748
rect 97794 13692 97804 13748
rect 97860 13692 98252 13748
rect 98308 13692 98318 13748
rect 99362 13692 99372 13748
rect 99428 13692 100268 13748
rect 100324 13692 102732 13748
rect 102788 13692 102798 13748
rect 71362 13580 71372 13636
rect 71428 13580 72492 13636
rect 72548 13580 75068 13636
rect 75124 13580 75134 13636
rect 77074 13580 77084 13636
rect 77140 13580 79324 13636
rect 79380 13580 79390 13636
rect 84550 13580 84588 13636
rect 84644 13580 84654 13636
rect 84924 13580 87500 13636
rect 87556 13580 87566 13636
rect 19058 13468 19068 13524
rect 19124 13468 19740 13524
rect 19796 13468 20412 13524
rect 20468 13468 20972 13524
rect 21028 13468 21038 13524
rect 21858 13468 21868 13524
rect 21924 13468 26908 13524
rect 34178 13468 34188 13524
rect 34244 13468 35084 13524
rect 35140 13468 35150 13524
rect 35746 13468 35756 13524
rect 35812 13468 37100 13524
rect 37156 13468 37166 13524
rect 37426 13468 37436 13524
rect 37492 13468 40684 13524
rect 40740 13468 40750 13524
rect 48066 13468 48076 13524
rect 48132 13468 51100 13524
rect 51156 13468 51166 13524
rect 58594 13468 58604 13524
rect 58660 13468 59332 13524
rect 60498 13468 60508 13524
rect 60564 13468 61628 13524
rect 61684 13468 61694 13524
rect 70242 13468 70252 13524
rect 70308 13468 72380 13524
rect 72436 13468 72446 13524
rect 74386 13468 74396 13524
rect 74452 13468 78204 13524
rect 78260 13468 78270 13524
rect 79090 13468 79100 13524
rect 79156 13468 81116 13524
rect 81172 13468 81182 13524
rect 81890 13468 81900 13524
rect 81956 13468 82796 13524
rect 82852 13468 82862 13524
rect 83906 13468 83916 13524
rect 83972 13468 87276 13524
rect 87332 13468 87342 13524
rect 59276 13412 59332 13468
rect 87724 13412 87780 13692
rect 87938 13580 87948 13636
rect 88004 13580 90524 13636
rect 90580 13580 90590 13636
rect 93090 13580 93100 13636
rect 93156 13580 95228 13636
rect 95284 13580 95294 13636
rect 104514 13580 104524 13636
rect 104580 13580 106204 13636
rect 106260 13580 107548 13636
rect 107604 13580 109004 13636
rect 109060 13580 109070 13636
rect 90850 13468 90860 13524
rect 90916 13468 91196 13524
rect 91252 13468 91262 13524
rect 94658 13468 94668 13524
rect 94724 13468 96180 13524
rect 98802 13468 98812 13524
rect 98868 13468 103964 13524
rect 104020 13468 104030 13524
rect 105634 13468 105644 13524
rect 105700 13468 108108 13524
rect 108164 13468 108174 13524
rect 110338 13468 110348 13524
rect 110404 13468 111132 13524
rect 111188 13468 111198 13524
rect 96124 13412 96180 13468
rect 27346 13356 27356 13412
rect 27412 13356 28252 13412
rect 28308 13356 28318 13412
rect 31714 13356 31724 13412
rect 31780 13356 32172 13412
rect 32228 13356 32238 13412
rect 45154 13356 45164 13412
rect 45220 13356 50988 13412
rect 51044 13356 51054 13412
rect 59266 13356 59276 13412
rect 59332 13356 59342 13412
rect 61058 13356 61068 13412
rect 61124 13356 61516 13412
rect 61572 13356 61582 13412
rect 67106 13356 67116 13412
rect 67172 13356 73948 13412
rect 83458 13356 83468 13412
rect 83524 13356 87780 13412
rect 89394 13356 89404 13412
rect 89460 13356 91084 13412
rect 91140 13356 91150 13412
rect 96124 13356 96348 13412
rect 96404 13356 96414 13412
rect 103170 13356 103180 13412
rect 103236 13356 103516 13412
rect 103572 13356 103582 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 73892 13300 73948 13356
rect 89404 13300 89460 13356
rect 96626 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96910 13356
rect 127346 13300 127356 13356
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127620 13300 127630 13356
rect 158066 13300 158076 13356
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158340 13300 158350 13356
rect 20066 13244 20076 13300
rect 20132 13244 21420 13300
rect 21476 13244 24220 13300
rect 24276 13244 26124 13300
rect 26180 13244 26684 13300
rect 26740 13244 31500 13300
rect 31556 13244 31566 13300
rect 59938 13244 59948 13300
rect 60004 13244 60732 13300
rect 60788 13244 60798 13300
rect 60946 13244 60956 13300
rect 61012 13244 61404 13300
rect 61460 13244 62748 13300
rect 62804 13244 62814 13300
rect 68786 13244 68796 13300
rect 68852 13244 72828 13300
rect 72884 13244 73724 13300
rect 73780 13244 73790 13300
rect 73892 13244 89460 13300
rect 98802 13244 98812 13300
rect 98868 13244 99596 13300
rect 99652 13244 102508 13300
rect 102564 13244 102574 13300
rect 103394 13244 103404 13300
rect 103460 13244 108668 13300
rect 108724 13244 108734 13300
rect 31938 13132 31948 13188
rect 32004 13132 32284 13188
rect 32340 13132 32350 13188
rect 38098 13132 38108 13188
rect 38164 13132 38780 13188
rect 38836 13132 48076 13188
rect 48132 13132 48142 13188
rect 49382 13132 49420 13188
rect 49476 13132 49486 13188
rect 60050 13132 60060 13188
rect 60116 13132 60620 13188
rect 60676 13132 60686 13188
rect 61730 13132 61740 13188
rect 61796 13132 69132 13188
rect 69188 13132 69198 13188
rect 84252 13132 85820 13188
rect 85876 13132 85886 13188
rect 88386 13132 88396 13188
rect 88452 13132 90076 13188
rect 90132 13132 90142 13188
rect 91746 13132 91756 13188
rect 91812 13132 91980 13188
rect 92036 13132 92046 13188
rect 97346 13132 97356 13188
rect 97412 13132 103292 13188
rect 103348 13132 103358 13188
rect 105298 13132 105308 13188
rect 105364 13132 108892 13188
rect 108948 13132 109116 13188
rect 109172 13132 109182 13188
rect 17826 13020 17836 13076
rect 17892 13020 19852 13076
rect 19908 13020 19918 13076
rect 24658 13020 24668 13076
rect 24724 13020 25452 13076
rect 25508 13020 25518 13076
rect 42802 13020 42812 13076
rect 42868 13020 43932 13076
rect 43988 13020 43998 13076
rect 49746 13020 49756 13076
rect 49812 13020 50316 13076
rect 50372 13020 50382 13076
rect 59490 13020 59500 13076
rect 59556 13020 63420 13076
rect 63476 13020 63868 13076
rect 63924 13020 64092 13076
rect 64148 13020 64158 13076
rect 70578 13020 70588 13076
rect 70644 13020 72268 13076
rect 72324 13020 72334 13076
rect 74162 13020 74172 13076
rect 74228 13020 79884 13076
rect 79940 13020 79950 13076
rect 81554 13020 81564 13076
rect 81620 13020 83804 13076
rect 83860 13020 83870 13076
rect 84252 12964 84308 13132
rect 88274 13020 88284 13076
rect 88340 13020 98644 13076
rect 107650 13020 107660 13076
rect 107716 13020 108220 13076
rect 108276 13020 110348 13076
rect 110404 13020 110414 13076
rect 98588 12964 98644 13020
rect 30818 12908 30828 12964
rect 30884 12908 32508 12964
rect 32564 12908 33964 12964
rect 34020 12908 34030 12964
rect 36642 12908 36652 12964
rect 36708 12908 38332 12964
rect 38388 12908 38398 12964
rect 49606 12908 49644 12964
rect 49700 12908 49710 12964
rect 52994 12908 53004 12964
rect 53060 12908 54348 12964
rect 54404 12908 55916 12964
rect 55972 12908 55982 12964
rect 59826 12908 59836 12964
rect 59892 12908 84252 12964
rect 84308 12908 84318 12964
rect 84802 12908 84812 12964
rect 84868 12908 86492 12964
rect 86548 12908 86558 12964
rect 88694 12908 88732 12964
rect 88788 12908 88798 12964
rect 88946 12908 88956 12964
rect 89012 12908 90076 12964
rect 90132 12908 90524 12964
rect 90580 12908 91308 12964
rect 91364 12908 91756 12964
rect 91812 12908 91822 12964
rect 93986 12908 93996 12964
rect 94052 12908 94062 12964
rect 96338 12908 96348 12964
rect 96404 12908 97804 12964
rect 97860 12908 97870 12964
rect 98588 12908 99708 12964
rect 99764 12908 100156 12964
rect 100212 12908 100222 12964
rect 100818 12908 100828 12964
rect 100884 12908 102844 12964
rect 102900 12908 102910 12964
rect 106530 12908 106540 12964
rect 106596 12908 109564 12964
rect 109620 12908 109630 12964
rect 110002 12908 110012 12964
rect 110068 12908 112140 12964
rect 112196 12908 112206 12964
rect 93996 12852 94052 12908
rect 29922 12796 29932 12852
rect 29988 12796 30940 12852
rect 30996 12796 31006 12852
rect 32834 12796 32844 12852
rect 32900 12796 34972 12852
rect 35028 12796 36988 12852
rect 37044 12796 37884 12852
rect 37940 12796 37950 12852
rect 44818 12796 44828 12852
rect 44884 12796 45836 12852
rect 45892 12796 49308 12852
rect 49364 12796 50876 12852
rect 50932 12796 50942 12852
rect 56802 12796 56812 12852
rect 56868 12796 57708 12852
rect 57764 12796 57774 12852
rect 60582 12796 60620 12852
rect 60676 12796 60686 12852
rect 66994 12796 67004 12852
rect 67060 12796 74508 12852
rect 74564 12796 78540 12852
rect 78596 12796 78606 12852
rect 82786 12796 82796 12852
rect 82852 12796 84476 12852
rect 84532 12796 84542 12852
rect 89282 12796 89292 12852
rect 89348 12796 89516 12852
rect 89572 12796 89582 12852
rect 90850 12796 90860 12852
rect 90916 12796 94052 12852
rect 100258 12796 100268 12852
rect 100324 12796 101276 12852
rect 101332 12796 101342 12852
rect 107660 12796 111692 12852
rect 111748 12796 111758 12852
rect 112690 12796 112700 12852
rect 112756 12796 121772 12852
rect 121828 12796 121838 12852
rect 107660 12740 107716 12796
rect 18610 12684 18620 12740
rect 18676 12684 19628 12740
rect 19684 12684 25004 12740
rect 25060 12684 25070 12740
rect 27122 12684 27132 12740
rect 27188 12684 28364 12740
rect 28420 12684 32060 12740
rect 32116 12684 33852 12740
rect 33908 12684 33918 12740
rect 47282 12684 47292 12740
rect 47348 12684 48524 12740
rect 48580 12684 49532 12740
rect 49588 12684 49598 12740
rect 57026 12684 57036 12740
rect 57092 12684 58828 12740
rect 58884 12684 58894 12740
rect 73938 12684 73948 12740
rect 74004 12684 74844 12740
rect 74900 12684 75292 12740
rect 75348 12684 75358 12740
rect 78082 12684 78092 12740
rect 78148 12684 80220 12740
rect 80276 12684 83244 12740
rect 83300 12684 83310 12740
rect 88274 12684 88284 12740
rect 88340 12684 89292 12740
rect 89348 12684 89358 12740
rect 89590 12684 89628 12740
rect 89684 12684 89694 12740
rect 91522 12684 91532 12740
rect 91588 12684 92204 12740
rect 92260 12684 92270 12740
rect 92866 12684 92876 12740
rect 92932 12684 93996 12740
rect 94052 12684 94062 12740
rect 96450 12684 96460 12740
rect 96516 12684 106428 12740
rect 106484 12684 106988 12740
rect 107044 12684 107054 12740
rect 107650 12684 107660 12740
rect 107716 12684 107726 12740
rect 107874 12684 107884 12740
rect 107940 12684 109676 12740
rect 109732 12684 109742 12740
rect 111234 12684 111244 12740
rect 111300 12684 113820 12740
rect 113876 12684 113886 12740
rect 29586 12572 29596 12628
rect 29652 12572 30604 12628
rect 30660 12572 35084 12628
rect 35140 12572 35150 12628
rect 52770 12572 52780 12628
rect 52836 12572 53452 12628
rect 53508 12572 54460 12628
rect 54516 12572 69692 12628
rect 69748 12572 69758 12628
rect 70130 12572 70140 12628
rect 70196 12572 79660 12628
rect 79716 12572 79726 12628
rect 88050 12572 88060 12628
rect 88116 12572 103628 12628
rect 103684 12572 103694 12628
rect 104850 12572 104860 12628
rect 104916 12572 110908 12628
rect 110964 12572 110974 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 81266 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81550 12572
rect 103628 12516 103684 12572
rect 111986 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112270 12572
rect 142706 12516 142716 12572
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142980 12516 142990 12572
rect 20188 12460 31052 12516
rect 31108 12460 31118 12516
rect 43138 12460 43148 12516
rect 43204 12460 45836 12516
rect 45892 12460 45902 12516
rect 46386 12460 46396 12516
rect 46452 12460 47180 12516
rect 47236 12460 47246 12516
rect 47506 12460 47516 12516
rect 47572 12460 50316 12516
rect 50372 12460 50382 12516
rect 53554 12460 53564 12516
rect 53620 12460 54684 12516
rect 54740 12460 58380 12516
rect 58436 12460 60508 12516
rect 60564 12460 60574 12516
rect 60834 12460 60844 12516
rect 60900 12460 61404 12516
rect 61460 12460 61516 12516
rect 61572 12460 61582 12516
rect 72818 12460 72828 12516
rect 72884 12460 73724 12516
rect 73780 12460 73790 12516
rect 87266 12460 87276 12516
rect 87332 12460 91868 12516
rect 91924 12460 92988 12516
rect 93044 12460 93054 12516
rect 103628 12460 110796 12516
rect 110852 12460 110862 12516
rect 20188 12404 20244 12460
rect 15586 12348 15596 12404
rect 15652 12348 18172 12404
rect 18228 12348 18956 12404
rect 19012 12348 20244 12404
rect 23314 12348 23324 12404
rect 23380 12348 23996 12404
rect 24052 12348 24062 12404
rect 24770 12348 24780 12404
rect 24836 12348 25788 12404
rect 25844 12348 29148 12404
rect 29204 12348 37324 12404
rect 37380 12348 37390 12404
rect 41794 12348 41804 12404
rect 41860 12348 43820 12404
rect 43876 12348 43886 12404
rect 45602 12348 45612 12404
rect 45668 12348 46956 12404
rect 47012 12348 47022 12404
rect 47954 12348 47964 12404
rect 48020 12348 50428 12404
rect 52210 12348 52220 12404
rect 52276 12348 53452 12404
rect 53508 12348 56028 12404
rect 56084 12348 57036 12404
rect 57092 12348 57102 12404
rect 57250 12348 57260 12404
rect 57316 12348 70756 12404
rect 21522 12236 21532 12292
rect 21588 12236 22428 12292
rect 22484 12236 22494 12292
rect 23996 12236 25564 12292
rect 25620 12236 26236 12292
rect 26292 12236 26302 12292
rect 29698 12236 29708 12292
rect 29764 12236 32844 12292
rect 32900 12236 32910 12292
rect 42354 12236 42364 12292
rect 42420 12236 48748 12292
rect 48804 12236 48814 12292
rect 49298 12236 49308 12292
rect 49364 12236 49756 12292
rect 49812 12236 49822 12292
rect 23996 12180 24052 12236
rect 50372 12180 50428 12348
rect 50754 12236 50764 12292
rect 50820 12236 51996 12292
rect 52052 12236 52062 12292
rect 55122 12236 55132 12292
rect 55188 12236 61292 12292
rect 61348 12236 61740 12292
rect 61796 12236 61806 12292
rect 17714 12124 17724 12180
rect 17780 12124 19628 12180
rect 19684 12124 19694 12180
rect 20962 12124 20972 12180
rect 21028 12124 21756 12180
rect 21812 12124 21822 12180
rect 22194 12124 22204 12180
rect 22260 12124 22876 12180
rect 22932 12124 24052 12180
rect 24546 12124 24556 12180
rect 24612 12124 25340 12180
rect 25396 12124 25406 12180
rect 27682 12124 27692 12180
rect 27748 12124 28812 12180
rect 28868 12124 30268 12180
rect 30324 12124 30334 12180
rect 30930 12124 30940 12180
rect 30996 12124 35532 12180
rect 35588 12124 35598 12180
rect 37650 12124 37660 12180
rect 37716 12124 39228 12180
rect 39284 12124 39294 12180
rect 40002 12124 40012 12180
rect 40068 12124 40908 12180
rect 40964 12124 40974 12180
rect 41906 12124 41916 12180
rect 41972 12124 46172 12180
rect 46228 12124 46238 12180
rect 46610 12124 46620 12180
rect 46676 12124 48860 12180
rect 48916 12124 49084 12180
rect 49140 12124 49868 12180
rect 49924 12124 50204 12180
rect 50260 12124 50270 12180
rect 50372 12124 51100 12180
rect 51156 12124 52892 12180
rect 52948 12124 52958 12180
rect 54898 12124 54908 12180
rect 54964 12124 54974 12180
rect 55906 12124 55916 12180
rect 55972 12124 56924 12180
rect 56980 12124 58716 12180
rect 58772 12124 58782 12180
rect 63074 12124 63084 12180
rect 63140 12124 70476 12180
rect 70532 12124 70542 12180
rect 18946 12012 18956 12068
rect 19012 12012 19964 12068
rect 20020 12012 20030 12068
rect 20972 11956 21028 12124
rect 41916 12068 41972 12124
rect 54908 12068 54964 12124
rect 70700 12068 70756 12348
rect 73724 12292 73780 12460
rect 83906 12348 83916 12404
rect 83972 12348 85708 12404
rect 85764 12348 85774 12404
rect 86482 12348 86492 12404
rect 86548 12348 88060 12404
rect 88116 12348 88126 12404
rect 90290 12348 90300 12404
rect 90356 12348 94556 12404
rect 94612 12348 94622 12404
rect 102498 12348 102508 12404
rect 102564 12348 103628 12404
rect 103684 12348 103694 12404
rect 105970 12348 105980 12404
rect 106036 12348 108668 12404
rect 108724 12348 108734 12404
rect 109330 12348 109340 12404
rect 109396 12348 112700 12404
rect 112756 12348 112766 12404
rect 73724 12236 75852 12292
rect 75908 12236 77196 12292
rect 77252 12236 77262 12292
rect 77410 12236 77420 12292
rect 77476 12236 78540 12292
rect 78596 12236 79436 12292
rect 79492 12236 79502 12292
rect 79650 12236 79660 12292
rect 79716 12236 82404 12292
rect 72706 12124 72716 12180
rect 72772 12124 74508 12180
rect 74564 12124 74574 12180
rect 78754 12124 78764 12180
rect 78820 12124 80108 12180
rect 80164 12124 80780 12180
rect 80836 12124 80846 12180
rect 82348 12068 82404 12236
rect 85652 12236 85820 12292
rect 85876 12236 85886 12292
rect 86146 12236 86156 12292
rect 86212 12236 88508 12292
rect 88564 12236 88574 12292
rect 94556 12236 95564 12292
rect 95620 12236 98140 12292
rect 98196 12236 98206 12292
rect 102582 12236 102620 12292
rect 102676 12236 102686 12292
rect 107986 12236 107996 12292
rect 108052 12236 108062 12292
rect 108546 12236 108556 12292
rect 108612 12236 112980 12292
rect 83234 12124 83244 12180
rect 83300 12124 84252 12180
rect 84308 12124 84318 12180
rect 25442 12012 25452 12068
rect 25508 12012 32060 12068
rect 32116 12012 32126 12068
rect 36530 12012 36540 12068
rect 36596 12012 41972 12068
rect 42700 12012 44044 12068
rect 44100 12012 54964 12068
rect 57026 12012 57036 12068
rect 57092 12012 59836 12068
rect 59892 12012 59902 12068
rect 65986 12012 65996 12068
rect 66052 12012 67116 12068
rect 67172 12012 67182 12068
rect 70700 12012 81564 12068
rect 81620 12012 81630 12068
rect 82348 12012 84700 12068
rect 84756 12012 84766 12068
rect 85110 12012 85148 12068
rect 85204 12012 85214 12068
rect 42700 11956 42756 12012
rect 65996 11956 66052 12012
rect 19170 11900 19180 11956
rect 19236 11900 21028 11956
rect 25218 11900 25228 11956
rect 25284 11900 26796 11956
rect 26852 11900 27132 11956
rect 27188 11900 27580 11956
rect 27636 11900 27646 11956
rect 30818 11900 30828 11956
rect 30884 11900 40180 11956
rect 40338 11900 40348 11956
rect 40404 11900 42756 11956
rect 42914 11900 42924 11956
rect 42980 11900 43708 11956
rect 43764 11900 43774 11956
rect 49298 11900 49308 11956
rect 49364 11900 49644 11956
rect 49700 11900 49710 11956
rect 52658 11900 52668 11956
rect 52724 11900 53564 11956
rect 53620 11900 53630 11956
rect 53890 11900 53900 11956
rect 53956 11900 58044 11956
rect 58100 11900 58110 11956
rect 65548 11900 66052 11956
rect 66882 11900 66892 11956
rect 66948 11900 66958 11956
rect 71922 11900 71932 11956
rect 71988 11900 83132 11956
rect 83188 11900 83198 11956
rect 83682 11900 83692 11956
rect 83748 11900 83804 11956
rect 83860 11900 83870 11956
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 19740 11732 19796 11900
rect 40124 11844 40180 11900
rect 21298 11788 21308 11844
rect 21364 11788 22204 11844
rect 22260 11788 22270 11844
rect 23874 11788 23884 11844
rect 23940 11788 24668 11844
rect 24724 11788 26460 11844
rect 26516 11788 26908 11844
rect 26964 11788 26974 11844
rect 27682 11788 27692 11844
rect 27748 11788 28364 11844
rect 28420 11788 28430 11844
rect 36978 11788 36988 11844
rect 37044 11788 37212 11844
rect 37268 11788 39564 11844
rect 39620 11788 39630 11844
rect 40124 11788 40404 11844
rect 42802 11788 42812 11844
rect 42868 11788 43092 11844
rect 43586 11788 43596 11844
rect 43652 11788 45612 11844
rect 45668 11788 45678 11844
rect 45826 11788 45836 11844
rect 45892 11788 62972 11844
rect 63028 11788 63038 11844
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 40328 11732 40348 11788
rect 40404 11732 40414 11788
rect 43036 11732 43092 11788
rect 65548 11732 65604 11900
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 19730 11676 19740 11732
rect 19796 11676 19806 11732
rect 21410 11676 21420 11732
rect 21476 11676 22540 11732
rect 22596 11676 24892 11732
rect 24948 11676 31836 11732
rect 31892 11676 31902 11732
rect 35644 11676 37548 11732
rect 37604 11676 40012 11732
rect 40068 11676 40078 11732
rect 43026 11676 43036 11732
rect 43092 11676 43102 11732
rect 47842 11676 47852 11732
rect 47908 11676 49084 11732
rect 49140 11676 50092 11732
rect 50148 11676 64652 11732
rect 64708 11676 64718 11732
rect 64866 11676 64876 11732
rect 64932 11676 65604 11732
rect 66322 11676 66332 11732
rect 66388 11676 66668 11732
rect 66724 11676 66734 11732
rect 35644 11620 35700 11676
rect 66892 11620 66948 11900
rect 85652 11844 85708 12236
rect 88508 12180 88564 12236
rect 94556 12180 94612 12236
rect 107996 12180 108052 12236
rect 88508 12124 94612 12180
rect 94770 12124 94780 12180
rect 94836 12124 95788 12180
rect 95844 12124 98812 12180
rect 98868 12124 98878 12180
rect 101266 12124 101276 12180
rect 101332 12124 103964 12180
rect 104020 12124 105644 12180
rect 105700 12124 107324 12180
rect 107380 12124 107390 12180
rect 107996 12124 109228 12180
rect 87266 12012 87276 12068
rect 87332 12012 89180 12068
rect 89236 12012 89246 12068
rect 89394 12012 89404 12068
rect 89460 12012 95228 12068
rect 95284 12012 95294 12068
rect 100146 12012 100156 12068
rect 100212 12012 108556 12068
rect 108612 12012 108622 12068
rect 109172 11956 109228 12124
rect 112924 12068 112980 12236
rect 109862 12012 109900 12068
rect 109956 12012 109966 12068
rect 112914 12012 112924 12068
rect 112980 12012 145516 12068
rect 145572 12012 145582 12068
rect 86930 11900 86940 11956
rect 86996 11900 96124 11956
rect 96180 11900 96190 11956
rect 98802 11900 98812 11956
rect 98868 11900 100044 11956
rect 100100 11900 100110 11956
rect 102396 11900 105308 11956
rect 105364 11900 105374 11956
rect 108098 11900 108108 11956
rect 108164 11900 108444 11956
rect 108500 11900 108510 11956
rect 109172 11900 112476 11956
rect 112532 11900 122668 11956
rect 122724 11900 122734 11956
rect 102396 11844 102452 11900
rect 108108 11844 108164 11900
rect 73378 11788 73388 11844
rect 73444 11788 76412 11844
rect 76468 11788 76478 11844
rect 79538 11788 79548 11844
rect 79604 11788 83468 11844
rect 83524 11788 84588 11844
rect 84644 11788 85708 11844
rect 92978 11788 92988 11844
rect 93044 11788 93548 11844
rect 93604 11788 93614 11844
rect 93762 11788 93772 11844
rect 93828 11788 94892 11844
rect 94948 11788 96460 11844
rect 96516 11788 96526 11844
rect 97794 11788 97804 11844
rect 97860 11788 102452 11844
rect 102610 11788 102620 11844
rect 102676 11788 102788 11844
rect 102946 11788 102956 11844
rect 103012 11788 103404 11844
rect 103460 11788 103470 11844
rect 103618 11788 103628 11844
rect 103684 11788 103964 11844
rect 104020 11788 108164 11844
rect 108658 11788 108668 11844
rect 108724 11788 110012 11844
rect 110068 11788 110078 11844
rect 96626 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96910 11788
rect 102722 11732 102732 11788
rect 102788 11732 102798 11788
rect 127346 11732 127356 11788
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127620 11732 127630 11788
rect 158066 11732 158076 11788
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158340 11732 158350 11788
rect 67554 11676 67564 11732
rect 67620 11676 84196 11732
rect 85474 11676 85484 11732
rect 85540 11676 86828 11732
rect 86884 11676 86894 11732
rect 89618 11676 89628 11732
rect 89684 11676 90076 11732
rect 90132 11676 90860 11732
rect 90916 11676 90926 11732
rect 94182 11676 94220 11732
rect 94276 11676 94286 11732
rect 95330 11676 95340 11732
rect 95396 11676 96180 11732
rect 97906 11676 97916 11732
rect 97972 11676 98364 11732
rect 98420 11676 98430 11732
rect 106418 11676 106428 11732
rect 106484 11676 109900 11732
rect 109956 11676 111580 11732
rect 111636 11676 111646 11732
rect 84140 11620 84196 11676
rect 96124 11620 96180 11676
rect 20290 11564 20300 11620
rect 20356 11564 21196 11620
rect 21252 11564 21262 11620
rect 28130 11564 28140 11620
rect 28196 11564 28476 11620
rect 28532 11564 30268 11620
rect 30324 11564 30334 11620
rect 32844 11564 34636 11620
rect 34692 11564 34702 11620
rect 35522 11564 35532 11620
rect 35588 11564 35700 11620
rect 40086 11564 40124 11620
rect 40180 11564 40190 11620
rect 42690 11564 42700 11620
rect 42756 11564 50428 11620
rect 52098 11564 52108 11620
rect 52164 11564 53788 11620
rect 53844 11564 53854 11620
rect 59826 11564 59836 11620
rect 59892 11564 64988 11620
rect 65044 11564 65054 11620
rect 65212 11564 66668 11620
rect 66724 11564 66734 11620
rect 66892 11564 71036 11620
rect 71092 11564 73500 11620
rect 73556 11564 75292 11620
rect 75348 11564 77196 11620
rect 77252 11564 77262 11620
rect 84102 11564 84140 11620
rect 84196 11564 84206 11620
rect 84466 11564 84476 11620
rect 84532 11564 86044 11620
rect 86100 11564 86110 11620
rect 92306 11564 92316 11620
rect 92372 11564 92382 11620
rect 94322 11564 94332 11620
rect 94388 11564 94556 11620
rect 94612 11564 96068 11620
rect 96124 11564 98476 11620
rect 98532 11564 99148 11620
rect 99204 11564 99214 11620
rect 100902 11564 100940 11620
rect 100996 11564 101006 11620
rect 104850 11564 104860 11620
rect 104916 11564 105196 11620
rect 105252 11564 105262 11620
rect 106306 11564 106316 11620
rect 106372 11564 116060 11620
rect 116116 11564 116126 11620
rect 32844 11508 32900 11564
rect 20066 11452 20076 11508
rect 20132 11452 20748 11508
rect 20804 11452 20814 11508
rect 28690 11452 28700 11508
rect 28756 11452 28924 11508
rect 28980 11452 32900 11508
rect 34412 11452 35980 11508
rect 36036 11452 36046 11508
rect 39442 11452 39452 11508
rect 39508 11452 40236 11508
rect 40292 11452 42812 11508
rect 42868 11452 42878 11508
rect 49410 11452 49420 11508
rect 49476 11452 49644 11508
rect 49700 11452 49710 11508
rect 20514 11340 20524 11396
rect 20580 11340 24332 11396
rect 24388 11340 24398 11396
rect 29922 11340 29932 11396
rect 29988 11340 30828 11396
rect 30884 11340 30894 11396
rect 34412 11284 34468 11452
rect 35410 11340 35420 11396
rect 35476 11340 37996 11396
rect 38052 11340 38556 11396
rect 38612 11340 40012 11396
rect 40068 11340 40078 11396
rect 40226 11340 40236 11396
rect 40292 11340 42476 11396
rect 42532 11340 42542 11396
rect 47618 11340 47628 11396
rect 47684 11340 48524 11396
rect 48580 11340 48590 11396
rect 50372 11284 50428 11564
rect 51762 11452 51772 11508
rect 51828 11452 52780 11508
rect 52836 11452 52846 11508
rect 58706 11452 58716 11508
rect 58772 11452 60060 11508
rect 60116 11452 60126 11508
rect 60722 11452 60732 11508
rect 60788 11452 61628 11508
rect 61684 11452 61694 11508
rect 61926 11452 61964 11508
rect 62020 11452 62030 11508
rect 65212 11396 65268 11564
rect 92316 11508 92372 11564
rect 96012 11508 96068 11564
rect 66210 11452 66220 11508
rect 66276 11452 68124 11508
rect 68180 11452 68190 11508
rect 68338 11452 68348 11508
rect 68404 11452 89404 11508
rect 89460 11452 89470 11508
rect 91970 11452 91980 11508
rect 92036 11452 94668 11508
rect 94724 11452 94734 11508
rect 95218 11452 95228 11508
rect 95284 11452 95788 11508
rect 95844 11452 95854 11508
rect 96012 11452 97916 11508
rect 97972 11452 97982 11508
rect 100594 11452 100604 11508
rect 100660 11452 101836 11508
rect 101892 11452 101902 11508
rect 105074 11452 105084 11508
rect 105140 11452 105420 11508
rect 105476 11452 105486 11508
rect 108780 11452 109452 11508
rect 109508 11452 109518 11508
rect 111010 11452 111020 11508
rect 111076 11452 112812 11508
rect 112868 11452 112878 11508
rect 51650 11340 51660 11396
rect 51716 11340 53004 11396
rect 53060 11340 53070 11396
rect 53900 11340 57484 11396
rect 57540 11340 57550 11396
rect 61842 11340 61852 11396
rect 61908 11340 61918 11396
rect 62066 11340 62076 11396
rect 62132 11340 64204 11396
rect 64260 11340 64270 11396
rect 64764 11340 65268 11396
rect 65426 11340 65436 11396
rect 65492 11340 70140 11396
rect 70196 11340 70206 11396
rect 71586 11340 71596 11396
rect 71652 11340 72156 11396
rect 72212 11340 72222 11396
rect 73042 11340 73052 11396
rect 73108 11340 74396 11396
rect 74452 11340 74462 11396
rect 74834 11340 74844 11396
rect 74900 11340 76076 11396
rect 76132 11340 76142 11396
rect 76290 11340 76300 11396
rect 76356 11340 76524 11396
rect 76580 11340 76972 11396
rect 77028 11340 77038 11396
rect 78194 11340 78204 11396
rect 78260 11340 83580 11396
rect 83636 11340 83646 11396
rect 84130 11340 84140 11396
rect 84196 11340 84364 11396
rect 84420 11340 84430 11396
rect 85026 11340 85036 11396
rect 85092 11340 86268 11396
rect 86324 11340 86334 11396
rect 88498 11340 88508 11396
rect 88564 11340 102956 11396
rect 103012 11340 104076 11396
rect 104132 11340 104142 11396
rect 53900 11284 53956 11340
rect 61852 11284 61908 11340
rect 18946 11228 18956 11284
rect 19012 11228 19404 11284
rect 19460 11228 21644 11284
rect 21700 11228 21710 11284
rect 29932 11228 34468 11284
rect 35074 11228 35084 11284
rect 35140 11228 37660 11284
rect 37716 11228 39004 11284
rect 39060 11228 39070 11284
rect 39330 11228 39340 11284
rect 39396 11228 41244 11284
rect 41300 11228 41310 11284
rect 42578 11228 42588 11284
rect 42644 11228 44940 11284
rect 44996 11228 45006 11284
rect 48178 11228 48188 11284
rect 48244 11228 48860 11284
rect 48916 11228 49532 11284
rect 49588 11228 49598 11284
rect 50372 11228 53956 11284
rect 54114 11228 54124 11284
rect 54180 11228 55580 11284
rect 55636 11228 55646 11284
rect 58258 11228 58268 11284
rect 58324 11228 60508 11284
rect 60564 11228 60574 11284
rect 61852 11228 64540 11284
rect 64596 11228 64606 11284
rect 29932 11172 29988 11228
rect 42588 11172 42644 11228
rect 64764 11172 64820 11340
rect 108780 11284 108836 11452
rect 109004 11340 112140 11396
rect 112196 11340 112206 11396
rect 64978 11228 64988 11284
rect 65044 11228 66556 11284
rect 66612 11228 66892 11284
rect 66948 11228 66958 11284
rect 70018 11228 70028 11284
rect 70084 11228 72380 11284
rect 72436 11228 73724 11284
rect 73780 11228 78988 11284
rect 79044 11228 79054 11284
rect 81554 11228 81564 11284
rect 81620 11228 84476 11284
rect 84532 11228 86380 11284
rect 86436 11228 86446 11284
rect 93090 11228 93100 11284
rect 93156 11228 93660 11284
rect 93716 11228 93726 11284
rect 102610 11228 102620 11284
rect 102676 11228 102844 11284
rect 102900 11228 102910 11284
rect 103394 11228 103404 11284
rect 103460 11228 106036 11284
rect 106194 11228 106204 11284
rect 106260 11228 107548 11284
rect 107604 11228 107614 11284
rect 108770 11228 108780 11284
rect 108836 11228 108846 11284
rect 105980 11172 106036 11228
rect 109004 11172 109060 11340
rect 111906 11228 111916 11284
rect 111972 11228 112364 11284
rect 112420 11228 112430 11284
rect 18162 11116 18172 11172
rect 18228 11116 20188 11172
rect 20244 11116 20254 11172
rect 22866 11116 22876 11172
rect 22932 11116 25340 11172
rect 25396 11116 29260 11172
rect 29316 11116 29326 11172
rect 29922 11116 29932 11172
rect 29988 11116 29998 11172
rect 34290 11116 34300 11172
rect 34356 11116 36092 11172
rect 36148 11116 36158 11172
rect 40226 11116 40236 11172
rect 40292 11116 42644 11172
rect 45154 11116 45164 11172
rect 45220 11116 45836 11172
rect 45892 11116 56700 11172
rect 56756 11116 59948 11172
rect 60004 11116 60014 11172
rect 61618 11116 61628 11172
rect 61684 11116 61964 11172
rect 62020 11116 62030 11172
rect 62132 11116 64820 11172
rect 65090 11116 65100 11172
rect 65156 11116 66444 11172
rect 66500 11116 66510 11172
rect 66658 11116 66668 11172
rect 66724 11116 67788 11172
rect 67844 11116 67854 11172
rect 69010 11116 69020 11172
rect 69076 11116 70924 11172
rect 70980 11116 71484 11172
rect 71540 11116 71550 11172
rect 71698 11116 71708 11172
rect 71764 11116 71802 11172
rect 71922 11116 71932 11172
rect 71988 11116 72716 11172
rect 72772 11116 75572 11172
rect 75702 11116 75740 11172
rect 75796 11116 75806 11172
rect 76178 11116 76188 11172
rect 76244 11116 76972 11172
rect 77028 11116 77038 11172
rect 79090 11116 79100 11172
rect 79156 11116 79772 11172
rect 79828 11116 79838 11172
rect 80434 11116 80444 11172
rect 80500 11116 84924 11172
rect 84980 11116 84990 11172
rect 88834 11116 88844 11172
rect 88900 11116 90636 11172
rect 90692 11116 90702 11172
rect 91634 11116 91644 11172
rect 91700 11116 92988 11172
rect 93044 11116 94220 11172
rect 94276 11116 94286 11172
rect 96338 11116 96348 11172
rect 96404 11116 97020 11172
rect 97076 11116 97086 11172
rect 99810 11116 99820 11172
rect 99876 11116 99886 11172
rect 102498 11116 102508 11172
rect 102564 11116 103180 11172
rect 103236 11116 103852 11172
rect 103908 11116 103918 11172
rect 104290 11116 104300 11172
rect 104356 11116 105364 11172
rect 105980 11116 109060 11172
rect 109172 11116 113036 11172
rect 113092 11116 113102 11172
rect 62132 11060 62188 11116
rect 20290 11004 20300 11060
rect 20356 11004 21420 11060
rect 21476 11004 21486 11060
rect 21634 11004 21644 11060
rect 21700 11004 22092 11060
rect 22148 11004 35756 11060
rect 35812 11004 35822 11060
rect 37538 11004 37548 11060
rect 37604 11004 43092 11060
rect 43894 11004 43932 11060
rect 43988 11004 43998 11060
rect 44146 11004 44156 11060
rect 44212 11004 44222 11060
rect 49494 11004 49532 11060
rect 49588 11004 49598 11060
rect 50278 11004 50316 11060
rect 50372 11004 50382 11060
rect 57138 11004 57148 11060
rect 57204 11004 57214 11060
rect 58818 11004 58828 11060
rect 58884 11004 62188 11060
rect 64306 11004 64316 11060
rect 64372 11004 67564 11060
rect 67620 11004 67630 11060
rect 67890 11004 67900 11060
rect 67956 11004 69468 11060
rect 69524 11004 70252 11060
rect 70308 11004 70318 11060
rect 71362 11004 71372 11060
rect 71428 11004 72828 11060
rect 72884 11004 72894 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 43036 10948 43092 11004
rect 28018 10892 28028 10948
rect 28084 10892 36988 10948
rect 37044 10892 38332 10948
rect 38388 10892 38398 10948
rect 38612 10892 38780 10948
rect 38836 10892 38846 10948
rect 40086 10892 40124 10948
rect 40180 10892 40190 10948
rect 43026 10892 43036 10948
rect 43092 10892 43102 10948
rect 38612 10836 38668 10892
rect 22978 10780 22988 10836
rect 23044 10780 23884 10836
rect 23940 10780 23950 10836
rect 26114 10780 26124 10836
rect 26180 10780 27244 10836
rect 27300 10780 30828 10836
rect 30884 10780 30894 10836
rect 31378 10780 31388 10836
rect 31444 10780 36540 10836
rect 36596 10780 36606 10836
rect 38444 10780 38668 10836
rect 40338 10780 40348 10836
rect 40404 10780 41916 10836
rect 41972 10780 42588 10836
rect 42644 10780 42654 10836
rect 16930 10668 16940 10724
rect 16996 10668 28924 10724
rect 28980 10668 28990 10724
rect 29922 10668 29932 10724
rect 29988 10668 31612 10724
rect 31668 10668 31678 10724
rect 32498 10668 32508 10724
rect 32564 10668 33404 10724
rect 33460 10668 33470 10724
rect 38444 10612 38500 10780
rect 44156 10724 44212 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 51538 10892 51548 10948
rect 51604 10892 55916 10948
rect 55972 10892 55982 10948
rect 46022 10780 46060 10836
rect 46116 10780 46126 10836
rect 49186 10780 49196 10836
rect 49252 10780 51996 10836
rect 52052 10780 52062 10836
rect 54002 10780 54012 10836
rect 54068 10780 54460 10836
rect 54516 10780 55468 10836
rect 55524 10780 56588 10836
rect 56644 10780 56654 10836
rect 57148 10724 57204 11004
rect 75516 10948 75572 11116
rect 75842 11004 75852 11060
rect 75908 11004 76748 11060
rect 76804 11004 77868 11060
rect 77924 11004 77934 11060
rect 85652 11004 86940 11060
rect 86996 11004 94108 11060
rect 94164 11004 94174 11060
rect 94332 11004 98252 11060
rect 98308 11004 98318 11060
rect 81266 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81550 11004
rect 85652 10948 85708 11004
rect 94332 10948 94388 11004
rect 99820 10948 99876 11116
rect 105308 11060 105364 11116
rect 109172 11060 109228 11116
rect 100940 11004 104748 11060
rect 104804 11004 104814 11060
rect 105308 11004 105532 11060
rect 105588 11004 109228 11060
rect 100940 10948 100996 11004
rect 111986 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112270 11004
rect 142706 10948 142716 11004
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142980 10948 142990 11004
rect 61926 10892 61964 10948
rect 62020 10892 62030 10948
rect 64642 10892 64652 10948
rect 64708 10892 65436 10948
rect 65492 10892 65502 10948
rect 68002 10892 68012 10948
rect 68068 10892 69356 10948
rect 69412 10892 69804 10948
rect 69860 10892 71932 10948
rect 71988 10892 71998 10948
rect 75516 10892 80444 10948
rect 80500 10892 80510 10948
rect 83570 10892 83580 10948
rect 83636 10892 85484 10948
rect 85540 10892 85708 10948
rect 87378 10892 87388 10948
rect 87444 10892 89628 10948
rect 89684 10892 90972 10948
rect 91028 10892 94388 10948
rect 94658 10892 94668 10948
rect 94724 10892 99876 10948
rect 100930 10892 100940 10948
rect 100996 10892 101006 10948
rect 102834 10892 102844 10948
rect 102900 10892 103292 10948
rect 103348 10892 110572 10948
rect 110628 10892 110638 10948
rect 59266 10780 59276 10836
rect 59332 10780 60844 10836
rect 60900 10780 60910 10836
rect 61068 10780 62412 10836
rect 62468 10780 62860 10836
rect 62916 10780 75740 10836
rect 75796 10780 75806 10836
rect 76962 10780 76972 10836
rect 77028 10780 78204 10836
rect 78260 10780 78270 10836
rect 78978 10780 78988 10836
rect 79044 10780 81452 10836
rect 81508 10780 81518 10836
rect 83878 10780 83916 10836
rect 83972 10780 83982 10836
rect 91522 10780 91532 10836
rect 91588 10780 92204 10836
rect 92260 10780 94556 10836
rect 94612 10780 94622 10836
rect 95330 10780 95340 10836
rect 95396 10780 96796 10836
rect 96852 10780 96862 10836
rect 99810 10780 99820 10836
rect 99876 10780 101164 10836
rect 101220 10780 101230 10836
rect 103842 10780 103852 10836
rect 103908 10780 106316 10836
rect 106372 10780 106382 10836
rect 110898 10780 110908 10836
rect 110964 10780 118300 10836
rect 118356 10780 118366 10836
rect 61068 10724 61124 10780
rect 39666 10668 39676 10724
rect 39732 10668 42140 10724
rect 42196 10668 44324 10724
rect 53778 10668 53788 10724
rect 53844 10668 56924 10724
rect 56980 10668 56990 10724
rect 57148 10668 61124 10724
rect 62178 10668 62188 10724
rect 62244 10668 62972 10724
rect 63028 10668 67228 10724
rect 67284 10668 67294 10724
rect 67890 10668 67900 10724
rect 67956 10668 71372 10724
rect 71428 10668 71438 10724
rect 44268 10612 44324 10668
rect 57260 10612 57316 10668
rect 76972 10612 77028 10780
rect 79650 10668 79660 10724
rect 79716 10668 83972 10724
rect 84914 10668 84924 10724
rect 84980 10668 84990 10724
rect 92082 10668 92092 10724
rect 92148 10668 92652 10724
rect 92708 10668 92718 10724
rect 94108 10668 94444 10724
rect 94500 10668 103908 10724
rect 106054 10668 106092 10724
rect 106148 10668 106158 10724
rect 106642 10668 106652 10724
rect 106708 10668 109452 10724
rect 109508 10668 109518 10724
rect 110002 10668 110012 10724
rect 110068 10668 117292 10724
rect 117348 10668 117358 10724
rect 83916 10612 83972 10668
rect 84924 10612 84980 10668
rect 94108 10612 94164 10668
rect 17490 10556 17500 10612
rect 17556 10556 18508 10612
rect 18564 10556 18574 10612
rect 20962 10556 20972 10612
rect 21028 10556 21420 10612
rect 21476 10556 22092 10612
rect 22148 10556 26572 10612
rect 26628 10556 28028 10612
rect 28084 10556 28094 10612
rect 30930 10556 30940 10612
rect 30996 10556 33068 10612
rect 33124 10556 33134 10612
rect 35074 10556 35084 10612
rect 35140 10556 38500 10612
rect 38658 10556 38668 10612
rect 38724 10556 41356 10612
rect 41412 10556 43596 10612
rect 43652 10556 43662 10612
rect 44258 10556 44268 10612
rect 44324 10556 44334 10612
rect 44566 10556 44604 10612
rect 44660 10556 44670 10612
rect 46722 10556 46732 10612
rect 46788 10556 49196 10612
rect 49252 10556 50204 10612
rect 50260 10556 50270 10612
rect 53666 10556 53676 10612
rect 53732 10556 54572 10612
rect 54628 10556 54638 10612
rect 56130 10556 56140 10612
rect 56196 10556 57260 10612
rect 57316 10556 57326 10612
rect 63074 10556 63084 10612
rect 63140 10556 63420 10612
rect 63476 10556 63486 10612
rect 63970 10556 63980 10612
rect 64036 10556 64876 10612
rect 64932 10556 66220 10612
rect 66276 10556 68348 10612
rect 68404 10556 68414 10612
rect 72482 10556 72492 10612
rect 72548 10556 77028 10612
rect 81218 10556 81228 10612
rect 81284 10556 82236 10612
rect 82292 10556 82908 10612
rect 82964 10556 82974 10612
rect 83906 10556 83916 10612
rect 83972 10556 83982 10612
rect 84924 10556 85820 10612
rect 85876 10556 85886 10612
rect 87826 10556 87836 10612
rect 87892 10556 88732 10612
rect 88788 10556 89180 10612
rect 89236 10556 89246 10612
rect 92194 10556 92204 10612
rect 92260 10556 94164 10612
rect 94322 10556 94332 10612
rect 94388 10556 97468 10612
rect 99026 10556 99036 10612
rect 99092 10556 101276 10612
rect 101332 10556 101342 10612
rect 101602 10556 101612 10612
rect 101668 10556 101678 10612
rect 102386 10556 102396 10612
rect 102452 10556 103628 10612
rect 103684 10556 103694 10612
rect 43596 10500 43652 10556
rect 23650 10444 23660 10500
rect 23716 10444 24444 10500
rect 24500 10444 24510 10500
rect 26226 10444 26236 10500
rect 26292 10444 27020 10500
rect 27076 10444 27086 10500
rect 31938 10444 31948 10500
rect 32004 10444 32956 10500
rect 33012 10444 34188 10500
rect 34244 10444 36316 10500
rect 36372 10444 36988 10500
rect 37044 10444 37054 10500
rect 40562 10444 40572 10500
rect 40628 10444 41132 10500
rect 41188 10444 42476 10500
rect 42532 10444 42542 10500
rect 43596 10444 44716 10500
rect 44772 10444 44782 10500
rect 50372 10444 51884 10500
rect 51940 10444 54796 10500
rect 54852 10444 54862 10500
rect 50372 10388 50428 10444
rect 56140 10388 56196 10556
rect 97412 10500 97468 10556
rect 101612 10500 101668 10556
rect 103852 10500 103908 10668
rect 104514 10556 104524 10612
rect 104580 10556 106204 10612
rect 106260 10556 106270 10612
rect 108770 10556 108780 10612
rect 108836 10556 109900 10612
rect 109956 10556 109966 10612
rect 110562 10556 110572 10612
rect 110628 10556 111580 10612
rect 111636 10556 111646 10612
rect 57922 10444 57932 10500
rect 57988 10444 59052 10500
rect 59108 10444 59118 10500
rect 64642 10444 64652 10500
rect 64708 10444 68572 10500
rect 68628 10444 72716 10500
rect 72772 10444 73612 10500
rect 73668 10444 73678 10500
rect 77522 10444 77532 10500
rect 77588 10444 84364 10500
rect 84420 10444 85372 10500
rect 85428 10444 85438 10500
rect 87266 10444 87276 10500
rect 87332 10444 90188 10500
rect 90244 10444 91308 10500
rect 91364 10444 91374 10500
rect 93090 10444 93100 10500
rect 93156 10444 93996 10500
rect 94052 10444 94062 10500
rect 94210 10444 94220 10500
rect 94276 10444 94286 10500
rect 96898 10444 96908 10500
rect 96964 10444 97244 10500
rect 97300 10444 97310 10500
rect 97412 10444 99820 10500
rect 99876 10444 101668 10500
rect 102582 10444 102620 10500
rect 102676 10444 102686 10500
rect 102834 10444 102844 10500
rect 102900 10444 103516 10500
rect 103572 10444 103582 10500
rect 103852 10444 114380 10500
rect 114436 10444 115500 10500
rect 115556 10444 115948 10500
rect 116004 10444 116014 10500
rect 94220 10388 94276 10444
rect 24210 10332 24220 10388
rect 24276 10332 25228 10388
rect 25284 10332 25294 10388
rect 25554 10332 25564 10388
rect 25620 10332 26796 10388
rect 26852 10332 26862 10388
rect 29698 10332 29708 10388
rect 29764 10332 35644 10388
rect 35700 10332 35710 10388
rect 40226 10332 40236 10388
rect 40292 10332 41580 10388
rect 41636 10332 41646 10388
rect 43138 10332 43148 10388
rect 43204 10332 46732 10388
rect 46788 10332 46798 10388
rect 47516 10332 50204 10388
rect 50260 10332 50428 10388
rect 53330 10332 53340 10388
rect 53396 10332 56196 10388
rect 57698 10332 57708 10388
rect 57764 10332 59276 10388
rect 59332 10332 59342 10388
rect 61282 10332 61292 10388
rect 61348 10332 62076 10388
rect 62132 10332 62142 10388
rect 65772 10332 65884 10388
rect 65940 10332 65950 10388
rect 67218 10332 67228 10388
rect 67284 10332 67788 10388
rect 67844 10332 67854 10388
rect 76402 10332 76412 10388
rect 76468 10332 78204 10388
rect 78260 10332 78270 10388
rect 83234 10332 83244 10388
rect 83300 10332 84476 10388
rect 84532 10332 84542 10388
rect 94220 10332 97804 10388
rect 97860 10332 97870 10388
rect 100370 10332 100380 10388
rect 100436 10332 104524 10388
rect 104580 10332 104590 10388
rect 104738 10332 104748 10388
rect 104804 10332 110348 10388
rect 110404 10332 110414 10388
rect 110786 10332 110796 10388
rect 110852 10332 114828 10388
rect 114884 10332 114894 10388
rect 47516 10276 47572 10332
rect 37436 10220 38444 10276
rect 38500 10220 38510 10276
rect 44146 10220 44156 10276
rect 44212 10220 47572 10276
rect 47730 10220 47740 10276
rect 47796 10220 48636 10276
rect 48692 10220 48702 10276
rect 50306 10220 50316 10276
rect 50372 10220 55132 10276
rect 55188 10220 55198 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 37436 10052 37492 10220
rect 42242 10108 42252 10164
rect 42308 10108 43036 10164
rect 43092 10108 43596 10164
rect 43652 10108 43662 10164
rect 43922 10108 43932 10164
rect 43988 10108 44604 10164
rect 44660 10108 44670 10164
rect 47954 10108 47964 10164
rect 48020 10108 48524 10164
rect 48580 10108 48590 10164
rect 48748 10108 50316 10164
rect 50372 10108 50382 10164
rect 53890 10108 53900 10164
rect 53956 10108 58716 10164
rect 58772 10108 58782 10164
rect 48748 10052 48804 10108
rect 65772 10052 65828 10332
rect 86034 10220 86044 10276
rect 86100 10220 88508 10276
rect 88564 10220 88574 10276
rect 93874 10220 93884 10276
rect 93940 10220 93950 10276
rect 98242 10220 98252 10276
rect 98308 10220 103852 10276
rect 103908 10220 103918 10276
rect 112130 10220 112140 10276
rect 112196 10220 115948 10276
rect 116004 10220 116014 10276
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 66994 10108 67004 10164
rect 67060 10108 70028 10164
rect 70084 10108 70094 10164
rect 73126 10108 73164 10164
rect 73220 10108 73230 10164
rect 73602 10108 73612 10164
rect 73668 10108 73948 10164
rect 80994 10108 81004 10164
rect 81060 10108 81452 10164
rect 81508 10108 81900 10164
rect 81956 10108 81966 10164
rect 82422 10108 82460 10164
rect 82516 10108 82526 10164
rect 73892 10052 73948 10108
rect 93884 10052 93940 10220
rect 96626 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96910 10220
rect 127346 10164 127356 10220
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127620 10164 127630 10220
rect 158066 10164 158076 10220
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158340 10164 158350 10220
rect 101126 10108 101164 10164
rect 101220 10108 102844 10164
rect 102900 10108 102910 10164
rect 103058 10108 103068 10164
rect 103124 10108 106092 10164
rect 106148 10108 106158 10164
rect 107986 10108 107996 10164
rect 108052 10108 108332 10164
rect 108388 10108 108398 10164
rect 111794 10108 111804 10164
rect 111860 10108 113148 10164
rect 113204 10108 113214 10164
rect 30482 9996 30492 10052
rect 30548 9996 35980 10052
rect 36036 9996 36046 10052
rect 37090 9996 37100 10052
rect 37156 9996 37492 10052
rect 39442 9996 39452 10052
rect 39508 9996 40796 10052
rect 40852 9996 40862 10052
rect 43810 9996 43820 10052
rect 43876 9996 44492 10052
rect 44548 9996 44716 10052
rect 44772 9996 44782 10052
rect 45490 9996 45500 10052
rect 45556 9996 46732 10052
rect 46788 9996 47628 10052
rect 47684 9996 48804 10052
rect 55010 9996 55020 10052
rect 55076 9996 56700 10052
rect 56756 9996 56766 10052
rect 57922 9996 57932 10052
rect 57988 9996 60396 10052
rect 60452 9996 65828 10052
rect 67788 9996 72436 10052
rect 72930 9996 72940 10052
rect 72996 9996 73006 10052
rect 73892 9996 82348 10052
rect 82404 9996 85484 10052
rect 85540 9996 85550 10052
rect 89618 9996 89628 10052
rect 89684 9996 93940 10052
rect 94546 9996 94556 10052
rect 94612 9996 95116 10052
rect 95172 9996 95182 10052
rect 95554 9996 95564 10052
rect 95620 9996 96460 10052
rect 96516 9996 96526 10052
rect 97010 9996 97020 10052
rect 97076 9996 99148 10052
rect 99204 9996 99214 10052
rect 103282 9996 103292 10052
rect 103348 9996 104188 10052
rect 104244 9996 104254 10052
rect 107090 9996 107100 10052
rect 107156 9996 109116 10052
rect 109172 9996 109182 10052
rect 110226 9996 110236 10052
rect 110292 9996 112028 10052
rect 112084 9996 112094 10052
rect 67788 9940 67844 9996
rect 72380 9940 72436 9996
rect 72940 9940 72996 9996
rect 95116 9940 95172 9996
rect 18834 9884 18844 9940
rect 18900 9884 21532 9940
rect 21588 9884 21598 9940
rect 25106 9884 25116 9940
rect 25172 9884 32284 9940
rect 32340 9884 32350 9940
rect 33394 9884 33404 9940
rect 33460 9884 40460 9940
rect 40516 9884 40526 9940
rect 40898 9884 40908 9940
rect 40964 9884 41356 9940
rect 41412 9884 41692 9940
rect 41748 9884 41758 9940
rect 44818 9884 44828 9940
rect 44884 9884 45164 9940
rect 45220 9884 45230 9940
rect 48962 9884 48972 9940
rect 49028 9884 52444 9940
rect 52500 9884 52510 9940
rect 55794 9884 55804 9940
rect 55860 9884 59388 9940
rect 59444 9884 59454 9940
rect 64530 9884 64540 9940
rect 64596 9884 67788 9940
rect 67844 9884 67854 9940
rect 70578 9884 70588 9940
rect 70644 9884 72324 9940
rect 72380 9884 74844 9940
rect 74900 9884 74910 9940
rect 79426 9884 79436 9940
rect 79492 9884 80668 9940
rect 80724 9884 80734 9940
rect 84550 9884 84588 9940
rect 84644 9884 84654 9940
rect 95116 9884 97468 9940
rect 100706 9884 100716 9940
rect 100772 9884 101836 9940
rect 101892 9884 101902 9940
rect 102834 9884 102844 9940
rect 102900 9884 106540 9940
rect 106596 9884 106606 9940
rect 29362 9772 29372 9828
rect 29428 9772 29932 9828
rect 29988 9772 29998 9828
rect 33506 9772 33516 9828
rect 33572 9772 38332 9828
rect 38388 9772 38398 9828
rect 38546 9772 38556 9828
rect 38612 9772 44156 9828
rect 44212 9772 44222 9828
rect 49186 9772 49196 9828
rect 49252 9772 49756 9828
rect 49812 9772 50540 9828
rect 50596 9772 50606 9828
rect 51436 9772 51884 9828
rect 51940 9772 51950 9828
rect 55682 9772 55692 9828
rect 55748 9772 58156 9828
rect 58212 9772 58222 9828
rect 51436 9716 51492 9772
rect 59388 9716 59444 9884
rect 72268 9828 72324 9884
rect 97412 9828 97468 9884
rect 59938 9772 59948 9828
rect 60004 9772 62524 9828
rect 62580 9772 63084 9828
rect 63140 9772 63420 9828
rect 63476 9772 63486 9828
rect 64754 9772 64764 9828
rect 64820 9772 65324 9828
rect 65380 9772 65390 9828
rect 67442 9772 67452 9828
rect 67508 9772 72212 9828
rect 72268 9772 73724 9828
rect 73780 9772 74956 9828
rect 75012 9772 75022 9828
rect 80322 9772 80332 9828
rect 80388 9772 82460 9828
rect 82516 9772 82526 9828
rect 83570 9772 83580 9828
rect 83636 9772 92652 9828
rect 92708 9772 92718 9828
rect 95218 9772 95228 9828
rect 95284 9772 96236 9828
rect 96292 9772 96302 9828
rect 97412 9772 103068 9828
rect 103124 9772 103134 9828
rect 105858 9772 105868 9828
rect 105924 9772 107996 9828
rect 108052 9772 108062 9828
rect 32946 9660 32956 9716
rect 33012 9660 35308 9716
rect 35364 9660 35374 9716
rect 37510 9660 37548 9716
rect 37604 9660 37614 9716
rect 37762 9660 37772 9716
rect 37828 9660 38668 9716
rect 38724 9660 38734 9716
rect 40002 9660 40012 9716
rect 40068 9660 40908 9716
rect 40964 9660 40974 9716
rect 45490 9660 45500 9716
rect 45556 9660 45948 9716
rect 46004 9660 46014 9716
rect 47506 9660 47516 9716
rect 47572 9660 51492 9716
rect 51650 9660 51660 9716
rect 51716 9660 55244 9716
rect 55300 9660 56028 9716
rect 56084 9660 56094 9716
rect 59388 9660 60844 9716
rect 60900 9660 60910 9716
rect 61058 9660 61068 9716
rect 61124 9660 61162 9716
rect 64194 9660 64204 9716
rect 64260 9660 65212 9716
rect 65268 9660 65278 9716
rect 66658 9660 66668 9716
rect 66724 9660 70140 9716
rect 70196 9660 70206 9716
rect 70466 9660 70476 9716
rect 70532 9660 70924 9716
rect 70980 9660 70990 9716
rect 51660 9604 51716 9660
rect 72156 9604 72212 9772
rect 109172 9716 109228 9940
rect 109284 9884 111468 9940
rect 111524 9884 111534 9940
rect 113698 9884 113708 9940
rect 113764 9884 114156 9940
rect 114212 9884 114222 9940
rect 111234 9772 111244 9828
rect 111300 9772 114492 9828
rect 114548 9772 115612 9828
rect 115668 9772 115678 9828
rect 73238 9660 73276 9716
rect 73332 9660 73342 9716
rect 79986 9660 79996 9716
rect 80052 9660 82908 9716
rect 82964 9660 82974 9716
rect 83906 9660 83916 9716
rect 83972 9660 85932 9716
rect 85988 9660 85998 9716
rect 86594 9660 86604 9716
rect 86660 9660 89068 9716
rect 89124 9660 89134 9716
rect 97234 9660 97244 9716
rect 97300 9660 97580 9716
rect 97636 9660 97646 9716
rect 99026 9660 99036 9716
rect 99092 9660 109228 9716
rect 113922 9660 113932 9716
rect 113988 9660 115948 9716
rect 116004 9660 116014 9716
rect 20738 9548 20748 9604
rect 20804 9548 26124 9604
rect 26180 9548 26190 9604
rect 30594 9548 30604 9604
rect 30660 9548 31052 9604
rect 31108 9548 34076 9604
rect 34132 9548 34142 9604
rect 35186 9548 35196 9604
rect 35252 9548 38556 9604
rect 38612 9548 38622 9604
rect 39330 9548 39340 9604
rect 39396 9548 49756 9604
rect 49812 9548 49822 9604
rect 50306 9548 50316 9604
rect 50372 9548 51716 9604
rect 52322 9548 52332 9604
rect 52388 9548 56140 9604
rect 56196 9548 56206 9604
rect 56354 9548 56364 9604
rect 56420 9548 56812 9604
rect 56868 9548 56878 9604
rect 58258 9548 58268 9604
rect 58324 9548 59052 9604
rect 59108 9548 59118 9604
rect 59714 9548 59724 9604
rect 59780 9548 61180 9604
rect 61236 9548 61246 9604
rect 62850 9548 62860 9604
rect 62916 9548 64316 9604
rect 64372 9548 64382 9604
rect 67106 9548 67116 9604
rect 67172 9548 69132 9604
rect 69188 9548 69198 9604
rect 69458 9548 69468 9604
rect 69524 9548 71260 9604
rect 71316 9548 71326 9604
rect 72146 9548 72156 9604
rect 72212 9548 72222 9604
rect 72706 9548 72716 9604
rect 72772 9548 75068 9604
rect 75124 9548 75134 9604
rect 82562 9548 82572 9604
rect 82628 9548 84812 9604
rect 84868 9548 84878 9604
rect 86482 9548 86492 9604
rect 86548 9548 88732 9604
rect 88788 9548 88798 9604
rect 92642 9548 92652 9604
rect 92708 9548 93436 9604
rect 93492 9548 93502 9604
rect 94098 9548 94108 9604
rect 94164 9548 94556 9604
rect 94612 9548 95228 9604
rect 95284 9548 95294 9604
rect 97346 9548 97356 9604
rect 97412 9548 97916 9604
rect 97972 9548 97982 9604
rect 101490 9548 101500 9604
rect 101556 9548 105308 9604
rect 105364 9548 109676 9604
rect 109732 9548 109742 9604
rect 110114 9548 110124 9604
rect 110180 9548 112476 9604
rect 112532 9548 113372 9604
rect 113428 9548 113438 9604
rect 115490 9548 115500 9604
rect 115556 9548 116396 9604
rect 116452 9548 116462 9604
rect 27906 9436 27916 9492
rect 27972 9436 28476 9492
rect 28532 9436 33068 9492
rect 33124 9436 33134 9492
rect 36418 9436 36428 9492
rect 36484 9436 36988 9492
rect 37044 9436 45836 9492
rect 45892 9436 47292 9492
rect 47348 9436 47358 9492
rect 50978 9436 50988 9492
rect 51044 9436 51054 9492
rect 51958 9436 51996 9492
rect 52052 9436 59836 9492
rect 59892 9436 59902 9492
rect 61964 9436 66444 9492
rect 66500 9436 71148 9492
rect 71204 9436 71708 9492
rect 71764 9436 72492 9492
rect 72548 9436 77868 9492
rect 77924 9436 77934 9492
rect 84130 9436 84140 9492
rect 84196 9436 84476 9492
rect 84532 9436 85708 9492
rect 85764 9436 85774 9492
rect 89170 9436 89180 9492
rect 89236 9436 89852 9492
rect 89908 9436 90860 9492
rect 90916 9436 90926 9492
rect 91522 9436 91532 9492
rect 91588 9436 94332 9492
rect 94388 9436 94398 9492
rect 96002 9436 96012 9492
rect 96068 9436 96684 9492
rect 96740 9436 96750 9492
rect 113138 9436 113148 9492
rect 113204 9436 113820 9492
rect 113876 9436 113886 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 50988 9380 51044 9436
rect 21970 9324 21980 9380
rect 22036 9324 44772 9380
rect 45490 9324 45500 9380
rect 45556 9324 46396 9380
rect 46452 9324 46462 9380
rect 49410 9324 49420 9380
rect 49476 9324 50428 9380
rect 50988 9324 61740 9380
rect 61796 9324 61806 9380
rect 20178 9212 20188 9268
rect 20244 9212 20972 9268
rect 21028 9212 23772 9268
rect 23828 9212 23838 9268
rect 34514 9212 34524 9268
rect 34580 9212 39676 9268
rect 39732 9212 39742 9268
rect 44716 9156 44772 9324
rect 50372 9268 50428 9324
rect 61964 9268 62020 9436
rect 81266 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81550 9436
rect 111986 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112270 9436
rect 142706 9380 142716 9436
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142980 9380 142990 9436
rect 66994 9324 67004 9380
rect 67060 9324 72716 9380
rect 72772 9324 74060 9380
rect 74116 9324 74126 9380
rect 74498 9324 74508 9380
rect 74564 9324 75964 9380
rect 76020 9324 77420 9380
rect 77476 9324 79772 9380
rect 79828 9324 80108 9380
rect 80164 9324 80174 9380
rect 85026 9324 85036 9380
rect 85092 9324 86940 9380
rect 86996 9324 87006 9380
rect 89964 9324 97692 9380
rect 97748 9324 97758 9380
rect 99138 9324 99148 9380
rect 99204 9324 99708 9380
rect 99764 9324 99774 9380
rect 103058 9324 103068 9380
rect 103124 9324 109900 9380
rect 109956 9324 109966 9380
rect 112886 9324 112924 9380
rect 112980 9324 112990 9380
rect 89964 9268 90020 9324
rect 45602 9212 45612 9268
rect 45668 9212 46564 9268
rect 48290 9212 48300 9268
rect 48356 9212 50092 9268
rect 50148 9212 50158 9268
rect 50372 9212 52108 9268
rect 52164 9212 52174 9268
rect 52546 9212 52556 9268
rect 52612 9212 61180 9268
rect 61236 9212 62020 9268
rect 62132 9212 62412 9268
rect 62468 9212 62478 9268
rect 65426 9212 65436 9268
rect 65492 9212 68180 9268
rect 71250 9212 71260 9268
rect 71316 9212 71708 9268
rect 71764 9212 72604 9268
rect 72660 9212 72940 9268
rect 72996 9212 73006 9268
rect 73602 9212 73612 9268
rect 73668 9212 73678 9268
rect 73938 9212 73948 9268
rect 74004 9212 87612 9268
rect 87668 9212 90020 9268
rect 94892 9212 97580 9268
rect 97636 9212 98252 9268
rect 98308 9212 98318 9268
rect 100370 9212 100380 9268
rect 100436 9212 106204 9268
rect 106260 9212 107436 9268
rect 107492 9212 107502 9268
rect 111682 9212 111692 9268
rect 111748 9212 112476 9268
rect 112532 9212 112542 9268
rect 112690 9212 112700 9268
rect 112756 9212 115388 9268
rect 115444 9212 115454 9268
rect 122658 9212 122668 9268
rect 122724 9212 137900 9268
rect 137956 9212 137966 9268
rect 46508 9156 46564 9212
rect 62132 9156 62188 9212
rect 68124 9156 68180 9212
rect 73612 9156 73668 9212
rect 94892 9156 94948 9212
rect 21746 9100 21756 9156
rect 21812 9100 22204 9156
rect 22260 9100 22428 9156
rect 22484 9100 22494 9156
rect 28886 9100 28924 9156
rect 28980 9100 28990 9156
rect 29250 9100 29260 9156
rect 29316 9100 34188 9156
rect 34244 9100 34254 9156
rect 38322 9100 38332 9156
rect 38388 9100 38668 9156
rect 38724 9100 38734 9156
rect 44706 9100 44716 9156
rect 44772 9100 46284 9156
rect 46340 9100 46350 9156
rect 46498 9100 46508 9156
rect 46564 9100 46574 9156
rect 48178 9100 48188 9156
rect 48244 9100 52220 9156
rect 52276 9100 54348 9156
rect 54404 9100 54414 9156
rect 55906 9100 55916 9156
rect 55972 9100 57148 9156
rect 57204 9100 59164 9156
rect 59220 9100 59230 9156
rect 60722 9100 60732 9156
rect 60788 9100 62188 9156
rect 64866 9100 64876 9156
rect 64932 9100 64942 9156
rect 65202 9100 65212 9156
rect 65268 9100 65716 9156
rect 66882 9100 66892 9156
rect 66948 9100 67900 9156
rect 67956 9100 67966 9156
rect 68124 9100 73668 9156
rect 77858 9100 77868 9156
rect 77924 9100 82460 9156
rect 82516 9100 82908 9156
rect 82964 9100 82974 9156
rect 84578 9100 84588 9156
rect 84644 9100 86492 9156
rect 86548 9100 86558 9156
rect 90626 9100 90636 9156
rect 90692 9100 91196 9156
rect 91252 9100 91262 9156
rect 92306 9100 92316 9156
rect 92372 9100 93324 9156
rect 93380 9100 93390 9156
rect 94882 9100 94892 9156
rect 94948 9100 94958 9156
rect 95890 9100 95900 9156
rect 95956 9100 96348 9156
rect 96404 9100 96414 9156
rect 97906 9100 97916 9156
rect 97972 9100 102844 9156
rect 102900 9100 102910 9156
rect 105746 9100 105756 9156
rect 105812 9100 107884 9156
rect 107940 9100 107950 9156
rect 111346 9100 111356 9156
rect 111412 9100 112644 9156
rect 114146 9100 114156 9156
rect 114212 9100 115276 9156
rect 115332 9100 115342 9156
rect 116162 9100 116172 9156
rect 116228 9100 126476 9156
rect 126532 9100 126542 9156
rect 64876 9044 64932 9100
rect 65660 9044 65716 9100
rect 112588 9044 112644 9100
rect 27010 8988 27020 9044
rect 27076 8988 29484 9044
rect 29540 8988 29550 9044
rect 30034 8988 30044 9044
rect 30100 8988 30716 9044
rect 30772 8988 30782 9044
rect 32498 8988 32508 9044
rect 32564 8988 34748 9044
rect 34804 8988 34814 9044
rect 43362 8988 43372 9044
rect 43428 8988 51212 9044
rect 51268 8988 51278 9044
rect 52098 8988 52108 9044
rect 52164 8988 52780 9044
rect 52836 8988 52846 9044
rect 56130 8988 56140 9044
rect 56196 8988 56364 9044
rect 56420 8988 56430 9044
rect 58772 8988 61852 9044
rect 61908 8988 61918 9044
rect 62066 8988 62076 9044
rect 62132 8988 62748 9044
rect 62804 8988 63420 9044
rect 63476 8988 63486 9044
rect 64876 8988 65436 9044
rect 65492 8988 65502 9044
rect 65660 8988 65772 9044
rect 65828 8988 66332 9044
rect 66388 8988 66398 9044
rect 67218 8988 67228 9044
rect 67284 8988 67844 9044
rect 71698 8988 71708 9044
rect 71764 8988 71774 9044
rect 72930 8988 72940 9044
rect 72996 8988 73276 9044
rect 73332 8988 73342 9044
rect 73602 8988 73612 9044
rect 73668 8988 74620 9044
rect 74676 8988 74686 9044
rect 75516 8988 77532 9044
rect 77588 8988 77598 9044
rect 83570 8988 83580 9044
rect 83636 8988 86268 9044
rect 86324 8988 86334 9044
rect 94098 8988 94108 9044
rect 94164 8988 99036 9044
rect 99092 8988 99102 9044
rect 105970 8988 105980 9044
rect 106036 8988 109004 9044
rect 109060 8988 112364 9044
rect 112420 8988 112430 9044
rect 112588 8988 113036 9044
rect 113092 8988 113102 9044
rect 113474 8988 113484 9044
rect 113540 8988 113932 9044
rect 113988 8988 113998 9044
rect 30044 8932 30100 8988
rect 20402 8876 20412 8932
rect 20468 8876 22316 8932
rect 22372 8876 22382 8932
rect 24434 8876 24444 8932
rect 24500 8876 26908 8932
rect 27122 8876 27132 8932
rect 27188 8876 27804 8932
rect 27860 8876 27870 8932
rect 28354 8876 28364 8932
rect 28420 8876 30100 8932
rect 49746 8876 49756 8932
rect 49812 8876 51548 8932
rect 51604 8876 55356 8932
rect 55412 8876 55422 8932
rect 26852 8820 26908 8876
rect 58772 8820 58828 8988
rect 63970 8876 63980 8932
rect 64036 8876 64876 8932
rect 64932 8876 64942 8932
rect 26852 8764 29260 8820
rect 29316 8764 30268 8820
rect 30324 8764 30334 8820
rect 31826 8764 31836 8820
rect 31892 8764 35868 8820
rect 35924 8764 37884 8820
rect 37940 8764 37950 8820
rect 51090 8764 51100 8820
rect 51156 8764 56588 8820
rect 56644 8764 58828 8820
rect 65538 8764 65548 8820
rect 65604 8764 67228 8820
rect 67284 8764 67294 8820
rect 67788 8708 67844 8988
rect 71708 8932 71764 8988
rect 75516 8932 75572 8988
rect 68674 8876 68684 8932
rect 68740 8876 69580 8932
rect 69636 8876 69646 8932
rect 71708 8876 75572 8932
rect 76626 8876 76636 8932
rect 76692 8876 78316 8932
rect 78372 8876 78382 8932
rect 81442 8876 81452 8932
rect 81508 8876 81518 8932
rect 95218 8876 95228 8932
rect 95284 8876 97916 8932
rect 97972 8876 97982 8932
rect 98130 8876 98140 8932
rect 98196 8876 102396 8932
rect 102452 8876 102462 8932
rect 110674 8876 110684 8932
rect 110740 8876 117628 8932
rect 117684 8876 117694 8932
rect 71596 8764 77084 8820
rect 77140 8764 77150 8820
rect 71596 8708 71652 8764
rect 81452 8708 81508 8876
rect 83122 8764 83132 8820
rect 83188 8764 91196 8820
rect 91252 8764 92092 8820
rect 92148 8764 92158 8820
rect 92866 8764 92876 8820
rect 92932 8764 94556 8820
rect 94612 8764 94622 8820
rect 95890 8764 95900 8820
rect 95956 8764 95966 8820
rect 96562 8764 96572 8820
rect 96628 8764 97468 8820
rect 98466 8764 98476 8820
rect 98532 8764 100828 8820
rect 100884 8764 100894 8820
rect 102834 8764 102844 8820
rect 102900 8764 105196 8820
rect 105252 8764 106428 8820
rect 106484 8764 106494 8820
rect 109890 8764 109900 8820
rect 109956 8764 116284 8820
rect 116340 8764 117180 8820
rect 117236 8764 117246 8820
rect 26002 8652 26012 8708
rect 26068 8652 29036 8708
rect 29092 8652 34468 8708
rect 39554 8652 39564 8708
rect 39620 8652 41356 8708
rect 41412 8652 41422 8708
rect 51314 8652 51324 8708
rect 51380 8652 51548 8708
rect 51604 8652 51884 8708
rect 51940 8652 62188 8708
rect 67788 8652 71652 8708
rect 72818 8652 72828 8708
rect 72884 8652 73612 8708
rect 73668 8652 81508 8708
rect 82292 8652 89292 8708
rect 89348 8652 92764 8708
rect 92820 8652 92830 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 25218 8540 25228 8596
rect 25284 8540 30884 8596
rect 30828 8484 30884 8540
rect 34412 8484 34468 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 62132 8596 62188 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 82292 8596 82348 8652
rect 38210 8540 38220 8596
rect 38276 8540 39004 8596
rect 39060 8540 39788 8596
rect 39844 8540 39854 8596
rect 55682 8540 55692 8596
rect 55748 8540 56812 8596
rect 56868 8540 56878 8596
rect 62132 8540 62300 8596
rect 62356 8540 62636 8596
rect 62692 8540 62702 8596
rect 67442 8540 67452 8596
rect 67508 8540 68460 8596
rect 68516 8540 68526 8596
rect 72258 8540 72268 8596
rect 72324 8540 73052 8596
rect 73108 8540 73118 8596
rect 78194 8540 78204 8596
rect 78260 8540 82348 8596
rect 83122 8540 83132 8596
rect 83188 8540 84084 8596
rect 84690 8540 84700 8596
rect 84756 8540 95116 8596
rect 95172 8540 95182 8596
rect 20178 8428 20188 8484
rect 20244 8428 21476 8484
rect 27794 8428 27804 8484
rect 27860 8428 30268 8484
rect 30324 8428 30334 8484
rect 30818 8428 30828 8484
rect 30884 8428 31612 8484
rect 31668 8428 31678 8484
rect 34412 8428 36988 8484
rect 37044 8428 37054 8484
rect 39106 8428 39116 8484
rect 39172 8428 40348 8484
rect 40404 8428 40414 8484
rect 45602 8428 45612 8484
rect 45668 8428 48412 8484
rect 48468 8428 48478 8484
rect 52294 8428 52332 8484
rect 52388 8428 52398 8484
rect 55234 8428 55244 8484
rect 55300 8428 55580 8484
rect 55636 8428 55646 8484
rect 55990 8428 56028 8484
rect 56084 8428 56094 8484
rect 56662 8428 56700 8484
rect 56756 8428 56766 8484
rect 56914 8428 56924 8484
rect 56980 8428 57596 8484
rect 57652 8428 57662 8484
rect 63970 8428 63980 8484
rect 64036 8428 64540 8484
rect 64596 8428 64606 8484
rect 69010 8428 69020 8484
rect 69076 8428 71932 8484
rect 71988 8428 74508 8484
rect 74564 8428 74574 8484
rect 79426 8428 79436 8484
rect 79492 8428 83804 8484
rect 83860 8428 83870 8484
rect 21420 8260 21476 8428
rect 84028 8372 84084 8540
rect 95900 8484 95956 8764
rect 96626 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96910 8652
rect 97412 8596 97468 8764
rect 98690 8652 98700 8708
rect 98756 8652 102508 8708
rect 102564 8652 102574 8708
rect 110562 8652 110572 8708
rect 110628 8652 112476 8708
rect 112532 8652 112542 8708
rect 127346 8596 127356 8652
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127620 8596 127630 8652
rect 158066 8596 158076 8652
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158340 8596 158350 8652
rect 97412 8540 104636 8596
rect 104692 8540 105644 8596
rect 105700 8540 105710 8596
rect 108770 8540 108780 8596
rect 108836 8540 110684 8596
rect 110740 8540 110750 8596
rect 110898 8540 110908 8596
rect 110964 8540 111356 8596
rect 111412 8540 111422 8596
rect 85446 8428 85484 8484
rect 85540 8428 85550 8484
rect 85698 8428 85708 8484
rect 85764 8428 86156 8484
rect 86212 8428 86222 8484
rect 86790 8428 86828 8484
rect 86884 8428 86894 8484
rect 90738 8428 90748 8484
rect 90804 8428 92876 8484
rect 92932 8428 92942 8484
rect 95638 8428 95676 8484
rect 95732 8428 95742 8484
rect 95900 8428 97468 8484
rect 97524 8428 97534 8484
rect 107426 8428 107436 8484
rect 107492 8428 107884 8484
rect 107940 8428 107950 8484
rect 109666 8428 109676 8484
rect 109732 8428 111132 8484
rect 111188 8428 111198 8484
rect 112354 8428 112364 8484
rect 112420 8428 115500 8484
rect 115556 8428 115566 8484
rect 21746 8316 21756 8372
rect 21812 8316 22540 8372
rect 22596 8316 28028 8372
rect 28084 8316 28094 8372
rect 28242 8316 28252 8372
rect 28308 8316 29484 8372
rect 29540 8316 29550 8372
rect 30482 8316 30492 8372
rect 30548 8316 32172 8372
rect 32228 8316 37100 8372
rect 37156 8316 37166 8372
rect 37650 8316 37660 8372
rect 37716 8316 39228 8372
rect 39284 8316 39294 8372
rect 43026 8316 43036 8372
rect 43092 8316 43820 8372
rect 43876 8316 45276 8372
rect 45332 8316 47068 8372
rect 47124 8316 48860 8372
rect 48916 8316 48926 8372
rect 49746 8316 49756 8372
rect 49812 8316 51548 8372
rect 51604 8316 51614 8372
rect 52444 8316 53228 8372
rect 53284 8316 53294 8372
rect 61730 8316 61740 8372
rect 61796 8316 63252 8372
rect 63410 8316 63420 8372
rect 63476 8316 65324 8372
rect 65380 8316 65390 8372
rect 67442 8316 67452 8372
rect 67508 8316 73164 8372
rect 73220 8316 73230 8372
rect 73490 8316 73500 8372
rect 73556 8316 75740 8372
rect 75796 8316 75806 8372
rect 77522 8316 77532 8372
rect 77588 8316 78540 8372
rect 78596 8316 79212 8372
rect 79268 8316 82236 8372
rect 82292 8316 82302 8372
rect 84018 8316 84028 8372
rect 84084 8316 84094 8372
rect 84466 8316 84476 8372
rect 84532 8316 85260 8372
rect 85316 8316 85326 8372
rect 86258 8316 86268 8372
rect 86324 8316 86716 8372
rect 86772 8316 86782 8372
rect 86930 8316 86940 8372
rect 86996 8316 87388 8372
rect 87444 8316 87454 8372
rect 91410 8316 91420 8372
rect 91476 8316 92988 8372
rect 93044 8316 94108 8372
rect 94164 8316 94174 8372
rect 96114 8316 96124 8372
rect 96180 8316 97916 8372
rect 97972 8316 97982 8372
rect 98354 8316 98364 8372
rect 98420 8316 100268 8372
rect 100324 8316 100334 8372
rect 100706 8316 100716 8372
rect 100772 8316 101948 8372
rect 102004 8316 102014 8372
rect 103954 8316 103964 8372
rect 104020 8316 105196 8372
rect 105252 8316 105262 8372
rect 106194 8316 106204 8372
rect 106260 8316 107660 8372
rect 107716 8316 107726 8372
rect 108518 8316 108556 8372
rect 108612 8316 108622 8372
rect 112914 8316 112924 8372
rect 112980 8316 113484 8372
rect 113540 8316 113550 8372
rect 114594 8316 114604 8372
rect 114660 8316 117516 8372
rect 117572 8316 117582 8372
rect 121762 8316 121772 8372
rect 121828 8316 128828 8372
rect 128884 8316 128894 8372
rect 28252 8260 28308 8316
rect 52444 8260 52500 8316
rect 63196 8260 63252 8316
rect 21410 8204 21420 8260
rect 21476 8204 21486 8260
rect 23426 8204 23436 8260
rect 23492 8204 23884 8260
rect 23940 8204 23950 8260
rect 25778 8204 25788 8260
rect 25844 8204 28308 8260
rect 29922 8204 29932 8260
rect 29988 8204 30716 8260
rect 30772 8204 30782 8260
rect 31388 8204 32620 8260
rect 32676 8204 33404 8260
rect 33460 8204 33470 8260
rect 35634 8204 35644 8260
rect 35700 8204 41356 8260
rect 41412 8204 42028 8260
rect 42084 8204 42094 8260
rect 44370 8204 44380 8260
rect 44436 8204 45052 8260
rect 45108 8204 45118 8260
rect 45714 8204 45724 8260
rect 45780 8204 46060 8260
rect 46116 8204 46126 8260
rect 49410 8204 49420 8260
rect 49476 8204 50540 8260
rect 50596 8204 52500 8260
rect 52770 8204 52780 8260
rect 52836 8204 61852 8260
rect 61908 8204 61918 8260
rect 63196 8204 64764 8260
rect 64820 8204 64830 8260
rect 64978 8204 64988 8260
rect 65044 8204 66668 8260
rect 66724 8204 66734 8260
rect 68226 8204 68236 8260
rect 68292 8204 72492 8260
rect 72548 8204 72558 8260
rect 72930 8204 72940 8260
rect 72996 8204 75404 8260
rect 75460 8204 75470 8260
rect 80994 8204 81004 8260
rect 81060 8204 85932 8260
rect 85988 8204 88620 8260
rect 88676 8204 88686 8260
rect 90514 8204 90524 8260
rect 90580 8204 92428 8260
rect 92484 8204 92494 8260
rect 93650 8204 93660 8260
rect 93716 8204 93996 8260
rect 94052 8204 94062 8260
rect 95666 8204 95676 8260
rect 95732 8204 96628 8260
rect 99138 8204 99148 8260
rect 99204 8204 101724 8260
rect 101780 8204 102956 8260
rect 103012 8204 103022 8260
rect 104850 8204 104860 8260
rect 104916 8204 110684 8260
rect 110740 8204 110750 8260
rect 111346 8204 111356 8260
rect 111412 8204 112140 8260
rect 112196 8204 112206 8260
rect 114258 8204 114268 8260
rect 114324 8204 115276 8260
rect 115332 8204 116732 8260
rect 116788 8204 118300 8260
rect 118356 8204 118748 8260
rect 118804 8204 118814 8260
rect 31388 8148 31444 8204
rect 96572 8148 96628 8204
rect 18050 8092 18060 8148
rect 18116 8092 20412 8148
rect 20468 8092 20478 8148
rect 28690 8092 28700 8148
rect 28756 8092 31444 8148
rect 32722 8092 32732 8148
rect 32788 8092 33516 8148
rect 33572 8092 33852 8148
rect 33908 8092 33918 8148
rect 34626 8092 34636 8148
rect 34692 8092 37212 8148
rect 37268 8092 39900 8148
rect 39956 8092 43708 8148
rect 43764 8092 43774 8148
rect 49522 8092 49532 8148
rect 49588 8092 53004 8148
rect 53060 8092 53070 8148
rect 53218 8092 53228 8148
rect 53284 8092 54684 8148
rect 54740 8092 54750 8148
rect 56018 8092 56028 8148
rect 56084 8092 59500 8148
rect 59556 8092 59566 8148
rect 62132 8092 68908 8148
rect 68964 8092 68974 8148
rect 69234 8092 69244 8148
rect 69300 8092 70364 8148
rect 70420 8092 70430 8148
rect 76962 8092 76972 8148
rect 77028 8092 81116 8148
rect 81172 8092 81452 8148
rect 81508 8092 81518 8148
rect 85026 8092 85036 8148
rect 85092 8092 86492 8148
rect 86548 8092 86558 8148
rect 88386 8092 88396 8148
rect 88452 8092 94668 8148
rect 94724 8092 94734 8148
rect 96572 8092 98364 8148
rect 98420 8092 98430 8148
rect 100370 8092 100380 8148
rect 100436 8092 111356 8148
rect 111412 8092 115612 8148
rect 115668 8092 115678 8148
rect 21522 7980 21532 8036
rect 21588 7980 22764 8036
rect 22820 7980 24668 8036
rect 24724 7980 24734 8036
rect 26562 7980 26572 8036
rect 26628 7980 28364 8036
rect 28420 7980 28430 8036
rect 42802 7980 42812 8036
rect 42868 7980 45276 8036
rect 45332 7980 45342 8036
rect 46946 7980 46956 8036
rect 47012 7980 48300 8036
rect 48356 7980 49756 8036
rect 49812 7980 49822 8036
rect 53106 7980 53116 8036
rect 53172 7980 54460 8036
rect 54516 7980 54526 8036
rect 21634 7868 21644 7924
rect 21700 7868 24332 7924
rect 24388 7868 30100 7924
rect 32162 7868 32172 7924
rect 32228 7868 39564 7924
rect 39620 7868 39630 7924
rect 51986 7868 51996 7924
rect 52052 7868 57036 7924
rect 57092 7868 57102 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 30044 7812 30100 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 62132 7812 62188 8092
rect 67442 7980 67452 8036
rect 67508 7980 71036 8036
rect 71092 7980 71102 8036
rect 75394 7980 75404 8036
rect 75460 7980 78092 8036
rect 78148 7980 78158 8036
rect 84354 7980 84364 8036
rect 84420 7980 85148 8036
rect 85204 7980 85214 8036
rect 85474 7980 85484 8036
rect 85540 7980 86044 8036
rect 86100 7980 86110 8036
rect 86594 7980 86604 8036
rect 86660 7980 87164 8036
rect 87220 7980 87230 8036
rect 90178 7980 90188 8036
rect 90244 7980 93100 8036
rect 93156 7980 93166 8036
rect 94770 7980 94780 8036
rect 94836 7980 94846 8036
rect 95778 7980 95788 8036
rect 95844 7980 100156 8036
rect 100212 7980 100222 8036
rect 100594 7980 100604 8036
rect 100660 7980 101612 8036
rect 101668 7980 101678 8036
rect 104290 7980 104300 8036
rect 104356 7980 106988 8036
rect 107044 7980 107054 8036
rect 107650 7980 107660 8036
rect 107716 7980 107726 8036
rect 107874 7980 107884 8036
rect 107940 7980 108892 8036
rect 108948 7980 108958 8036
rect 111010 7980 111020 8036
rect 111076 7980 113540 8036
rect 113810 7980 113820 8036
rect 113876 7980 114828 8036
rect 114884 7980 114894 8036
rect 117282 7980 117292 8036
rect 117348 7980 120988 8036
rect 94780 7924 94836 7980
rect 107660 7924 107716 7980
rect 113484 7924 113540 7980
rect 64754 7868 64764 7924
rect 64820 7868 65660 7924
rect 65716 7868 65726 7924
rect 66434 7868 66444 7924
rect 66500 7868 67228 7924
rect 67284 7868 67294 7924
rect 82674 7868 82684 7924
rect 82740 7868 86828 7924
rect 86884 7868 86894 7924
rect 87378 7868 87388 7924
rect 87444 7868 87454 7924
rect 89842 7868 89852 7924
rect 89908 7868 93212 7924
rect 93268 7868 94836 7924
rect 95666 7868 95676 7924
rect 95732 7868 107716 7924
rect 110870 7868 110908 7924
rect 110964 7868 110974 7924
rect 113484 7868 114604 7924
rect 114660 7868 114670 7924
rect 81266 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81550 7868
rect 87388 7812 87444 7868
rect 111986 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112270 7868
rect 120932 7812 120988 7980
rect 142706 7812 142716 7868
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142980 7812 142990 7868
rect 15922 7756 15932 7812
rect 15988 7756 16940 7812
rect 16996 7756 17006 7812
rect 25554 7756 25564 7812
rect 25620 7756 26236 7812
rect 26292 7756 28700 7812
rect 28756 7756 28766 7812
rect 30034 7756 30044 7812
rect 30100 7756 31388 7812
rect 31444 7756 31454 7812
rect 34066 7756 34076 7812
rect 34132 7756 50316 7812
rect 50372 7756 50382 7812
rect 51996 7756 62188 7812
rect 62514 7756 62524 7812
rect 62580 7756 63532 7812
rect 63588 7756 63598 7812
rect 86482 7756 86492 7812
rect 86548 7756 87444 7812
rect 94546 7756 94556 7812
rect 94612 7756 97020 7812
rect 97076 7756 97086 7812
rect 97906 7756 97916 7812
rect 97972 7756 108444 7812
rect 108500 7756 108510 7812
rect 114034 7756 114044 7812
rect 114100 7756 120148 7812
rect 120932 7756 121324 7812
rect 121380 7756 121390 7812
rect 24546 7644 24556 7700
rect 24612 7644 25788 7700
rect 25844 7644 28812 7700
rect 28868 7644 28878 7700
rect 40226 7644 40236 7700
rect 40292 7644 41132 7700
rect 41188 7644 41198 7700
rect 44930 7644 44940 7700
rect 44996 7644 46732 7700
rect 46788 7644 50652 7700
rect 50708 7644 50718 7700
rect 51996 7588 52052 7756
rect 52182 7644 52220 7700
rect 52276 7644 52286 7700
rect 55990 7644 56028 7700
rect 56084 7644 56094 7700
rect 56466 7644 56476 7700
rect 56532 7644 57092 7700
rect 57250 7644 57260 7700
rect 57316 7644 58716 7700
rect 58772 7644 58782 7700
rect 59826 7644 59836 7700
rect 59892 7644 62188 7700
rect 62850 7644 62860 7700
rect 62916 7644 64428 7700
rect 64484 7644 64494 7700
rect 67106 7644 67116 7700
rect 67172 7644 67788 7700
rect 67844 7644 67854 7700
rect 72146 7644 72156 7700
rect 72212 7644 75964 7700
rect 76020 7644 84476 7700
rect 84532 7644 85260 7700
rect 85316 7644 85326 7700
rect 86706 7644 86716 7700
rect 86772 7644 95788 7700
rect 95844 7644 95854 7700
rect 100258 7644 100268 7700
rect 100324 7644 101388 7700
rect 101444 7644 101454 7700
rect 101724 7644 103068 7700
rect 103124 7644 103964 7700
rect 104020 7644 104030 7700
rect 57036 7588 57092 7644
rect 62132 7588 62188 7644
rect 101724 7588 101780 7644
rect 114044 7588 114100 7756
rect 120092 7700 120148 7756
rect 118738 7644 118748 7700
rect 118804 7644 119868 7700
rect 119924 7644 119934 7700
rect 120092 7644 120988 7700
rect 120932 7588 120988 7644
rect 125972 7644 141036 7700
rect 141092 7644 141102 7700
rect 125972 7588 126028 7644
rect 24658 7532 24668 7588
rect 24724 7532 25900 7588
rect 25956 7532 25966 7588
rect 26852 7532 27244 7588
rect 27300 7532 27310 7588
rect 31042 7532 31052 7588
rect 31108 7532 32284 7588
rect 32340 7532 32350 7588
rect 43698 7532 43708 7588
rect 43764 7532 48188 7588
rect 48244 7532 48254 7588
rect 49084 7532 52052 7588
rect 53890 7532 53900 7588
rect 53956 7532 56588 7588
rect 56644 7532 56654 7588
rect 57036 7532 60284 7588
rect 60340 7532 61292 7588
rect 61348 7532 61358 7588
rect 61926 7532 61964 7588
rect 62020 7532 62030 7588
rect 62132 7532 64316 7588
rect 64372 7532 64382 7588
rect 65212 7532 66668 7588
rect 66724 7532 66734 7588
rect 72258 7532 72268 7588
rect 72324 7532 74060 7588
rect 74116 7532 74126 7588
rect 77298 7532 77308 7588
rect 77364 7532 77980 7588
rect 78036 7532 78046 7588
rect 78978 7532 78988 7588
rect 79044 7532 79772 7588
rect 79828 7532 90076 7588
rect 90132 7532 90142 7588
rect 92082 7532 92092 7588
rect 92148 7532 93996 7588
rect 94052 7532 94062 7588
rect 94546 7532 94556 7588
rect 94612 7532 95452 7588
rect 95508 7532 97468 7588
rect 100146 7532 100156 7588
rect 100212 7532 101052 7588
rect 101108 7532 101780 7588
rect 105074 7532 105084 7588
rect 105140 7532 114100 7588
rect 115714 7532 115724 7588
rect 115780 7532 116396 7588
rect 116452 7532 120316 7588
rect 120372 7532 120382 7588
rect 120932 7532 126028 7588
rect 26852 7476 26908 7532
rect 49084 7476 49140 7532
rect 22306 7420 22316 7476
rect 22372 7420 23212 7476
rect 23268 7420 23278 7476
rect 24556 7420 25676 7476
rect 25732 7420 26908 7476
rect 28466 7420 28476 7476
rect 28532 7420 29148 7476
rect 29204 7420 29214 7476
rect 32610 7420 32620 7476
rect 32676 7420 39900 7476
rect 39956 7420 41356 7476
rect 41412 7420 41422 7476
rect 41570 7420 41580 7476
rect 41636 7420 43932 7476
rect 43988 7420 49140 7476
rect 49298 7420 49308 7476
rect 49364 7420 49756 7476
rect 49812 7420 52556 7476
rect 52612 7420 52622 7476
rect 54002 7420 54012 7476
rect 54068 7420 54078 7476
rect 55682 7420 55692 7476
rect 55748 7420 64652 7476
rect 64708 7420 64718 7476
rect 24556 7364 24612 7420
rect 20514 7308 20524 7364
rect 20580 7308 22876 7364
rect 22932 7308 22942 7364
rect 24546 7308 24556 7364
rect 24612 7308 24622 7364
rect 47618 7308 47628 7364
rect 47684 7308 48188 7364
rect 48244 7308 49868 7364
rect 49924 7308 49934 7364
rect 51874 7308 51884 7364
rect 51940 7308 52332 7364
rect 52388 7308 52398 7364
rect 52994 7308 53004 7364
rect 53060 7308 53452 7364
rect 53508 7308 53518 7364
rect 54012 7252 54068 7420
rect 54674 7308 54684 7364
rect 54740 7308 56140 7364
rect 56196 7308 56206 7364
rect 60834 7308 60844 7364
rect 60900 7308 61068 7364
rect 61124 7308 63308 7364
rect 63364 7308 63374 7364
rect 65212 7252 65268 7532
rect 65426 7420 65436 7476
rect 65492 7420 67116 7476
rect 67172 7420 67182 7476
rect 71250 7420 71260 7476
rect 71316 7420 72212 7476
rect 72370 7420 72380 7476
rect 72436 7420 72828 7476
rect 72884 7420 73948 7476
rect 74004 7420 82124 7476
rect 82180 7420 82684 7476
rect 82740 7420 82750 7476
rect 86706 7420 86716 7476
rect 86772 7420 89964 7476
rect 90020 7420 90030 7476
rect 92194 7420 92204 7476
rect 92260 7420 95004 7476
rect 95060 7420 95070 7476
rect 72156 7364 72212 7420
rect 66210 7308 66220 7364
rect 66276 7308 66286 7364
rect 70466 7308 70476 7364
rect 70532 7308 71148 7364
rect 71204 7308 71214 7364
rect 72156 7308 73444 7364
rect 75506 7308 75516 7364
rect 75572 7308 76748 7364
rect 76804 7308 77196 7364
rect 77252 7308 77262 7364
rect 80658 7308 80668 7364
rect 80724 7308 85820 7364
rect 85876 7308 86156 7364
rect 86212 7308 86222 7364
rect 86818 7308 86828 7364
rect 86884 7308 87948 7364
rect 88004 7308 88014 7364
rect 89506 7308 89516 7364
rect 89572 7308 90860 7364
rect 90916 7308 94892 7364
rect 94948 7308 94958 7364
rect 21298 7196 21308 7252
rect 21364 7196 24780 7252
rect 24836 7196 25452 7252
rect 25508 7196 31220 7252
rect 31378 7196 31388 7252
rect 31444 7196 39228 7252
rect 39284 7196 39294 7252
rect 40002 7196 40012 7252
rect 40068 7196 41020 7252
rect 41076 7196 41086 7252
rect 47170 7196 47180 7252
rect 47236 7196 54068 7252
rect 60844 7196 65268 7252
rect 66220 7252 66276 7308
rect 66220 7196 66500 7252
rect 66658 7196 66668 7252
rect 66724 7196 72044 7252
rect 72100 7196 72604 7252
rect 72660 7196 72670 7252
rect 31164 7140 31220 7196
rect 60844 7140 60900 7196
rect 22530 7084 22540 7140
rect 22596 7084 29484 7140
rect 29540 7084 31108 7140
rect 31164 7084 34076 7140
rect 34132 7084 34142 7140
rect 38994 7084 39004 7140
rect 39060 7084 39340 7140
rect 39396 7084 39406 7140
rect 45826 7084 45836 7140
rect 45892 7084 47292 7140
rect 47348 7084 47358 7140
rect 52322 7084 52332 7140
rect 52388 7084 55468 7140
rect 55524 7084 55534 7140
rect 56802 7084 56812 7140
rect 56868 7084 60508 7140
rect 60564 7084 60574 7140
rect 60834 7084 60844 7140
rect 60900 7084 60910 7140
rect 61506 7084 61516 7140
rect 61572 7084 61852 7140
rect 61908 7084 61918 7140
rect 62132 7084 63420 7140
rect 63476 7084 63486 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 31052 7028 31108 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 62132 7028 62188 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 66444 7028 66500 7196
rect 73388 7140 73444 7308
rect 97412 7252 97468 7532
rect 101490 7420 101500 7476
rect 101556 7420 102508 7476
rect 102564 7420 102574 7476
rect 102946 7420 102956 7476
rect 103012 7420 105532 7476
rect 105588 7420 105598 7476
rect 109554 7420 109564 7476
rect 109620 7420 110572 7476
rect 110628 7420 110638 7476
rect 114706 7420 114716 7476
rect 114772 7420 122668 7476
rect 122724 7420 122734 7476
rect 110226 7308 110236 7364
rect 110292 7308 115612 7364
rect 115668 7308 115678 7364
rect 117394 7308 117404 7364
rect 117460 7308 117740 7364
rect 117796 7308 117806 7364
rect 118178 7308 118188 7364
rect 118244 7308 118254 7364
rect 118188 7252 118244 7308
rect 73602 7196 73612 7252
rect 73668 7196 76300 7252
rect 76356 7196 76366 7252
rect 77308 7196 84476 7252
rect 84532 7196 84542 7252
rect 86706 7196 86716 7252
rect 86772 7196 86828 7252
rect 86884 7196 86894 7252
rect 87042 7196 87052 7252
rect 87108 7196 87724 7252
rect 87780 7196 87790 7252
rect 94210 7196 94220 7252
rect 94276 7196 96572 7252
rect 96628 7196 96638 7252
rect 97412 7196 118244 7252
rect 77308 7140 77364 7196
rect 72818 7084 72828 7140
rect 72884 7084 73164 7140
rect 73220 7084 73230 7140
rect 73388 7084 77364 7140
rect 79398 7084 79436 7140
rect 79492 7084 79502 7140
rect 82562 7084 82572 7140
rect 82628 7084 83916 7140
rect 83972 7084 83982 7140
rect 86146 7084 86156 7140
rect 86212 7084 86492 7140
rect 86548 7084 86558 7140
rect 108434 7084 108444 7140
rect 108500 7084 109004 7140
rect 109060 7084 109070 7140
rect 115014 7084 115052 7140
rect 115108 7084 115118 7140
rect 96626 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96910 7084
rect 127346 7028 127356 7084
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127620 7028 127630 7084
rect 158066 7028 158076 7084
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158340 7028 158350 7084
rect 17378 6972 17388 7028
rect 17444 6972 18508 7028
rect 18564 6972 20076 7028
rect 20132 6972 22764 7028
rect 22820 6972 23436 7028
rect 23492 6972 24332 7028
rect 24388 6972 24398 7028
rect 28802 6972 28812 7028
rect 28868 6972 29260 7028
rect 29316 6972 29326 7028
rect 29586 6972 29596 7028
rect 29652 6972 30492 7028
rect 30548 6972 30558 7028
rect 31052 6972 33852 7028
rect 33908 6972 33918 7028
rect 39554 6972 39564 7028
rect 39620 6972 41020 7028
rect 41076 6972 41086 7028
rect 44930 6972 44940 7028
rect 44996 6972 46284 7028
rect 46340 6972 46350 7028
rect 56690 6972 56700 7028
rect 56756 6972 57036 7028
rect 57092 6972 57102 7028
rect 57260 6972 62188 7028
rect 66444 6972 81004 7028
rect 81060 6972 90524 7028
rect 90580 6972 90590 7028
rect 102498 6972 102508 7028
rect 102564 6972 104860 7028
rect 104916 6972 104926 7028
rect 106194 6972 106204 7028
rect 106260 6972 112028 7028
rect 112084 6972 117964 7028
rect 118020 6972 118030 7028
rect 57260 6916 57316 6972
rect 28578 6860 28588 6916
rect 28644 6860 29484 6916
rect 29540 6860 30156 6916
rect 30212 6860 30604 6916
rect 30660 6860 31724 6916
rect 31780 6860 31790 6916
rect 38994 6860 39004 6916
rect 39060 6860 39340 6916
rect 39396 6860 40572 6916
rect 40628 6860 40638 6916
rect 48850 6860 48860 6916
rect 48916 6860 50092 6916
rect 50148 6860 50158 6916
rect 51538 6860 51548 6916
rect 51604 6860 57316 6916
rect 61058 6860 61068 6916
rect 61124 6860 64204 6916
rect 64260 6860 64270 6916
rect 65426 6860 65436 6916
rect 65492 6860 65502 6916
rect 69906 6860 69916 6916
rect 69972 6860 70588 6916
rect 70644 6860 70654 6916
rect 71138 6860 71148 6916
rect 71204 6860 76076 6916
rect 76132 6860 76142 6916
rect 77298 6860 77308 6916
rect 77364 6860 83300 6916
rect 83458 6860 83468 6916
rect 83524 6860 84476 6916
rect 84532 6860 84542 6916
rect 85698 6860 85708 6916
rect 85764 6860 92484 6916
rect 93202 6860 93212 6916
rect 93268 6860 99708 6916
rect 99764 6860 99774 6916
rect 105746 6860 105756 6916
rect 105812 6860 105822 6916
rect 106530 6860 106540 6916
rect 106596 6860 116284 6916
rect 116340 6860 116350 6916
rect 22642 6748 22652 6804
rect 22708 6748 26236 6804
rect 26292 6748 26302 6804
rect 29250 6748 29260 6804
rect 29316 6748 30828 6804
rect 30884 6748 30894 6804
rect 34626 6748 34636 6804
rect 34692 6748 34702 6804
rect 36418 6748 36428 6804
rect 36484 6748 37660 6804
rect 37716 6748 37726 6804
rect 39666 6748 39676 6804
rect 39732 6748 39844 6804
rect 44370 6748 44380 6804
rect 44436 6748 45052 6804
rect 45108 6748 45118 6804
rect 47842 6748 47852 6804
rect 47908 6748 48636 6804
rect 48692 6748 48702 6804
rect 50978 6748 50988 6804
rect 51044 6748 51054 6804
rect 52098 6748 52108 6804
rect 52164 6748 52892 6804
rect 52948 6748 53340 6804
rect 53396 6748 53406 6804
rect 57698 6748 57708 6804
rect 57764 6748 58380 6804
rect 58436 6748 61740 6804
rect 61796 6748 63196 6804
rect 63252 6748 63262 6804
rect 34636 6692 34692 6748
rect 39788 6692 39844 6748
rect 50988 6692 51044 6748
rect 57708 6692 57764 6748
rect 65436 6692 65492 6860
rect 71148 6804 71204 6860
rect 83244 6804 83300 6860
rect 67666 6748 67676 6804
rect 67732 6748 71204 6804
rect 72482 6748 72492 6804
rect 72548 6748 73388 6804
rect 73444 6748 73454 6804
rect 81106 6748 81116 6804
rect 81172 6748 82348 6804
rect 82404 6748 82414 6804
rect 83244 6748 84364 6804
rect 84420 6748 84430 6804
rect 85362 6748 85372 6804
rect 85428 6748 85484 6804
rect 85540 6748 85550 6804
rect 87714 6748 87724 6804
rect 87780 6748 88172 6804
rect 88228 6748 92204 6804
rect 92260 6748 92270 6804
rect 82348 6692 82404 6748
rect 18610 6636 18620 6692
rect 18676 6636 22540 6692
rect 22596 6636 22606 6692
rect 24780 6636 28140 6692
rect 28196 6636 30492 6692
rect 30548 6636 34692 6692
rect 37538 6636 37548 6692
rect 37604 6636 38556 6692
rect 38612 6636 39564 6692
rect 39620 6636 39630 6692
rect 39788 6636 41132 6692
rect 41188 6636 41198 6692
rect 41542 6636 41580 6692
rect 41636 6636 41646 6692
rect 41794 6636 41804 6692
rect 41860 6636 43708 6692
rect 43764 6636 43774 6692
rect 45938 6636 45948 6692
rect 46004 6636 46060 6692
rect 46116 6636 46126 6692
rect 46386 6636 46396 6692
rect 46452 6636 47292 6692
rect 47348 6636 47358 6692
rect 49186 6636 49196 6692
rect 49252 6636 52668 6692
rect 52724 6636 52734 6692
rect 54338 6636 54348 6692
rect 54404 6636 57764 6692
rect 60722 6636 60732 6692
rect 60788 6636 65492 6692
rect 67554 6636 67564 6692
rect 67620 6636 68236 6692
rect 68292 6636 71708 6692
rect 71764 6636 71774 6692
rect 73154 6636 73164 6692
rect 73220 6636 76412 6692
rect 76468 6636 77196 6692
rect 77252 6636 77262 6692
rect 77420 6636 81396 6692
rect 82348 6636 85260 6692
rect 85316 6636 85326 6692
rect 85652 6636 87276 6692
rect 87332 6636 87342 6692
rect 87826 6636 87836 6692
rect 87892 6636 89516 6692
rect 89572 6636 89582 6692
rect 16818 6524 16828 6580
rect 16884 6524 20412 6580
rect 20468 6524 20478 6580
rect 20860 6524 21756 6580
rect 21812 6524 21822 6580
rect 22866 6524 22876 6580
rect 22932 6524 23436 6580
rect 23492 6524 23502 6580
rect 23650 6524 23660 6580
rect 23716 6524 23996 6580
rect 24052 6524 24062 6580
rect 20860 6468 20916 6524
rect 24780 6468 24836 6636
rect 39788 6580 39844 6636
rect 25890 6524 25900 6580
rect 25956 6524 29932 6580
rect 29988 6524 29998 6580
rect 30594 6524 30604 6580
rect 30660 6524 33180 6580
rect 33236 6524 38108 6580
rect 38164 6524 38174 6580
rect 38994 6524 39004 6580
rect 39060 6524 39844 6580
rect 41132 6580 41188 6636
rect 77420 6580 77476 6636
rect 81340 6580 81396 6636
rect 85652 6580 85708 6636
rect 92428 6580 92484 6860
rect 97412 6748 100268 6804
rect 100324 6748 100334 6804
rect 102050 6748 102060 6804
rect 102116 6748 102732 6804
rect 102788 6748 102798 6804
rect 104822 6748 104860 6804
rect 104916 6748 104926 6804
rect 92754 6636 92764 6692
rect 92820 6636 93884 6692
rect 93940 6636 94668 6692
rect 94724 6636 94734 6692
rect 97412 6580 97468 6748
rect 105756 6692 105812 6860
rect 110226 6748 110236 6804
rect 110292 6748 110628 6804
rect 114258 6748 114268 6804
rect 114324 6748 117852 6804
rect 117908 6748 117918 6804
rect 102386 6636 102396 6692
rect 102452 6636 105420 6692
rect 105476 6636 105486 6692
rect 105756 6636 110348 6692
rect 110404 6636 110414 6692
rect 41132 6524 42252 6580
rect 42308 6524 42318 6580
rect 43138 6524 43148 6580
rect 43204 6524 44156 6580
rect 44212 6524 44222 6580
rect 44370 6524 44380 6580
rect 44436 6524 45388 6580
rect 45444 6524 45454 6580
rect 48850 6524 48860 6580
rect 48916 6524 49644 6580
rect 49700 6524 49710 6580
rect 49970 6524 49980 6580
rect 50036 6524 54124 6580
rect 54180 6524 54190 6580
rect 55794 6524 55804 6580
rect 55860 6524 57484 6580
rect 57540 6524 57550 6580
rect 61170 6524 61180 6580
rect 61236 6524 66332 6580
rect 66388 6524 66398 6580
rect 66882 6524 66892 6580
rect 66948 6524 72268 6580
rect 72324 6524 72334 6580
rect 72818 6524 72828 6580
rect 72884 6524 73724 6580
rect 73780 6524 73790 6580
rect 73892 6524 74172 6580
rect 74228 6524 77476 6580
rect 80098 6524 80108 6580
rect 80164 6524 81116 6580
rect 81172 6524 81182 6580
rect 81340 6524 84140 6580
rect 84196 6524 84206 6580
rect 84466 6524 84476 6580
rect 84532 6524 85708 6580
rect 85922 6524 85932 6580
rect 85988 6524 87724 6580
rect 87780 6524 87790 6580
rect 92428 6524 97468 6580
rect 100930 6524 100940 6580
rect 100996 6524 103404 6580
rect 103460 6524 103470 6580
rect 104178 6524 104188 6580
rect 104244 6524 107212 6580
rect 107268 6524 107278 6580
rect 73892 6468 73948 6524
rect 110572 6468 110628 6748
rect 112354 6524 112364 6580
rect 112420 6524 112924 6580
rect 112980 6524 113708 6580
rect 113764 6524 113774 6580
rect 114706 6524 114716 6580
rect 114772 6524 115500 6580
rect 115556 6524 115566 6580
rect 19618 6412 19628 6468
rect 19684 6412 20916 6468
rect 21074 6412 21084 6468
rect 21140 6412 24780 6468
rect 24836 6412 24846 6468
rect 26898 6412 26908 6468
rect 26964 6412 27580 6468
rect 27636 6412 27646 6468
rect 28354 6412 28364 6468
rect 28420 6412 29148 6468
rect 29204 6412 29214 6468
rect 37426 6412 37436 6468
rect 37492 6412 39228 6468
rect 39284 6412 40124 6468
rect 40180 6412 40190 6468
rect 43922 6412 43932 6468
rect 43988 6412 44268 6468
rect 44324 6412 44604 6468
rect 44660 6412 44670 6468
rect 50530 6412 50540 6468
rect 50596 6412 52108 6468
rect 52164 6412 52174 6468
rect 52434 6412 52444 6468
rect 52500 6412 53340 6468
rect 53396 6412 53406 6468
rect 56018 6412 56028 6468
rect 56084 6412 58492 6468
rect 58548 6412 58558 6468
rect 61730 6412 61740 6468
rect 61796 6412 62188 6468
rect 62244 6412 63084 6468
rect 63140 6412 63150 6468
rect 68450 6412 68460 6468
rect 68516 6412 73948 6468
rect 76402 6412 76412 6468
rect 76468 6412 81788 6468
rect 81844 6412 81854 6468
rect 84690 6412 84700 6468
rect 84756 6412 84766 6468
rect 86930 6412 86940 6468
rect 86996 6412 88060 6468
rect 88116 6412 88126 6468
rect 89058 6412 89068 6468
rect 89124 6412 90860 6468
rect 90916 6412 90926 6468
rect 93426 6412 93436 6468
rect 93492 6412 94892 6468
rect 94948 6412 94958 6468
rect 95218 6412 95228 6468
rect 95284 6412 97244 6468
rect 97300 6412 97310 6468
rect 100482 6412 100492 6468
rect 100548 6412 103516 6468
rect 103572 6412 103582 6468
rect 106642 6412 106652 6468
rect 106708 6412 107436 6468
rect 107492 6412 109228 6468
rect 109284 6412 109294 6468
rect 110572 6412 114380 6468
rect 114436 6412 114446 6468
rect 117282 6412 117292 6468
rect 117348 6412 118636 6468
rect 118692 6412 134092 6468
rect 134148 6412 134158 6468
rect 27580 6356 27636 6412
rect 84700 6356 84756 6412
rect 23100 6300 26460 6356
rect 26516 6300 27356 6356
rect 27412 6300 27422 6356
rect 27580 6300 28924 6356
rect 28980 6300 28990 6356
rect 34178 6300 34188 6356
rect 34244 6300 39452 6356
rect 39508 6300 39518 6356
rect 42354 6300 42364 6356
rect 42420 6300 44044 6356
rect 44100 6300 48748 6356
rect 48804 6300 48814 6356
rect 51650 6300 51660 6356
rect 51716 6300 54684 6356
rect 54740 6300 55580 6356
rect 55636 6300 55646 6356
rect 70690 6300 70700 6356
rect 70756 6300 72044 6356
rect 72100 6300 72110 6356
rect 72230 6300 72268 6356
rect 72324 6300 72334 6356
rect 77634 6300 77644 6356
rect 77700 6300 81172 6356
rect 84130 6300 84140 6356
rect 84196 6300 84756 6356
rect 85026 6300 85036 6356
rect 85092 6300 85596 6356
rect 85652 6300 86604 6356
rect 86660 6300 86670 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 23100 6132 23156 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 26674 6188 26684 6244
rect 26740 6188 32060 6244
rect 32116 6188 34076 6244
rect 34132 6188 34142 6244
rect 37314 6188 37324 6244
rect 37380 6188 45388 6244
rect 45444 6188 45454 6244
rect 61954 6188 61964 6244
rect 62020 6188 62188 6244
rect 64754 6188 64764 6244
rect 64820 6188 73948 6244
rect 62132 6132 62188 6188
rect 18386 6076 18396 6132
rect 18452 6076 23156 6132
rect 23314 6076 23324 6132
rect 23380 6076 24388 6132
rect 26786 6076 26796 6132
rect 26852 6076 29820 6132
rect 29876 6076 29886 6132
rect 39106 6076 39116 6132
rect 39172 6076 40236 6132
rect 40292 6076 40684 6132
rect 40740 6076 41468 6132
rect 41524 6076 41534 6132
rect 48290 6076 48300 6132
rect 48356 6076 52556 6132
rect 52612 6076 52622 6132
rect 62132 6076 68460 6132
rect 68516 6076 68526 6132
rect 24332 6020 24388 6076
rect 73892 6020 73948 6188
rect 81116 6132 81172 6300
rect 81266 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81550 6300
rect 86940 6244 86996 6412
rect 93436 6356 93492 6412
rect 88946 6300 88956 6356
rect 89012 6300 93492 6356
rect 93548 6300 94556 6356
rect 94612 6300 94622 6356
rect 96226 6300 96236 6356
rect 96292 6300 109228 6356
rect 112354 6300 112364 6356
rect 112420 6300 113484 6356
rect 113540 6300 113550 6356
rect 93548 6244 93604 6300
rect 84914 6188 84924 6244
rect 84980 6188 86996 6244
rect 87154 6188 87164 6244
rect 87220 6188 89292 6244
rect 89348 6188 89358 6244
rect 90514 6188 90524 6244
rect 90580 6188 93100 6244
rect 93156 6188 93604 6244
rect 102834 6188 102844 6244
rect 102900 6188 106092 6244
rect 106148 6188 106158 6244
rect 109172 6132 109228 6300
rect 111986 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112270 6300
rect 142706 6244 142716 6300
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142980 6244 142990 6300
rect 78418 6076 78428 6132
rect 78484 6076 79436 6132
rect 79492 6076 79502 6132
rect 81116 6076 85820 6132
rect 85876 6076 88116 6132
rect 93314 6076 93324 6132
rect 93380 6076 94220 6132
rect 94276 6076 94286 6132
rect 95218 6076 95228 6132
rect 95284 6076 97916 6132
rect 97972 6076 97982 6132
rect 106866 6076 106876 6132
rect 106932 6076 108780 6132
rect 108836 6076 108846 6132
rect 109172 6076 114268 6132
rect 114324 6076 114334 6132
rect 115154 6076 115164 6132
rect 115220 6076 117628 6132
rect 117684 6076 117694 6132
rect 24332 5964 27244 6020
rect 27300 5964 27310 6020
rect 28886 5964 28924 6020
rect 28980 5964 28990 6020
rect 29586 5964 29596 6020
rect 29652 5964 30044 6020
rect 30100 5964 32060 6020
rect 32116 5964 32126 6020
rect 34626 5964 34636 6020
rect 34692 5964 37548 6020
rect 37604 5964 38220 6020
rect 38276 5964 38286 6020
rect 41010 5964 41020 6020
rect 41076 5964 41916 6020
rect 41972 5964 43372 6020
rect 43428 5964 43438 6020
rect 51874 5964 51884 6020
rect 51940 5964 52780 6020
rect 52836 5964 52846 6020
rect 53330 5964 53340 6020
rect 53396 5964 56812 6020
rect 56868 5964 56878 6020
rect 60274 5964 60284 6020
rect 60340 5964 60620 6020
rect 60676 5964 62188 6020
rect 66322 5964 66332 6020
rect 66388 5964 68012 6020
rect 68068 5964 72940 6020
rect 72996 5964 73006 6020
rect 73154 5964 73164 6020
rect 73220 5964 73388 6020
rect 73444 5964 73454 6020
rect 73892 5964 75292 6020
rect 75348 5964 76972 6020
rect 77028 5964 77038 6020
rect 78306 5964 78316 6020
rect 78372 5964 82348 6020
rect 62132 5908 62188 5964
rect 21858 5852 21868 5908
rect 21924 5852 23212 5908
rect 23268 5852 23278 5908
rect 26338 5852 26348 5908
rect 26404 5852 26908 5908
rect 27346 5852 27356 5908
rect 27412 5852 35756 5908
rect 35812 5852 35822 5908
rect 38322 5852 38332 5908
rect 38388 5852 39900 5908
rect 39956 5852 39966 5908
rect 40226 5852 40236 5908
rect 40292 5852 40908 5908
rect 40964 5852 40974 5908
rect 41570 5852 41580 5908
rect 41636 5852 41646 5908
rect 45266 5852 45276 5908
rect 45332 5852 48860 5908
rect 48916 5852 48926 5908
rect 52658 5852 52668 5908
rect 52724 5852 54236 5908
rect 54292 5852 54302 5908
rect 62132 5852 63868 5908
rect 63924 5852 63934 5908
rect 67554 5852 67564 5908
rect 67620 5852 69132 5908
rect 69188 5852 69198 5908
rect 72370 5852 72380 5908
rect 72436 5852 78652 5908
rect 78708 5852 78718 5908
rect 26852 5796 26908 5852
rect 41580 5796 41636 5852
rect 26852 5740 31500 5796
rect 31556 5740 36988 5796
rect 37044 5740 37054 5796
rect 37314 5740 37324 5796
rect 37380 5740 38444 5796
rect 38500 5740 38510 5796
rect 40236 5740 41636 5796
rect 42802 5740 42812 5796
rect 42868 5740 49644 5796
rect 49700 5740 51548 5796
rect 51604 5740 51614 5796
rect 57698 5740 57708 5796
rect 57764 5740 64092 5796
rect 64148 5740 64876 5796
rect 64932 5740 64942 5796
rect 67106 5740 67116 5796
rect 67172 5740 68460 5796
rect 68516 5740 69244 5796
rect 69300 5740 69310 5796
rect 40236 5684 40292 5740
rect 82292 5684 82348 5964
rect 88060 5908 88116 6076
rect 115164 6020 115220 6076
rect 91858 5964 91868 6020
rect 91924 5964 92652 6020
rect 92708 5964 92718 6020
rect 95078 5964 95116 6020
rect 95172 5964 95182 6020
rect 104850 5964 104860 6020
rect 104916 5964 107884 6020
rect 107940 5964 109228 6020
rect 110674 5964 110684 6020
rect 110740 5964 111356 6020
rect 111412 5964 111422 6020
rect 112690 5964 112700 6020
rect 112756 5964 115220 6020
rect 116834 5964 116844 6020
rect 116900 5964 119084 6020
rect 119140 5964 119150 6020
rect 85782 5852 85820 5908
rect 85876 5852 85886 5908
rect 86482 5852 86492 5908
rect 86548 5852 87836 5908
rect 87892 5852 87902 5908
rect 88060 5852 94108 5908
rect 94182 5852 94220 5908
rect 94276 5852 95004 5908
rect 95060 5852 95070 5908
rect 95554 5852 95564 5908
rect 95620 5852 100940 5908
rect 100996 5852 101006 5908
rect 94052 5796 94108 5852
rect 109172 5796 109228 5964
rect 111570 5852 111580 5908
rect 111636 5852 112924 5908
rect 112980 5852 112990 5908
rect 117842 5852 117852 5908
rect 117908 5852 119644 5908
rect 119700 5852 119710 5908
rect 82786 5740 82796 5796
rect 82852 5740 86268 5796
rect 86324 5740 86334 5796
rect 86706 5740 86716 5796
rect 86772 5740 87052 5796
rect 87108 5740 88284 5796
rect 88340 5740 88350 5796
rect 94052 5740 103740 5796
rect 103796 5740 103806 5796
rect 109172 5740 117068 5796
rect 117124 5740 117134 5796
rect 117628 5740 119420 5796
rect 119476 5740 119486 5796
rect 117628 5684 117684 5740
rect 19058 5628 19068 5684
rect 19124 5628 25228 5684
rect 25284 5628 25900 5684
rect 25956 5628 25966 5684
rect 36754 5628 36764 5684
rect 36820 5628 40012 5684
rect 40068 5628 40078 5684
rect 40226 5628 40236 5684
rect 40292 5628 40302 5684
rect 42914 5628 42924 5684
rect 42980 5628 49196 5684
rect 49252 5628 49262 5684
rect 72034 5628 72044 5684
rect 72100 5628 80668 5684
rect 80724 5628 80734 5684
rect 82292 5628 87164 5684
rect 87220 5628 87230 5684
rect 88498 5628 88508 5684
rect 88564 5628 91868 5684
rect 91924 5628 91934 5684
rect 115938 5628 115948 5684
rect 116004 5628 117628 5684
rect 117684 5628 117694 5684
rect 118626 5628 118636 5684
rect 118692 5628 127148 5684
rect 127204 5628 127214 5684
rect 17490 5516 17500 5572
rect 17556 5516 31836 5572
rect 31892 5516 31902 5572
rect 45378 5516 45388 5572
rect 45444 5516 56476 5572
rect 56532 5516 56542 5572
rect 86258 5516 86268 5572
rect 86324 5516 89404 5572
rect 89460 5516 89470 5572
rect 97794 5516 97804 5572
rect 97860 5516 100492 5572
rect 100548 5516 100558 5572
rect 101602 5516 101612 5572
rect 101668 5516 102844 5572
rect 102900 5516 104748 5572
rect 104804 5516 109564 5572
rect 109620 5516 109630 5572
rect 111234 5516 111244 5572
rect 111300 5516 116396 5572
rect 116452 5516 117852 5572
rect 117908 5516 117918 5572
rect 118514 5516 118524 5572
rect 118580 5516 121660 5572
rect 121716 5516 121726 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 96626 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96910 5516
rect 127346 5460 127356 5516
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127620 5460 127630 5516
rect 158066 5460 158076 5516
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158340 5460 158350 5516
rect 21522 5404 21532 5460
rect 21588 5404 22316 5460
rect 22372 5404 22382 5460
rect 52770 5404 52780 5460
rect 52836 5404 57036 5460
rect 57092 5404 57102 5460
rect 69346 5404 69356 5460
rect 69412 5404 92484 5460
rect 97234 5404 97244 5460
rect 97300 5404 111860 5460
rect 120306 5404 120316 5460
rect 120372 5404 122892 5460
rect 122948 5404 122958 5460
rect 138898 5404 138908 5460
rect 138964 5404 142940 5460
rect 142996 5404 143006 5460
rect 19170 5292 19180 5348
rect 19236 5292 20300 5348
rect 20356 5292 21868 5348
rect 21924 5292 21934 5348
rect 32946 5292 32956 5348
rect 33012 5292 41132 5348
rect 41188 5292 42980 5348
rect 45602 5292 45612 5348
rect 45668 5292 47740 5348
rect 47796 5292 47806 5348
rect 53330 5292 53340 5348
rect 53396 5292 57260 5348
rect 57316 5292 57326 5348
rect 66770 5292 66780 5348
rect 66836 5292 68460 5348
rect 68516 5292 68526 5348
rect 69458 5292 69468 5348
rect 69524 5292 72604 5348
rect 72660 5292 73052 5348
rect 73108 5292 73118 5348
rect 77074 5292 77084 5348
rect 77140 5292 77644 5348
rect 77700 5292 77710 5348
rect 82908 5292 87052 5348
rect 87108 5292 87118 5348
rect 42924 5236 42980 5292
rect 15092 5180 16380 5236
rect 16436 5180 16446 5236
rect 16594 5180 16604 5236
rect 16660 5180 19292 5236
rect 19348 5180 19358 5236
rect 21746 5180 21756 5236
rect 21812 5180 23548 5236
rect 23604 5180 23614 5236
rect 34178 5180 34188 5236
rect 34244 5180 35308 5236
rect 35364 5180 35374 5236
rect 37202 5180 37212 5236
rect 37268 5180 38332 5236
rect 38388 5180 38398 5236
rect 38882 5180 38892 5236
rect 38948 5180 39900 5236
rect 39956 5180 41244 5236
rect 41300 5180 41310 5236
rect 42914 5180 42924 5236
rect 42980 5180 43260 5236
rect 43316 5180 43326 5236
rect 43698 5180 43708 5236
rect 43764 5180 48748 5236
rect 48804 5180 48814 5236
rect 56578 5180 56588 5236
rect 56644 5180 57036 5236
rect 57092 5180 57102 5236
rect 68796 5180 70700 5236
rect 70756 5180 70766 5236
rect 73490 5180 73500 5236
rect 73556 5180 74172 5236
rect 74228 5180 74238 5236
rect 15092 5124 15148 5180
rect 68796 5124 68852 5180
rect 82908 5124 82964 5292
rect 92428 5236 92484 5404
rect 111804 5348 111860 5404
rect 98690 5292 98700 5348
rect 98756 5292 101724 5348
rect 101780 5292 101790 5348
rect 108546 5292 108556 5348
rect 108612 5292 111636 5348
rect 111794 5292 111804 5348
rect 111860 5292 136220 5348
rect 136276 5292 136286 5348
rect 142034 5292 142044 5348
rect 142100 5292 147868 5348
rect 147924 5292 147934 5348
rect 111580 5236 111636 5292
rect 89618 5180 89628 5236
rect 89684 5180 91980 5236
rect 92036 5180 92046 5236
rect 92418 5180 92428 5236
rect 92484 5180 92494 5236
rect 94780 5180 100044 5236
rect 100100 5180 100110 5236
rect 110086 5180 110124 5236
rect 110180 5180 110190 5236
rect 111318 5180 111356 5236
rect 111412 5180 111422 5236
rect 111580 5180 112364 5236
rect 112420 5180 112430 5236
rect 137330 5180 137340 5236
rect 137396 5180 140140 5236
rect 140196 5180 140206 5236
rect 142146 5180 142156 5236
rect 142212 5180 142940 5236
rect 142996 5180 143006 5236
rect 94780 5124 94836 5180
rect 11330 5068 11340 5124
rect 11396 5068 15148 5124
rect 17042 5068 17052 5124
rect 17108 5068 21308 5124
rect 21364 5068 21374 5124
rect 29474 5068 29484 5124
rect 29540 5068 40236 5124
rect 40292 5068 40302 5124
rect 41346 5068 41356 5124
rect 41412 5068 42252 5124
rect 42308 5068 42318 5124
rect 53666 5068 53676 5124
rect 53732 5068 54908 5124
rect 54964 5068 54974 5124
rect 59938 5068 59948 5124
rect 60004 5068 61964 5124
rect 62020 5068 62030 5124
rect 65202 5068 65212 5124
rect 65268 5068 67788 5124
rect 67844 5068 67854 5124
rect 68674 5068 68684 5124
rect 68740 5068 68852 5124
rect 69010 5068 69020 5124
rect 69076 5068 71596 5124
rect 71652 5068 71662 5124
rect 72230 5068 72268 5124
rect 72324 5068 75740 5124
rect 75796 5068 75806 5124
rect 76178 5068 76188 5124
rect 76244 5068 82908 5124
rect 82964 5068 82974 5124
rect 83234 5068 83244 5124
rect 83300 5068 86380 5124
rect 86436 5068 86446 5124
rect 88610 5068 88620 5124
rect 88676 5068 94836 5124
rect 94994 5068 95004 5124
rect 95060 5068 95564 5124
rect 95620 5068 95630 5124
rect 98242 5068 98252 5124
rect 98308 5068 98924 5124
rect 98980 5068 98990 5124
rect 104514 5068 104524 5124
rect 104580 5068 111916 5124
rect 111972 5068 119308 5124
rect 119364 5068 119374 5124
rect 135762 5068 135772 5124
rect 135828 5068 138236 5124
rect 138292 5068 138302 5124
rect 141698 5068 141708 5124
rect 141764 5068 144732 5124
rect 144788 5068 144798 5124
rect 147634 5068 147644 5124
rect 147700 5068 148092 5124
rect 148148 5068 148158 5124
rect 21308 5012 21364 5068
rect 17826 4956 17836 5012
rect 17892 4956 18844 5012
rect 18900 4956 20300 5012
rect 20356 4956 20366 5012
rect 21308 4956 23212 5012
rect 23268 4956 23278 5012
rect 25666 4956 25676 5012
rect 25732 4956 28812 5012
rect 28868 4956 28878 5012
rect 30706 4956 30716 5012
rect 30772 4956 33180 5012
rect 33236 4956 33246 5012
rect 36082 4956 36092 5012
rect 36148 4956 37436 5012
rect 37492 4956 37502 5012
rect 42578 4956 42588 5012
rect 42644 4956 43596 5012
rect 43652 4956 43662 5012
rect 47394 4956 47404 5012
rect 47460 4956 48076 5012
rect 48132 4956 50876 5012
rect 50932 4956 50942 5012
rect 52770 4956 52780 5012
rect 52836 4956 55020 5012
rect 55076 4956 57148 5012
rect 57204 4956 57214 5012
rect 58930 4956 58940 5012
rect 58996 4956 60396 5012
rect 60452 4956 60462 5012
rect 61702 4956 61740 5012
rect 61796 4956 61806 5012
rect 65762 4956 65772 5012
rect 65828 4956 66556 5012
rect 66612 4956 67228 5012
rect 67284 4956 67294 5012
rect 67666 4956 67676 5012
rect 67732 4956 71148 5012
rect 71204 4956 71214 5012
rect 72706 4956 72716 5012
rect 72772 4956 76524 5012
rect 76580 4956 76590 5012
rect 80210 4956 80220 5012
rect 80276 4956 86940 5012
rect 86996 4956 87006 5012
rect 96002 4956 96012 5012
rect 96068 4956 99036 5012
rect 99092 4956 99102 5012
rect 102162 4956 102172 5012
rect 102228 4956 103740 5012
rect 103796 4956 103806 5012
rect 106754 4956 106764 5012
rect 106820 4956 107660 5012
rect 107716 4956 107726 5012
rect 111804 4956 120988 5012
rect 124786 4956 124796 5012
rect 124852 4956 125580 5012
rect 125636 4956 128044 5012
rect 128100 4956 128110 5012
rect 137732 4956 149772 5012
rect 149828 4956 149838 5012
rect 111804 4900 111860 4956
rect 120932 4900 120988 4956
rect 137732 4900 137788 4956
rect 18610 4844 18620 4900
rect 18676 4844 20468 4900
rect 20626 4844 20636 4900
rect 20692 4844 32060 4900
rect 32116 4844 32126 4900
rect 36866 4844 36876 4900
rect 36932 4844 40796 4900
rect 40852 4844 40862 4900
rect 41458 4844 41468 4900
rect 41524 4844 50428 4900
rect 52994 4844 53004 4900
rect 53060 4844 56588 4900
rect 56644 4844 56654 4900
rect 63634 4844 63644 4900
rect 63700 4844 76412 4900
rect 76468 4844 76478 4900
rect 80434 4844 80444 4900
rect 80500 4844 82348 4900
rect 82404 4844 83692 4900
rect 83748 4844 83758 4900
rect 87154 4844 87164 4900
rect 87220 4844 91756 4900
rect 91812 4844 91822 4900
rect 96226 4844 96236 4900
rect 96292 4844 101780 4900
rect 103618 4844 103628 4900
rect 103684 4844 107324 4900
rect 107380 4844 107390 4900
rect 111794 4844 111804 4900
rect 111860 4844 111870 4900
rect 112578 4844 112588 4900
rect 112644 4844 113260 4900
rect 113316 4844 113326 4900
rect 115910 4844 115948 4900
rect 116004 4844 116956 4900
rect 117012 4844 117022 4900
rect 117842 4844 117852 4900
rect 117908 4844 117918 4900
rect 120932 4844 137788 4900
rect 138338 4844 138348 4900
rect 138404 4844 141484 4900
rect 141540 4844 141550 4900
rect 142706 4844 142716 4900
rect 142772 4844 143948 4900
rect 144004 4844 144014 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 20412 4676 20468 4844
rect 28018 4732 28028 4788
rect 28084 4732 28700 4788
rect 28756 4732 29820 4788
rect 29876 4732 29886 4788
rect 31826 4732 31836 4788
rect 31892 4732 34636 4788
rect 34692 4732 34702 4788
rect 34850 4732 34860 4788
rect 34916 4732 34926 4788
rect 39442 4732 39452 4788
rect 39508 4732 43932 4788
rect 43988 4732 47964 4788
rect 48020 4732 48030 4788
rect 34860 4676 34916 4732
rect 20412 4620 26460 4676
rect 26516 4620 28140 4676
rect 28196 4620 28206 4676
rect 28364 4620 34916 4676
rect 39106 4620 39116 4676
rect 39172 4620 47180 4676
rect 47236 4620 47246 4676
rect 28364 4564 28420 4620
rect 50372 4564 50428 4844
rect 51538 4732 51548 4788
rect 51604 4732 64596 4788
rect 68898 4732 68908 4788
rect 68964 4732 69468 4788
rect 69524 4732 71036 4788
rect 71092 4732 71102 4788
rect 95330 4732 95340 4788
rect 95396 4732 96124 4788
rect 96180 4732 96190 4788
rect 97234 4732 97244 4788
rect 97300 4732 100716 4788
rect 100772 4732 100782 4788
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 64540 4676 64596 4732
rect 81266 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81550 4732
rect 101724 4676 101780 4844
rect 117852 4788 117908 4844
rect 101938 4732 101948 4788
rect 102004 4732 103740 4788
rect 103796 4732 103806 4788
rect 104178 4732 104188 4788
rect 104244 4732 104254 4788
rect 107426 4732 107436 4788
rect 107492 4732 110012 4788
rect 110068 4732 110078 4788
rect 117852 4732 131180 4788
rect 131236 4732 131246 4788
rect 104188 4676 104244 4732
rect 111986 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112270 4732
rect 142706 4676 142716 4732
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142980 4676 142990 4732
rect 61506 4620 61516 4676
rect 61572 4620 64316 4676
rect 64372 4620 64382 4676
rect 64530 4620 64540 4676
rect 64596 4620 64606 4676
rect 74274 4620 74284 4676
rect 74340 4620 76412 4676
rect 76468 4620 79100 4676
rect 79156 4620 79166 4676
rect 83122 4620 83132 4676
rect 83188 4620 85036 4676
rect 85092 4620 85102 4676
rect 85474 4620 85484 4676
rect 85540 4620 100156 4676
rect 100212 4620 100222 4676
rect 101724 4620 104244 4676
rect 105634 4620 105644 4676
rect 105700 4620 108556 4676
rect 108612 4620 110124 4676
rect 110180 4620 110190 4676
rect 116722 4620 116732 4676
rect 116788 4620 118748 4676
rect 118804 4620 118814 4676
rect 122546 4620 122556 4676
rect 122612 4620 125244 4676
rect 125300 4620 125310 4676
rect 23314 4508 23324 4564
rect 23380 4508 25676 4564
rect 25732 4508 25742 4564
rect 28252 4508 28420 4564
rect 29708 4508 33964 4564
rect 34020 4508 34030 4564
rect 34850 4508 34860 4564
rect 34916 4508 39340 4564
rect 39396 4508 39406 4564
rect 42578 4508 42588 4564
rect 42644 4508 46508 4564
rect 46564 4508 46574 4564
rect 50372 4508 65548 4564
rect 65604 4508 65614 4564
rect 75506 4508 75516 4564
rect 75572 4508 76972 4564
rect 77028 4508 77038 4564
rect 85586 4508 85596 4564
rect 85652 4508 86044 4564
rect 86100 4508 86110 4564
rect 86482 4508 86492 4564
rect 86548 4508 91196 4564
rect 91252 4508 91262 4564
rect 105858 4508 105868 4564
rect 105924 4508 110908 4564
rect 110964 4508 110974 4564
rect 111346 4508 111356 4564
rect 111412 4508 113036 4564
rect 113092 4508 113820 4564
rect 113876 4508 113886 4564
rect 126130 4508 126140 4564
rect 126196 4508 132524 4564
rect 132580 4508 132590 4564
rect 13794 4396 13804 4452
rect 13860 4396 15484 4452
rect 15540 4396 15550 4452
rect 16818 4396 16828 4452
rect 16884 4396 18956 4452
rect 19012 4396 19022 4452
rect 22866 4396 22876 4452
rect 22932 4396 27132 4452
rect 27188 4396 27198 4452
rect 28252 4340 28308 4508
rect 29708 4452 29764 4508
rect 28466 4396 28476 4452
rect 28532 4396 29148 4452
rect 29204 4396 29214 4452
rect 29596 4396 29764 4452
rect 32050 4396 32060 4452
rect 32116 4396 34636 4452
rect 34692 4396 34702 4452
rect 41458 4396 41468 4452
rect 41524 4396 44604 4452
rect 44660 4396 44670 4452
rect 49298 4396 49308 4452
rect 49364 4396 51212 4452
rect 51268 4396 51278 4452
rect 56690 4396 56700 4452
rect 56756 4396 62524 4452
rect 62580 4396 62590 4452
rect 68012 4396 79436 4452
rect 79492 4396 81116 4452
rect 81172 4396 81182 4452
rect 84466 4396 84476 4452
rect 84532 4396 86604 4452
rect 86660 4396 89964 4452
rect 90020 4396 90030 4452
rect 93874 4396 93884 4452
rect 93940 4396 94556 4452
rect 94612 4396 94622 4452
rect 99026 4396 99036 4452
rect 99092 4396 105756 4452
rect 105812 4396 105822 4452
rect 121202 4396 121212 4452
rect 121268 4396 122780 4452
rect 122836 4396 122846 4452
rect 124562 4396 124572 4452
rect 124628 4396 127260 4452
rect 127316 4396 127326 4452
rect 127922 4396 127932 4452
rect 127988 4396 129948 4452
rect 130004 4396 130014 4452
rect 136882 4396 136892 4452
rect 136948 4396 137676 4452
rect 137732 4396 137742 4452
rect 22082 4284 22092 4340
rect 22148 4284 24108 4340
rect 24164 4284 24174 4340
rect 24434 4284 24444 4340
rect 24500 4284 28308 4340
rect 24108 4228 24164 4284
rect 29596 4228 29652 4396
rect 68012 4340 68068 4396
rect 29810 4284 29820 4340
rect 29876 4284 34972 4340
rect 35028 4284 35038 4340
rect 47618 4284 47628 4340
rect 47684 4284 48748 4340
rect 48804 4284 48814 4340
rect 51874 4284 51884 4340
rect 51940 4284 51996 4340
rect 52052 4284 52062 4340
rect 55682 4284 55692 4340
rect 55748 4284 68068 4340
rect 69234 4284 69244 4340
rect 69300 4284 73164 4340
rect 73220 4284 73230 4340
rect 76514 4284 76524 4340
rect 76580 4284 77196 4340
rect 77252 4284 77262 4340
rect 85474 4284 85484 4340
rect 85540 4284 86156 4340
rect 86212 4284 86222 4340
rect 92530 4284 92540 4340
rect 92596 4284 96236 4340
rect 96292 4284 96302 4340
rect 108098 4284 108108 4340
rect 108164 4284 110572 4340
rect 110628 4284 110638 4340
rect 113250 4284 113260 4340
rect 113316 4284 115388 4340
rect 115444 4284 115454 4340
rect 131506 4284 131516 4340
rect 131572 4284 132300 4340
rect 132356 4284 132748 4340
rect 132804 4284 132814 4340
rect 139010 4284 139020 4340
rect 139076 4284 141932 4340
rect 141988 4284 141998 4340
rect 143042 4284 143052 4340
rect 143108 4284 144284 4340
rect 144340 4284 144350 4340
rect 24108 4172 25228 4228
rect 25284 4172 25294 4228
rect 27794 4172 27804 4228
rect 27860 4172 29652 4228
rect 30594 4172 30604 4228
rect 30660 4172 32172 4228
rect 32228 4172 32238 4228
rect 33730 4172 33740 4228
rect 33796 4172 36316 4228
rect 36372 4172 36382 4228
rect 41682 4172 41692 4228
rect 41748 4172 43708 4228
rect 43764 4172 43774 4228
rect 15474 4060 15484 4116
rect 15540 4060 17836 4116
rect 17892 4060 17902 4116
rect 26226 4060 26236 4116
rect 26292 4060 33404 4116
rect 33460 4060 39004 4116
rect 39060 4060 39070 4116
rect 51884 4004 51940 4284
rect 72790 4172 72828 4228
rect 72884 4172 77252 4228
rect 79762 4172 79772 4228
rect 79828 4172 85596 4228
rect 85652 4172 85662 4228
rect 89618 4172 89628 4228
rect 89684 4172 93548 4228
rect 93604 4172 93614 4228
rect 102946 4172 102956 4228
rect 103012 4172 107548 4228
rect 107604 4172 107614 4228
rect 111682 4172 111692 4228
rect 111748 4172 112252 4228
rect 112308 4172 112318 4228
rect 115042 4172 115052 4228
rect 115108 4172 115164 4228
rect 115220 4172 115230 4228
rect 120754 4172 120764 4228
rect 120820 4172 122892 4228
rect 122948 4172 122958 4228
rect 129154 4172 129164 4228
rect 129220 4172 130732 4228
rect 130788 4172 130798 4228
rect 142594 4172 142604 4228
rect 142660 4172 143612 4228
rect 143668 4172 143678 4228
rect 144946 4172 144956 4228
rect 145012 4172 147532 4228
rect 147588 4172 148876 4228
rect 148932 4172 148942 4228
rect 77196 4116 77252 4172
rect 63298 4060 63308 4116
rect 63364 4060 73948 4116
rect 77186 4060 77196 4116
rect 77252 4060 77262 4116
rect 79090 4060 79100 4116
rect 79156 4060 82460 4116
rect 82516 4060 82526 4116
rect 87154 4060 87164 4116
rect 87220 4060 92764 4116
rect 92820 4060 92830 4116
rect 93874 4060 93884 4116
rect 93940 4060 96012 4116
rect 96068 4060 96078 4116
rect 105970 4060 105980 4116
rect 106036 4060 107212 4116
rect 107268 4060 107278 4116
rect 118402 4060 118412 4116
rect 118468 4060 119756 4116
rect 119812 4060 119822 4116
rect 24658 3948 24668 4004
rect 24724 3948 28924 4004
rect 28980 3948 33180 4004
rect 33236 3948 33246 4004
rect 42130 3948 42140 4004
rect 42196 3948 51940 4004
rect 73892 4004 73948 4060
rect 73892 3948 85484 4004
rect 85540 3948 85550 4004
rect 91186 3948 91196 4004
rect 91252 3948 94108 4004
rect 94164 3948 94174 4004
rect 103282 3948 103292 4004
rect 103348 3948 104636 4004
rect 104692 3948 116620 4004
rect 116676 3948 116686 4004
rect 119410 3948 119420 4004
rect 119476 3948 122108 4004
rect 122164 3948 122174 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 96626 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96910 3948
rect 127346 3892 127356 3948
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127620 3892 127630 3948
rect 158066 3892 158076 3948
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158340 3892 158350 3948
rect 23762 3836 23772 3892
rect 23828 3836 31276 3892
rect 31332 3836 31342 3892
rect 97010 3836 97020 3892
rect 97076 3836 108332 3892
rect 108388 3836 108398 3892
rect 109666 3836 109676 3892
rect 109732 3836 122332 3892
rect 122388 3836 122398 3892
rect 65874 3724 65884 3780
rect 65940 3724 77980 3780
rect 78036 3724 78046 3780
rect 92306 3724 92316 3780
rect 92372 3724 103964 3780
rect 104020 3724 104030 3780
rect 110114 3724 110124 3780
rect 110180 3724 121884 3780
rect 121940 3724 121950 3780
rect 140914 3724 140924 3780
rect 140980 3724 142492 3780
rect 142548 3724 142558 3780
rect 11890 3612 11900 3668
rect 11956 3612 13356 3668
rect 13412 3612 13422 3668
rect 16146 3612 16156 3668
rect 16212 3612 17052 3668
rect 17108 3612 17118 3668
rect 17938 3612 17948 3668
rect 18004 3612 18732 3668
rect 18788 3612 18798 3668
rect 20178 3612 20188 3668
rect 20244 3612 20972 3668
rect 21028 3612 21038 3668
rect 36194 3612 36204 3668
rect 36260 3612 40796 3668
rect 40852 3612 40862 3668
rect 57586 3612 57596 3668
rect 57652 3612 59052 3668
rect 59108 3612 59118 3668
rect 64866 3612 64876 3668
rect 64932 3612 65660 3668
rect 65716 3612 65726 3668
rect 66882 3612 66892 3668
rect 66948 3612 68572 3668
rect 68628 3612 68638 3668
rect 69682 3612 69692 3668
rect 69748 3612 70476 3668
rect 70532 3612 70542 3668
rect 77746 3612 77756 3668
rect 77812 3612 78988 3668
rect 79044 3612 79054 3668
rect 81778 3612 81788 3668
rect 81844 3612 83020 3668
rect 83076 3612 83086 3668
rect 91074 3612 91084 3668
rect 91140 3612 96908 3668
rect 96964 3612 96974 3668
rect 110450 3612 110460 3668
rect 110516 3612 112924 3668
rect 112980 3612 112990 3668
rect 118066 3612 118076 3668
rect 118132 3612 120988 3668
rect 121044 3612 121054 3668
rect 122098 3612 122108 3668
rect 122164 3612 124572 3668
rect 124628 3612 124638 3668
rect 126130 3612 126140 3668
rect 126196 3612 128380 3668
rect 128436 3612 128446 3668
rect 134194 3612 134204 3668
rect 134260 3612 136108 3668
rect 136164 3612 136174 3668
rect 138338 3612 138348 3668
rect 138404 3612 139804 3668
rect 139860 3612 139870 3668
rect 142258 3612 142268 3668
rect 142324 3612 143612 3668
rect 143668 3612 143678 3668
rect 150322 3612 150332 3668
rect 150388 3612 151564 3668
rect 151620 3612 151630 3668
rect 28690 3500 28700 3556
rect 28756 3500 31052 3556
rect 31108 3500 31118 3556
rect 34962 3500 34972 3556
rect 35028 3500 35980 3556
rect 36036 3500 36046 3556
rect 38546 3500 38556 3556
rect 38612 3500 42924 3556
rect 42980 3500 42990 3556
rect 76962 3500 76972 3556
rect 77028 3500 85484 3556
rect 85540 3500 85550 3556
rect 94098 3500 94108 3556
rect 94164 3500 102620 3556
rect 102676 3500 102686 3556
rect 103954 3500 103964 3556
rect 104020 3500 109228 3556
rect 109284 3500 109294 3556
rect 120642 3500 120652 3556
rect 120708 3500 123564 3556
rect 123620 3500 123630 3556
rect 128818 3500 128828 3556
rect 128884 3500 130396 3556
rect 130452 3500 131740 3556
rect 131796 3500 131806 3556
rect 137732 3500 139244 3556
rect 139300 3500 139310 3556
rect 139570 3500 139580 3556
rect 139636 3500 143052 3556
rect 143108 3500 143118 3556
rect 145842 3500 145852 3556
rect 145908 3500 147756 3556
rect 147812 3500 147822 3556
rect 149762 3500 149772 3556
rect 149828 3500 150556 3556
rect 150612 3500 150622 3556
rect 14578 3388 14588 3444
rect 14644 3388 16268 3444
rect 16324 3388 17500 3444
rect 17556 3388 17566 3444
rect 18050 3388 18060 3444
rect 18116 3388 19740 3444
rect 19796 3388 21308 3444
rect 21364 3388 21374 3444
rect 38770 3388 38780 3444
rect 38836 3388 41804 3444
rect 41860 3388 41870 3444
rect 51510 3388 51548 3444
rect 51604 3388 51614 3444
rect 53106 3388 53116 3444
rect 53172 3388 61740 3444
rect 61796 3388 61806 3444
rect 76066 3388 76076 3444
rect 76132 3388 77644 3444
rect 77700 3388 77710 3444
rect 85922 3388 85932 3444
rect 85988 3388 87052 3444
rect 87108 3388 87118 3444
rect 96562 3388 96572 3444
rect 96628 3388 99036 3444
rect 99092 3388 99102 3444
rect 100594 3388 100604 3444
rect 100660 3388 106876 3444
rect 106932 3388 106942 3444
rect 114034 3388 114044 3444
rect 114100 3388 117628 3444
rect 117684 3388 117694 3444
rect 118850 3388 118860 3444
rect 118916 3388 119532 3444
rect 119588 3388 119598 3444
rect 120754 3388 120764 3444
rect 120820 3388 122556 3444
rect 122612 3388 122622 3444
rect 130162 3388 130172 3444
rect 130228 3388 132748 3444
rect 132804 3388 132814 3444
rect 137732 3332 137788 3500
rect 141026 3388 141036 3444
rect 141092 3388 141708 3444
rect 141764 3388 141774 3444
rect 146290 3388 146300 3444
rect 146356 3388 147532 3444
rect 147588 3388 147598 3444
rect 24882 3276 24892 3332
rect 24948 3276 43148 3332
rect 43204 3276 43214 3332
rect 44594 3276 44604 3332
rect 44660 3276 61068 3332
rect 61124 3276 61134 3332
rect 84018 3276 84028 3332
rect 84084 3276 107548 3332
rect 107604 3276 107614 3332
rect 114594 3276 114604 3332
rect 114660 3276 137788 3332
rect 24546 3164 24556 3220
rect 24612 3164 33292 3220
rect 33348 3164 33358 3220
rect 53778 3164 53788 3220
rect 53844 3164 69468 3220
rect 69524 3164 69534 3220
rect 99362 3164 99372 3220
rect 99428 3164 109676 3220
rect 109732 3164 109742 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 81266 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81550 3164
rect 111986 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112270 3164
rect 142706 3108 142716 3164
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142980 3108 142990 3164
rect 23538 3052 23548 3108
rect 23604 3052 33628 3108
rect 33684 3052 33694 3108
rect 113362 3052 113372 3108
rect 113428 3052 142380 3108
rect 142436 3052 142446 3108
rect 23090 2940 23100 2996
rect 23156 2940 48076 2996
rect 48132 2940 48142 2996
rect 63074 2940 63084 2996
rect 63140 2940 89068 2996
rect 89124 2940 89134 2996
rect 90850 2940 90860 2996
rect 90916 2940 111468 2996
rect 111524 2940 111534 2996
rect 115490 2940 115500 2996
rect 115556 2940 134988 2996
rect 135044 2940 135054 2996
rect 15698 2828 15708 2884
rect 15764 2828 40460 2884
rect 40516 2828 40526 2884
rect 51986 2828 51996 2884
rect 52052 2828 70700 2884
rect 70756 2828 70766 2884
rect 79762 2828 79772 2884
rect 79828 2828 80556 2884
rect 80612 2828 104412 2884
rect 104468 2828 104478 2884
rect 106866 2828 106876 2884
rect 106932 2828 120876 2884
rect 120932 2828 120942 2884
rect 49410 2716 49420 2772
rect 49476 2716 71708 2772
rect 71764 2716 71774 2772
rect 84354 2716 84364 2772
rect 84420 2716 105644 2772
rect 105700 2716 105710 2772
rect 113922 2716 113932 2772
rect 113988 2716 145964 2772
rect 146020 2716 146030 2772
rect 33506 2604 33516 2660
rect 33572 2604 87948 2660
rect 88004 2604 88014 2660
rect 92418 2604 92428 2660
rect 92484 2604 115052 2660
rect 115108 2604 115118 2660
rect 17826 2492 17836 2548
rect 17892 2492 38444 2548
rect 38500 2492 38510 2548
rect 61394 2492 61404 2548
rect 61460 2492 74284 2548
rect 74340 2492 74350 2548
rect 74508 2492 97132 2548
rect 97188 2492 97198 2548
rect 74508 2436 74564 2492
rect 70242 2380 70252 2436
rect 70308 2380 74564 2436
rect 75618 2380 75628 2436
rect 75684 2380 101164 2436
rect 101220 2380 101230 2436
rect 42466 2268 42476 2324
rect 42532 2268 90524 2324
rect 90580 2268 90590 2324
rect 31602 1596 31612 1652
rect 31668 1596 52332 1652
rect 52388 1596 52398 1652
rect 59378 1596 59388 1652
rect 59444 1596 89180 1652
rect 89236 1596 89246 1652
rect 103170 1596 103180 1652
rect 103236 1596 149660 1652
rect 149716 1596 149726 1652
rect 48850 1484 48860 1540
rect 48916 1484 94108 1540
rect 94164 1484 94174 1540
rect 52770 1372 52780 1428
rect 52836 1372 94780 1428
rect 94836 1372 94846 1428
rect 56130 1260 56140 1316
rect 56196 1260 94444 1316
rect 94500 1260 94510 1316
rect 59266 1148 59276 1204
rect 59332 1148 95676 1204
rect 95732 1148 95742 1204
rect 35746 1036 35756 1092
rect 35812 1036 72268 1092
rect 72324 1036 72334 1092
rect 42242 924 42252 980
rect 42308 924 80556 980
rect 80612 924 80622 980
rect 31602 812 31612 868
rect 31668 812 91644 868
rect 91700 812 91710 868
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 81276 56420 81332 56476
rect 81380 56420 81436 56476
rect 81484 56420 81540 56476
rect 111996 56420 112052 56476
rect 112100 56420 112156 56476
rect 112204 56420 112260 56476
rect 142716 56420 142772 56476
rect 142820 56420 142876 56476
rect 142924 56420 142980 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 96636 55636 96692 55692
rect 96740 55636 96796 55692
rect 96844 55636 96900 55692
rect 127356 55636 127412 55692
rect 127460 55636 127516 55692
rect 127564 55636 127620 55692
rect 158076 55636 158132 55692
rect 158180 55636 158236 55692
rect 158284 55636 158340 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 81276 54852 81332 54908
rect 81380 54852 81436 54908
rect 81484 54852 81540 54908
rect 111996 54852 112052 54908
rect 112100 54852 112156 54908
rect 112204 54852 112260 54908
rect 142716 54852 142772 54908
rect 142820 54852 142876 54908
rect 142924 54852 142980 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 96636 54068 96692 54124
rect 96740 54068 96796 54124
rect 96844 54068 96900 54124
rect 127356 54068 127412 54124
rect 127460 54068 127516 54124
rect 127564 54068 127620 54124
rect 158076 54068 158132 54124
rect 158180 54068 158236 54124
rect 158284 54068 158340 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 81276 53284 81332 53340
rect 81380 53284 81436 53340
rect 81484 53284 81540 53340
rect 111996 53284 112052 53340
rect 112100 53284 112156 53340
rect 112204 53284 112260 53340
rect 142716 53284 142772 53340
rect 142820 53284 142876 53340
rect 142924 53284 142980 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 96636 52500 96692 52556
rect 96740 52500 96796 52556
rect 96844 52500 96900 52556
rect 127356 52500 127412 52556
rect 127460 52500 127516 52556
rect 127564 52500 127620 52556
rect 158076 52500 158132 52556
rect 158180 52500 158236 52556
rect 158284 52500 158340 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 81276 51716 81332 51772
rect 81380 51716 81436 51772
rect 81484 51716 81540 51772
rect 111996 51716 112052 51772
rect 112100 51716 112156 51772
rect 112204 51716 112260 51772
rect 142716 51716 142772 51772
rect 142820 51716 142876 51772
rect 142924 51716 142980 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 96636 50932 96692 50988
rect 96740 50932 96796 50988
rect 96844 50932 96900 50988
rect 127356 50932 127412 50988
rect 127460 50932 127516 50988
rect 127564 50932 127620 50988
rect 158076 50932 158132 50988
rect 158180 50932 158236 50988
rect 158284 50932 158340 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 81276 50148 81332 50204
rect 81380 50148 81436 50204
rect 81484 50148 81540 50204
rect 111996 50148 112052 50204
rect 112100 50148 112156 50204
rect 112204 50148 112260 50204
rect 142716 50148 142772 50204
rect 142820 50148 142876 50204
rect 142924 50148 142980 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 96636 49364 96692 49420
rect 96740 49364 96796 49420
rect 96844 49364 96900 49420
rect 127356 49364 127412 49420
rect 127460 49364 127516 49420
rect 127564 49364 127620 49420
rect 158076 49364 158132 49420
rect 158180 49364 158236 49420
rect 158284 49364 158340 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 81276 48580 81332 48636
rect 81380 48580 81436 48636
rect 81484 48580 81540 48636
rect 111996 48580 112052 48636
rect 112100 48580 112156 48636
rect 112204 48580 112260 48636
rect 142716 48580 142772 48636
rect 142820 48580 142876 48636
rect 142924 48580 142980 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 96636 47796 96692 47852
rect 96740 47796 96796 47852
rect 96844 47796 96900 47852
rect 127356 47796 127412 47852
rect 127460 47796 127516 47852
rect 127564 47796 127620 47852
rect 158076 47796 158132 47852
rect 158180 47796 158236 47852
rect 158284 47796 158340 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 81276 47012 81332 47068
rect 81380 47012 81436 47068
rect 81484 47012 81540 47068
rect 111996 47012 112052 47068
rect 112100 47012 112156 47068
rect 112204 47012 112260 47068
rect 142716 47012 142772 47068
rect 142820 47012 142876 47068
rect 142924 47012 142980 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 96636 46228 96692 46284
rect 96740 46228 96796 46284
rect 96844 46228 96900 46284
rect 127356 46228 127412 46284
rect 127460 46228 127516 46284
rect 127564 46228 127620 46284
rect 158076 46228 158132 46284
rect 158180 46228 158236 46284
rect 158284 46228 158340 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 81276 45444 81332 45500
rect 81380 45444 81436 45500
rect 81484 45444 81540 45500
rect 111996 45444 112052 45500
rect 112100 45444 112156 45500
rect 112204 45444 112260 45500
rect 142716 45444 142772 45500
rect 142820 45444 142876 45500
rect 142924 45444 142980 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 96636 44660 96692 44716
rect 96740 44660 96796 44716
rect 96844 44660 96900 44716
rect 127356 44660 127412 44716
rect 127460 44660 127516 44716
rect 127564 44660 127620 44716
rect 158076 44660 158132 44716
rect 158180 44660 158236 44716
rect 158284 44660 158340 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 81276 43876 81332 43932
rect 81380 43876 81436 43932
rect 81484 43876 81540 43932
rect 111996 43876 112052 43932
rect 112100 43876 112156 43932
rect 112204 43876 112260 43932
rect 142716 43876 142772 43932
rect 142820 43876 142876 43932
rect 142924 43876 142980 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 96636 43092 96692 43148
rect 96740 43092 96796 43148
rect 96844 43092 96900 43148
rect 127356 43092 127412 43148
rect 127460 43092 127516 43148
rect 127564 43092 127620 43148
rect 158076 43092 158132 43148
rect 158180 43092 158236 43148
rect 158284 43092 158340 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 81276 42308 81332 42364
rect 81380 42308 81436 42364
rect 81484 42308 81540 42364
rect 111996 42308 112052 42364
rect 112100 42308 112156 42364
rect 112204 42308 112260 42364
rect 142716 42308 142772 42364
rect 142820 42308 142876 42364
rect 142924 42308 142980 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 96636 41524 96692 41580
rect 96740 41524 96796 41580
rect 96844 41524 96900 41580
rect 127356 41524 127412 41580
rect 127460 41524 127516 41580
rect 127564 41524 127620 41580
rect 158076 41524 158132 41580
rect 158180 41524 158236 41580
rect 158284 41524 158340 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 81276 40740 81332 40796
rect 81380 40740 81436 40796
rect 81484 40740 81540 40796
rect 111996 40740 112052 40796
rect 112100 40740 112156 40796
rect 112204 40740 112260 40796
rect 142716 40740 142772 40796
rect 142820 40740 142876 40796
rect 142924 40740 142980 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 96636 39956 96692 40012
rect 96740 39956 96796 40012
rect 96844 39956 96900 40012
rect 127356 39956 127412 40012
rect 127460 39956 127516 40012
rect 127564 39956 127620 40012
rect 158076 39956 158132 40012
rect 158180 39956 158236 40012
rect 158284 39956 158340 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 81276 39172 81332 39228
rect 81380 39172 81436 39228
rect 81484 39172 81540 39228
rect 111996 39172 112052 39228
rect 112100 39172 112156 39228
rect 112204 39172 112260 39228
rect 142716 39172 142772 39228
rect 142820 39172 142876 39228
rect 142924 39172 142980 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 96636 38388 96692 38444
rect 96740 38388 96796 38444
rect 96844 38388 96900 38444
rect 127356 38388 127412 38444
rect 127460 38388 127516 38444
rect 127564 38388 127620 38444
rect 158076 38388 158132 38444
rect 158180 38388 158236 38444
rect 158284 38388 158340 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 81276 37604 81332 37660
rect 81380 37604 81436 37660
rect 81484 37604 81540 37660
rect 111996 37604 112052 37660
rect 112100 37604 112156 37660
rect 112204 37604 112260 37660
rect 142716 37604 142772 37660
rect 142820 37604 142876 37660
rect 142924 37604 142980 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 96636 36820 96692 36876
rect 96740 36820 96796 36876
rect 96844 36820 96900 36876
rect 127356 36820 127412 36876
rect 127460 36820 127516 36876
rect 127564 36820 127620 36876
rect 158076 36820 158132 36876
rect 158180 36820 158236 36876
rect 158284 36820 158340 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 81276 36036 81332 36092
rect 81380 36036 81436 36092
rect 81484 36036 81540 36092
rect 111996 36036 112052 36092
rect 112100 36036 112156 36092
rect 112204 36036 112260 36092
rect 142716 36036 142772 36092
rect 142820 36036 142876 36092
rect 142924 36036 142980 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 96636 35252 96692 35308
rect 96740 35252 96796 35308
rect 96844 35252 96900 35308
rect 127356 35252 127412 35308
rect 127460 35252 127516 35308
rect 127564 35252 127620 35308
rect 158076 35252 158132 35308
rect 158180 35252 158236 35308
rect 158284 35252 158340 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 81276 34468 81332 34524
rect 81380 34468 81436 34524
rect 81484 34468 81540 34524
rect 111996 34468 112052 34524
rect 112100 34468 112156 34524
rect 112204 34468 112260 34524
rect 142716 34468 142772 34524
rect 142820 34468 142876 34524
rect 142924 34468 142980 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 96636 33684 96692 33740
rect 96740 33684 96796 33740
rect 96844 33684 96900 33740
rect 127356 33684 127412 33740
rect 127460 33684 127516 33740
rect 127564 33684 127620 33740
rect 158076 33684 158132 33740
rect 158180 33684 158236 33740
rect 158284 33684 158340 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 81276 32900 81332 32956
rect 81380 32900 81436 32956
rect 81484 32900 81540 32956
rect 111996 32900 112052 32956
rect 112100 32900 112156 32956
rect 112204 32900 112260 32956
rect 142716 32900 142772 32956
rect 142820 32900 142876 32956
rect 142924 32900 142980 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 96636 32116 96692 32172
rect 96740 32116 96796 32172
rect 96844 32116 96900 32172
rect 127356 32116 127412 32172
rect 127460 32116 127516 32172
rect 127564 32116 127620 32172
rect 158076 32116 158132 32172
rect 158180 32116 158236 32172
rect 158284 32116 158340 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 81276 31332 81332 31388
rect 81380 31332 81436 31388
rect 81484 31332 81540 31388
rect 111996 31332 112052 31388
rect 112100 31332 112156 31388
rect 112204 31332 112260 31388
rect 142716 31332 142772 31388
rect 142820 31332 142876 31388
rect 142924 31332 142980 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 96636 30548 96692 30604
rect 96740 30548 96796 30604
rect 96844 30548 96900 30604
rect 127356 30548 127412 30604
rect 127460 30548 127516 30604
rect 127564 30548 127620 30604
rect 158076 30548 158132 30604
rect 158180 30548 158236 30604
rect 158284 30548 158340 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 81276 29764 81332 29820
rect 81380 29764 81436 29820
rect 81484 29764 81540 29820
rect 111996 29764 112052 29820
rect 112100 29764 112156 29820
rect 112204 29764 112260 29820
rect 142716 29764 142772 29820
rect 142820 29764 142876 29820
rect 142924 29764 142980 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 96636 28980 96692 29036
rect 96740 28980 96796 29036
rect 96844 28980 96900 29036
rect 127356 28980 127412 29036
rect 127460 28980 127516 29036
rect 127564 28980 127620 29036
rect 158076 28980 158132 29036
rect 158180 28980 158236 29036
rect 158284 28980 158340 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 81276 28196 81332 28252
rect 81380 28196 81436 28252
rect 81484 28196 81540 28252
rect 111996 28196 112052 28252
rect 112100 28196 112156 28252
rect 112204 28196 112260 28252
rect 142716 28196 142772 28252
rect 142820 28196 142876 28252
rect 142924 28196 142980 28252
rect 51100 28028 51156 28084
rect 51324 27692 51380 27748
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 96636 27412 96692 27468
rect 96740 27412 96796 27468
rect 96844 27412 96900 27468
rect 127356 27412 127412 27468
rect 127460 27412 127516 27468
rect 127564 27412 127620 27468
rect 158076 27412 158132 27468
rect 158180 27412 158236 27468
rect 158284 27412 158340 27468
rect 49756 27244 49812 27300
rect 51996 27244 52052 27300
rect 35644 26908 35700 26964
rect 51436 26796 51492 26852
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 81276 26628 81332 26684
rect 81380 26628 81436 26684
rect 81484 26628 81540 26684
rect 111996 26628 112052 26684
rect 112100 26628 112156 26684
rect 112204 26628 112260 26684
rect 142716 26628 142772 26684
rect 142820 26628 142876 26684
rect 142924 26628 142980 26684
rect 49756 26572 49812 26628
rect 51212 26012 51268 26068
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 96636 25844 96692 25900
rect 96740 25844 96796 25900
rect 96844 25844 96900 25900
rect 127356 25844 127412 25900
rect 127460 25844 127516 25900
rect 127564 25844 127620 25900
rect 158076 25844 158132 25900
rect 158180 25844 158236 25900
rect 158284 25844 158340 25900
rect 50092 25452 50148 25508
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 51324 25004 51380 25060
rect 81276 25060 81332 25116
rect 81380 25060 81436 25116
rect 81484 25060 81540 25116
rect 111996 25060 112052 25116
rect 112100 25060 112156 25116
rect 112204 25060 112260 25116
rect 142716 25060 142772 25116
rect 142820 25060 142876 25116
rect 142924 25060 142980 25116
rect 66668 24892 66724 24948
rect 35644 24780 35700 24836
rect 51324 24668 51380 24724
rect 66668 24444 66724 24500
rect 55356 24332 55412 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 96636 24276 96692 24332
rect 96740 24276 96796 24332
rect 96844 24276 96900 24332
rect 127356 24276 127412 24332
rect 127460 24276 127516 24332
rect 127564 24276 127620 24332
rect 158076 24276 158132 24332
rect 158180 24276 158236 24332
rect 158284 24276 158340 24332
rect 53676 23996 53732 24052
rect 51212 23660 51268 23716
rect 51996 23660 52052 23716
rect 51100 23548 51156 23604
rect 51436 23548 51492 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 81276 23492 81332 23548
rect 81380 23492 81436 23548
rect 81484 23492 81540 23548
rect 111996 23492 112052 23548
rect 112100 23492 112156 23548
rect 112204 23492 112260 23548
rect 142716 23492 142772 23548
rect 142820 23492 142876 23548
rect 142924 23492 142980 23548
rect 52668 23324 52724 23380
rect 53676 23324 53732 23380
rect 75180 22876 75236 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 96636 22708 96692 22764
rect 96740 22708 96796 22764
rect 96844 22708 96900 22764
rect 127356 22708 127412 22764
rect 127460 22708 127516 22764
rect 127564 22708 127620 22764
rect 158076 22708 158132 22764
rect 158180 22708 158236 22764
rect 158284 22708 158340 22764
rect 50092 22540 50148 22596
rect 51548 22428 51604 22484
rect 90972 22204 91028 22260
rect 50092 22092 50148 22148
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 81276 21924 81332 21980
rect 81380 21924 81436 21980
rect 81484 21924 81540 21980
rect 111996 21924 112052 21980
rect 112100 21924 112156 21980
rect 112204 21924 112260 21980
rect 142716 21924 142772 21980
rect 142820 21924 142876 21980
rect 142924 21924 142980 21980
rect 51996 21756 52052 21812
rect 52668 21756 52724 21812
rect 55356 21644 55412 21700
rect 60620 21308 60676 21364
rect 89628 21308 89684 21364
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 96636 21140 96692 21196
rect 96740 21140 96796 21196
rect 96844 21140 96900 21196
rect 127356 21140 127412 21196
rect 127460 21140 127516 21196
rect 127564 21140 127620 21196
rect 158076 21140 158132 21196
rect 158180 21140 158236 21196
rect 158284 21140 158340 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 81276 20356 81332 20412
rect 81380 20356 81436 20412
rect 81484 20356 81540 20412
rect 111996 20356 112052 20412
rect 112100 20356 112156 20412
rect 112204 20356 112260 20412
rect 142716 20356 142772 20412
rect 142820 20356 142876 20412
rect 142924 20356 142980 20412
rect 74620 20300 74676 20356
rect 74620 20076 74676 20132
rect 87948 19964 88004 20020
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 110124 19740 110180 19796
rect 94892 19628 94948 19684
rect 44716 19516 44772 19572
rect 68236 19516 68292 19572
rect 96636 19572 96692 19628
rect 96740 19572 96796 19628
rect 96844 19572 96900 19628
rect 127356 19572 127412 19628
rect 127460 19572 127516 19628
rect 127564 19572 127620 19628
rect 158076 19572 158132 19628
rect 158180 19572 158236 19628
rect 158284 19572 158340 19628
rect 68012 19292 68068 19348
rect 68012 18956 68068 19012
rect 85484 18956 85540 19012
rect 68236 18844 68292 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 44716 18732 44772 18788
rect 81276 18788 81332 18844
rect 81380 18788 81436 18844
rect 81484 18788 81540 18844
rect 111996 18788 112052 18844
rect 112100 18788 112156 18844
rect 112204 18788 112260 18844
rect 88732 18732 88788 18788
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 90972 18396 91028 18452
rect 142716 18788 142772 18844
rect 142820 18788 142876 18844
rect 142924 18788 142980 18844
rect 94444 18284 94500 18340
rect 75180 18172 75236 18228
rect 51548 18060 51604 18116
rect 77196 18060 77252 18116
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 96636 18004 96692 18060
rect 96740 18004 96796 18060
rect 96844 18004 96900 18060
rect 127356 18004 127412 18060
rect 127460 18004 127516 18060
rect 127564 18004 127620 18060
rect 158076 18004 158132 18060
rect 158180 18004 158236 18060
rect 158284 18004 158340 18060
rect 51548 17724 51604 17780
rect 87948 17612 88004 17668
rect 57148 17388 57204 17444
rect 84364 17388 84420 17444
rect 85148 17388 85204 17444
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 89292 17276 89348 17332
rect 81276 17220 81332 17276
rect 81380 17220 81436 17276
rect 81484 17220 81540 17276
rect 111996 17220 112052 17276
rect 112100 17220 112156 17276
rect 112204 17220 112260 17276
rect 142716 17220 142772 17276
rect 142820 17220 142876 17276
rect 142924 17220 142980 17276
rect 85484 16828 85540 16884
rect 92428 16828 92484 16884
rect 95004 16716 95060 16772
rect 77196 16604 77252 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 96636 16436 96692 16492
rect 96740 16436 96796 16492
rect 96844 16436 96900 16492
rect 127356 16436 127412 16492
rect 127460 16436 127516 16492
rect 127564 16436 127620 16492
rect 158076 16436 158132 16492
rect 158180 16436 158236 16492
rect 158284 16436 158340 16492
rect 83132 15820 83188 15876
rect 83580 15820 83636 15876
rect 84476 15820 84532 15876
rect 94892 15820 94948 15876
rect 105756 15820 105812 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 81276 15652 81332 15708
rect 81380 15652 81436 15708
rect 81484 15652 81540 15708
rect 111996 15652 112052 15708
rect 112100 15652 112156 15708
rect 112204 15652 112260 15708
rect 142716 15652 142772 15708
rect 142820 15652 142876 15708
rect 142924 15652 142980 15708
rect 31836 15484 31892 15540
rect 41356 15372 41412 15428
rect 57148 15372 57204 15428
rect 39340 15148 39396 15204
rect 83020 15036 83076 15092
rect 94444 15036 94500 15092
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 96636 14868 96692 14924
rect 96740 14868 96796 14924
rect 96844 14868 96900 14924
rect 127356 14868 127412 14924
rect 127460 14868 127516 14924
rect 127564 14868 127620 14924
rect 158076 14868 158132 14924
rect 158180 14868 158236 14924
rect 158284 14868 158340 14924
rect 49756 14476 49812 14532
rect 61404 14476 61460 14532
rect 83692 14140 83748 14196
rect 83916 14140 83972 14196
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 81276 14084 81332 14140
rect 81380 14084 81436 14140
rect 81484 14084 81540 14140
rect 30492 14028 30548 14084
rect 49532 13916 49588 13972
rect 83020 13916 83076 13972
rect 83580 13916 83636 13972
rect 50316 13692 50372 13748
rect 30492 13580 30548 13636
rect 111996 14084 112052 14140
rect 112100 14084 112156 14140
rect 112204 14084 112260 14140
rect 142716 14084 142772 14140
rect 142820 14084 142876 14140
rect 142924 14084 142980 14140
rect 95004 13804 95060 13860
rect 84588 13580 84644 13636
rect 87276 13468 87332 13524
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 96636 13300 96692 13356
rect 96740 13300 96796 13356
rect 96844 13300 96900 13356
rect 127356 13300 127412 13356
rect 127460 13300 127516 13356
rect 127564 13300 127620 13356
rect 158076 13300 158132 13356
rect 158180 13300 158236 13356
rect 158284 13300 158340 13356
rect 72828 13244 72884 13300
rect 103404 13244 103460 13300
rect 49420 13132 49476 13188
rect 72268 13020 72324 13076
rect 49644 12908 49700 12964
rect 88732 12908 88788 12964
rect 60620 12796 60676 12852
rect 89292 12796 89348 12852
rect 89628 12684 89684 12740
rect 96460 12684 96516 12740
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 81276 12516 81332 12572
rect 81380 12516 81436 12572
rect 81484 12516 81540 12572
rect 111996 12516 112052 12572
rect 112100 12516 112156 12572
rect 112204 12516 112260 12572
rect 142716 12516 142772 12572
rect 142820 12516 142876 12572
rect 142924 12516 142980 12572
rect 50316 12460 50372 12516
rect 61404 12460 61460 12516
rect 87276 12460 87332 12516
rect 49756 12236 49812 12292
rect 51996 12236 52052 12292
rect 102620 12236 102676 12292
rect 85148 12012 85204 12068
rect 30828 11900 30884 11956
rect 49644 11900 49700 11956
rect 83692 11900 83748 11956
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 40348 11732 40404 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 31836 11676 31892 11732
rect 37548 11676 37604 11732
rect 40012 11676 40068 11732
rect 64652 11676 64708 11732
rect 109900 12012 109956 12068
rect 94892 11788 94948 11844
rect 96460 11788 96516 11844
rect 102620 11788 102676 11844
rect 103404 11788 103460 11844
rect 96636 11732 96692 11788
rect 96740 11732 96796 11788
rect 96844 11732 96900 11788
rect 127356 11732 127412 11788
rect 127460 11732 127516 11788
rect 127564 11732 127620 11788
rect 158076 11732 158132 11788
rect 158180 11732 158236 11788
rect 158284 11732 158340 11788
rect 94220 11676 94276 11732
rect 40124 11564 40180 11620
rect 66668 11564 66724 11620
rect 84140 11564 84196 11620
rect 100940 11564 100996 11620
rect 104860 11564 104916 11620
rect 49420 11452 49476 11508
rect 40236 11340 40292 11396
rect 61964 11452 62020 11508
rect 102620 11228 102676 11284
rect 112364 11228 112420 11284
rect 56700 11116 56756 11172
rect 66668 11116 66724 11172
rect 71708 11116 71764 11172
rect 75740 11116 75796 11172
rect 103180 11116 103236 11172
rect 43932 11004 43988 11060
rect 49532 11004 49588 11060
rect 50316 11004 50372 11060
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 40124 10892 40180 10948
rect 30828 10780 30884 10836
rect 40348 10780 40404 10836
rect 31612 10668 31668 10724
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 46060 10780 46116 10836
rect 81276 10948 81332 11004
rect 81380 10948 81436 11004
rect 81484 10948 81540 11004
rect 104748 11004 104804 11060
rect 111996 10948 112052 11004
rect 112100 10948 112156 11004
rect 112204 10948 112260 11004
rect 142716 10948 142772 11004
rect 142820 10948 142876 11004
rect 142924 10948 142980 11004
rect 61964 10892 62020 10948
rect 85484 10892 85540 10948
rect 100940 10892 100996 10948
rect 75740 10780 75796 10836
rect 83916 10780 83972 10836
rect 106092 10668 106148 10724
rect 44604 10556 44660 10612
rect 64652 10444 64708 10500
rect 102620 10444 102676 10500
rect 104748 10332 104804 10388
rect 50316 10220 50372 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 44604 10108 44660 10164
rect 115948 10220 116004 10276
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 73164 10108 73220 10164
rect 73612 10108 73668 10164
rect 82460 10108 82516 10164
rect 96636 10164 96692 10220
rect 96740 10164 96796 10220
rect 96844 10164 96900 10220
rect 127356 10164 127412 10220
rect 127460 10164 127516 10220
rect 127564 10164 127620 10220
rect 158076 10164 158132 10220
rect 158180 10164 158236 10220
rect 158284 10164 158340 10220
rect 101164 10108 101220 10164
rect 84588 9884 84644 9940
rect 37548 9660 37604 9716
rect 61068 9660 61124 9716
rect 73276 9660 73332 9716
rect 56364 9548 56420 9604
rect 51996 9436 52052 9492
rect 84140 9436 84196 9492
rect 85708 9436 85764 9492
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 81276 9380 81332 9436
rect 81380 9380 81436 9436
rect 81484 9380 81540 9436
rect 111996 9380 112052 9436
rect 112100 9380 112156 9436
rect 112204 9380 112260 9436
rect 142716 9380 142772 9436
rect 142820 9380 142876 9436
rect 142924 9380 142980 9436
rect 109900 9324 109956 9380
rect 112924 9324 112980 9380
rect 52108 9212 52164 9268
rect 72940 9212 72996 9268
rect 73612 9212 73668 9268
rect 28924 9100 28980 9156
rect 34188 9100 34244 9156
rect 52220 9100 52276 9156
rect 82460 9100 82516 9156
rect 97916 9100 97972 9156
rect 52108 8988 52164 9044
rect 52780 8988 52836 9044
rect 56364 8988 56420 9044
rect 71708 8988 71764 9044
rect 73276 8988 73332 9044
rect 51548 8876 51604 8932
rect 97916 8876 97972 8932
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 83132 8540 83188 8596
rect 95116 8540 95172 8596
rect 52332 8428 52388 8484
rect 56028 8428 56084 8484
rect 56700 8428 56756 8484
rect 96636 8596 96692 8652
rect 96740 8596 96796 8652
rect 96844 8596 96900 8652
rect 127356 8596 127412 8652
rect 127460 8596 127516 8652
rect 127564 8596 127620 8652
rect 158076 8596 158132 8652
rect 158180 8596 158236 8652
rect 158284 8596 158340 8652
rect 110908 8540 110964 8596
rect 85484 8428 85540 8484
rect 85708 8428 85764 8484
rect 86828 8428 86884 8484
rect 95676 8428 95732 8484
rect 86716 8316 86772 8372
rect 108556 8316 108612 8372
rect 112924 8316 112980 8372
rect 46060 8204 46116 8260
rect 72940 8204 72996 8260
rect 92428 8204 92484 8260
rect 111356 8204 111412 8260
rect 43708 8092 43764 8148
rect 56028 8092 56084 8148
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 84364 7980 84420 8036
rect 85484 7980 85540 8036
rect 95676 7868 95732 7924
rect 110908 7868 110964 7924
rect 81276 7812 81332 7868
rect 81380 7812 81436 7868
rect 81484 7812 81540 7868
rect 111996 7812 112052 7868
rect 112100 7812 112156 7868
rect 112204 7812 112260 7868
rect 142716 7812 142772 7868
rect 142820 7812 142876 7868
rect 142924 7812 142980 7868
rect 50316 7756 50372 7812
rect 52220 7644 52276 7700
rect 56028 7644 56084 7700
rect 84476 7644 84532 7700
rect 86716 7644 86772 7700
rect 61964 7532 62020 7588
rect 41356 7420 41412 7476
rect 43932 7420 43988 7476
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 86828 7196 86884 7252
rect 79436 7084 79492 7140
rect 115052 7084 115108 7140
rect 96636 7028 96692 7084
rect 96740 7028 96796 7084
rect 96844 7028 96900 7084
rect 127356 7028 127412 7084
rect 127460 7028 127516 7084
rect 127564 7028 127620 7084
rect 158076 7028 158132 7084
rect 158180 7028 158236 7084
rect 158284 7028 158340 7084
rect 61740 6748 61796 6804
rect 84364 6748 84420 6804
rect 85372 6748 85428 6804
rect 41580 6636 41636 6692
rect 46060 6636 46116 6692
rect 73164 6636 73220 6692
rect 104860 6748 104916 6804
rect 34188 6300 34244 6356
rect 72268 6300 72324 6356
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 61964 6188 62020 6244
rect 81276 6244 81332 6300
rect 81380 6244 81436 6300
rect 81484 6244 81540 6300
rect 112364 6300 112420 6356
rect 106092 6188 106148 6244
rect 111996 6244 112052 6300
rect 112100 6244 112156 6300
rect 112204 6244 112260 6300
rect 142716 6244 142772 6300
rect 142820 6244 142876 6300
rect 142924 6244 142980 6300
rect 85820 6076 85876 6132
rect 28924 5964 28980 6020
rect 73164 5964 73220 6020
rect 41580 5852 41636 5908
rect 95116 5964 95172 6020
rect 85820 5852 85876 5908
rect 94220 5852 94276 5908
rect 100940 5852 100996 5908
rect 115948 5628 116004 5684
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 96636 5460 96692 5516
rect 96740 5460 96796 5516
rect 96844 5460 96900 5516
rect 127356 5460 127412 5516
rect 127460 5460 127516 5516
rect 127564 5460 127620 5516
rect 158076 5460 158132 5516
rect 158180 5460 158236 5516
rect 158284 5460 158340 5516
rect 34188 5180 34244 5236
rect 43708 5180 43764 5236
rect 110124 5180 110180 5236
rect 111356 5180 111412 5236
rect 72268 5068 72324 5124
rect 61740 4956 61796 5012
rect 115948 4844 116004 4900
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 81276 4676 81332 4732
rect 81380 4676 81436 4732
rect 81484 4676 81540 4732
rect 111996 4676 112052 4732
rect 112100 4676 112156 4732
rect 112204 4676 112260 4732
rect 142716 4676 142772 4732
rect 142820 4676 142876 4732
rect 142924 4676 142980 4732
rect 108556 4620 108612 4676
rect 39340 4508 39396 4564
rect 79436 4396 79492 4452
rect 105756 4396 105812 4452
rect 51996 4284 52052 4340
rect 72828 4172 72884 4228
rect 115052 4172 115108 4228
rect 85484 3948 85540 4004
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 96636 3892 96692 3948
rect 96740 3892 96796 3948
rect 96844 3892 96900 3948
rect 127356 3892 127412 3948
rect 127460 3892 127516 3948
rect 127564 3892 127620 3948
rect 158076 3892 158132 3948
rect 158180 3892 158236 3948
rect 158284 3892 158340 3948
rect 102620 3500 102676 3556
rect 51548 3388 51604 3444
rect 44604 3276 44660 3332
rect 61068 3276 61124 3332
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 81276 3108 81332 3164
rect 81380 3108 81436 3164
rect 81484 3108 81540 3164
rect 111996 3108 112052 3164
rect 112100 3108 112156 3164
rect 112204 3108 112260 3164
rect 142716 3108 142772 3164
rect 142820 3108 142876 3164
rect 142924 3108 142980 3164
rect 71708 2716 71764 2772
rect 84364 2716 84420 2772
rect 92428 2604 92484 2660
rect 101164 2380 101220 2436
rect 52332 1596 52388 1652
rect 103180 1596 103236 1652
rect 52780 1372 52836 1428
rect 95676 1148 95732 1204
rect 72268 1036 72324 1092
rect 31612 812 31668 868
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 49756 27300 49812 27310
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35644 26964 35700 26974
rect 35644 24836 35700 26908
rect 49756 26628 49812 27244
rect 49756 26562 49812 26572
rect 50528 26684 50848 28196
rect 65888 55692 66208 56508
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 35644 24770 35700 24780
rect 50092 25508 50148 25518
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 50092 22596 50148 25452
rect 50092 22148 50148 22540
rect 50092 22082 50148 22092
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 51100 28084 51156 28094
rect 51100 23604 51156 28028
rect 51324 27748 51380 27758
rect 51212 26068 51268 26078
rect 51212 23716 51268 26012
rect 51324 25060 51380 27692
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 51996 27300 52052 27310
rect 51324 24724 51380 25004
rect 51324 24658 51380 24668
rect 51436 26852 51492 26862
rect 51212 23650 51268 23660
rect 51100 23538 51156 23548
rect 51436 23604 51492 26796
rect 51996 23716 52052 27244
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 55356 24388 55412 24398
rect 51996 23650 52052 23660
rect 53676 24052 53732 24062
rect 51436 23538 51492 23548
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 50528 21980 50848 23492
rect 52668 23380 52724 23390
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 35168 18060 35488 19572
rect 44716 19572 44772 19582
rect 44716 18788 44772 19516
rect 44716 18722 44772 18732
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 31836 15540 31892 15550
rect 19808 12572 20128 14084
rect 30492 14084 30548 14094
rect 30492 13636 30548 14028
rect 30492 13570 30548 13580
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 30828 11956 30884 11966
rect 30828 10836 30884 11900
rect 31836 11732 31892 15484
rect 31836 11666 31892 11676
rect 35168 14924 35488 16436
rect 50528 17276 50848 18788
rect 51548 22484 51604 22494
rect 51548 18116 51604 22428
rect 51548 17780 51604 18060
rect 51548 17714 51604 17724
rect 51996 21812 52052 21822
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 41356 15428 41412 15438
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 39340 15204 39396 15214
rect 30828 10770 30884 10780
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 31612 10724 31668 10734
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 28924 9156 28980 9166
rect 28924 6020 28980 9100
rect 28924 5954 28980 5964
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 31612 868 31668 10668
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 34188 9156 34244 9166
rect 34188 6356 34244 9100
rect 34188 5236 34244 6300
rect 34188 5170 34244 5180
rect 35168 8652 35488 10164
rect 37548 11732 37604 11742
rect 37548 9716 37604 11676
rect 37548 9650 37604 9660
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 39340 4564 39396 15148
rect 40348 11788 40404 11798
rect 40012 11732 40292 11788
rect 40012 11666 40068 11676
rect 40124 11620 40180 11630
rect 40124 10948 40180 11564
rect 40236 11396 40292 11732
rect 40236 11330 40292 11340
rect 40124 10882 40180 10892
rect 40348 10836 40404 11732
rect 40348 10770 40404 10780
rect 41356 7476 41412 15372
rect 49756 14532 49812 14542
rect 49532 13972 49588 13982
rect 49420 13188 49476 13198
rect 49420 11508 49476 13132
rect 49420 11442 49476 11452
rect 43932 11060 43988 11070
rect 41356 7410 41412 7420
rect 43708 8148 43764 8158
rect 41580 6692 41636 6702
rect 41580 5908 41636 6636
rect 41580 5842 41636 5852
rect 43708 5236 43764 8092
rect 43932 7476 43988 11004
rect 49532 11060 49588 13916
rect 49644 12964 49700 12974
rect 49644 11956 49700 12908
rect 49756 12292 49812 14476
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 49756 12226 49812 12236
rect 50316 13748 50372 13758
rect 50316 12516 50372 13692
rect 49644 11890 49700 11900
rect 49532 10994 49588 11004
rect 50316 11060 50372 12460
rect 50316 10994 50372 11004
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 51996 12292 52052 21756
rect 52668 21812 52724 23324
rect 53676 23380 53732 23996
rect 53676 23314 53732 23324
rect 52668 21746 52724 21756
rect 55356 21700 55412 24332
rect 55356 21634 55412 21644
rect 65888 24332 66208 25844
rect 81248 56476 81568 56508
rect 81248 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81568 56476
rect 81248 54908 81568 56420
rect 81248 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81568 54908
rect 81248 53340 81568 54852
rect 81248 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81568 53340
rect 81248 51772 81568 53284
rect 81248 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81568 51772
rect 81248 50204 81568 51716
rect 81248 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81568 50204
rect 81248 48636 81568 50148
rect 81248 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81568 48636
rect 81248 47068 81568 48580
rect 81248 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81568 47068
rect 81248 45500 81568 47012
rect 81248 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81568 45500
rect 81248 43932 81568 45444
rect 81248 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81568 43932
rect 81248 42364 81568 43876
rect 81248 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81568 42364
rect 81248 40796 81568 42308
rect 81248 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81568 40796
rect 81248 39228 81568 40740
rect 81248 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81568 39228
rect 81248 37660 81568 39172
rect 81248 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81568 37660
rect 81248 36092 81568 37604
rect 81248 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81568 36092
rect 81248 34524 81568 36036
rect 81248 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81568 34524
rect 81248 32956 81568 34468
rect 81248 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81568 32956
rect 81248 31388 81568 32900
rect 81248 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81568 31388
rect 81248 29820 81568 31332
rect 81248 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81568 29820
rect 81248 28252 81568 29764
rect 81248 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81568 28252
rect 81248 26684 81568 28196
rect 81248 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81568 26684
rect 81248 25116 81568 26628
rect 81248 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81568 25116
rect 66668 24948 66724 24958
rect 66668 24500 66724 24892
rect 66668 24434 66724 24444
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 81248 23548 81568 25060
rect 81248 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81568 23548
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 60620 21364 60676 21374
rect 57148 17444 57204 17454
rect 57148 15428 57204 17388
rect 57148 15362 57204 15372
rect 60620 12852 60676 21308
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 75180 22932 75236 22942
rect 74620 20356 74676 20366
rect 74620 20132 74676 20300
rect 74620 20066 74676 20076
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 68236 19572 68292 19582
rect 68012 19348 68068 19358
rect 68012 19012 68068 19292
rect 68012 18946 68068 18956
rect 68236 18900 68292 19516
rect 68236 18834 68292 18844
rect 75180 18228 75236 22876
rect 75180 18162 75236 18172
rect 81248 21980 81568 23492
rect 96608 55692 96928 56508
rect 96608 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96928 55692
rect 96608 54124 96928 55636
rect 96608 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96928 54124
rect 96608 52556 96928 54068
rect 96608 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96928 52556
rect 96608 50988 96928 52500
rect 96608 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96928 50988
rect 96608 49420 96928 50932
rect 96608 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96928 49420
rect 96608 47852 96928 49364
rect 96608 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96928 47852
rect 96608 46284 96928 47796
rect 96608 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96928 46284
rect 96608 44716 96928 46228
rect 96608 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96928 44716
rect 96608 43148 96928 44660
rect 96608 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96928 43148
rect 96608 41580 96928 43092
rect 96608 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96928 41580
rect 96608 40012 96928 41524
rect 96608 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96928 40012
rect 96608 38444 96928 39956
rect 96608 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96928 38444
rect 96608 36876 96928 38388
rect 96608 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96928 36876
rect 96608 35308 96928 36820
rect 96608 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96928 35308
rect 96608 33740 96928 35252
rect 96608 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96928 33740
rect 96608 32172 96928 33684
rect 96608 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96928 32172
rect 96608 30604 96928 32116
rect 96608 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96928 30604
rect 96608 29036 96928 30548
rect 96608 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96928 29036
rect 96608 27468 96928 28980
rect 96608 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96928 27468
rect 96608 25900 96928 27412
rect 96608 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96928 25900
rect 96608 24332 96928 25844
rect 96608 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96928 24332
rect 96608 22764 96928 24276
rect 96608 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96928 22764
rect 81248 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81568 21980
rect 81248 20412 81568 21924
rect 90972 22260 91028 22270
rect 81248 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81568 20412
rect 81248 18844 81568 20356
rect 89628 21364 89684 21374
rect 87948 20020 88004 20030
rect 81248 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81568 18844
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 77196 18116 77252 18126
rect 77196 16660 77252 18060
rect 77196 16594 77252 16604
rect 81248 17276 81568 18788
rect 85484 19012 85540 19022
rect 81248 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81568 17276
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 60620 12786 60676 12796
rect 61404 14532 61460 14542
rect 61404 12516 61460 14476
rect 61404 12450 61460 12460
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 81248 15708 81568 17220
rect 84364 17444 84420 17454
rect 81248 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81568 15708
rect 81248 14140 81568 15652
rect 83132 15876 83188 15886
rect 81248 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81568 14140
rect 51996 12226 52052 12236
rect 65888 11788 66208 13300
rect 72828 13300 72884 13310
rect 64652 11732 64708 11742
rect 61964 11508 62020 11518
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 46060 10836 46116 10846
rect 43932 7410 43988 7420
rect 44604 10612 44660 10622
rect 44604 10164 44660 10556
rect 43708 5170 43764 5180
rect 39340 4498 39396 4508
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 44604 3332 44660 10108
rect 46060 8260 46116 10780
rect 46060 6692 46116 8204
rect 50316 10276 50372 10286
rect 50316 7812 50372 10220
rect 50316 7746 50372 7756
rect 50528 9436 50848 10948
rect 56700 11172 56756 11182
rect 56364 9604 56420 9614
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 51996 9492 52052 9502
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 46060 6626 46116 6636
rect 44604 3266 44660 3276
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 51548 8932 51604 8942
rect 51548 3444 51604 8876
rect 51996 4340 52052 9436
rect 52108 9268 52164 9278
rect 52108 9044 52164 9212
rect 52108 8978 52164 8988
rect 52220 9156 52276 9166
rect 52220 7700 52276 9100
rect 52780 9044 52836 9054
rect 52220 7634 52276 7644
rect 52332 8484 52388 8494
rect 51996 4274 52052 4284
rect 51548 3378 51604 3388
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 52332 1652 52388 8428
rect 52332 1586 52388 1596
rect 52780 1428 52836 8988
rect 56364 9044 56420 9548
rect 56364 8978 56420 8988
rect 56028 8484 56084 8494
rect 56028 8148 56084 8428
rect 56700 8484 56756 11116
rect 61964 10948 62020 11452
rect 61964 10882 62020 10892
rect 64652 10500 64708 11676
rect 64652 10434 64708 10444
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 72268 13076 72324 13086
rect 66668 11620 66724 11630
rect 66668 11172 66724 11564
rect 66668 11106 66724 11116
rect 71708 11172 71764 11182
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 56700 8418 56756 8428
rect 61068 9716 61124 9726
rect 56028 7700 56084 8092
rect 56028 7634 56084 7644
rect 61068 3332 61124 9660
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 61964 7588 62020 7598
rect 61740 6804 61796 6814
rect 61740 5012 61796 6748
rect 61964 6244 62020 7532
rect 61964 6178 62020 6188
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 61740 4946 61796 4956
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 61068 3266 61124 3276
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
rect 71708 9044 71764 11116
rect 71708 2772 71764 8988
rect 72268 6356 72324 13020
rect 72268 6290 72324 6300
rect 71708 2706 71764 2716
rect 72268 5124 72324 5134
rect 52780 1362 52836 1372
rect 72268 1092 72324 5068
rect 72828 4228 72884 13244
rect 81248 12572 81568 14084
rect 83020 15092 83076 15102
rect 83020 13972 83076 15036
rect 83020 13906 83076 13916
rect 81248 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81568 12572
rect 75740 11172 75796 11182
rect 75740 10836 75796 11116
rect 75740 10770 75796 10780
rect 81248 11004 81568 12516
rect 81248 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81568 11004
rect 73164 10164 73220 10174
rect 72940 9268 72996 9278
rect 72940 8260 72996 9212
rect 72940 8194 72996 8204
rect 73164 6692 73220 10108
rect 73612 10164 73668 10174
rect 73276 9716 73332 9726
rect 73276 9044 73332 9660
rect 73612 9268 73668 10108
rect 73612 9202 73668 9212
rect 81248 9436 81568 10948
rect 81248 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81568 9436
rect 73276 8978 73332 8988
rect 81248 7868 81568 9380
rect 82460 10164 82516 10174
rect 82460 9156 82516 10108
rect 82460 9090 82516 9100
rect 83132 8596 83188 15820
rect 83580 15876 83636 15886
rect 83580 13972 83636 15820
rect 83580 13906 83636 13916
rect 83692 14196 83748 14206
rect 83692 11956 83748 14140
rect 83692 11890 83748 11900
rect 83916 14196 83972 14206
rect 83916 10836 83972 14140
rect 83916 10770 83972 10780
rect 84140 11620 84196 11630
rect 84140 9492 84196 11564
rect 84140 9426 84196 9436
rect 83132 8530 83188 8540
rect 84364 8036 84420 17388
rect 85148 17444 85204 17454
rect 84364 7970 84420 7980
rect 84476 15876 84532 15886
rect 81248 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81568 7868
rect 73164 6020 73220 6636
rect 73164 5954 73220 5964
rect 79436 7140 79492 7150
rect 79436 4452 79492 7084
rect 79436 4386 79492 4396
rect 81248 6300 81568 7812
rect 84476 7700 84532 15820
rect 84588 13636 84644 13646
rect 84588 9940 84644 13580
rect 85148 12068 85204 17388
rect 85484 17038 85540 18956
rect 87948 17668 88004 19964
rect 87948 17602 88004 17612
rect 88732 18788 88788 18798
rect 85148 12002 85204 12012
rect 85372 16982 85540 17038
rect 84588 9874 84644 9884
rect 84476 7634 84532 7644
rect 81248 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81568 6300
rect 81248 4732 81568 6244
rect 81248 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81568 4732
rect 72828 4162 72884 4172
rect 81248 3164 81568 4676
rect 81248 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81568 3164
rect 81248 3076 81568 3108
rect 84364 6804 84420 6814
rect 84364 2772 84420 6748
rect 85372 6804 85428 16982
rect 85484 16884 85540 16894
rect 85484 15148 85540 16828
rect 85484 15092 85652 15148
rect 85484 10948 85540 10958
rect 85484 8484 85540 10892
rect 85484 8418 85540 8428
rect 85372 6738 85428 6748
rect 85484 8036 85540 8046
rect 85596 8036 85652 15092
rect 87276 13524 87332 13534
rect 87276 12516 87332 13468
rect 88732 12964 88788 18732
rect 88732 12898 88788 12908
rect 89292 17332 89348 17342
rect 89292 12852 89348 17276
rect 89292 12786 89348 12796
rect 89628 12740 89684 21308
rect 90972 18452 91028 22204
rect 96608 21196 96928 22708
rect 96608 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96928 21196
rect 90972 18386 91028 18396
rect 94892 19684 94948 19694
rect 94444 18340 94500 18350
rect 89628 12674 89684 12684
rect 92428 16884 92484 16894
rect 87276 12450 87332 12460
rect 85708 9492 85764 9502
rect 85708 8484 85764 9436
rect 85708 8418 85764 8428
rect 86828 8484 86884 8494
rect 85540 7980 85652 8036
rect 86716 8372 86772 8382
rect 85484 4004 85540 7980
rect 86716 7700 86772 8316
rect 86716 7634 86772 7644
rect 86828 7252 86884 8428
rect 86828 7186 86884 7196
rect 92428 8260 92484 16828
rect 94444 15092 94500 18284
rect 94444 15026 94500 15036
rect 94892 15876 94948 19628
rect 96608 19628 96928 21140
rect 111968 56476 112288 56508
rect 111968 56420 111996 56476
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 112260 56420 112288 56476
rect 111968 54908 112288 56420
rect 111968 54852 111996 54908
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 112260 54852 112288 54908
rect 111968 53340 112288 54852
rect 111968 53284 111996 53340
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 112260 53284 112288 53340
rect 111968 51772 112288 53284
rect 111968 51716 111996 51772
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 112260 51716 112288 51772
rect 111968 50204 112288 51716
rect 111968 50148 111996 50204
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 112260 50148 112288 50204
rect 111968 48636 112288 50148
rect 111968 48580 111996 48636
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 112260 48580 112288 48636
rect 111968 47068 112288 48580
rect 111968 47012 111996 47068
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 112260 47012 112288 47068
rect 111968 45500 112288 47012
rect 111968 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112288 45500
rect 111968 43932 112288 45444
rect 111968 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112288 43932
rect 111968 42364 112288 43876
rect 111968 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112288 42364
rect 111968 40796 112288 42308
rect 111968 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112288 40796
rect 111968 39228 112288 40740
rect 111968 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112288 39228
rect 111968 37660 112288 39172
rect 111968 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112288 37660
rect 111968 36092 112288 37604
rect 111968 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112288 36092
rect 111968 34524 112288 36036
rect 111968 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112288 34524
rect 111968 32956 112288 34468
rect 111968 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112288 32956
rect 111968 31388 112288 32900
rect 111968 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112288 31388
rect 111968 29820 112288 31332
rect 111968 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112288 29820
rect 111968 28252 112288 29764
rect 111968 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112288 28252
rect 111968 26684 112288 28196
rect 111968 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112288 26684
rect 111968 25116 112288 26628
rect 111968 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112288 25116
rect 111968 23548 112288 25060
rect 111968 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112288 23548
rect 111968 21980 112288 23492
rect 111968 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112288 21980
rect 111968 20412 112288 21924
rect 111968 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112288 20412
rect 96608 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96928 19628
rect 96608 18060 96928 19572
rect 96608 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96928 18060
rect 94892 11844 94948 15820
rect 95004 16772 95060 16782
rect 95004 13860 95060 16716
rect 95004 13794 95060 13804
rect 96608 16492 96928 18004
rect 96608 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96928 16492
rect 96608 14924 96928 16436
rect 110124 19796 110180 19806
rect 96608 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96928 14924
rect 96608 13356 96928 14868
rect 96608 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96928 13356
rect 105756 15876 105812 15886
rect 94892 11778 94948 11788
rect 96460 12740 96516 12750
rect 96460 11844 96516 12684
rect 96460 11778 96516 11788
rect 96608 11788 96928 13300
rect 103404 13300 103460 13310
rect 85820 6132 85876 6142
rect 85820 5908 85876 6076
rect 85820 5842 85876 5852
rect 85484 3938 85540 3948
rect 84364 2706 84420 2716
rect 92428 2660 92484 8204
rect 94220 11732 94276 11742
rect 94220 5908 94276 11676
rect 96608 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96928 11788
rect 102620 12292 102676 12302
rect 102620 11844 102676 12236
rect 102620 11778 102676 11788
rect 103404 11844 103460 13244
rect 103404 11778 103460 11788
rect 96608 10220 96928 11732
rect 96608 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96928 10220
rect 96608 8652 96928 10164
rect 100940 11620 100996 11630
rect 100940 10948 100996 11564
rect 104860 11620 104916 11630
rect 97916 9156 97972 9166
rect 97916 8932 97972 9100
rect 97916 8866 97972 8876
rect 95116 8596 95172 8606
rect 95116 6020 95172 8540
rect 96608 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96928 8652
rect 95116 5954 95172 5964
rect 95676 8484 95732 8494
rect 95676 7924 95732 8428
rect 94220 5842 94276 5852
rect 92428 2594 92484 2604
rect 95676 1204 95732 7868
rect 96608 7084 96928 8596
rect 96608 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96928 7084
rect 96608 5516 96928 7028
rect 100940 5908 100996 10892
rect 102620 11284 102676 11294
rect 102620 10500 102676 11228
rect 100940 5842 100996 5852
rect 101164 10164 101220 10174
rect 96608 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96928 5516
rect 96608 3948 96928 5460
rect 96608 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96928 3948
rect 96608 3076 96928 3892
rect 101164 2436 101220 10108
rect 102620 3556 102676 10444
rect 102620 3490 102676 3500
rect 103180 11172 103236 11182
rect 101164 2370 101220 2380
rect 103180 1652 103236 11116
rect 104748 11060 104804 11070
rect 104748 10388 104804 11004
rect 104748 10322 104804 10332
rect 104860 6804 104916 11564
rect 104860 6738 104916 6748
rect 105756 4452 105812 15820
rect 109900 12068 109956 12078
rect 106092 10724 106148 10734
rect 106092 6244 106148 10668
rect 109900 9380 109956 12012
rect 109900 9314 109956 9324
rect 106092 6178 106148 6188
rect 108556 8372 108612 8382
rect 108556 4676 108612 8316
rect 110124 5236 110180 19740
rect 111968 18844 112288 20356
rect 111968 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112288 18844
rect 111968 17276 112288 18788
rect 111968 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112288 17276
rect 111968 15708 112288 17220
rect 111968 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112288 15708
rect 111968 14140 112288 15652
rect 111968 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112288 14140
rect 111968 12572 112288 14084
rect 111968 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112288 12572
rect 111968 11004 112288 12516
rect 127328 55692 127648 56508
rect 127328 55636 127356 55692
rect 127412 55636 127460 55692
rect 127516 55636 127564 55692
rect 127620 55636 127648 55692
rect 127328 54124 127648 55636
rect 127328 54068 127356 54124
rect 127412 54068 127460 54124
rect 127516 54068 127564 54124
rect 127620 54068 127648 54124
rect 127328 52556 127648 54068
rect 127328 52500 127356 52556
rect 127412 52500 127460 52556
rect 127516 52500 127564 52556
rect 127620 52500 127648 52556
rect 127328 50988 127648 52500
rect 127328 50932 127356 50988
rect 127412 50932 127460 50988
rect 127516 50932 127564 50988
rect 127620 50932 127648 50988
rect 127328 49420 127648 50932
rect 127328 49364 127356 49420
rect 127412 49364 127460 49420
rect 127516 49364 127564 49420
rect 127620 49364 127648 49420
rect 127328 47852 127648 49364
rect 127328 47796 127356 47852
rect 127412 47796 127460 47852
rect 127516 47796 127564 47852
rect 127620 47796 127648 47852
rect 127328 46284 127648 47796
rect 127328 46228 127356 46284
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127620 46228 127648 46284
rect 127328 44716 127648 46228
rect 127328 44660 127356 44716
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127620 44660 127648 44716
rect 127328 43148 127648 44660
rect 127328 43092 127356 43148
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127620 43092 127648 43148
rect 127328 41580 127648 43092
rect 127328 41524 127356 41580
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127620 41524 127648 41580
rect 127328 40012 127648 41524
rect 127328 39956 127356 40012
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127620 39956 127648 40012
rect 127328 38444 127648 39956
rect 127328 38388 127356 38444
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127620 38388 127648 38444
rect 127328 36876 127648 38388
rect 127328 36820 127356 36876
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127620 36820 127648 36876
rect 127328 35308 127648 36820
rect 127328 35252 127356 35308
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127620 35252 127648 35308
rect 127328 33740 127648 35252
rect 127328 33684 127356 33740
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127620 33684 127648 33740
rect 127328 32172 127648 33684
rect 127328 32116 127356 32172
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127620 32116 127648 32172
rect 127328 30604 127648 32116
rect 127328 30548 127356 30604
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127620 30548 127648 30604
rect 127328 29036 127648 30548
rect 127328 28980 127356 29036
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127620 28980 127648 29036
rect 127328 27468 127648 28980
rect 127328 27412 127356 27468
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127620 27412 127648 27468
rect 127328 25900 127648 27412
rect 127328 25844 127356 25900
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127620 25844 127648 25900
rect 127328 24332 127648 25844
rect 127328 24276 127356 24332
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127620 24276 127648 24332
rect 127328 22764 127648 24276
rect 127328 22708 127356 22764
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127620 22708 127648 22764
rect 127328 21196 127648 22708
rect 127328 21140 127356 21196
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127620 21140 127648 21196
rect 127328 19628 127648 21140
rect 127328 19572 127356 19628
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127620 19572 127648 19628
rect 127328 18060 127648 19572
rect 127328 18004 127356 18060
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127620 18004 127648 18060
rect 127328 16492 127648 18004
rect 127328 16436 127356 16492
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127620 16436 127648 16492
rect 127328 14924 127648 16436
rect 127328 14868 127356 14924
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127620 14868 127648 14924
rect 127328 13356 127648 14868
rect 127328 13300 127356 13356
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127620 13300 127648 13356
rect 127328 11788 127648 13300
rect 127328 11732 127356 11788
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127620 11732 127648 11788
rect 111968 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112288 11004
rect 111968 9436 112288 10948
rect 111968 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112288 9436
rect 110908 8596 110964 8606
rect 110908 7924 110964 8540
rect 110908 7858 110964 7868
rect 111356 8260 111412 8270
rect 110124 5170 110180 5180
rect 111356 5236 111412 8204
rect 111356 5170 111412 5180
rect 111968 7868 112288 9380
rect 111968 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112288 7868
rect 111968 6300 112288 7812
rect 111968 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112288 6300
rect 112364 11284 112420 11294
rect 112364 6356 112420 11228
rect 115948 10276 116004 10286
rect 112924 9380 112980 9390
rect 112924 8372 112980 9324
rect 112924 8306 112980 8316
rect 112364 6290 112420 6300
rect 115052 7140 115108 7150
rect 108556 4610 108612 4620
rect 111968 4732 112288 6244
rect 111968 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112288 4732
rect 105756 4386 105812 4396
rect 111968 3164 112288 4676
rect 115052 4228 115108 7084
rect 115948 5684 116004 10220
rect 115948 4900 116004 5628
rect 115948 4834 116004 4844
rect 127328 10220 127648 11732
rect 127328 10164 127356 10220
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127620 10164 127648 10220
rect 127328 8652 127648 10164
rect 127328 8596 127356 8652
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127620 8596 127648 8652
rect 127328 7084 127648 8596
rect 127328 7028 127356 7084
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127620 7028 127648 7084
rect 127328 5516 127648 7028
rect 127328 5460 127356 5516
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127620 5460 127648 5516
rect 115052 4162 115108 4172
rect 111968 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112288 3164
rect 111968 3076 112288 3108
rect 127328 3948 127648 5460
rect 127328 3892 127356 3948
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127620 3892 127648 3948
rect 127328 3076 127648 3892
rect 142688 56476 143008 56508
rect 142688 56420 142716 56476
rect 142772 56420 142820 56476
rect 142876 56420 142924 56476
rect 142980 56420 143008 56476
rect 142688 54908 143008 56420
rect 142688 54852 142716 54908
rect 142772 54852 142820 54908
rect 142876 54852 142924 54908
rect 142980 54852 143008 54908
rect 142688 53340 143008 54852
rect 142688 53284 142716 53340
rect 142772 53284 142820 53340
rect 142876 53284 142924 53340
rect 142980 53284 143008 53340
rect 142688 51772 143008 53284
rect 142688 51716 142716 51772
rect 142772 51716 142820 51772
rect 142876 51716 142924 51772
rect 142980 51716 143008 51772
rect 142688 50204 143008 51716
rect 142688 50148 142716 50204
rect 142772 50148 142820 50204
rect 142876 50148 142924 50204
rect 142980 50148 143008 50204
rect 142688 48636 143008 50148
rect 142688 48580 142716 48636
rect 142772 48580 142820 48636
rect 142876 48580 142924 48636
rect 142980 48580 143008 48636
rect 142688 47068 143008 48580
rect 142688 47012 142716 47068
rect 142772 47012 142820 47068
rect 142876 47012 142924 47068
rect 142980 47012 143008 47068
rect 142688 45500 143008 47012
rect 142688 45444 142716 45500
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142980 45444 143008 45500
rect 142688 43932 143008 45444
rect 142688 43876 142716 43932
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142980 43876 143008 43932
rect 142688 42364 143008 43876
rect 142688 42308 142716 42364
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142980 42308 143008 42364
rect 142688 40796 143008 42308
rect 142688 40740 142716 40796
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142980 40740 143008 40796
rect 142688 39228 143008 40740
rect 142688 39172 142716 39228
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142980 39172 143008 39228
rect 142688 37660 143008 39172
rect 142688 37604 142716 37660
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142980 37604 143008 37660
rect 142688 36092 143008 37604
rect 142688 36036 142716 36092
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142980 36036 143008 36092
rect 142688 34524 143008 36036
rect 142688 34468 142716 34524
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142980 34468 143008 34524
rect 142688 32956 143008 34468
rect 142688 32900 142716 32956
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142980 32900 143008 32956
rect 142688 31388 143008 32900
rect 142688 31332 142716 31388
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142980 31332 143008 31388
rect 142688 29820 143008 31332
rect 142688 29764 142716 29820
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142980 29764 143008 29820
rect 142688 28252 143008 29764
rect 142688 28196 142716 28252
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142980 28196 143008 28252
rect 142688 26684 143008 28196
rect 142688 26628 142716 26684
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142980 26628 143008 26684
rect 142688 25116 143008 26628
rect 142688 25060 142716 25116
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142980 25060 143008 25116
rect 142688 23548 143008 25060
rect 142688 23492 142716 23548
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142980 23492 143008 23548
rect 142688 21980 143008 23492
rect 142688 21924 142716 21980
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142980 21924 143008 21980
rect 142688 20412 143008 21924
rect 142688 20356 142716 20412
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142980 20356 143008 20412
rect 142688 18844 143008 20356
rect 142688 18788 142716 18844
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142980 18788 143008 18844
rect 142688 17276 143008 18788
rect 142688 17220 142716 17276
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142980 17220 143008 17276
rect 142688 15708 143008 17220
rect 142688 15652 142716 15708
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142980 15652 143008 15708
rect 142688 14140 143008 15652
rect 142688 14084 142716 14140
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142980 14084 143008 14140
rect 142688 12572 143008 14084
rect 142688 12516 142716 12572
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142980 12516 143008 12572
rect 142688 11004 143008 12516
rect 142688 10948 142716 11004
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142980 10948 143008 11004
rect 142688 9436 143008 10948
rect 142688 9380 142716 9436
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142980 9380 143008 9436
rect 142688 7868 143008 9380
rect 142688 7812 142716 7868
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142980 7812 143008 7868
rect 142688 6300 143008 7812
rect 142688 6244 142716 6300
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142980 6244 143008 6300
rect 142688 4732 143008 6244
rect 142688 4676 142716 4732
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142980 4676 143008 4732
rect 142688 3164 143008 4676
rect 142688 3108 142716 3164
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142980 3108 143008 3164
rect 142688 3076 143008 3108
rect 158048 55692 158368 56508
rect 158048 55636 158076 55692
rect 158132 55636 158180 55692
rect 158236 55636 158284 55692
rect 158340 55636 158368 55692
rect 158048 54124 158368 55636
rect 158048 54068 158076 54124
rect 158132 54068 158180 54124
rect 158236 54068 158284 54124
rect 158340 54068 158368 54124
rect 158048 52556 158368 54068
rect 158048 52500 158076 52556
rect 158132 52500 158180 52556
rect 158236 52500 158284 52556
rect 158340 52500 158368 52556
rect 158048 50988 158368 52500
rect 158048 50932 158076 50988
rect 158132 50932 158180 50988
rect 158236 50932 158284 50988
rect 158340 50932 158368 50988
rect 158048 49420 158368 50932
rect 158048 49364 158076 49420
rect 158132 49364 158180 49420
rect 158236 49364 158284 49420
rect 158340 49364 158368 49420
rect 158048 47852 158368 49364
rect 158048 47796 158076 47852
rect 158132 47796 158180 47852
rect 158236 47796 158284 47852
rect 158340 47796 158368 47852
rect 158048 46284 158368 47796
rect 158048 46228 158076 46284
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158340 46228 158368 46284
rect 158048 44716 158368 46228
rect 158048 44660 158076 44716
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158340 44660 158368 44716
rect 158048 43148 158368 44660
rect 158048 43092 158076 43148
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158340 43092 158368 43148
rect 158048 41580 158368 43092
rect 158048 41524 158076 41580
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158340 41524 158368 41580
rect 158048 40012 158368 41524
rect 158048 39956 158076 40012
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158340 39956 158368 40012
rect 158048 38444 158368 39956
rect 158048 38388 158076 38444
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158340 38388 158368 38444
rect 158048 36876 158368 38388
rect 158048 36820 158076 36876
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158340 36820 158368 36876
rect 158048 35308 158368 36820
rect 158048 35252 158076 35308
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158340 35252 158368 35308
rect 158048 33740 158368 35252
rect 158048 33684 158076 33740
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158340 33684 158368 33740
rect 158048 32172 158368 33684
rect 158048 32116 158076 32172
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158340 32116 158368 32172
rect 158048 30604 158368 32116
rect 158048 30548 158076 30604
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158340 30548 158368 30604
rect 158048 29036 158368 30548
rect 158048 28980 158076 29036
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158340 28980 158368 29036
rect 158048 27468 158368 28980
rect 158048 27412 158076 27468
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158340 27412 158368 27468
rect 158048 25900 158368 27412
rect 158048 25844 158076 25900
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158340 25844 158368 25900
rect 158048 24332 158368 25844
rect 158048 24276 158076 24332
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158340 24276 158368 24332
rect 158048 22764 158368 24276
rect 158048 22708 158076 22764
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158340 22708 158368 22764
rect 158048 21196 158368 22708
rect 158048 21140 158076 21196
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158340 21140 158368 21196
rect 158048 19628 158368 21140
rect 158048 19572 158076 19628
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158340 19572 158368 19628
rect 158048 18060 158368 19572
rect 158048 18004 158076 18060
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158340 18004 158368 18060
rect 158048 16492 158368 18004
rect 158048 16436 158076 16492
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158340 16436 158368 16492
rect 158048 14924 158368 16436
rect 158048 14868 158076 14924
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158340 14868 158368 14924
rect 158048 13356 158368 14868
rect 158048 13300 158076 13356
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158340 13300 158368 13356
rect 158048 11788 158368 13300
rect 158048 11732 158076 11788
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158340 11732 158368 11788
rect 158048 10220 158368 11732
rect 158048 10164 158076 10220
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158340 10164 158368 10220
rect 158048 8652 158368 10164
rect 158048 8596 158076 8652
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158340 8596 158368 8652
rect 158048 7084 158368 8596
rect 158048 7028 158076 7084
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158340 7028 158368 7084
rect 158048 5516 158368 7028
rect 158048 5460 158076 5516
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158340 5460 158368 5516
rect 158048 3948 158368 5460
rect 158048 3892 158076 3948
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158340 3892 158368 3948
rect 158048 3076 158368 3892
rect 103180 1586 103236 1596
rect 95676 1138 95732 1148
rect 72268 1026 72324 1036
rect 31612 802 31668 812
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _0972_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19824 0 -1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0973_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 72576 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0974_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 73696 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0975_
timestamp 1698431365
transform -1 0 73136 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0976_
timestamp 1698431365
transform -1 0 28784 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0977_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 54768 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0978_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 53760 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0979_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 55552 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0980_
timestamp 1698431365
transform 1 0 55552 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0981_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 55552 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0982_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 53760 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0983_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28672 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0984_
timestamp 1698431365
transform 1 0 54880 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0985_
timestamp 1698431365
transform 1 0 58352 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0986_
timestamp 1698431365
transform 1 0 59248 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0987_
timestamp 1698431365
transform 1 0 60368 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0988_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 59248 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0989_
timestamp 1698431365
transform 1 0 60368 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0990_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 59136 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0991_
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0992_
timestamp 1698431365
transform 1 0 55104 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0993_
timestamp 1698431365
transform 1 0 57568 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0994_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 61488 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0995_
timestamp 1698431365
transform -1 0 61488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0996_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 62720 0 -1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0997_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15232 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0998_
timestamp 1698431365
transform 1 0 38304 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0999_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 138096 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1000_
timestamp 1698431365
transform 1 0 138768 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1001_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 142352 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1002_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 126784 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1003_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 90384 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1004_
timestamp 1698431365
transform 1 0 91056 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1005_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 94640 0 -1 7840
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1006_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 93408 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1007_
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1008_
timestamp 1698431365
transform 1 0 47824 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1009_
timestamp 1698431365
transform 1 0 47712 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1010_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15232 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1011_
timestamp 1698431365
transform 1 0 38640 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1012_
timestamp 1698431365
transform 1 0 92960 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1013_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 93296 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1014_
timestamp 1698431365
transform 1 0 91056 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1015_
timestamp 1698431365
transform -1 0 95424 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1016_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 95984 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1017_
timestamp 1698431365
transform -1 0 40544 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _1018_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44464 0 1 4704
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1019_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29344 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1020_
timestamp 1698431365
transform -1 0 42560 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1021_
timestamp 1698431365
transform 1 0 33712 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1022_
timestamp 1698431365
transform 1 0 38080 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1023_
timestamp 1698431365
transform 1 0 68208 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1024_
timestamp 1698431365
transform -1 0 67984 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1025_
timestamp 1698431365
transform -1 0 66192 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1026_
timestamp 1698431365
transform 1 0 64288 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1027_
timestamp 1698431365
transform 1 0 39424 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1028_
timestamp 1698431365
transform -1 0 38640 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1029_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37520 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1030_
timestamp 1698431365
transform -1 0 36624 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1031_
timestamp 1698431365
transform 1 0 33040 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1032_
timestamp 1698431365
transform 1 0 31360 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1033_
timestamp 1698431365
transform -1 0 38304 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1034_
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1035_
timestamp 1698431365
transform -1 0 53648 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1036_
timestamp 1698431365
transform -1 0 73920 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1037_
timestamp 1698431365
transform -1 0 68432 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1038_
timestamp 1698431365
transform -1 0 52304 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1039_
timestamp 1698431365
transform 1 0 27888 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1040_
timestamp 1698431365
transform -1 0 33600 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1041_
timestamp 1698431365
transform -1 0 39424 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1042_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 93520 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1043_
timestamp 1698431365
transform -1 0 95648 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1044_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 91280 0 -1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1045_
timestamp 1698431365
transform 1 0 89600 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1046_
timestamp 1698431365
transform -1 0 91280 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1047_
timestamp 1698431365
transform -1 0 39312 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1048_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40544 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1049_
timestamp 1698431365
transform -1 0 38080 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1050_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41552 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1051_
timestamp 1698431365
transform -1 0 40880 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1052_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34720 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1053_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 103488 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1054_
timestamp 1698431365
transform -1 0 37744 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1055_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33040 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1056_
timestamp 1698431365
transform 1 0 29120 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1057_
timestamp 1698431365
transform 1 0 29568 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1058_
timestamp 1698431365
transform 1 0 35840 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1059_
timestamp 1698431365
transform -1 0 91728 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1060_
timestamp 1698431365
transform 1 0 30128 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1061_
timestamp 1698431365
transform -1 0 38416 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1062_
timestamp 1698431365
transform -1 0 38192 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1063_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30240 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1064_
timestamp 1698431365
transform -1 0 34384 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1065_
timestamp 1698431365
transform 1 0 27440 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1066_
timestamp 1698431365
transform -1 0 92736 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1067_
timestamp 1698431365
transform 1 0 30128 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1068_
timestamp 1698431365
transform 1 0 29232 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1069_
timestamp 1698431365
transform -1 0 32144 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1070_
timestamp 1698431365
transform 1 0 29344 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1071_
timestamp 1698431365
transform 1 0 88592 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1072_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30240 0 1 7840
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1073_
timestamp 1698431365
transform 1 0 34832 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1074_
timestamp 1698431365
transform -1 0 36512 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1075_
timestamp 1698431365
transform 1 0 38864 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1076_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 50736 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1077_
timestamp 1698431365
transform -1 0 49504 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1078_
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1079_
timestamp 1698431365
transform -1 0 43904 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1080_
timestamp 1698431365
transform -1 0 42448 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1081_
timestamp 1698431365
transform 1 0 45808 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1082_
timestamp 1698431365
transform 1 0 45696 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1083_
timestamp 1698431365
transform -1 0 47152 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1084_
timestamp 1698431365
transform 1 0 48160 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1085_
timestamp 1698431365
transform -1 0 49840 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1086_
timestamp 1698431365
transform 1 0 49168 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1087_
timestamp 1698431365
transform 1 0 49840 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1088_
timestamp 1698431365
transform -1 0 75152 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1089_
timestamp 1698431365
transform 1 0 72128 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1090_
timestamp 1698431365
transform -1 0 77952 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1091_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 76832 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1092_
timestamp 1698431365
transform 1 0 73920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1093_
timestamp 1698431365
transform -1 0 78960 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1094_
timestamp 1698431365
transform 1 0 77952 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1095_
timestamp 1698431365
transform 1 0 76272 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1096_
timestamp 1698431365
transform -1 0 79296 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1097_
timestamp 1698431365
transform -1 0 79968 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1098_
timestamp 1698431365
transform 1 0 77952 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1099_
timestamp 1698431365
transform 1 0 81312 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1100_
timestamp 1698431365
transform -1 0 86016 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1101_
timestamp 1698431365
transform 1 0 81760 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1102_
timestamp 1698431365
transform -1 0 80416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1103_
timestamp 1698431365
transform -1 0 77952 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1104_
timestamp 1698431365
transform -1 0 82880 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1105_
timestamp 1698431365
transform -1 0 82768 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1106_
timestamp 1698431365
transform 1 0 84112 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1107_
timestamp 1698431365
transform 1 0 101024 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1108_
timestamp 1698431365
transform 1 0 102368 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1109_
timestamp 1698431365
transform -1 0 86128 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1110_
timestamp 1698431365
transform 1 0 98000 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1111_
timestamp 1698431365
transform 1 0 102368 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1112_
timestamp 1698431365
transform -1 0 103488 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1113_
timestamp 1698431365
transform 1 0 103488 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1114_
timestamp 1698431365
transform 1 0 97552 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1115_
timestamp 1698431365
transform 1 0 100576 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1116_
timestamp 1698431365
transform 1 0 98112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1117_
timestamp 1698431365
transform 1 0 99568 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1118_
timestamp 1698431365
transform 1 0 98896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1119_
timestamp 1698431365
transform 1 0 105168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1120_
timestamp 1698431365
transform 1 0 108976 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1121_
timestamp 1698431365
transform 1 0 102816 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1122_
timestamp 1698431365
transform 1 0 111328 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1123_
timestamp 1698431365
transform -1 0 106960 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1124_
timestamp 1698431365
transform 1 0 105392 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1125_
timestamp 1698431365
transform -1 0 108976 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1126_
timestamp 1698431365
transform -1 0 105392 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1127_
timestamp 1698431365
transform -1 0 106848 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1128_
timestamp 1698431365
transform 1 0 105168 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1129_
timestamp 1698431365
transform 1 0 110656 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1130_
timestamp 1698431365
transform -1 0 118720 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1131_
timestamp 1698431365
transform 1 0 114800 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1132_
timestamp 1698431365
transform 1 0 111440 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1133_
timestamp 1698431365
transform -1 0 120736 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1134_
timestamp 1698431365
transform 1 0 113904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1135_
timestamp 1698431365
transform -1 0 118944 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1136_
timestamp 1698431365
transform 1 0 115472 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1137_
timestamp 1698431365
transform -1 0 118160 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1138_
timestamp 1698431365
transform 1 0 112224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1139_
timestamp 1698431365
transform 1 0 109312 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1140_
timestamp 1698431365
transform -1 0 117152 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1141_
timestamp 1698431365
transform 1 0 110544 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1142_
timestamp 1698431365
transform 1 0 111328 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1143_
timestamp 1698431365
transform -1 0 114912 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1144_
timestamp 1698431365
transform 1 0 111328 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1145_
timestamp 1698431365
transform -1 0 115024 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1146_
timestamp 1698431365
transform 1 0 110096 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1147_
timestamp 1698431365
transform -1 0 114240 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1148_
timestamp 1698431365
transform 1 0 107632 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1149_
timestamp 1698431365
transform -1 0 112112 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1150_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 93072 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1151_
timestamp 1698431365
transform -1 0 63952 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1152_
timestamp 1698431365
transform 1 0 56896 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1153_
timestamp 1698431365
transform -1 0 64064 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1154_
timestamp 1698431365
transform -1 0 67312 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1155_
timestamp 1698431365
transform -1 0 61600 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1156_
timestamp 1698431365
transform -1 0 62384 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1157_
timestamp 1698431365
transform 1 0 61712 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1158_
timestamp 1698431365
transform 1 0 81200 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1159_
timestamp 1698431365
transform 1 0 86016 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1160_
timestamp 1698431365
transform 1 0 58688 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1161_
timestamp 1698431365
transform 1 0 60592 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1162_
timestamp 1698431365
transform 1 0 77728 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1163_
timestamp 1698431365
transform 1 0 86688 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1164_
timestamp 1698431365
transform -1 0 57568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1165_
timestamp 1698431365
transform 1 0 61824 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1166_
timestamp 1698431365
transform -1 0 61824 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1167_
timestamp 1698431365
transform 1 0 56112 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1168_
timestamp 1698431365
transform 1 0 57232 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1169_
timestamp 1698431365
transform 1 0 60480 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1170_
timestamp 1698431365
transform 1 0 61264 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1171_
timestamp 1698431365
transform -1 0 66304 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1172_
timestamp 1698431365
transform 1 0 65184 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1173_
timestamp 1698431365
transform 1 0 57456 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1174_
timestamp 1698431365
transform 1 0 58912 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1175_
timestamp 1698431365
transform -1 0 91504 0 1 9408
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1176_
timestamp 1698431365
transform 1 0 60368 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1177_
timestamp 1698431365
transform 1 0 61264 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1178_
timestamp 1698431365
transform -1 0 85008 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1179_
timestamp 1698431365
transform 1 0 64512 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1180_
timestamp 1698431365
transform -1 0 61264 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1181_
timestamp 1698431365
transform 1 0 64176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1182_
timestamp 1698431365
transform 1 0 65408 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1183_
timestamp 1698431365
transform -1 0 68432 0 -1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1184_
timestamp 1698431365
transform -1 0 77728 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1185_
timestamp 1698431365
transform 1 0 76048 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1186_
timestamp 1698431365
transform 1 0 74368 0 -1 12544
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1187_
timestamp 1698431365
transform -1 0 54880 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1188_
timestamp 1698431365
transform -1 0 57568 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1189_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 54992 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1190_
timestamp 1698431365
transform 1 0 60592 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1191_
timestamp 1698431365
transform 1 0 91952 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1192_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 86576 0 1 15680
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1193_
timestamp 1698431365
transform 1 0 57568 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1194_
timestamp 1698431365
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1195_
timestamp 1698431365
transform -1 0 92400 0 -1 10976
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1196_
timestamp 1698431365
transform -1 0 75712 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1197_
timestamp 1698431365
transform 1 0 75040 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1198_
timestamp 1698431365
transform 1 0 74592 0 -1 14112
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1199_
timestamp 1698431365
transform 1 0 86464 0 1 14112
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1200_
timestamp 1698431365
transform 1 0 95424 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1201_
timestamp 1698431365
transform 1 0 94304 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1202_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 60704 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1203_
timestamp 1698431365
transform 1 0 95648 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1204_
timestamp 1698431365
transform 1 0 95648 0 -1 10976
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1205_
timestamp 1698431365
transform 1 0 56784 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1206_
timestamp 1698431365
transform -1 0 82880 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1207_
timestamp 1698431365
transform -1 0 77616 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1208_
timestamp 1698431365
transform -1 0 79520 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1209_
timestamp 1698431365
transform -1 0 81312 0 1 14112
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1210_
timestamp 1698431365
transform 1 0 92736 0 1 14112
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1211_
timestamp 1698431365
transform 1 0 58240 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1212_
timestamp 1698431365
transform 1 0 82096 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1213_
timestamp 1698431365
transform 1 0 76832 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1214_
timestamp 1698431365
transform 1 0 83888 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1215_
timestamp 1698431365
transform 1 0 83888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1216_
timestamp 1698431365
transform -1 0 88592 0 1 12544
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1217_
timestamp 1698431365
transform -1 0 90608 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1218_
timestamp 1698431365
transform 1 0 88480 0 -1 14112
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1219_
timestamp 1698431365
transform 1 0 93744 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1220_
timestamp 1698431365
transform -1 0 85904 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1221_
timestamp 1698431365
transform 1 0 84784 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1222_
timestamp 1698431365
transform -1 0 88816 0 1 10976
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1223_
timestamp 1698431365
transform -1 0 90832 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1224_
timestamp 1698431365
transform 1 0 94192 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1225_
timestamp 1698431365
transform 1 0 94192 0 1 12544
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1226_
timestamp 1698431365
transform 1 0 66080 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1227_
timestamp 1698431365
transform 1 0 97104 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1228_
timestamp 1698431365
transform 1 0 96096 0 -1 9408
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1229_
timestamp 1698431365
transform -1 0 67088 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1230_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 80976 0 -1 14112
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1231_
timestamp 1698431365
transform 1 0 95648 0 -1 12544
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1232_
timestamp 1698431365
transform -1 0 86912 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1233_
timestamp 1698431365
transform 1 0 95648 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1234_
timestamp 1698431365
transform 1 0 94864 0 1 9408
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1235_
timestamp 1698431365
transform 1 0 64288 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1236_
timestamp 1698431365
transform 1 0 79968 0 -1 12544
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1237_
timestamp 1698431365
transform 1 0 95648 0 -1 15680
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1238_
timestamp 1698431365
transform -1 0 85232 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1239_
timestamp 1698431365
transform 1 0 94976 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1240_
timestamp 1698431365
transform 1 0 96096 0 -1 7840
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1241_
timestamp 1698431365
transform -1 0 43344 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1242_
timestamp 1698431365
transform -1 0 38864 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1243_
timestamp 1698431365
transform 1 0 43344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1244_
timestamp 1698431365
transform 1 0 78400 0 1 12544
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1245_
timestamp 1698431365
transform 1 0 95648 0 -1 14112
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1246_
timestamp 1698431365
transform 1 0 49840 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_4  _1247_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 49728 0 -1 7840
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1248_
timestamp 1698431365
transform 1 0 60368 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1249_
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1250_
timestamp 1698431365
transform 1 0 57568 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1251_
timestamp 1698431365
transform -1 0 73472 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1252_
timestamp 1698431365
transform 1 0 63840 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1253_
timestamp 1698431365
transform -1 0 71904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1254_
timestamp 1698431365
transform 1 0 65184 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1255_
timestamp 1698431365
transform 1 0 64512 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1256_
timestamp 1698431365
transform -1 0 73808 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1257_
timestamp 1698431365
transform 1 0 67312 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1258_
timestamp 1698431365
transform 1 0 66864 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1259_
timestamp 1698431365
transform 1 0 68208 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1260_
timestamp 1698431365
transform 1 0 57456 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1261_
timestamp 1698431365
transform -1 0 74592 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1262_
timestamp 1698431365
transform 1 0 72464 0 1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1263_
timestamp 1698431365
transform 1 0 108528 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1264_
timestamp 1698431365
transform -1 0 54544 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1265_
timestamp 1698431365
transform -1 0 54880 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1266_
timestamp 1698431365
transform 1 0 64288 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1267_
timestamp 1698431365
transform -1 0 77952 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1268_
timestamp 1698431365
transform 1 0 73472 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1269_
timestamp 1698431365
transform 1 0 108080 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1270_
timestamp 1698431365
transform 1 0 73136 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1271_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 112784 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1272_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 113680 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1273_
timestamp 1698431365
transform -1 0 78400 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1274_
timestamp 1698431365
transform 1 0 109648 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1275_
timestamp 1698431365
transform 1 0 108752 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1276_
timestamp 1698431365
transform 1 0 87472 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1277_
timestamp 1698431365
transform -1 0 90048 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1278_
timestamp 1698431365
transform 1 0 112560 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1279_
timestamp 1698431365
transform 1 0 111664 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1280_
timestamp 1698431365
transform -1 0 101584 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1281_
timestamp 1698431365
transform 1 0 105952 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1282_
timestamp 1698431365
transform -1 0 110096 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1283_
timestamp 1698431365
transform 1 0 108864 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1284_
timestamp 1698431365
transform -1 0 106400 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1285_
timestamp 1698431365
transform -1 0 107184 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1286_
timestamp 1698431365
transform 1 0 106288 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1287_
timestamp 1698431365
transform 1 0 108640 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1288_
timestamp 1698431365
transform 1 0 106288 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1289_
timestamp 1698431365
transform -1 0 108416 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1290_
timestamp 1698431365
transform 1 0 107744 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1291_
timestamp 1698431365
transform -1 0 108640 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1292_
timestamp 1698431365
transform -1 0 87248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1293_
timestamp 1698431365
transform -1 0 106736 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1294_
timestamp 1698431365
transform 1 0 107408 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1295_
timestamp 1698431365
transform 1 0 106064 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1296_
timestamp 1698431365
transform -1 0 105728 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1297_
timestamp 1698431365
transform -1 0 104720 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1298_
timestamp 1698431365
transform -1 0 106288 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1299_
timestamp 1698431365
transform 1 0 104496 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1300_
timestamp 1698431365
transform 1 0 72464 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1301_
timestamp 1698431365
transform 1 0 68656 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1302_
timestamp 1698431365
transform 1 0 74032 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1303_
timestamp 1698431365
transform -1 0 75376 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1304_
timestamp 1698431365
transform -1 0 87136 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1305_
timestamp 1698431365
transform 1 0 86688 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1306_
timestamp 1698431365
transform 1 0 93632 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1307_
timestamp 1698431365
transform 1 0 92848 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1308_
timestamp 1698431365
transform 1 0 92624 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1309_
timestamp 1698431365
transform 1 0 91728 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1310_
timestamp 1698431365
transform 1 0 91728 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1311_
timestamp 1698431365
transform 1 0 90496 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1312_
timestamp 1698431365
transform 1 0 76608 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1313_
timestamp 1698431365
transform -1 0 87584 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1314_
timestamp 1698431365
transform -1 0 88704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1315_
timestamp 1698431365
transform 1 0 86240 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1316_
timestamp 1698431365
transform -1 0 86688 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1317_
timestamp 1698431365
transform 1 0 86800 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1318_
timestamp 1698431365
transform 1 0 86016 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1319_
timestamp 1698431365
transform -1 0 86128 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1320_
timestamp 1698431365
transform -1 0 88256 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1321_
timestamp 1698431365
transform -1 0 88480 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1322_
timestamp 1698431365
transform 1 0 86464 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1323_
timestamp 1698431365
transform 1 0 85904 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1324_
timestamp 1698431365
transform -1 0 93296 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1325_
timestamp 1698431365
transform 1 0 91392 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1326_
timestamp 1698431365
transform 1 0 90608 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1327_
timestamp 1698431365
transform 1 0 69104 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1328_
timestamp 1698431365
transform 1 0 68880 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1329_
timestamp 1698431365
transform -1 0 73696 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1330_
timestamp 1698431365
transform -1 0 76048 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1331_
timestamp 1698431365
transform 1 0 95648 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1332_
timestamp 1698431365
transform 1 0 95872 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1333_
timestamp 1698431365
transform -1 0 98448 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1334_
timestamp 1698431365
transform 1 0 97664 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1335_
timestamp 1698431365
transform 1 0 97216 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1336_
timestamp 1698431365
transform 1 0 96320 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1337_
timestamp 1698431365
transform 1 0 96544 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1338_
timestamp 1698431365
transform 1 0 95648 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1339_
timestamp 1698431365
transform 1 0 93744 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1340_
timestamp 1698431365
transform 1 0 97216 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1341_
timestamp 1698431365
transform 1 0 96320 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1342_
timestamp 1698431365
transform 1 0 99904 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1343_
timestamp 1698431365
transform 1 0 99680 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1344_
timestamp 1698431365
transform 1 0 100464 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1345_
timestamp 1698431365
transform 1 0 99904 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1346_
timestamp 1698431365
transform -1 0 101920 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1347_
timestamp 1698431365
transform 1 0 103488 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1348_
timestamp 1698431365
transform 1 0 101920 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1349_
timestamp 1698431365
transform 1 0 101248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1350_
timestamp 1698431365
transform 1 0 92400 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1351_
timestamp 1698431365
transform -1 0 101248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1352_
timestamp 1698431365
transform -1 0 102144 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1353_
timestamp 1698431365
transform -1 0 46816 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1354_
timestamp 1698431365
transform -1 0 46032 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1355_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40992 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1356_
timestamp 1698431365
transform -1 0 57904 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1357_
timestamp 1698431365
transform 1 0 45024 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1358_
timestamp 1698431365
transform -1 0 48384 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1359_
timestamp 1698431365
transform 1 0 48384 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1360_
timestamp 1698431365
transform 1 0 73472 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1361_
timestamp 1698431365
transform -1 0 75488 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1362_
timestamp 1698431365
transform -1 0 71568 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1363_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48272 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1364_
timestamp 1698431365
transform 1 0 50400 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1365_
timestamp 1698431365
transform 1 0 61600 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1366_
timestamp 1698431365
transform -1 0 62944 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1367_
timestamp 1698431365
transform 1 0 61488 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1368_
timestamp 1698431365
transform -1 0 69888 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1369_
timestamp 1698431365
transform -1 0 69216 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1370_
timestamp 1698431365
transform 1 0 65744 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1371_
timestamp 1698431365
transform 1 0 69104 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1372_
timestamp 1698431365
transform 1 0 61152 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1373_
timestamp 1698431365
transform 1 0 63056 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1374_
timestamp 1698431365
transform 1 0 49504 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1375_
timestamp 1698431365
transform -1 0 88480 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1376_
timestamp 1698431365
transform 1 0 76048 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1377_
timestamp 1698431365
transform 1 0 72912 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1378_
timestamp 1698431365
transform 1 0 76832 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1379_
timestamp 1698431365
transform 1 0 74928 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1380_
timestamp 1698431365
transform -1 0 72688 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1381_
timestamp 1698431365
transform -1 0 63616 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1382_
timestamp 1698431365
transform 1 0 63168 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1383_
timestamp 1698431365
transform -1 0 70672 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1384_
timestamp 1698431365
transform -1 0 71232 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1385_
timestamp 1698431365
transform 1 0 63280 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1386_
timestamp 1698431365
transform 1 0 67984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1387_
timestamp 1698431365
transform 1 0 49840 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1388_
timestamp 1698431365
transform 1 0 62384 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1389_
timestamp 1698431365
transform -1 0 66976 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1390_
timestamp 1698431365
transform -1 0 60144 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1391_
timestamp 1698431365
transform 1 0 64848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1392_
timestamp 1698431365
transform -1 0 65184 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1393_
timestamp 1698431365
transform 1 0 62384 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1394_
timestamp 1698431365
transform -1 0 65632 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1395_
timestamp 1698431365
transform 1 0 64288 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1396_
timestamp 1698431365
transform 1 0 66752 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1397_
timestamp 1698431365
transform 1 0 65184 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1398_
timestamp 1698431365
transform 1 0 65632 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1399_
timestamp 1698431365
transform 1 0 65856 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1400_
timestamp 1698431365
transform -1 0 65968 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1401_
timestamp 1698431365
transform -1 0 64400 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1402_
timestamp 1698431365
transform 1 0 64624 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1403_
timestamp 1698431365
transform -1 0 73024 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1404_
timestamp 1698431365
transform 1 0 71232 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1405_
timestamp 1698431365
transform -1 0 69664 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1406_
timestamp 1698431365
transform 1 0 65072 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1407_
timestamp 1698431365
transform -1 0 67424 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1408_
timestamp 1698431365
transform -1 0 71456 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1409_
timestamp 1698431365
transform 1 0 66192 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1410_
timestamp 1698431365
transform 1 0 70000 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1411_
timestamp 1698431365
transform 1 0 70000 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1412_
timestamp 1698431365
transform 1 0 75264 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1413_
timestamp 1698431365
transform 1 0 74032 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1414_
timestamp 1698431365
transform 1 0 79968 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1415_
timestamp 1698431365
transform 1 0 71792 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1416_
timestamp 1698431365
transform 1 0 73024 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1417_
timestamp 1698431365
transform 1 0 72464 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1418_
timestamp 1698431365
transform -1 0 67984 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1419_
timestamp 1698431365
transform 1 0 73024 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1420_
timestamp 1698431365
transform 1 0 77728 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1421_
timestamp 1698431365
transform -1 0 76608 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1422_
timestamp 1698431365
transform 1 0 72576 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1423_
timestamp 1698431365
transform 1 0 74368 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1424_
timestamp 1698431365
transform -1 0 89488 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1425_
timestamp 1698431365
transform 1 0 85680 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1426_
timestamp 1698431365
transform 1 0 71680 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1427_
timestamp 1698431365
transform 1 0 79968 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1428_
timestamp 1698431365
transform 1 0 86128 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1429_
timestamp 1698431365
transform 1 0 90496 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1430_
timestamp 1698431365
transform 1 0 89264 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1431_
timestamp 1698431365
transform -1 0 93296 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1432_
timestamp 1698431365
transform 1 0 89712 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1433_
timestamp 1698431365
transform -1 0 93856 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1434_
timestamp 1698431365
transform -1 0 92736 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1435_
timestamp 1698431365
transform -1 0 92960 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1436_
timestamp 1698431365
transform -1 0 93296 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1437_
timestamp 1698431365
transform -1 0 92624 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1438_
timestamp 1698431365
transform 1 0 82768 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1439_
timestamp 1698431365
transform -1 0 86016 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1440_
timestamp 1698431365
transform 1 0 99568 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1441_
timestamp 1698431365
transform -1 0 86128 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1442_
timestamp 1698431365
transform -1 0 84784 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1443_
timestamp 1698431365
transform -1 0 93184 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1444_
timestamp 1698431365
transform 1 0 79072 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1445_
timestamp 1698431365
transform -1 0 83664 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1446_
timestamp 1698431365
transform -1 0 87472 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1447_
timestamp 1698431365
transform 1 0 78736 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1448_
timestamp 1698431365
transform -1 0 81312 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1449_
timestamp 1698431365
transform -1 0 80864 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1450_
timestamp 1698431365
transform -1 0 79744 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1451_
timestamp 1698431365
transform 1 0 83664 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1452_
timestamp 1698431365
transform -1 0 79744 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1453_
timestamp 1698431365
transform -1 0 81760 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1454_
timestamp 1698431365
transform 1 0 80192 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1455_
timestamp 1698431365
transform 1 0 48720 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1456_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 62048 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1457_
timestamp 1698431365
transform 1 0 64288 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1458_
timestamp 1698431365
transform 1 0 64288 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1459_
timestamp 1698431365
transform 1 0 77056 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1460_
timestamp 1698431365
transform -1 0 76160 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1461_
timestamp 1698431365
transform 1 0 74928 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1462_
timestamp 1698431365
transform 1 0 73920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1463_
timestamp 1698431365
transform 1 0 63504 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1464_
timestamp 1698431365
transform -1 0 66416 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1465_
timestamp 1698431365
transform -1 0 69664 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1466_
timestamp 1698431365
transform -1 0 65184 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1467_
timestamp 1698431365
transform 1 0 59248 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1468_
timestamp 1698431365
transform -1 0 58800 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1469_
timestamp 1698431365
transform -1 0 49504 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1470_
timestamp 1698431365
transform 1 0 50624 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1471_
timestamp 1698431365
transform 1 0 61488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1472_
timestamp 1698431365
transform -1 0 48384 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1473_
timestamp 1698431365
transform 1 0 45024 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1474_
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1475_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26208 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1476_
timestamp 1698431365
transform -1 0 70896 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1477_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 62384 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1478_
timestamp 1698431365
transform 1 0 68768 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1479_
timestamp 1698431365
transform -1 0 59808 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1480_
timestamp 1698431365
transform 1 0 73472 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1481_
timestamp 1698431365
transform 1 0 75152 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1482_
timestamp 1698431365
transform 1 0 74928 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1483_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 73472 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1484_
timestamp 1698431365
transform -1 0 72464 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1485_
timestamp 1698431365
transform 1 0 70560 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1486_
timestamp 1698431365
transform 1 0 67424 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1487_
timestamp 1698431365
transform 1 0 69776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1488_
timestamp 1698431365
transform 1 0 70224 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1489_
timestamp 1698431365
transform -1 0 71456 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1490_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 71344 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1491_
timestamp 1698431365
transform -1 0 70224 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1492_
timestamp 1698431365
transform -1 0 65968 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1493_
timestamp 1698431365
transform 1 0 37968 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1494_
timestamp 1698431365
transform -1 0 41664 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1495_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40432 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1496_
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1497_
timestamp 1698431365
transform 1 0 72128 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1498_
timestamp 1698431365
transform -1 0 75152 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1499_
timestamp 1698431365
transform -1 0 77056 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1500_
timestamp 1698431365
transform 1 0 76384 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1501_
timestamp 1698431365
transform 1 0 74368 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1502_
timestamp 1698431365
transform -1 0 76496 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1503_
timestamp 1698431365
transform 1 0 74368 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1504_
timestamp 1698431365
transform 1 0 73696 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1505_
timestamp 1698431365
transform 1 0 76384 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1506_
timestamp 1698431365
transform 1 0 78176 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1507_
timestamp 1698431365
transform 1 0 77280 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1508_
timestamp 1698431365
transform 1 0 78064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1509_
timestamp 1698431365
transform 1 0 78400 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1510_
timestamp 1698431365
transform 1 0 80416 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1511_
timestamp 1698431365
transform 1 0 80640 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1512_
timestamp 1698431365
transform -1 0 82432 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1513_
timestamp 1698431365
transform 1 0 82880 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1514_
timestamp 1698431365
transform -1 0 81984 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1515_
timestamp 1698431365
transform -1 0 82880 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1516_
timestamp 1698431365
transform 1 0 76160 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1517_
timestamp 1698431365
transform -1 0 81536 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1518_
timestamp 1698431365
transform -1 0 82432 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1519_
timestamp 1698431365
transform 1 0 81984 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1520_
timestamp 1698431365
transform 1 0 81088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1521_
timestamp 1698431365
transform -1 0 49504 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1522_
timestamp 1698431365
transform -1 0 33936 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1523_
timestamp 1698431365
transform -1 0 32704 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1524_
timestamp 1698431365
transform -1 0 26992 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1525_
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1526_
timestamp 1698431365
transform 1 0 33264 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1527_
timestamp 1698431365
transform -1 0 32032 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1528_
timestamp 1698431365
transform 1 0 30576 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1529_
timestamp 1698431365
transform 1 0 32368 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1530_
timestamp 1698431365
transform 1 0 33712 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1531_
timestamp 1698431365
transform -1 0 33824 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1532_
timestamp 1698431365
transform 1 0 31696 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1533_
timestamp 1698431365
transform 1 0 32480 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1534_
timestamp 1698431365
transform -1 0 24864 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1535_
timestamp 1698431365
transform -1 0 26544 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1536_
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1537_
timestamp 1698431365
transform -1 0 24752 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1538_
timestamp 1698431365
transform -1 0 24304 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1539_
timestamp 1698431365
transform 1 0 31808 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1540_
timestamp 1698431365
transform -1 0 34384 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1541_
timestamp 1698431365
transform 1 0 30576 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1542_
timestamp 1698431365
transform -1 0 69888 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1543_
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1544_
timestamp 1698431365
transform -1 0 30128 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1545_
timestamp 1698431365
transform -1 0 30240 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1546_
timestamp 1698431365
transform -1 0 33712 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1547_
timestamp 1698431365
transform -1 0 36176 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1548_
timestamp 1698431365
transform -1 0 32704 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1549_
timestamp 1698431365
transform 1 0 34496 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1550_
timestamp 1698431365
transform 1 0 29792 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1551_
timestamp 1698431365
transform -1 0 29680 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1552_
timestamp 1698431365
transform 1 0 30464 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1553_
timestamp 1698431365
transform 1 0 31584 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1554_
timestamp 1698431365
transform 1 0 27552 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1555_
timestamp 1698431365
transform -1 0 27440 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1556_
timestamp 1698431365
transform 1 0 27328 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1557_
timestamp 1698431365
transform -1 0 27664 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1558_
timestamp 1698431365
transform 1 0 30016 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1559_
timestamp 1698431365
transform 1 0 31136 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1560_
timestamp 1698431365
transform 1 0 27776 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1561_
timestamp 1698431365
transform -1 0 28784 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1562_
timestamp 1698431365
transform -1 0 31920 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1563_
timestamp 1698431365
transform -1 0 30576 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1564_
timestamp 1698431365
transform 1 0 30912 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1565_
timestamp 1698431365
transform 1 0 38192 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1566_
timestamp 1698431365
transform 1 0 33936 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1567_
timestamp 1698431365
transform 1 0 35504 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1568_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1569_
timestamp 1698431365
transform -1 0 38304 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1570_
timestamp 1698431365
transform 1 0 36064 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1571_
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1572_
timestamp 1698431365
transform -1 0 29456 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1573_
timestamp 1698431365
transform -1 0 29568 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1574_
timestamp 1698431365
transform 1 0 27552 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1575_
timestamp 1698431365
transform 1 0 34384 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1576_
timestamp 1698431365
transform 1 0 40096 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1577_
timestamp 1698431365
transform 1 0 37856 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1578_
timestamp 1698431365
transform -1 0 70784 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1579_
timestamp 1698431365
transform -1 0 43344 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1580_
timestamp 1698431365
transform 1 0 41552 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1581_
timestamp 1698431365
transform 1 0 40880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1582_
timestamp 1698431365
transform -1 0 39760 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1583_
timestamp 1698431365
transform -1 0 25536 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1584_
timestamp 1698431365
transform -1 0 26320 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1585_
timestamp 1698431365
transform -1 0 25424 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1586_
timestamp 1698431365
transform 1 0 30464 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1587_
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1588_
timestamp 1698431365
transform -1 0 43904 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1589_
timestamp 1698431365
transform 1 0 40880 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1590_
timestamp 1698431365
transform 1 0 29680 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1591_
timestamp 1698431365
transform 1 0 40656 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1592_
timestamp 1698431365
transform 1 0 45136 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1593_
timestamp 1698431365
transform 1 0 26656 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1594_
timestamp 1698431365
transform 1 0 26320 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1595_
timestamp 1698431365
transform -1 0 27104 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1596_
timestamp 1698431365
transform -1 0 39200 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1597_
timestamp 1698431365
transform 1 0 35616 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1598_
timestamp 1698431365
transform 1 0 36960 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1599_
timestamp 1698431365
transform -1 0 23072 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1600_
timestamp 1698431365
transform -1 0 25648 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1601_
timestamp 1698431365
transform -1 0 24304 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1602_
timestamp 1698431365
transform -1 0 24080 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1603_
timestamp 1698431365
transform -1 0 22960 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1604_
timestamp 1698431365
transform 1 0 22960 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1605_
timestamp 1698431365
transform -1 0 23632 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1606_
timestamp 1698431365
transform -1 0 24304 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1607_
timestamp 1698431365
transform -1 0 23520 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1608_
timestamp 1698431365
transform 1 0 18816 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1609_
timestamp 1698431365
transform -1 0 20608 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1610_
timestamp 1698431365
transform -1 0 61040 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1611_
timestamp 1698431365
transform -1 0 54992 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1612_
timestamp 1698431365
transform -1 0 54096 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1613_
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1614_
timestamp 1698431365
transform 1 0 23520 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1615_
timestamp 1698431365
transform -1 0 76384 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1616_
timestamp 1698431365
transform 1 0 55328 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1617_
timestamp 1698431365
transform 1 0 53424 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1618_
timestamp 1698431365
transform -1 0 61376 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1619_
timestamp 1698431365
transform 1 0 55664 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1620_
timestamp 1698431365
transform 1 0 30240 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1621_
timestamp 1698431365
transform 1 0 55888 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1622_
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1623_
timestamp 1698431365
transform 1 0 56448 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1624_
timestamp 1698431365
transform -1 0 27888 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1625_
timestamp 1698431365
transform -1 0 26880 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1626_
timestamp 1698431365
transform 1 0 56560 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1627_
timestamp 1698431365
transform -1 0 58464 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1628_
timestamp 1698431365
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1629_
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1630_
timestamp 1698431365
transform 1 0 54544 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1631_
timestamp 1698431365
transform 1 0 43680 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1632_
timestamp 1698431365
transform 1 0 61824 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1633_
timestamp 1698431365
transform 1 0 60592 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1634_
timestamp 1698431365
transform -1 0 59584 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1635_
timestamp 1698431365
transform 1 0 55104 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1636_
timestamp 1698431365
transform 1 0 56896 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1637_
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1638_
timestamp 1698431365
transform 1 0 61264 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1639_
timestamp 1698431365
transform 1 0 60368 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1640_
timestamp 1698431365
transform 1 0 51744 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1641_
timestamp 1698431365
transform -1 0 77616 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1642_
timestamp 1698431365
transform -1 0 59024 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1643_
timestamp 1698431365
transform -1 0 53984 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1644_
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1645_
timestamp 1698431365
transform 1 0 52864 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1646_
timestamp 1698431365
transform 1 0 56672 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1647_
timestamp 1698431365
transform 1 0 72576 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1648_
timestamp 1698431365
transform -1 0 73024 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1649_
timestamp 1698431365
transform -1 0 60928 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1650_
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1651_
timestamp 1698431365
transform -1 0 62160 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1652_
timestamp 1698431365
transform 1 0 60368 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1653_
timestamp 1698431365
transform -1 0 71792 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1654_
timestamp 1698431365
transform 1 0 67088 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1655_
timestamp 1698431365
transform 1 0 67312 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1656_
timestamp 1698431365
transform 1 0 71904 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1657_
timestamp 1698431365
transform 1 0 83888 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1658_
timestamp 1698431365
transform -1 0 77504 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1659_
timestamp 1698431365
transform -1 0 76832 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1660_
timestamp 1698431365
transform -1 0 73696 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1661_
timestamp 1698431365
transform 1 0 66304 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1662_
timestamp 1698431365
transform -1 0 73024 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1663_
timestamp 1698431365
transform -1 0 67088 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1664_
timestamp 1698431365
transform 1 0 86912 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1665_
timestamp 1698431365
transform -1 0 88368 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1666_
timestamp 1698431365
transform 1 0 85344 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1667_
timestamp 1698431365
transform 1 0 75712 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1668_
timestamp 1698431365
transform 1 0 86016 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1669_
timestamp 1698431365
transform -1 0 87696 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1670_
timestamp 1698431365
transform -1 0 86800 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1671_
timestamp 1698431365
transform -1 0 83664 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1672_
timestamp 1698431365
transform -1 0 92288 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1673_
timestamp 1698431365
transform 1 0 105840 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1674_
timestamp 1698431365
transform -1 0 87584 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1675_
timestamp 1698431365
transform -1 0 87584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1676_
timestamp 1698431365
transform -1 0 95200 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1677_
timestamp 1698431365
transform -1 0 91168 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1678_
timestamp 1698431365
transform -1 0 88928 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1679_
timestamp 1698431365
transform 1 0 105168 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1680_
timestamp 1698431365
transform -1 0 101472 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1681_
timestamp 1698431365
transform -1 0 103936 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1682_
timestamp 1698431365
transform 1 0 70784 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1683_
timestamp 1698431365
transform -1 0 106736 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1684_
timestamp 1698431365
transform -1 0 101024 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1685_
timestamp 1698431365
transform -1 0 100464 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1686_
timestamp 1698431365
transform -1 0 104048 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1687_
timestamp 1698431365
transform -1 0 100912 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1688_
timestamp 1698431365
transform 1 0 103824 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1689_
timestamp 1698431365
transform 1 0 105392 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1690_
timestamp 1698431365
transform -1 0 111216 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1691_
timestamp 1698431365
transform -1 0 105168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1692_
timestamp 1698431365
transform 1 0 107184 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1693_
timestamp 1698431365
transform -1 0 111104 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1694_
timestamp 1698431365
transform -1 0 108304 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1695_
timestamp 1698431365
transform 1 0 110432 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1696_
timestamp 1698431365
transform 1 0 111328 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1697_
timestamp 1698431365
transform 1 0 110544 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1698_
timestamp 1698431365
transform 1 0 109648 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1699_
timestamp 1698431365
transform 1 0 112896 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1700_
timestamp 1698431365
transform -1 0 115920 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1701_
timestamp 1698431365
transform 1 0 114464 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1702_
timestamp 1698431365
transform -1 0 113232 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1703_
timestamp 1698431365
transform -1 0 115808 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1704_
timestamp 1698431365
transform 1 0 108304 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1705_
timestamp 1698431365
transform 1 0 117040 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1706_
timestamp 1698431365
transform -1 0 114688 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1707_
timestamp 1698431365
transform -1 0 114688 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1708_
timestamp 1698431365
transform -1 0 116480 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1709_
timestamp 1698431365
transform -1 0 114128 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1710_
timestamp 1698431365
transform 1 0 102816 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1711_
timestamp 1698431365
transform -1 0 109312 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1712_
timestamp 1698431365
transform -1 0 109648 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1713_
timestamp 1698431365
transform -1 0 107184 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1714_
timestamp 1698431365
transform -1 0 107184 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1715_
timestamp 1698431365
transform 1 0 107408 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1716_
timestamp 1698431365
transform 1 0 117040 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1717_
timestamp 1698431365
transform -1 0 110208 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1718_
timestamp 1698431365
transform 1 0 104384 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1719_
timestamp 1698431365
transform 1 0 103488 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1720_
timestamp 1698431365
transform -1 0 108304 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1721_
timestamp 1698431365
transform -1 0 105952 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1722_
timestamp 1698431365
transform -1 0 106400 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1723_
timestamp 1698431365
transform -1 0 105392 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1724_
timestamp 1698431365
transform 1 0 102368 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1725_
timestamp 1698431365
transform 1 0 94304 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1726_
timestamp 1698431365
transform -1 0 97104 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1727_
timestamp 1698431365
transform 1 0 108304 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1728_
timestamp 1698431365
transform -1 0 93856 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1729_
timestamp 1698431365
transform -1 0 95984 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1730_
timestamp 1698431365
transform 1 0 98784 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1731_
timestamp 1698431365
transform -1 0 102816 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1732_
timestamp 1698431365
transform 1 0 102144 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1733_
timestamp 1698431365
transform 1 0 52640 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1734_
timestamp 1698431365
transform -1 0 45360 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1735_
timestamp 1698431365
transform -1 0 39648 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1736_
timestamp 1698431365
transform 1 0 53984 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1737_
timestamp 1698431365
transform 1 0 49056 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1738_
timestamp 1698431365
transform 1 0 47824 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1739_
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1740_
timestamp 1698431365
transform -1 0 47824 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1741_
timestamp 1698431365
transform 1 0 43904 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1742_
timestamp 1698431365
transform -1 0 47488 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1743_
timestamp 1698431365
transform 1 0 45360 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1744_
timestamp 1698431365
transform -1 0 46928 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1745_
timestamp 1698431365
transform 1 0 43904 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1746_
timestamp 1698431365
transform 1 0 45024 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1747_
timestamp 1698431365
transform -1 0 49168 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1748_
timestamp 1698431365
transform -1 0 53536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1749_
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1750_
timestamp 1698431365
transform 1 0 45696 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1751_
timestamp 1698431365
transform 1 0 47824 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1752_
timestamp 1698431365
transform -1 0 50064 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1753_
timestamp 1698431365
transform -1 0 48160 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1754_
timestamp 1698431365
transform -1 0 59024 0 1 26656
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1755_
timestamp 1698431365
transform 1 0 53984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1756_
timestamp 1698431365
transform -1 0 53312 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1757_
timestamp 1698431365
transform -1 0 53424 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1758_
timestamp 1698431365
transform 1 0 50064 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1759_
timestamp 1698431365
transform 1 0 62048 0 1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1760_
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1761_
timestamp 1698431365
transform -1 0 57008 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1762_
timestamp 1698431365
transform -1 0 58800 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1763_
timestamp 1698431365
transform -1 0 56224 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1764_
timestamp 1698431365
transform -1 0 57344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1698431365
transform -1 0 56224 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1766_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 57904 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1767_
timestamp 1698431365
transform -1 0 55552 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1768_
timestamp 1698431365
transform -1 0 54320 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1769_
timestamp 1698431365
transform -1 0 52976 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1770_
timestamp 1698431365
transform -1 0 57456 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1771_
timestamp 1698431365
transform -1 0 53536 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1772_
timestamp 1698431365
transform -1 0 52304 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1773_
timestamp 1698431365
transform -1 0 56224 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1774_
timestamp 1698431365
transform -1 0 46592 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1775_
timestamp 1698431365
transform -1 0 57568 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1776_
timestamp 1698431365
transform 1 0 49056 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1777_
timestamp 1698431365
transform -1 0 43568 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1778_
timestamp 1698431365
transform -1 0 43120 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1779_
timestamp 1698431365
transform 1 0 43120 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1780_
timestamp 1698431365
transform 1 0 44128 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1781_
timestamp 1698431365
transform 1 0 47152 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1782_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47600 0 1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1783_
timestamp 1698431365
transform 1 0 49392 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1784_
timestamp 1698431365
transform 1 0 49504 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1785_
timestamp 1698431365
transform -1 0 53312 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1786_
timestamp 1698431365
transform 1 0 48944 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1787_
timestamp 1698431365
transform 1 0 51296 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1788_
timestamp 1698431365
transform -1 0 51408 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1789_
timestamp 1698431365
transform 1 0 47488 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1790_
timestamp 1698431365
transform 1 0 50064 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1791_
timestamp 1698431365
transform -1 0 49168 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1792_
timestamp 1698431365
transform 1 0 48720 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1793_
timestamp 1698431365
transform -1 0 45472 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1794_
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1795_
timestamp 1698431365
transform 1 0 54656 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1796_
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1797_
timestamp 1698431365
transform 1 0 50512 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1798_
timestamp 1698431365
transform -1 0 51296 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1799_
timestamp 1698431365
transform -1 0 56672 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1800_
timestamp 1698431365
transform 1 0 56672 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1801_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 54320 0 1 23520
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1802_
timestamp 1698431365
transform 1 0 54768 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1803_
timestamp 1698431365
transform 1 0 44912 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1804_
timestamp 1698431365
transform 1 0 49952 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1805_
timestamp 1698431365
transform 1 0 49728 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1806_
timestamp 1698431365
transform 1 0 50960 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1807_
timestamp 1698431365
transform -1 0 69104 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1808_
timestamp 1698431365
transform 1 0 53536 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1809_
timestamp 1698431365
transform -1 0 54432 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1810_
timestamp 1698431365
transform -1 0 54656 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1811_
timestamp 1698431365
transform -1 0 53760 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1812_
timestamp 1698431365
transform 1 0 52304 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1813_
timestamp 1698431365
transform -1 0 58912 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1814_
timestamp 1698431365
transform -1 0 44128 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1815_
timestamp 1698431365
transform -1 0 42224 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1816_
timestamp 1698431365
transform 1 0 23184 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1817_
timestamp 1698431365
transform -1 0 39872 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1818_
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1819_
timestamp 1698431365
transform 1 0 40432 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1820_
timestamp 1698431365
transform -1 0 41664 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1821_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1822_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44352 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1823_
timestamp 1698431365
transform 1 0 45248 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1824_
timestamp 1698431365
transform 1 0 44912 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1825_
timestamp 1698431365
transform 1 0 47040 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1826_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45808 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1827_
timestamp 1698431365
transform 1 0 46256 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1828_
timestamp 1698431365
transform -1 0 49616 0 1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1829_
timestamp 1698431365
transform -1 0 49280 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1830_
timestamp 1698431365
transform -1 0 47824 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1831_
timestamp 1698431365
transform -1 0 47040 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1832_
timestamp 1698431365
transform 1 0 47264 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1833_
timestamp 1698431365
transform -1 0 50624 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1834_
timestamp 1698431365
transform 1 0 49616 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1835_
timestamp 1698431365
transform 1 0 62384 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1836_
timestamp 1698431365
transform 1 0 69216 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1837_
timestamp 1698431365
transform 1 0 69888 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1838_
timestamp 1698431365
transform -1 0 59472 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1839_
timestamp 1698431365
transform 1 0 30688 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1840_
timestamp 1698431365
transform -1 0 40432 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1841_
timestamp 1698431365
transform 1 0 39648 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1842_
timestamp 1698431365
transform -1 0 39648 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1843_
timestamp 1698431365
transform 1 0 39872 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1844_
timestamp 1698431365
transform 1 0 40880 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1845_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41440 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1846_
timestamp 1698431365
transform 1 0 43008 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1847_
timestamp 1698431365
transform 1 0 51184 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1848_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 50064 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1849_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 50288 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1850_
timestamp 1698431365
transform 1 0 50512 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1851_
timestamp 1698431365
transform -1 0 52192 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1852_
timestamp 1698431365
transform 1 0 52528 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1853_
timestamp 1698431365
transform 1 0 41328 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1854_
timestamp 1698431365
transform -1 0 51408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1855_
timestamp 1698431365
transform -1 0 58128 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1856_
timestamp 1698431365
transform -1 0 53312 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1857_
timestamp 1698431365
transform -1 0 48384 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1858_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 52304 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1859_
timestamp 1698431365
transform 1 0 52416 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1860_
timestamp 1698431365
transform -1 0 56224 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1861_
timestamp 1698431365
transform -1 0 55552 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1862_
timestamp 1698431365
transform -1 0 51072 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1863_
timestamp 1698431365
transform 1 0 59360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1864_
timestamp 1698431365
transform -1 0 61376 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1865_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 52304 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1866_
timestamp 1698431365
transform -1 0 37744 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1867_
timestamp 1698431365
transform 1 0 33712 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1868_
timestamp 1698431365
transform 1 0 34160 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1869_
timestamp 1698431365
transform 1 0 37184 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1870_
timestamp 1698431365
transform 1 0 35728 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1871_
timestamp 1698431365
transform 1 0 38192 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1872_
timestamp 1698431365
transform 1 0 38080 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1873_
timestamp 1698431365
transform 1 0 39200 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1874_
timestamp 1698431365
transform 1 0 43120 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1875_
timestamp 1698431365
transform 1 0 41552 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1876_
timestamp 1698431365
transform -1 0 43008 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1877_
timestamp 1698431365
transform 1 0 46256 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1878_
timestamp 1698431365
transform 1 0 47488 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1879_
timestamp 1698431365
transform -1 0 48384 0 -1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1880_
timestamp 1698431365
transform -1 0 47600 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1881_
timestamp 1698431365
transform 1 0 51184 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1882_
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1883_
timestamp 1698431365
transform 1 0 66192 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1884_
timestamp 1698431365
transform -1 0 64736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1885_
timestamp 1698431365
transform 1 0 58912 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1886_
timestamp 1698431365
transform -1 0 61712 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1887_
timestamp 1698431365
transform -1 0 60144 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1888_
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1889_
timestamp 1698431365
transform 1 0 41552 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1890_
timestamp 1698431365
transform 1 0 43120 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1891_
timestamp 1698431365
transform 1 0 45248 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1892_
timestamp 1698431365
transform 1 0 59920 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1893_
timestamp 1698431365
transform 1 0 33824 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1894_
timestamp 1698431365
transform -1 0 31584 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1895_
timestamp 1698431365
transform 1 0 30800 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1896_
timestamp 1698431365
transform 1 0 34496 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1897_
timestamp 1698431365
transform -1 0 36960 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1898_
timestamp 1698431365
transform 1 0 35392 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1899_
timestamp 1698431365
transform 1 0 35392 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1900_
timestamp 1698431365
transform 1 0 49504 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1901_
timestamp 1698431365
transform 1 0 63280 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1902_
timestamp 1698431365
transform -1 0 59920 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1903_
timestamp 1698431365
transform 1 0 59584 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1904_
timestamp 1698431365
transform 1 0 60816 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1905_
timestamp 1698431365
transform 1 0 31584 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1906_
timestamp 1698431365
transform -1 0 35728 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1907_
timestamp 1698431365
transform 1 0 34832 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1908_
timestamp 1698431365
transform -1 0 43120 0 1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1909_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1910_
timestamp 1698431365
transform 1 0 51408 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1911_
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1912_
timestamp 1698431365
transform -1 0 44800 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1913_
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1914_
timestamp 1698431365
transform 1 0 60368 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1915_
timestamp 1698431365
transform 1 0 30464 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1916_
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1917_
timestamp 1698431365
transform 1 0 34496 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1918_
timestamp 1698431365
transform 1 0 18928 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1919_
timestamp 1698431365
transform -1 0 19600 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1920_
timestamp 1698431365
transform -1 0 19376 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1921_
timestamp 1698431365
transform 1 0 20496 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1922_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1923_
timestamp 1698431365
transform -1 0 24976 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1924_
timestamp 1698431365
transform 1 0 19376 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1925_
timestamp 1698431365
transform -1 0 20608 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1926_
timestamp 1698431365
transform 1 0 19600 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1927_
timestamp 1698431365
transform 1 0 21168 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1928_
timestamp 1698431365
transform 1 0 21728 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1929_
timestamp 1698431365
transform -1 0 22624 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1930_
timestamp 1698431365
transform -1 0 21840 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1931_
timestamp 1698431365
transform 1 0 19600 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1932_
timestamp 1698431365
transform 1 0 20832 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1933_
timestamp 1698431365
transform 1 0 20496 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1934_
timestamp 1698431365
transform -1 0 32704 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1935_
timestamp 1698431365
transform 1 0 30016 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1936_
timestamp 1698431365
transform -1 0 28000 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1937_
timestamp 1698431365
transform -1 0 27328 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1938_
timestamp 1698431365
transform -1 0 25760 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1939_
timestamp 1698431365
transform -1 0 24864 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1940_
timestamp 1698431365
transform 1 0 26992 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1941_
timestamp 1698431365
transform 1 0 27888 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1942_
timestamp 1698431365
transform 1 0 26320 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1943_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1944_
timestamp 1698431365
transform 1 0 23744 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1945_
timestamp 1698431365
transform 1 0 27440 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1946_
timestamp 1698431365
transform 1 0 26768 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1947_
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1948_
timestamp 1698431365
transform -1 0 37184 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1949_
timestamp 1698431365
transform -1 0 37520 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1950_
timestamp 1698431365
transform 1 0 34832 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1951_
timestamp 1698431365
transform -1 0 34832 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1952_
timestamp 1698431365
transform -1 0 33040 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1953_
timestamp 1698431365
transform 1 0 31248 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1954_
timestamp 1698431365
transform -1 0 29904 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1955_
timestamp 1698431365
transform -1 0 30576 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1956_
timestamp 1698431365
transform 1 0 39200 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1957_
timestamp 1698431365
transform 1 0 39648 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1958_
timestamp 1698431365
transform -1 0 40544 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1959_
timestamp 1698431365
transform 1 0 38192 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1960_
timestamp 1698431365
transform -1 0 42336 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1961_
timestamp 1698431365
transform 1 0 42448 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1962_
timestamp 1698431365
transform -1 0 44464 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1963_
timestamp 1698431365
transform 1 0 44912 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1964_
timestamp 1698431365
transform 1 0 44128 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1965_
timestamp 1698431365
transform -1 0 38080 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1966_
timestamp 1698431365
transform -1 0 38528 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1967_
timestamp 1698431365
transform 1 0 45360 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1968_
timestamp 1698431365
transform 1 0 44688 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1969_
timestamp 1698431365
transform -1 0 29904 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1970_
timestamp 1698431365
transform -1 0 26768 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1971_
timestamp 1698431365
transform -1 0 28560 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1972_
timestamp 1698431365
transform -1 0 22176 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1973_
timestamp 1698431365
transform 1 0 16576 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1974_
timestamp 1698431365
transform -1 0 22288 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1975_
timestamp 1698431365
transform -1 0 31024 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1976_
timestamp 1698431365
transform -1 0 24864 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1977_
timestamp 1698431365
transform -1 0 24192 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1978_
timestamp 1698431365
transform 1 0 23744 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1979_
timestamp 1698431365
transform -1 0 26096 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1980_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1981_
timestamp 1698431365
transform -1 0 25536 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1982_
timestamp 1698431365
transform 1 0 28000 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1983_
timestamp 1698431365
transform 1 0 28560 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1984_
timestamp 1698431365
transform -1 0 21728 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1985_
timestamp 1698431365
transform 1 0 21280 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1986_
timestamp 1698431365
transform -1 0 20944 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1987_
timestamp 1698431365
transform 1 0 22624 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1988_
timestamp 1698431365
transform -1 0 22624 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1989_
timestamp 1698431365
transform -1 0 23408 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1990_
timestamp 1698431365
transform 1 0 39424 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1991_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 111664 0 1 20384
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1992_
timestamp 1698431365
transform 1 0 108192 0 1 20384
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1993_
timestamp 1698431365
transform 1 0 112112 0 -1 17248
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1994_
timestamp 1698431365
transform 1 0 109088 0 1 17248
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1995_
timestamp 1698431365
transform 1 0 107408 0 1 14112
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1996_
timestamp 1698431365
transform 1 0 107408 0 -1 14112
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1997_
timestamp 1698431365
transform 1 0 105616 0 -1 17248
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1998_
timestamp 1698431365
transform 1 0 103488 0 1 20384
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1999_
timestamp 1698431365
transform -1 0 96208 0 1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2000_
timestamp 1698431365
transform 1 0 90272 0 -1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2001_
timestamp 1698431365
transform 1 0 89488 0 -1 23520
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2002_
timestamp 1698431365
transform 1 0 85456 0 1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2003_
timestamp 1698431365
transform -1 0 87136 0 -1 17248
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2004_
timestamp 1698431365
transform -1 0 91168 0 -1 18816
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2005_
timestamp 1698431365
transform -1 0 88480 0 1 20384
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2006_
timestamp 1698431365
transform 1 0 90048 0 -1 20384
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2007_
timestamp 1698431365
transform -1 0 101584 0 -1 20384
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2008_
timestamp 1698431365
transform 1 0 95536 0 1 20384
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2009_
timestamp 1698431365
transform 1 0 94080 0 1 17248
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2010_
timestamp 1698431365
transform 1 0 95648 0 1 15680
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2011_
timestamp 1698431365
transform 1 0 99568 0 1 14112
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2012_
timestamp 1698431365
transform 1 0 102928 0 1 14112
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2013_
timestamp 1698431365
transform 1 0 103488 0 -1 15680
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2014_
timestamp 1698431365
transform 1 0 101248 0 1 15680
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2015_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42784 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2016_
timestamp 1698431365
transform 1 0 68768 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2017_
timestamp 1698431365
transform 1 0 72240 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2018_
timestamp 1698431365
transform 1 0 74928 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2019_
timestamp 1698431365
transform 1 0 69664 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2020_
timestamp 1698431365
transform 1 0 68208 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2021_
timestamp 1698431365
transform 1 0 64288 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2022_
timestamp 1698431365
transform 1 0 63056 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2023_
timestamp 1698431365
transform -1 0 69104 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2024_
timestamp 1698431365
transform 1 0 63616 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2025_
timestamp 1698431365
transform 1 0 66864 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2026_
timestamp 1698431365
transform 1 0 68656 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2027_
timestamp 1698431365
transform 1 0 73696 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2028_
timestamp 1698431365
transform 1 0 72016 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2029_
timestamp 1698431365
transform 1 0 73472 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2030_
timestamp 1698431365
transform 1 0 87808 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2031_
timestamp 1698431365
transform 1 0 88480 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2032_
timestamp 1698431365
transform -1 0 94976 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2033_
timestamp 1698431365
transform -1 0 94304 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2034_
timestamp 1698431365
transform -1 0 87024 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2035_
timestamp 1698431365
transform 1 0 82432 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2036_
timestamp 1698431365
transform -1 0 81200 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2037_
timestamp 1698431365
transform -1 0 81648 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2038_
timestamp 1698431365
transform 1 0 79968 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2039_
timestamp 1698431365
transform -1 0 65744 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2040_
timestamp 1698431365
transform -1 0 71456 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2041_
timestamp 1698431365
transform 1 0 62832 0 1 28224
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2042_
timestamp 1698431365
transform -1 0 26656 0 1 25088
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2043_
timestamp 1698431365
transform -1 0 79408 0 1 26656
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_2  _2044_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 70448 0 -1 28224
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2045_
timestamp 1698431365
transform 1 0 64624 0 1 23520
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2046_
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2047_
timestamp 1698431365
transform 1 0 72240 0 -1 23520
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2048_
timestamp 1698431365
transform 1 0 72016 0 1 20384
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2049_
timestamp 1698431365
transform 1 0 76384 0 -1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2050_
timestamp 1698431365
transform 1 0 77280 0 1 25088
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2051_
timestamp 1698431365
transform -1 0 83664 0 1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2052_
timestamp 1698431365
transform -1 0 84672 0 -1 25088
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2053_
timestamp 1698431365
transform 1 0 79968 0 1 17248
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2054_
timestamp 1698431365
transform 1 0 80304 0 -1 18816
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2055_
timestamp 1698431365
transform 1 0 33376 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2056_
timestamp 1698431365
transform 1 0 30912 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2057_
timestamp 1698431365
transform 1 0 20944 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2058_
timestamp 1698431365
transform 1 0 31136 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2059_
timestamp 1698431365
transform 1 0 29568 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2060_
timestamp 1698431365
transform 1 0 26656 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2061_
timestamp 1698431365
transform 1 0 26992 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2062_
timestamp 1698431365
transform 1 0 27664 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2063_
timestamp 1698431365
transform 1 0 34944 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2064_
timestamp 1698431365
transform -1 0 40096 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2065_
timestamp 1698431365
transform 1 0 26544 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2066_
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2067_
timestamp 1698431365
transform 1 0 37184 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2068_
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2069_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25312 0 1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2070_
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2071_
timestamp 1698431365
transform 1 0 21616 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2072_
timestamp 1698431365
transform 1 0 21280 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2073_
timestamp 1698431365
transform 1 0 18928 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2074_
timestamp 1698431365
transform 1 0 50848 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2075_
timestamp 1698431365
transform 1 0 52640 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2076_
timestamp 1698431365
transform 1 0 54096 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2077_
timestamp 1698431365
transform 1 0 56672 0 -1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2078_
timestamp 1698431365
transform 1 0 54096 0 1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2079_
timestamp 1698431365
transform 1 0 59920 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2080_
timestamp 1698431365
transform 1 0 57792 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2081_
timestamp 1698431365
transform 1 0 59136 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2082_
timestamp 1698431365
transform 1 0 53984 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2083_
timestamp 1698431365
transform -1 0 58128 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2084_
timestamp 1698431365
transform -1 0 62048 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2085_
timestamp 1698431365
transform 1 0 68208 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2086_
timestamp 1698431365
transform 1 0 73024 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2087_
timestamp 1698431365
transform -1 0 69552 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2088_
timestamp 1698431365
transform 1 0 81872 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2089_
timestamp 1698431365
transform 1 0 82768 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2090_
timestamp 1698431365
transform 1 0 86464 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2091_
timestamp 1698431365
transform 1 0 87808 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2092_
timestamp 1698431365
transform -1 0 102816 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2093_
timestamp 1698431365
transform -1 0 102816 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2094_
timestamp 1698431365
transform -1 0 106064 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2095_
timestamp 1698431365
transform -1 0 109312 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2096_
timestamp 1698431365
transform -1 0 112336 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2097_
timestamp 1698431365
transform -1 0 114464 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2098_
timestamp 1698431365
transform -1 0 115584 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2099_
timestamp 1698431365
transform 1 0 112448 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2100_
timestamp 1698431365
transform 1 0 105392 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2101_
timestamp 1698431365
transform -1 0 110656 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2102_
timestamp 1698431365
transform -1 0 103376 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2103_
timestamp 1698431365
transform 1 0 101584 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2104_
timestamp 1698431365
transform -1 0 99344 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2105_
timestamp 1698431365
transform -1 0 99120 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2106_
timestamp 1698431365
transform 1 0 49056 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2107_
timestamp 1698431365
transform -1 0 52864 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2108_
timestamp 1698431365
transform 1 0 45136 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2109_
timestamp 1698431365
transform 1 0 41888 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2110_
timestamp 1698431365
transform 1 0 45136 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2111_
timestamp 1698431365
transform -1 0 53984 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2112_
timestamp 1698431365
transform 1 0 45808 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2113_
timestamp 1698431365
transform 1 0 50848 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2114_
timestamp 1698431365
transform 1 0 49056 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_2  _2115_
timestamp 1698431365
transform -1 0 47040 0 -1 29792
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2116_
timestamp 1698431365
transform 1 0 52640 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2117_
timestamp 1698431365
transform -1 0 71568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2118_
timestamp 1698431365
transform 1 0 55216 0 1 17248
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2119_
timestamp 1698431365
transform -1 0 68096 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2120_
timestamp 1698431365
transform -1 0 67536 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2121_
timestamp 1698431365
transform 1 0 60032 0 -1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2122_
timestamp 1698431365
transform -1 0 18704 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2123_
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2124_
timestamp 1698431365
transform 1 0 21504 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2125_
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2126_
timestamp 1698431365
transform 1 0 17696 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2127_
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2128_
timestamp 1698431365
transform 1 0 25424 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2129_
timestamp 1698431365
transform 1 0 22400 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2130_
timestamp 1698431365
transform 1 0 25312 0 1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2131_
timestamp 1698431365
transform 1 0 33376 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2132_
timestamp 1698431365
transform 1 0 30912 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2133_
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2134_
timestamp 1698431365
transform -1 0 41664 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2135_
timestamp 1698431365
transform 1 0 40880 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2136_
timestamp 1698431365
transform 1 0 43568 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2137_
timestamp 1698431365
transform 1 0 37296 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2138_
timestamp 1698431365
transform -1 0 47936 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2139_
timestamp 1698431365
transform -1 0 22512 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2140_
timestamp 1698431365
transform 1 0 22736 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2141_
timestamp 1698431365
transform 1 0 24192 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2142_
timestamp 1698431365
transform -1 0 30128 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2143_
timestamp 1698431365
transform 1 0 17136 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2144_
timestamp 1698431365
transform 1 0 19600 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2145_
timestamp 1698431365
transform -1 0 35280 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2150_
timestamp 1698431365
transform 1 0 69888 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2151_
timestamp 1698431365
transform 1 0 81312 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2152_
timestamp 1698431365
transform 1 0 92736 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2153_
timestamp 1698431365
transform 1 0 104160 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2154_
timestamp 1698431365
transform 1 0 115584 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2155_
timestamp 1698431365
transform 1 0 127008 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2156_
timestamp 1698431365
transform 1 0 138768 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__A1 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__A2
timestamp 1698431365
transform -1 0 19376 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__I
timestamp 1698431365
transform -1 0 72576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0975__I
timestamp 1698431365
transform 1 0 73136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__I
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__A1
timestamp 1698431365
transform 1 0 27888 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__A2
timestamp 1698431365
transform -1 0 29456 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A1
timestamp 1698431365
transform -1 0 60816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A2
timestamp 1698431365
transform 1 0 61488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0996__A1
timestamp 1698431365
transform -1 0 60704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0996__A2
timestamp 1698431365
transform 1 0 62720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__I
timestamp 1698431365
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A1
timestamp 1698431365
transform -1 0 92848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A2
timestamp 1698431365
transform -1 0 90944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A3
timestamp 1698431365
transform -1 0 97552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1005__B
timestamp 1698431365
transform -1 0 94864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1006__A1
timestamp 1698431365
transform -1 0 94976 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1006__A2
timestamp 1698431365
transform 1 0 100800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__I
timestamp 1698431365
transform -1 0 50288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1011__A2
timestamp 1698431365
transform 1 0 34608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__I
timestamp 1698431365
transform -1 0 93632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A2
timestamp 1698431365
transform -1 0 94416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A3
timestamp 1698431365
transform -1 0 98896 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__I
timestamp 1698431365
transform -1 0 29568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1018__A2
timestamp 1698431365
transform -1 0 33040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__A1
timestamp 1698431365
transform 1 0 25424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__A2
timestamp 1698431365
transform -1 0 29680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A2
timestamp 1698431365
transform -1 0 70224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A3
timestamp 1698431365
transform -1 0 69776 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A1
timestamp 1698431365
transform 1 0 51520 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A2
timestamp 1698431365
transform 1 0 51520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A3
timestamp 1698431365
transform 1 0 51968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A1
timestamp 1698431365
transform 1 0 43120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A2
timestamp 1698431365
transform -1 0 44240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A4
timestamp 1698431365
transform 1 0 44464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1028__A1
timestamp 1698431365
transform 1 0 37520 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1033__A2
timestamp 1698431365
transform 1 0 35280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A1
timestamp 1698431365
transform -1 0 49504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A2
timestamp 1698431365
transform -1 0 47488 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A3
timestamp 1698431365
transform 1 0 49728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A4
timestamp 1698431365
transform -1 0 54656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__A3
timestamp 1698431365
transform 1 0 70784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__A4
timestamp 1698431365
transform -1 0 66192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__A3
timestamp 1698431365
transform -1 0 51968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__I
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A1
timestamp 1698431365
transform 1 0 111776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A2
timestamp 1698431365
transform 1 0 114352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__A1
timestamp 1698431365
transform 1 0 93520 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__A2
timestamp 1698431365
transform -1 0 93296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__B
timestamp 1698431365
transform -1 0 93744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1045__I
timestamp 1698431365
transform 1 0 93520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__A2
timestamp 1698431365
transform -1 0 39984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__I0
timestamp 1698431365
transform 1 0 31360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__I1
timestamp 1698431365
transform -1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__S
timestamp 1698431365
transform -1 0 32256 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A1
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A2
timestamp 1698431365
transform 1 0 22512 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__A1
timestamp 1698431365
transform -1 0 41216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__B2
timestamp 1698431365
transform 1 0 30240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__I
timestamp 1698431365
transform 1 0 112112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__I
timestamp 1698431365
transform -1 0 36848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__C
timestamp 1698431365
transform -1 0 32256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__C
timestamp 1698431365
transform -1 0 30128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1072__C
timestamp 1698431365
transform -1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__B2
timestamp 1698431365
transform 1 0 34832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A1
timestamp 1698431365
transform 1 0 39648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__I
timestamp 1698431365
transform 1 0 50736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A1
timestamp 1698431365
transform 1 0 49728 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__B2
timestamp 1698431365
transform 1 0 39872 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__I
timestamp 1698431365
transform 1 0 43008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__A1
timestamp 1698431365
transform -1 0 47264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__B2
timestamp 1698431365
transform 1 0 46256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__A1
timestamp 1698431365
transform 1 0 49168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__A1
timestamp 1698431365
transform 1 0 50400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1089__I
timestamp 1698431365
transform 1 0 70336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__I
timestamp 1698431365
transform 1 0 71680 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__A1
timestamp 1698431365
transform -1 0 73024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__A2
timestamp 1698431365
transform -1 0 70672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A2
timestamp 1698431365
transform 1 0 73808 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__A2
timestamp 1698431365
transform 1 0 76272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__I
timestamp 1698431365
transform -1 0 79072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__I
timestamp 1698431365
transform 1 0 103712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__I
timestamp 1698431365
transform -1 0 103040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1109__A2
timestamp 1698431365
transform -1 0 85568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1111__I
timestamp 1698431365
transform 1 0 108640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1113__A2
timestamp 1698431365
transform 1 0 113008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__A2
timestamp 1698431365
transform 1 0 105280 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__A2
timestamp 1698431365
transform 1 0 104160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A1
timestamp 1698431365
transform 1 0 122304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1130__A1
timestamp 1698431365
transform 1 0 121632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A2
timestamp 1698431365
transform 1 0 119392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__I
timestamp 1698431365
transform 1 0 92848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__I
timestamp 1698431365
transform 1 0 64512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__A2
timestamp 1698431365
transform 1 0 60368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__I
timestamp 1698431365
transform 1 0 82096 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__I
timestamp 1698431365
transform 1 0 88480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__A1
timestamp 1698431365
transform 1 0 59472 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__I
timestamp 1698431365
transform 1 0 73696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__I
timestamp 1698431365
transform 1 0 94080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1168__I
timestamp 1698431365
transform -1 0 57232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A2
timestamp 1698431365
transform 1 0 59920 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__I
timestamp 1698431365
transform -1 0 63616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__B2
timestamp 1698431365
transform -1 0 91728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__C
timestamp 1698431365
transform 1 0 93520 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1177__I
timestamp 1698431365
transform 1 0 61040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1178__I
timestamp 1698431365
transform 1 0 85232 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1184__A2
timestamp 1698431365
transform -1 0 72576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1184__B1
timestamp 1698431365
transform 1 0 71008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1186__A2
timestamp 1698431365
transform 1 0 73472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1191__I
timestamp 1698431365
transform -1 0 92176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__B2
timestamp 1698431365
transform -1 0 94640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__C
timestamp 1698431365
transform 1 0 93968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1196__A2
timestamp 1698431365
transform 1 0 67760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1196__B1
timestamp 1698431365
transform 1 0 74256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1198__A2
timestamp 1698431365
transform 1 0 74368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1200__I
timestamp 1698431365
transform 1 0 97776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1201__I
timestamp 1698431365
transform 1 0 98336 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1203__I
timestamp 1698431365
transform 1 0 107632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__I
timestamp 1698431365
transform 1 0 55888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__I
timestamp 1698431365
transform 1 0 83104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__A2
timestamp 1698431365
transform 1 0 72800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__B1
timestamp 1698431365
transform 1 0 73248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1209__A2
timestamp 1698431365
transform -1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__I
timestamp 1698431365
transform 1 0 85456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1213__I
timestamp 1698431365
transform 1 0 73696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1214__A1
timestamp 1698431365
transform 1 0 84560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1214__B2
timestamp 1698431365
transform -1 0 83216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A1
timestamp 1698431365
transform -1 0 85904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A2
timestamp 1698431365
transform 1 0 86464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1217__A1
timestamp 1698431365
transform 1 0 95200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__I
timestamp 1698431365
transform 1 0 93520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1220__A1
timestamp 1698431365
transform -1 0 85232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1220__B1
timestamp 1698431365
transform -1 0 83664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1220__B2
timestamp 1698431365
transform 1 0 101360 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__A1
timestamp 1698431365
transform 1 0 86352 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__A2
timestamp 1698431365
transform 1 0 88032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1223__A1
timestamp 1698431365
transform 1 0 91056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1224__I
timestamp 1698431365
transform 1 0 93968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1226__A2
timestamp 1698431365
transform 1 0 64288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__I
timestamp 1698431365
transform 1 0 98784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1230__A1
timestamp 1698431365
transform 1 0 80304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1230__C2
timestamp 1698431365
transform 1 0 80752 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1232__A1
timestamp 1698431365
transform -1 0 85568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1232__A2
timestamp 1698431365
transform -1 0 85120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1235__I
timestamp 1698431365
transform 1 0 65408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__A1
timestamp 1698431365
transform -1 0 79520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__C1
timestamp 1698431365
transform 1 0 79072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__C2
timestamp 1698431365
transform -1 0 78848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__A1
timestamp 1698431365
transform 1 0 86912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__A2
timestamp 1698431365
transform 1 0 84112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1241__I
timestamp 1698431365
transform 1 0 43568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1244__C1
timestamp 1698431365
transform 1 0 74144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1244__C2
timestamp 1698431365
transform 1 0 74592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__I
timestamp 1698431365
transform 1 0 49616 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1247__S0
timestamp 1698431365
transform -1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1247__S1
timestamp 1698431365
transform -1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1248__A1
timestamp 1698431365
transform 1 0 61712 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1248__A2
timestamp 1698431365
transform 1 0 59920 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1252__A2
timestamp 1698431365
transform 1 0 63168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__A1
timestamp 1698431365
transform 1 0 63616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1261__A2
timestamp 1698431365
transform 1 0 72352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__I
timestamp 1698431365
transform 1 0 108304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__I
timestamp 1698431365
transform 1 0 76832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__A1
timestamp 1698431365
transform 1 0 73360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1269__I
timestamp 1698431365
transform 1 0 107856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__I
timestamp 1698431365
transform 1 0 73584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__B
timestamp 1698431365
transform 1 0 110880 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1272__A2
timestamp 1698431365
transform 1 0 113904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__A1
timestamp 1698431365
transform 1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__B
timestamp 1698431365
transform 1 0 109424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1275__A2
timestamp 1698431365
transform -1 0 108752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1276__I
timestamp 1698431365
transform 1 0 87248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1277__A1
timestamp 1698431365
transform 1 0 90272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1277__A2
timestamp 1698431365
transform -1 0 89040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1278__B
timestamp 1698431365
transform 1 0 112336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1279__A2
timestamp 1698431365
transform -1 0 111104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A1
timestamp 1698431365
transform 1 0 101808 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A2
timestamp 1698431365
transform -1 0 100576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1281__I
timestamp 1698431365
transform 1 0 105728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1283__A2
timestamp 1698431365
transform 1 0 108640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1284__I
timestamp 1698431365
transform 1 0 104944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1285__A1
timestamp 1698431365
transform -1 0 107408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1285__A2
timestamp 1698431365
transform -1 0 106176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__I
timestamp 1698431365
transform 1 0 107184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1288__A2
timestamp 1698431365
transform 1 0 107520 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1289__A1
timestamp 1698431365
transform 1 0 108640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1289__A2
timestamp 1698431365
transform -1 0 107632 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__A2
timestamp 1698431365
transform 1 0 108864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1292__I
timestamp 1698431365
transform 1 0 86128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1293__A1
timestamp 1698431365
transform -1 0 107184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1293__A2
timestamp 1698431365
transform 1 0 105504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__A2
timestamp 1698431365
transform 1 0 106960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A1
timestamp 1698431365
transform 1 0 105728 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A2
timestamp 1698431365
transform 1 0 104496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__I
timestamp 1698431365
transform 1 0 103040 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1299__A2
timestamp 1698431365
transform 1 0 105392 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1302__A2
timestamp 1698431365
transform 1 0 74704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1307__A1
timestamp 1698431365
transform 1 0 92624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1309__A1
timestamp 1698431365
transform 1 0 91280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1311__A1
timestamp 1698431365
transform 1 0 90272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1313__I
timestamp 1698431365
transform 1 0 87136 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1315__A1
timestamp 1698431365
transform 1 0 87360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__A1
timestamp 1698431365
transform 1 0 85792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1319__A1
timestamp 1698431365
transform 1 0 86352 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__A1
timestamp 1698431365
transform -1 0 88704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1321__A1
timestamp 1698431365
transform 1 0 88704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__A1
timestamp 1698431365
transform 1 0 86240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1323__A1
timestamp 1698431365
transform 1 0 85680 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1324__I
timestamp 1698431365
transform 1 0 92176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1325__A1
timestamp 1698431365
transform 1 0 92400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1326__A1
timestamp 1698431365
transform 1 0 91952 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1331__I
timestamp 1698431365
transform 1 0 95200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1332__I
timestamp 1698431365
transform 1 0 95200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1334__A1
timestamp 1698431365
transform 1 0 97440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1336__A1
timestamp 1698431365
transform -1 0 95872 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A1
timestamp 1698431365
transform -1 0 95424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1339__I
timestamp 1698431365
transform -1 0 93744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1341__A1
timestamp 1698431365
transform -1 0 96320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__I
timestamp 1698431365
transform 1 0 99680 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__I
timestamp 1698431365
transform -1 0 99680 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__A1
timestamp 1698431365
transform 1 0 100800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1347__A1
timestamp 1698431365
transform -1 0 107296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__A1
timestamp 1698431365
transform -1 0 102592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1350__I
timestamp 1698431365
transform -1 0 92400 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__B
timestamp 1698431365
transform 1 0 100240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1352__A1
timestamp 1698431365
transform -1 0 102592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1353__I
timestamp 1698431365
transform 1 0 45920 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1355__A1
timestamp 1698431365
transform 1 0 42112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1355__A3
timestamp 1698431365
transform -1 0 42784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A2
timestamp 1698431365
transform 1 0 44912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A3
timestamp 1698431365
transform -1 0 46480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__A2
timestamp 1698431365
transform 1 0 48160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1360__I
timestamp 1698431365
transform -1 0 73472 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1361__I
timestamp 1698431365
transform 1 0 73920 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A2
timestamp 1698431365
transform -1 0 47824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1365__I
timestamp 1698431365
transform -1 0 60816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1367__A1
timestamp 1698431365
transform 1 0 61264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__I
timestamp 1698431365
transform 1 0 67760 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__I
timestamp 1698431365
transform 1 0 62720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__I
timestamp 1698431365
transform 1 0 88032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A2
timestamp 1698431365
transform 1 0 77168 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__B
timestamp 1698431365
transform 1 0 77616 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1377__A1
timestamp 1698431365
transform -1 0 72128 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1377__A2
timestamp 1698431365
transform 1 0 72464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__A2
timestamp 1698431365
transform 1 0 77952 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__B
timestamp 1698431365
transform 1 0 78400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__A1
timestamp 1698431365
transform -1 0 74928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__A2
timestamp 1698431365
transform 1 0 74256 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1382__A1
timestamp 1698431365
transform 1 0 62944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A1
timestamp 1698431365
transform 1 0 63392 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1387__I
timestamp 1698431365
transform -1 0 47936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1388__I
timestamp 1698431365
transform 1 0 62272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1390__A1
timestamp 1698431365
transform -1 0 59584 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A1
timestamp 1698431365
transform -1 0 64064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1393__A1
timestamp 1698431365
transform 1 0 63280 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1396__A1
timestamp 1698431365
transform -1 0 64960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__A1
timestamp 1698431365
transform 1 0 66192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__I
timestamp 1698431365
transform -1 0 67088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__I
timestamp 1698431365
transform 1 0 66416 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1405__A1
timestamp 1698431365
transform -1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1413__I
timestamp 1698431365
transform -1 0 74032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__I
timestamp 1698431365
transform 1 0 75600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A2
timestamp 1698431365
transform 1 0 69328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1418__A2
timestamp 1698431365
transform 1 0 68096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__I
timestamp 1698431365
transform 1 0 71680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__A2
timestamp 1698431365
transform -1 0 73472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1422__A1
timestamp 1698431365
transform 1 0 71232 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1422__A2
timestamp 1698431365
transform 1 0 69776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1424__A2
timestamp 1698431365
transform 1 0 98672 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__A1
timestamp 1698431365
transform 1 0 92400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__A2
timestamp 1698431365
transform -1 0 85232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1428__B
timestamp 1698431365
transform 1 0 85904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A2
timestamp 1698431365
transform 1 0 90384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__B
timestamp 1698431365
transform 1 0 91952 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1430__A2
timestamp 1698431365
transform 1 0 89040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A2
timestamp 1698431365
transform -1 0 95312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1432__I
timestamp 1698431365
transform 1 0 90048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1434__B
timestamp 1698431365
transform 1 0 92400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__A2
timestamp 1698431365
transform 1 0 99120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__B
timestamp 1698431365
transform 1 0 99792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__I
timestamp 1698431365
transform -1 0 82768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__B
timestamp 1698431365
transform 1 0 87360 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1443__A1
timestamp 1698431365
transform 1 0 95312 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1447__I
timestamp 1698431365
transform -1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1448__A1
timestamp 1698431365
transform -1 0 66304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1448__A2
timestamp 1698431365
transform -1 0 79072 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__A1
timestamp 1698431365
transform -1 0 86352 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__A2
timestamp 1698431365
transform 1 0 83440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A1
timestamp 1698431365
transform 1 0 62608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A2
timestamp 1698431365
transform -1 0 60368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A3
timestamp 1698431365
transform 1 0 64512 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A1
timestamp 1698431365
transform 1 0 66640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1458__A1
timestamp 1698431365
transform 1 0 63840 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__A1
timestamp 1698431365
transform 1 0 74256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__A2
timestamp 1698431365
transform -1 0 74928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__A1
timestamp 1698431365
transform 1 0 73696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__A2
timestamp 1698431365
transform 1 0 74144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__A2
timestamp 1698431365
transform 1 0 63280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1464__A1
timestamp 1698431365
transform 1 0 66416 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__B
timestamp 1698431365
transform -1 0 65408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1471__A2
timestamp 1698431365
transform 1 0 62384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__A1
timestamp 1698431365
transform -1 0 46144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__A2
timestamp 1698431365
transform -1 0 46592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1474__A2
timestamp 1698431365
transform -1 0 24304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A1
timestamp 1698431365
transform -1 0 26432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A2
timestamp 1698431365
transform 1 0 27104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__C
timestamp 1698431365
transform 1 0 26656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1480__A1
timestamp 1698431365
transform 1 0 71232 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A1
timestamp 1698431365
transform 1 0 71680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1485__A1
timestamp 1698431365
transform -1 0 71120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__B
timestamp 1698431365
transform 1 0 68432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__A1
timestamp 1698431365
transform 1 0 71680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__A1
timestamp 1698431365
transform 1 0 72016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__A2
timestamp 1698431365
transform 1 0 71568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__A1
timestamp 1698431365
transform 1 0 65072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__A1
timestamp 1698431365
transform -1 0 41888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__A3
timestamp 1698431365
transform 1 0 42560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__A1
timestamp 1698431365
transform 1 0 41664 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__A1
timestamp 1698431365
transform 1 0 75600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__A1
timestamp 1698431365
transform 1 0 75376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__A1
timestamp 1698431365
transform 1 0 79296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1509__A1
timestamp 1698431365
transform 1 0 79520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__A1
timestamp 1698431365
transform 1 0 84448 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1515__A1
timestamp 1698431365
transform 1 0 84000 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__B
timestamp 1698431365
transform 1 0 79968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1518__A1
timestamp 1698431365
transform -1 0 83328 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__B
timestamp 1698431365
transform 1 0 80864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A1
timestamp 1698431365
transform 1 0 81984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A1
timestamp 1698431365
transform 1 0 31808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A2
timestamp 1698431365
transform -1 0 36288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A1
timestamp 1698431365
transform -1 0 34160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A2
timestamp 1698431365
transform -1 0 35056 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__B
timestamp 1698431365
transform 1 0 34832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1533__B
timestamp 1698431365
transform 1 0 33376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1538__C
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__B
timestamp 1698431365
transform -1 0 34384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1545__B
timestamp 1698431365
transform 1 0 24304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1549__B
timestamp 1698431365
transform 1 0 35616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__I
timestamp 1698431365
transform -1 0 30128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__B
timestamp 1698431365
transform -1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1565__A1
timestamp 1698431365
transform 1 0 38976 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__B
timestamp 1698431365
transform 1 0 37968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__B
timestamp 1698431365
transform 1 0 38528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__A1
timestamp 1698431365
transform 1 0 29792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__I
timestamp 1698431365
transform 1 0 43568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__A1
timestamp 1698431365
transform 1 0 25200 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__A2
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__A1
timestamp 1698431365
transform -1 0 29680 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__I
timestamp 1698431365
transform 1 0 46256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__A1
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A1
timestamp 1698431365
transform -1 0 35616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__I
timestamp 1698431365
transform 1 0 23296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A1
timestamp 1698431365
transform -1 0 22400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1604__A1
timestamp 1698431365
transform 1 0 24528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A1
timestamp 1698431365
transform 1 0 23520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__A1
timestamp 1698431365
transform -1 0 24528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__I
timestamp 1698431365
transform 1 0 51856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__B
timestamp 1698431365
transform -1 0 54544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A1
timestamp 1698431365
transform 1 0 51632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__B
timestamp 1698431365
transform -1 0 52976 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__A1
timestamp 1698431365
transform 1 0 52080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__I
timestamp 1698431365
transform -1 0 52640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__A1
timestamp 1698431365
transform 1 0 52304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__A2
timestamp 1698431365
transform 1 0 51632 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__I
timestamp 1698431365
transform -1 0 51296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A1
timestamp 1698431365
transform -1 0 53872 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__B
timestamp 1698431365
transform -1 0 53424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A1
timestamp 1698431365
transform -1 0 57568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__I
timestamp 1698431365
transform 1 0 39424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1629__A1
timestamp 1698431365
transform 1 0 57568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1629__B
timestamp 1698431365
transform 1 0 58016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__I
timestamp 1698431365
transform -1 0 44352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__B
timestamp 1698431365
transform 1 0 62944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__A1
timestamp 1698431365
transform -1 0 58688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__A1
timestamp 1698431365
transform 1 0 49728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__A2
timestamp 1698431365
transform -1 0 50400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1638__A1
timestamp 1698431365
transform -1 0 62608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1638__B
timestamp 1698431365
transform 1 0 62832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__A1
timestamp 1698431365
transform -1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__I
timestamp 1698431365
transform -1 0 69104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__A2
timestamp 1698431365
transform 1 0 56000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A2
timestamp 1698431365
transform -1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__I
timestamp 1698431365
transform -1 0 68656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__I
timestamp 1698431365
transform -1 0 73248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A2
timestamp 1698431365
transform -1 0 57120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I
timestamp 1698431365
transform 1 0 63728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A1
timestamp 1698431365
transform -1 0 69104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A2
timestamp 1698431365
transform 1 0 67648 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A1
timestamp 1698431365
transform -1 0 67536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1698431365
transform 1 0 68432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__I
timestamp 1698431365
transform -1 0 78288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A2
timestamp 1698431365
transform 1 0 74256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A2
timestamp 1698431365
transform -1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__I
timestamp 1698431365
transform 1 0 97776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A2
timestamp 1698431365
transform -1 0 85120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__I
timestamp 1698431365
transform 1 0 74816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A2
timestamp 1698431365
transform 1 0 93072 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__I
timestamp 1698431365
transform 1 0 109984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A2
timestamp 1698431365
transform -1 0 89376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A2
timestamp 1698431365
transform 1 0 98224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__I
timestamp 1698431365
transform 1 0 109088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A2
timestamp 1698431365
transform 1 0 116032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__I
timestamp 1698431365
transform 1 0 112560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A2
timestamp 1698431365
transform 1 0 117152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__I
timestamp 1698431365
transform 1 0 121856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__I
timestamp 1698431365
transform 1 0 117600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__I
timestamp 1698431365
transform 1 0 113344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__A1
timestamp 1698431365
transform 1 0 116368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__I
timestamp 1698431365
transform 1 0 112112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A1
timestamp 1698431365
transform 1 0 115920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__I
timestamp 1698431365
transform 1 0 109872 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__A1
timestamp 1698431365
transform -1 0 112784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__I
timestamp 1698431365
transform 1 0 111552 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__A1
timestamp 1698431365
transform 1 0 111664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__A1
timestamp 1698431365
transform -1 0 118720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__A1
timestamp 1698431365
transform 1 0 106624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__I
timestamp 1698431365
transform 1 0 110768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__A1
timestamp 1698431365
transform 1 0 112448 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A1
timestamp 1698431365
transform -1 0 114128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__I
timestamp 1698431365
transform -1 0 95088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__A2
timestamp 1698431365
transform 1 0 98224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A1
timestamp 1698431365
transform 1 0 112896 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__I
timestamp 1698431365
transform 1 0 94864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__B
timestamp 1698431365
transform -1 0 94528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__A2
timestamp 1698431365
transform 1 0 100240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__A1
timestamp 1698431365
transform -1 0 103936 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__B
timestamp 1698431365
transform 1 0 109536 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__A2
timestamp 1698431365
transform 1 0 49280 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__I
timestamp 1698431365
transform -1 0 43904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__A1
timestamp 1698431365
transform -1 0 39088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__A2
timestamp 1698431365
transform -1 0 47264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__B
timestamp 1698431365
transform -1 0 49504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A2
timestamp 1698431365
transform 1 0 49616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__A1
timestamp 1698431365
transform -1 0 47824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__B
timestamp 1698431365
transform 1 0 51184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A2
timestamp 1698431365
transform 1 0 47488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__A1
timestamp 1698431365
transform -1 0 43792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1744__A2
timestamp 1698431365
transform -1 0 45584 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A1
timestamp 1698431365
transform 1 0 49392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__A1
timestamp 1698431365
transform 1 0 48832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__A1
timestamp 1698431365
transform -1 0 54208 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__A2
timestamp 1698431365
transform 1 0 55104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A1
timestamp 1698431365
transform -1 0 51856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A2
timestamp 1698431365
transform 1 0 53536 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A3
timestamp 1698431365
transform -1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__I
timestamp 1698431365
transform 1 0 49840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__A1
timestamp 1698431365
transform 1 0 57792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__A1
timestamp 1698431365
transform 1 0 57792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__A1
timestamp 1698431365
transform 1 0 54320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__I
timestamp 1698431365
transform -1 0 43120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A2
timestamp 1698431365
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__A1
timestamp 1698431365
transform 1 0 46816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A1
timestamp 1698431365
transform -1 0 51856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__B1
timestamp 1698431365
transform -1 0 51184 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A2
timestamp 1698431365
transform -1 0 48720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__A1
timestamp 1698431365
transform 1 0 49840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A1
timestamp 1698431365
transform 1 0 44128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A2
timestamp 1698431365
transform 1 0 45696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A1
timestamp 1698431365
transform 1 0 52304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A2
timestamp 1698431365
transform 1 0 51856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__A2
timestamp 1698431365
transform 1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A1
timestamp 1698431365
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A2
timestamp 1698431365
transform 1 0 49504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__C
timestamp 1698431365
transform -1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__B2
timestamp 1698431365
transform 1 0 53984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__A2
timestamp 1698431365
transform -1 0 43568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__I
timestamp 1698431365
transform 1 0 38976 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__A2
timestamp 1698431365
transform -1 0 40432 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A4
timestamp 1698431365
transform 1 0 44576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__B
timestamp 1698431365
transform 1 0 48160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__A1
timestamp 1698431365
transform 1 0 51296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A1
timestamp 1698431365
transform -1 0 70784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A2
timestamp 1698431365
transform 1 0 68992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__A1
timestamp 1698431365
transform 1 0 50288 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__B2
timestamp 1698431365
transform 1 0 52752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__A1
timestamp 1698431365
transform 1 0 51744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__C
timestamp 1698431365
transform 1 0 51632 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A1
timestamp 1698431365
transform 1 0 52304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A1
timestamp 1698431365
transform 1 0 53648 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__A1
timestamp 1698431365
transform -1 0 50960 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A1
timestamp 1698431365
transform -1 0 54768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A2
timestamp 1698431365
transform 1 0 59360 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__B2
timestamp 1698431365
transform 1 0 52752 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A1
timestamp 1698431365
transform 1 0 37968 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__B
timestamp 1698431365
transform -1 0 40544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__B
timestamp 1698431365
transform 1 0 43008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A2
timestamp 1698431365
transform 1 0 48832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__A1
timestamp 1698431365
transform 1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__C
timestamp 1698431365
transform 1 0 67536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__A2
timestamp 1698431365
transform 1 0 58240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A1
timestamp 1698431365
transform -1 0 58912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A1
timestamp 1698431365
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__I
timestamp 1698431365
transform 1 0 33600 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A1
timestamp 1698431365
transform -1 0 50064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A3
timestamp 1698431365
transform 1 0 49280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A1
timestamp 1698431365
transform 1 0 45024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A1
timestamp 1698431365
transform -1 0 59472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__B
timestamp 1698431365
transform 1 0 59360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A1
timestamp 1698431365
transform 1 0 31584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A3
timestamp 1698431365
transform 1 0 25536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A4
timestamp 1698431365
transform -1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A1
timestamp 1698431365
transform -1 0 26096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A3
timestamp 1698431365
transform -1 0 39536 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__I
timestamp 1698431365
transform -1 0 19824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__I
timestamp 1698431365
transform 1 0 19600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A1
timestamp 1698431365
transform -1 0 18256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__I
timestamp 1698431365
transform 1 0 20272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__I
timestamp 1698431365
transform 1 0 35728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__A1
timestamp 1698431365
transform -1 0 18704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__A2
timestamp 1698431365
transform -1 0 21056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A1
timestamp 1698431365
transform -1 0 21504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__I
timestamp 1698431365
transform 1 0 22064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__A1
timestamp 1698431365
transform 1 0 22848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A1
timestamp 1698431365
transform 1 0 22512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A2
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__A1
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A1
timestamp 1698431365
transform -1 0 21952 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__A2
timestamp 1698431365
transform -1 0 21168 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1939__A1
timestamp 1698431365
transform 1 0 23520 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1941__I
timestamp 1698431365
transform 1 0 26544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__A1
timestamp 1698431365
transform 1 0 26096 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__A1
timestamp 1698431365
transform 1 0 26208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A1
timestamp 1698431365
transform 1 0 26096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A3
timestamp 1698431365
transform -1 0 39088 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__A1
timestamp 1698431365
transform 1 0 33488 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__A1
timestamp 1698431365
transform -1 0 31248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__I
timestamp 1698431365
transform -1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A1
timestamp 1698431365
transform 1 0 42560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__A1
timestamp 1698431365
transform -1 0 39424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__A1
timestamp 1698431365
transform 1 0 38752 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__A1
timestamp 1698431365
transform 1 0 45808 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A1
timestamp 1698431365
transform -1 0 19712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__I
timestamp 1698431365
transform 1 0 16352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__A1
timestamp 1698431365
transform -1 0 19152 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A1
timestamp 1698431365
transform 1 0 20944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A1
timestamp 1698431365
transform 1 0 22400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__A1
timestamp 1698431365
transform 1 0 22848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A1
timestamp 1698431365
transform -1 0 22064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__A1
timestamp 1698431365
transform 1 0 40992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__CLKN
timestamp 1698431365
transform 1 0 111552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__CLKN
timestamp 1698431365
transform 1 0 107968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__CLKN
timestamp 1698431365
transform 1 0 111888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__CLKN
timestamp 1698431365
transform 1 0 108864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__CLKN
timestamp 1698431365
transform 1 0 106960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__CLKN
timestamp 1698431365
transform 1 0 109760 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__CLKN
timestamp 1698431365
transform 1 0 104944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__CLKN
timestamp 1698431365
transform 1 0 103264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1999__CLKN
timestamp 1698431365
transform 1 0 96432 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__CLKN
timestamp 1698431365
transform 1 0 93744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__CLKN
timestamp 1698431365
transform -1 0 93296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__CLKN
timestamp 1698431365
transform 1 0 85232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__CLKN
timestamp 1698431365
transform 1 0 87360 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__CLKN
timestamp 1698431365
transform 1 0 91168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__CLKN
timestamp 1698431365
transform 1 0 88704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__CLKN
timestamp 1698431365
transform 1 0 93632 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__CLKN
timestamp 1698431365
transform 1 0 101808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__CLKN
timestamp 1698431365
transform 1 0 99120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2009__CLKN
timestamp 1698431365
transform 1 0 98672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__CLKN
timestamp 1698431365
transform 1 0 99792 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__CLKN
timestamp 1698431365
transform 1 0 103040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__CLKN
timestamp 1698431365
transform 1 0 106288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__CLKN
timestamp 1698431365
transform 1 0 107072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__CLKN
timestamp 1698431365
transform 1 0 104832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__CLK
timestamp 1698431365
transform 1 0 46032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__CLK
timestamp 1698431365
transform -1 0 72464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__CLK
timestamp 1698431365
transform 1 0 75712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__CLK
timestamp 1698431365
transform 1 0 78400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__CLK
timestamp 1698431365
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__CLK
timestamp 1698431365
transform 1 0 71456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__CLK
timestamp 1698431365
transform 1 0 64064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__CLK
timestamp 1698431365
transform 1 0 63280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__CLK
timestamp 1698431365
transform 1 0 69104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__CLK
timestamp 1698431365
transform 1 0 63392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__CLK
timestamp 1698431365
transform 1 0 64848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__CLK
timestamp 1698431365
transform 1 0 69552 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2027__CLK
timestamp 1698431365
transform 1 0 68432 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__CLK
timestamp 1698431365
transform 1 0 74704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__CLK
timestamp 1698431365
transform 1 0 72352 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__CLK
timestamp 1698431365
transform 1 0 89600 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__CLK
timestamp 1698431365
transform -1 0 88480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__CLK
timestamp 1698431365
transform 1 0 98784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2033__CLK
timestamp 1698431365
transform 1 0 98672 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2034__CLK
timestamp 1698431365
transform 1 0 87248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__CLK
timestamp 1698431365
transform 1 0 83552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__CLK
timestamp 1698431365
transform -1 0 86016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__CLK
timestamp 1698431365
transform 1 0 81872 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__CLK
timestamp 1698431365
transform 1 0 79520 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2039__CLK
timestamp 1698431365
transform 1 0 62832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__CLK
timestamp 1698431365
transform 1 0 71680 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__CLKN
timestamp 1698431365
transform 1 0 62608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__CLKN
timestamp 1698431365
transform 1 0 26880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__CLKN
timestamp 1698431365
transform 1 0 79632 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2044__CLKN
timestamp 1698431365
transform -1 0 70672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__CLKN
timestamp 1698431365
transform 1 0 64400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__CLK
timestamp 1698431365
transform -1 0 39536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__CLKN
timestamp 1698431365
transform 1 0 75600 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2048__CLKN
timestamp 1698431365
transform 1 0 75600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__CLKN
timestamp 1698431365
transform 1 0 80192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__CLKN
timestamp 1698431365
transform 1 0 80864 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2051__CLKN
timestamp 1698431365
transform 1 0 84112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__CLKN
timestamp 1698431365
transform 1 0 84896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__CLKN
timestamp 1698431365
transform 1 0 79296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2054__CLKN
timestamp 1698431365
transform 1 0 79744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__CLK
timestamp 1698431365
transform 1 0 36624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__CLK
timestamp 1698431365
transform 1 0 34384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2057__CLK
timestamp 1698431365
transform 1 0 24528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__CLK
timestamp 1698431365
transform -1 0 35504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__CLK
timestamp 1698431365
transform 1 0 33040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2060__CLK
timestamp 1698431365
transform 1 0 30128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__CLK
timestamp 1698431365
transform 1 0 30464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__CLK
timestamp 1698431365
transform -1 0 30688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__CLK
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__CLK
timestamp 1698431365
transform 1 0 40320 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__CLK
timestamp 1698431365
transform 1 0 30016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2066__CLK
timestamp 1698431365
transform 1 0 44240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2067__CLK
timestamp 1698431365
transform 1 0 36960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2068__CLK
timestamp 1698431365
transform 1 0 44240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2069__CLK
timestamp 1698431365
transform 1 0 28784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2070__CLK
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__CLK
timestamp 1698431365
transform 1 0 25872 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__CLK
timestamp 1698431365
transform 1 0 22400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__CLK
timestamp 1698431365
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2075__CLK
timestamp 1698431365
transform 1 0 55888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__CLK
timestamp 1698431365
transform 1 0 50624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__CLK
timestamp 1698431365
transform 1 0 59472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__CLK
timestamp 1698431365
transform 1 0 58688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__CLK
timestamp 1698431365
transform 1 0 54096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__CLK
timestamp 1698431365
transform 1 0 57792 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2081__CLK
timestamp 1698431365
transform 1 0 58912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2082__CLK
timestamp 1698431365
transform 1 0 48832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2083__CLK
timestamp 1698431365
transform -1 0 58352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__CLK
timestamp 1698431365
transform -1 0 58800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__CLK
timestamp 1698431365
transform -1 0 60816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2086__CLK
timestamp 1698431365
transform 1 0 65408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__CLK
timestamp 1698431365
transform 1 0 69104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__CLK
timestamp 1698431365
transform 1 0 84448 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2089__CLK
timestamp 1698431365
transform -1 0 85456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__CLK
timestamp 1698431365
transform 1 0 84000 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__CLK
timestamp 1698431365
transform 1 0 90832 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2092__CLK
timestamp 1698431365
transform 1 0 110320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2093__CLK
timestamp 1698431365
transform 1 0 108192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2094__CLK
timestamp 1698431365
transform 1 0 111216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__CLK
timestamp 1698431365
transform 1 0 114800 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2096__CLK
timestamp 1698431365
transform 1 0 114352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2097__CLK
timestamp 1698431365
transform 1 0 118720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__CLK
timestamp 1698431365
transform 1 0 119840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2099__CLK
timestamp 1698431365
transform 1 0 113792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__CLK
timestamp 1698431365
transform 1 0 118272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2101__CLK
timestamp 1698431365
transform 1 0 118720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__CLK
timestamp 1698431365
transform 1 0 116704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2103__CLK
timestamp 1698431365
transform 1 0 113456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2104__CLK
timestamp 1698431365
transform -1 0 100016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2105__CLK
timestamp 1698431365
transform -1 0 99344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2106__CLK
timestamp 1698431365
transform 1 0 47152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2107__CLK
timestamp 1698431365
transform 1 0 51072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2108__CLK
timestamp 1698431365
transform 1 0 47712 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2109__CLK
timestamp 1698431365
transform 1 0 42112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__CLK
timestamp 1698431365
transform -1 0 48720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2111__CLK
timestamp 1698431365
transform 1 0 53984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2112__CLK
timestamp 1698431365
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2113__CLK
timestamp 1698431365
transform 1 0 54096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__CLK
timestamp 1698431365
transform 1 0 52752 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__CLKN
timestamp 1698431365
transform 1 0 47264 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2116__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__CLK
timestamp 1698431365
transform 1 0 71568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__CLK
timestamp 1698431365
transform 1 0 58688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__CLK
timestamp 1698431365
transform 1 0 68320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2120__CLK
timestamp 1698431365
transform 1 0 67760 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2121__CLK
timestamp 1698431365
transform 1 0 59808 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__CLK
timestamp 1698431365
transform -1 0 18928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__CLK
timestamp 1698431365
transform 1 0 20384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__CLK
timestamp 1698431365
transform -1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__CLK
timestamp 1698431365
transform -1 0 20496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__CLK
timestamp 1698431365
transform 1 0 25312 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__CLK
timestamp 1698431365
transform -1 0 28896 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__CLK
timestamp 1698431365
transform 1 0 25648 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__CLK
timestamp 1698431365
transform 1 0 29232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__CLK
timestamp 1698431365
transform 1 0 34384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2133__CLK
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2134__CLK
timestamp 1698431365
transform 1 0 38416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2135__CLK
timestamp 1698431365
transform 1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2136__CLK
timestamp 1698431365
transform 1 0 46816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__CLK
timestamp 1698431365
transform 1 0 37072 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__CLK
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__CLK
timestamp 1698431365
transform -1 0 18592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__CLK
timestamp 1698431365
transform 1 0 20048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2141__CLK
timestamp 1698431365
transform 1 0 23408 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__CLK
timestamp 1698431365
transform 1 0 23856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2143__CLK
timestamp 1698431365
transform 1 0 20384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2144__CLK
timestamp 1698431365
transform 1 0 22848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__CLK
timestamp 1698431365
transform 1 0 35728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__I
timestamp 1698431365
transform 1 0 71456 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2151__I
timestamp 1698431365
transform 1 0 81088 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2152__I
timestamp 1698431365
transform 1 0 92512 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__I
timestamp 1698431365
transform 1 0 103936 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__I
timestamp 1698431365
transform -1 0 116704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2155__I
timestamp 1698431365
transform 1 0 126784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__I
timestamp 1698431365
transform 1 0 138320 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 66304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 36176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 55104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 36064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 53984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 81312 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 102704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 76608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 94752 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout138_I
timestamp 1698431365
transform -1 0 69888 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout139_I
timestamp 1698431365
transform -1 0 115808 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold22_I
timestamp 1698431365
transform -1 0 17920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold27_I
timestamp 1698431365
transform -1 0 20720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold38_I
timestamp 1698431365
transform 1 0 130368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold41_I
timestamp 1698431365
transform -1 0 48272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold42_I
timestamp 1698431365
transform -1 0 67648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold44_I
timestamp 1698431365
transform -1 0 133616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold45_I
timestamp 1698431365
transform -1 0 30016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold48_I
timestamp 1698431365
transform -1 0 26656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold49_I
timestamp 1698431365
transform -1 0 17920 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold51_I
timestamp 1698431365
transform -1 0 26096 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold52_I
timestamp 1698431365
transform -1 0 137536 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold53_I
timestamp 1698431365
transform -1 0 47040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold54_I
timestamp 1698431365
transform -1 0 29232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold55_I
timestamp 1698431365
transform -1 0 142800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold56_I
timestamp 1698431365
transform -1 0 149296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold57_I
timestamp 1698431365
transform -1 0 18704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold58_I
timestamp 1698431365
transform 1 0 147504 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold59_I
timestamp 1698431365
transform -1 0 45136 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold60_I
timestamp 1698431365
transform -1 0 38864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold61_I
timestamp 1698431365
transform -1 0 40432 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold62_I
timestamp 1698431365
transform -1 0 18144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold63_I
timestamp 1698431365
transform 1 0 121632 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold65_I
timestamp 1698431365
transform 1 0 68880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold66_I
timestamp 1698431365
transform 1 0 120288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold67_I
timestamp 1698431365
transform -1 0 143920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold69_I
timestamp 1698431365
transform 1 0 116480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold70_I
timestamp 1698431365
transform -1 0 51632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold71_I
timestamp 1698431365
transform 1 0 117824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold72_I
timestamp 1698431365
transform 1 0 96880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold73_I
timestamp 1698431365
transform -1 0 47488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold74_I
timestamp 1698431365
transform -1 0 68656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold75_I
timestamp 1698431365
transform -1 0 23520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold76_I
timestamp 1698431365
transform 1 0 85904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold77_I
timestamp 1698431365
transform -1 0 90832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold78_I
timestamp 1698431365
transform -1 0 85680 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold79_I
timestamp 1698431365
transform 1 0 43456 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold80_I
timestamp 1698431365
transform -1 0 45696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold81_I
timestamp 1698431365
transform -1 0 62720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold82_I
timestamp 1698431365
transform 1 0 61712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold83_I
timestamp 1698431365
transform -1 0 99344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold84_I
timestamp 1698431365
transform 1 0 112000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold87_I
timestamp 1698431365
transform -1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold88_I
timestamp 1698431365
transform -1 0 28784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold89_I
timestamp 1698431365
transform 1 0 113008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold90_I
timestamp 1698431365
transform -1 0 26208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold91_I
timestamp 1698431365
transform -1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold92_I
timestamp 1698431365
transform 1 0 118048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold93_I
timestamp 1698431365
transform -1 0 67312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold94_I
timestamp 1698431365
transform 1 0 85792 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold95_I
timestamp 1698431365
transform -1 0 122640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold96_I
timestamp 1698431365
transform -1 0 51744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold97_I
timestamp 1698431365
transform 1 0 116928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold98_I
timestamp 1698431365
transform 1 0 63840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold99_I
timestamp 1698431365
transform -1 0 86576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold100_I
timestamp 1698431365
transform 1 0 92624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold101_I
timestamp 1698431365
transform -1 0 74368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold102_I
timestamp 1698431365
transform -1 0 127792 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold104_I
timestamp 1698431365
transform 1 0 106960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold105_I
timestamp 1698431365
transform 1 0 112000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold106_I
timestamp 1698431365
transform -1 0 125888 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold107_I
timestamp 1698431365
transform -1 0 68656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold108_I
timestamp 1698431365
transform 1 0 119168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold109_I
timestamp 1698431365
transform 1 0 105728 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold110_I
timestamp 1698431365
transform 1 0 120848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 123760 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 135184 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 146832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 55216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 66640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 78064 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 89488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 100912 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 112336 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 10640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 123872 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 132384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 135968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 144144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 147728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 13328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1698431365
transform 1 0 17472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1698431365
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output85_I
timestamp 1698431365
transform -1 0 149856 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output86_I
timestamp 1698431365
transform 1 0 62160 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output92_I
timestamp 1698431365
transform -1 0 21056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output93_I
timestamp 1698431365
transform 1 0 131152 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output94_I
timestamp 1698431365
transform 1 0 142576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output95_I
timestamp 1698431365
transform 1 0 154000 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output97_I
timestamp 1698431365
transform -1 0 43904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output100_I
timestamp 1698431365
transform 1 0 77168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output101_I
timestamp 1698431365
transform 1 0 88592 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output102_I
timestamp 1698431365
transform 1 0 96880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output103_I
timestamp 1698431365
transform 1 0 108304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output104_I
timestamp 1698431365
transform 1 0 119728 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output105_I
timestamp 1698431365
transform 1 0 15008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output125_I
timestamp 1698431365
transform 1 0 135072 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output126_I
timestamp 1698431365
transform 1 0 139552 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output127_I
timestamp 1698431365
transform 1 0 143584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output129_I
timestamp 1698431365
transform 1 0 146160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output130_I
timestamp 1698431365
transform -1 0 149856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 66304 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_3_0_0_wb_clk_i asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36176 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_3_1_0_wb_clk_i
timestamp 1698431365
transform 1 0 51968 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_3_2_0_wb_clk_i
timestamp 1698431365
transform -1 0 35840 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_3_3_0_wb_clk_i
timestamp 1698431365
transform -1 0 52304 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_3_4_0_wb_clk_i
timestamp 1698431365
transform -1 0 83664 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_3_5_0_wb_clk_i
timestamp 1698431365
transform 1 0 99568 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_3_6_0_wb_clk_i
timestamp 1698431365
transform -1 0 79744 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_3_7_0_wb_clk_i
timestamp 1698431365
transform 1 0 96544 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_0__f_wb_clk_i
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_1__f_wb_clk_i
timestamp 1698431365
transform -1 0 36064 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_2__f_wb_clk_i
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 54432 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_4__f_wb_clk_i
timestamp 1698431365
transform -1 0 35280 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_5__f_wb_clk_i
timestamp 1698431365
transform 1 0 30688 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_6__f_wb_clk_i
timestamp 1698431365
transform -1 0 51184 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_7__f_wb_clk_i
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_8__f_wb_clk_i
timestamp 1698431365
transform 1 0 79968 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_9__f_wb_clk_i
timestamp 1698431365
transform -1 0 83552 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_10__f_wb_clk_i
timestamp 1698431365
transform 1 0 103488 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_11__f_wb_clk_i
timestamp 1698431365
transform 1 0 101360 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_12__f_wb_clk_i
timestamp 1698431365
transform 1 0 76048 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_13__f_wb_clk_i
timestamp 1698431365
transform 1 0 78064 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_14__f_wb_clk_i
timestamp 1698431365
transform 1 0 99568 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_4_15__f_wb_clk_i
timestamp 1698431365
transform 1 0 99568 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout138
timestamp 1698431365
transform -1 0 71232 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout139
timestamp 1698431365
transform 1 0 115808 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_70 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_78 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_80 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10304 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_91
timestamp 1698431365
transform 1 0 11536 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_99
timestamp 1698431365
transform 1 0 12432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142
timestamp 1698431365
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_146
timestamp 1698431365
transform 1 0 17696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_150
timestamp 1698431365
transform 1 0 18144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_337
timestamp 1698431365
transform 1 0 39088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_507
timestamp 1698431365
transform 1 0 58128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_509
timestamp 1698431365
transform 1 0 58352 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_609
timestamp 1698431365
transform 1 0 69552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_611
timestamp 1698431365
transform 1 0 69776 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_682
timestamp 1698431365
transform 1 0 77728 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_716
timestamp 1698431365
transform 1 0 81536 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_718
timestamp 1698431365
transform 1 0 81760 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_745
timestamp 1698431365
transform 1 0 84784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_747
timestamp 1698431365
transform 1 0 85008 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_781
timestamp 1698431365
transform 1 0 88816 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_848
timestamp 1698431365
transform 1 0 96320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_951
timestamp 1698431365
transform 1 0 107856 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1150
timestamp 1698431365
transform 1 0 130144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1154
timestamp 1698431365
transform 1 0 130592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1294
timestamp 1698431365
transform 1 0 146272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1321
timestamp 1698431365
transform 1 0 149296 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1323
timestamp 1698431365
transform 1 0 149520 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1328
timestamp 1698431365
transform 1 0 150080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1330
timestamp 1698431365
transform 1 0 150304 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1357
timestamp 1698431365
transform 1 0 153328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1359
timestamp 1698431365
transform 1 0 153552 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1362
timestamp 1698431365
transform 1 0 153888 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1396 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 157696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1400
timestamp 1698431365
transform 1 0 158144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_104
timestamp 1698431365
transform 1 0 12992 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_113
timestamp 1698431365
transform 1 0 14000 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_121
timestamp 1698431365
transform 1 0 14896 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_133
timestamp 1698431365
transform 1 0 16240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_189
timestamp 1698431365
transform 1 0 22512 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_257
timestamp 1698431365
transform 1 0 30128 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_259
timestamp 1698431365
transform 1 0 30352 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_483
timestamp 1698431365
transform 1 0 55440 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_542
timestamp 1698431365
transform 1 0 62048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_632
timestamp 1698431365
transform 1 0 72128 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_634
timestamp 1698431365
transform 1 0 72352 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_674
timestamp 1698431365
transform 1 0 76832 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_838
timestamp 1698431365
transform 1 0 95200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_909
timestamp 1698431365
transform 1 0 103152 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_912
timestamp 1698431365
transform 1 0 103488 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1048
timestamp 1698431365
transform 1 0 118720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1074
timestamp 1698431365
transform 1 0 121632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1078
timestamp 1698431365
transform 1 0 122080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1082
timestamp 1698431365
transform 1 0 122528 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1122
timestamp 1698431365
transform 1 0 127008 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1176
timestamp 1698431365
transform 1 0 133056 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1184
timestamp 1698431365
transform 1 0 133952 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1188
timestamp 1698431365
transform 1 0 134400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1192
timestamp 1698431365
transform 1 0 134848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1232
timestamp 1698431365
transform 1 0 139328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1236
timestamp 1698431365
transform 1 0 139776 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1244
timestamp 1698431365
transform 1 0 140672 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1248
timestamp 1698431365
transform 1 0 141120 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1259
timestamp 1698431365
transform 1 0 142352 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1268
timestamp 1698431365
transform 1 0 143360 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1272
timestamp 1698431365
transform 1 0 143808 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1289
timestamp 1698431365
transform 1 0 145712 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1295
timestamp 1698431365
transform 1 0 146384 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1303
timestamp 1698431365
transform 1 0 147280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1329
timestamp 1698431365
transform 1 0 150192 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1332
timestamp 1698431365
transform 1 0 150528 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1396
timestamp 1698431365
transform 1 0 157696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_123
timestamp 1698431365
transform 1 0 15120 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_132
timestamp 1698431365
transform 1 0 16128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_150
timestamp 1698431365
transform 1 0 18144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_152
timestamp 1698431365
transform 1 0 18368 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_155
timestamp 1698431365
transform 1 0 18704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_187
timestamp 1698431365
transform 1 0 22288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_220
timestamp 1698431365
transform 1 0 25984 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_249
timestamp 1698431365
transform 1 0 29232 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_277
timestamp 1698431365
transform 1 0 32368 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_389
timestamp 1698431365
transform 1 0 44912 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_499
timestamp 1698431365
transform 1 0 57232 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_648
timestamp 1698431365
transform 1 0 73920 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_693
timestamp 1698431365
transform 1 0 78960 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_757
timestamp 1698431365
transform 1 0 86128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_759
timestamp 1698431365
transform 1 0 86352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_812
timestamp 1698431365
transform 1 0 92288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_877
timestamp 1698431365
transform 1 0 99568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_942
timestamp 1698431365
transform 1 0 106848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_944
timestamp 1698431365
transform 1 0 107072 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1084
timestamp 1698431365
transform 1 0 122752 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1143
timestamp 1698431365
transform 1 0 129360 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1151
timestamp 1698431365
transform 1 0 130256 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1157
timestamp 1698431365
transform 1 0 130928 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1165
timestamp 1698431365
transform 1 0 131824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1167
timestamp 1698431365
transform 1 0 132048 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1170
timestamp 1698431365
transform 1 0 132384 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1178
timestamp 1698431365
transform 1 0 133280 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1197
timestamp 1698431365
transform 1 0 135408 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1201
timestamp 1698431365
transform 1 0 135856 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1204
timestamp 1698431365
transform 1 0 136192 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1212
timestamp 1698431365
transform 1 0 137088 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1216
timestamp 1698431365
transform 1 0 137536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1220
timestamp 1698431365
transform 1 0 137984 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1227
timestamp 1698431365
transform 1 0 138768 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1235
timestamp 1698431365
transform 1 0 139664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1237
timestamp 1698431365
transform 1 0 139888 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1254
timestamp 1698431365
transform 1 0 141792 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1258
timestamp 1698431365
transform 1 0 142240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1260
timestamp 1698431365
transform 1 0 142464 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1285
timestamp 1698431365
transform 1 0 145264 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1293
timestamp 1698431365
transform 1 0 146160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1297
timestamp 1698431365
transform 1 0 146608 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1313
timestamp 1698431365
transform 1 0 148400 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1317
timestamp 1698431365
transform 1 0 148848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_1337
timestamp 1698431365
transform 1 0 151088 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1353
timestamp 1698431365
transform 1 0 152880 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1361
timestamp 1698431365
transform 1 0 153776 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_1367
timestamp 1698431365
transform 1 0 154448 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1399
timestamp 1698431365
transform 1 0 158032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1401
timestamp 1698431365
transform 1 0 158256 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_164
timestamp 1698431365
transform 1 0 19712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_166
timestamp 1698431365
transform 1 0 19936 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_169
timestamp 1698431365
transform 1 0 20272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_173
timestamp 1698431365
transform 1 0 20720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_185
timestamp 1698431365
transform 1 0 22064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_187
timestamp 1698431365
transform 1 0 22288 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_237
timestamp 1698431365
transform 1 0 27888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_255
timestamp 1698431365
transform 1 0 29904 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_418
timestamp 1698431365
transform 1 0 48160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_430
timestamp 1698431365
transform 1 0 49504 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_588
timestamp 1698431365
transform 1 0 67200 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_626
timestamp 1698431365
transform 1 0 71456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_646
timestamp 1698431365
transform 1 0 73696 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_698
timestamp 1698431365
transform 1 0 79520 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_702
timestamp 1698431365
transform 1 0 79968 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_769
timestamp 1698431365
transform 1 0 87472 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_777
timestamp 1698431365
transform 1 0 88368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_842
timestamp 1698431365
transform 1 0 95648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_844
timestamp 1698431365
transform 1 0 95872 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_912
timestamp 1698431365
transform 1 0 103488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_957
timestamp 1698431365
transform 1 0 108528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1007
timestamp 1698431365
transform 1 0 114128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1072
timestamp 1698431365
transform 1 0 121408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1076
timestamp 1698431365
transform 1 0 121856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1100
timestamp 1698431365
transform 1 0 124544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1122
timestamp 1698431365
transform 1 0 127008 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1126
timestamp 1698431365
transform 1 0 127456 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_1129
timestamp 1698431365
transform 1 0 127792 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_1161
timestamp 1698431365
transform 1 0 131376 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_1177
timestamp 1698431365
transform 1 0 133168 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1185
timestamp 1698431365
transform 1 0 134064 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1189
timestamp 1698431365
transform 1 0 134512 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_1192
timestamp 1698431365
transform 1 0 134848 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1224
timestamp 1698431365
transform 1 0 138432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1226
timestamp 1698431365
transform 1 0 138656 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_1231
timestamp 1698431365
transform 1 0 139216 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_1247
timestamp 1698431365
transform 1 0 141008 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1255
timestamp 1698431365
transform 1 0 141904 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1259
timestamp 1698431365
transform 1 0 142352 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_1262
timestamp 1698431365
transform 1 0 142688 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1270
timestamp 1698431365
transform 1 0 143584 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1273
timestamp 1698431365
transform 1 0 143920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_1277
timestamp 1698431365
transform 1 0 144368 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_1309
timestamp 1698431365
transform 1 0 147952 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1325
timestamp 1698431365
transform 1 0 149744 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1329
timestamp 1698431365
transform 1 0 150192 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1332
timestamp 1698431365
transform 1 0 150528 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1396
timestamp 1698431365
transform 1 0 157696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_139
timestamp 1698431365
transform 1 0 16912 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_143
timestamp 1698431365
transform 1 0 17360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_145
timestamp 1698431365
transform 1 0 17584 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_148
timestamp 1698431365
transform 1 0 17920 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_160
timestamp 1698431365
transform 1 0 19264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_179
timestamp 1698431365
transform 1 0 21392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_202
timestamp 1698431365
transform 1 0 23968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_265
timestamp 1698431365
transform 1 0 31024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_267
timestamp 1698431365
transform 1 0 31248 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_288
timestamp 1698431365
transform 1 0 33600 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_339
timestamp 1698431365
transform 1 0 39312 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_377
timestamp 1698431365
transform 1 0 43568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_379
timestamp 1698431365
transform 1 0 43792 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_507
timestamp 1698431365
transform 1 0 58128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_527
timestamp 1698431365
transform 1 0 60368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_597
timestamp 1698431365
transform 1 0 68208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_667
timestamp 1698431365
transform 1 0 76048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_695
timestamp 1698431365
transform 1 0 79184 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_732
timestamp 1698431365
transform 1 0 83328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_734
timestamp 1698431365
transform 1 0 83552 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_784
timestamp 1698431365
transform 1 0 89152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_807
timestamp 1698431365
transform 1 0 91728 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_842
timestamp 1698431365
transform 1 0 95648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_873
timestamp 1698431365
transform 1 0 99120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_942
timestamp 1698431365
transform 1 0 106848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_944
timestamp 1698431365
transform 1 0 107072 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_984
timestamp 1698431365
transform 1 0 111552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1013
timestamp 1698431365
transform 1 0 114800 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1038
timestamp 1698431365
transform 1 0 117600 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1065
timestamp 1698431365
transform 1 0 120624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1069
timestamp 1698431365
transform 1 0 121072 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1073
timestamp 1698431365
transform 1 0 121520 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1076
timestamp 1698431365
transform 1 0 121856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1080
timestamp 1698431365
transform 1 0 122304 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1083
timestamp 1698431365
transform 1 0 122640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1087
timestamp 1698431365
transform 1 0 123088 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1091
timestamp 1698431365
transform 1 0 123536 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_1094
timestamp 1698431365
transform 1 0 123872 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_1112
timestamp 1698431365
transform 1 0 125888 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_1144
timestamp 1698431365
transform 1 0 129472 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1152
timestamp 1698431365
transform 1 0 130368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1154
timestamp 1698431365
transform 1 0 130592 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1157
timestamp 1698431365
transform 1 0 130928 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1221
timestamp 1698431365
transform 1 0 138096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1227
timestamp 1698431365
transform 1 0 138768 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1291
timestamp 1698431365
transform 1 0 145936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1297
timestamp 1698431365
transform 1 0 146608 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1361
timestamp 1698431365
transform 1 0 153776 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_1367
timestamp 1698431365
transform 1 0 154448 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1399
timestamp 1698431365
transform 1 0 158032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1401
timestamp 1698431365
transform 1 0 158256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_158
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_162
timestamp 1698431365
transform 1 0 19488 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_197
timestamp 1698431365
transform 1 0 23408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_199
timestamp 1698431365
transform 1 0 23632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_214
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_217
timestamp 1698431365
transform 1 0 25648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_269
timestamp 1698431365
transform 1 0 31472 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_273
timestamp 1698431365
transform 1 0 31920 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_333
timestamp 1698431365
transform 1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_360
timestamp 1698431365
transform 1 0 41664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_431
timestamp 1698431365
transform 1 0 49616 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_478
timestamp 1698431365
transform 1 0 54880 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_487
timestamp 1698431365
transform 1 0 55888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_489
timestamp 1698431365
transform 1 0 56112 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_533
timestamp 1698431365
transform 1 0 61040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_576
timestamp 1698431365
transform 1 0 65856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_699
timestamp 1698431365
transform 1 0 79632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_752
timestamp 1698431365
transform 1 0 85568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_811
timestamp 1698431365
transform 1 0 92176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_813
timestamp 1698431365
transform 1 0 92400 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_838
timestamp 1698431365
transform 1 0 95200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_926
timestamp 1698431365
transform 1 0 105056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_928
timestamp 1698431365
transform 1 0 105280 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_990
timestamp 1698431365
transform 1 0 112224 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1020
timestamp 1698431365
transform 1 0 115584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1046
timestamp 1698431365
transform 1 0 118496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1052
timestamp 1698431365
transform 1 0 119168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1056
timestamp 1698431365
transform 1 0 119616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1060
timestamp 1698431365
transform 1 0 120064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_1064
timestamp 1698431365
transform 1 0 120512 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_1096
timestamp 1698431365
transform 1 0 124096 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_1112
timestamp 1698431365
transform 1 0 125888 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1122
timestamp 1698431365
transform 1 0 127008 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1186
timestamp 1698431365
transform 1 0 134176 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1192
timestamp 1698431365
transform 1 0 134848 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1256
timestamp 1698431365
transform 1 0 142016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1262
timestamp 1698431365
transform 1 0 142688 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1326
timestamp 1698431365
transform 1 0 149856 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1332
timestamp 1698431365
transform 1 0 150528 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1396
timestamp 1698431365
transform 1 0 157696 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_195
timestamp 1698431365
transform 1 0 23184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_199
timestamp 1698431365
transform 1 0 23632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_203
timestamp 1698431365
transform 1 0 24080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_207
timestamp 1698431365
transform 1 0 24528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_389
timestamp 1698431365
transform 1 0 44912 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_419
timestamp 1698431365
transform 1 0 48272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_423
timestamp 1698431365
transform 1 0 48720 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_426
timestamp 1698431365
transform 1 0 49056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_446
timestamp 1698431365
transform 1 0 51296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_580
timestamp 1698431365
transform 1 0 66304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_630
timestamp 1698431365
transform 1 0 71904 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_667
timestamp 1698431365
transform 1 0 76048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_669
timestamp 1698431365
transform 1 0 76272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_733
timestamp 1698431365
transform 1 0 83440 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_764
timestamp 1698431365
transform 1 0 86912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_771
timestamp 1698431365
transform 1 0 87696 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_773
timestamp 1698431365
transform 1 0 87920 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_787
timestamp 1698431365
transform 1 0 89488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_845
timestamp 1698431365
transform 1 0 95984 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_891
timestamp 1698431365
transform 1 0 101136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_943
timestamp 1698431365
transform 1 0 106960 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_947
timestamp 1698431365
transform 1 0 107408 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1038
timestamp 1698431365
transform 1 0 117600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1042
timestamp 1698431365
transform 1 0 118048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1046
timestamp 1698431365
transform 1 0 118496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1050
timestamp 1698431365
transform 1 0 118944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_1054
timestamp 1698431365
transform 1 0 119392 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1070
timestamp 1698431365
transform 1 0 121184 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1078
timestamp 1698431365
transform 1 0 122080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1082
timestamp 1698431365
transform 1 0 122528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1084
timestamp 1698431365
transform 1 0 122752 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1087
timestamp 1698431365
transform 1 0 123088 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1151
timestamp 1698431365
transform 1 0 130256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1157
timestamp 1698431365
transform 1 0 130928 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1221
timestamp 1698431365
transform 1 0 138096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1227
timestamp 1698431365
transform 1 0 138768 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1291
timestamp 1698431365
transform 1 0 145936 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1297
timestamp 1698431365
transform 1 0 146608 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1361
timestamp 1698431365
transform 1 0 153776 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_1367
timestamp 1698431365
transform 1 0 154448 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1399
timestamp 1698431365
transform 1 0 158032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1401
timestamp 1698431365
transform 1 0 158256 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_158
timestamp 1698431365
transform 1 0 19040 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_166
timestamp 1698431365
transform 1 0 19936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_172
timestamp 1698431365
transform 1 0 20608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_174
timestamp 1698431365
transform 1 0 20832 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_177
timestamp 1698431365
transform 1 0 21168 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_186
timestamp 1698431365
transform 1 0 22176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_190
timestamp 1698431365
transform 1 0 22624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_194
timestamp 1698431365
transform 1 0 23072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_204
timestamp 1698431365
transform 1 0 24192 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_218
timestamp 1698431365
transform 1 0 25760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_222
timestamp 1698431365
transform 1 0 26208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_266
timestamp 1698431365
transform 1 0 31136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_348
timestamp 1698431365
transform 1 0 40320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_359
timestamp 1698431365
transform 1 0 41552 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_376
timestamp 1698431365
transform 1 0 43456 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_406
timestamp 1698431365
transform 1 0 46816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_415
timestamp 1698431365
transform 1 0 47824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_417
timestamp 1698431365
transform 1 0 48048 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_426
timestamp 1698431365
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_430
timestamp 1698431365
transform 1 0 49504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_434
timestamp 1698431365
transform 1 0 49952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_438
timestamp 1698431365
transform 1 0 50400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_442
timestamp 1698431365
transform 1 0 50848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_446
timestamp 1698431365
transform 1 0 51296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_450
timestamp 1698431365
transform 1 0 51744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_454
timestamp 1698431365
transform 1 0 52192 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_479
timestamp 1698431365
transform 1 0 54992 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_536
timestamp 1698431365
transform 1 0 61376 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_556
timestamp 1698431365
transform 1 0 63616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_570
timestamp 1698431365
transform 1 0 65184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_584
timestamp 1698431365
transform 1 0 66752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_586
timestamp 1698431365
transform 1 0 66976 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_632
timestamp 1698431365
transform 1 0 72128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_698
timestamp 1698431365
transform 1 0 79520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_710
timestamp 1698431365
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_722
timestamp 1698431365
transform 1 0 82208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_763
timestamp 1698431365
transform 1 0 86800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_838
timestamp 1698431365
transform 1 0 95200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_908
timestamp 1698431365
transform 1 0 103040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_934
timestamp 1698431365
transform 1 0 105952 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_978
timestamp 1698431365
transform 1 0 110880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1028
timestamp 1698431365
transform 1 0 116480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1032
timestamp 1698431365
transform 1 0 116928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1036
timestamp 1698431365
transform 1 0 117376 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1040
timestamp 1698431365
transform 1 0 117824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1044
timestamp 1698431365
transform 1 0 118272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1048
timestamp 1698431365
transform 1 0 118720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1052
timestamp 1698431365
transform 1 0 119168 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1116
timestamp 1698431365
transform 1 0 126336 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1122
timestamp 1698431365
transform 1 0 127008 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1186
timestamp 1698431365
transform 1 0 134176 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1192
timestamp 1698431365
transform 1 0 134848 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1256
timestamp 1698431365
transform 1 0 142016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1262
timestamp 1698431365
transform 1 0 142688 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1326
timestamp 1698431365
transform 1 0 149856 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1332
timestamp 1698431365
transform 1 0 150528 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1396
timestamp 1698431365
transform 1 0 157696 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_139
timestamp 1698431365
transform 1 0 16912 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_157
timestamp 1698431365
transform 1 0 18928 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_161
timestamp 1698431365
transform 1 0 19376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_165
timestamp 1698431365
transform 1 0 19824 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_181
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_298
timestamp 1698431365
transform 1 0 34720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_300
timestamp 1698431365
transform 1 0 34944 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_395
timestamp 1698431365
transform 1 0 45584 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_401
timestamp 1698431365
transform 1 0 46256 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_407
timestamp 1698431365
transform 1 0 46928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_411
timestamp 1698431365
transform 1 0 47376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_415
timestamp 1698431365
transform 1 0 47824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_429
timestamp 1698431365
transform 1 0 49392 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_444
timestamp 1698431365
transform 1 0 51072 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_448
timestamp 1698431365
transform 1 0 51520 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_451
timestamp 1698431365
transform 1 0 51856 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_500
timestamp 1698431365
transform 1 0 57344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_511
timestamp 1698431365
transform 1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_513
timestamp 1698431365
transform 1 0 58800 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_527
timestamp 1698431365
transform 1 0 60368 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_543
timestamp 1698431365
transform 1 0 62160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_550
timestamp 1698431365
transform 1 0 62944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_552
timestamp 1698431365
transform 1 0 63168 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_563
timestamp 1698431365
transform 1 0 64400 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_574
timestamp 1698431365
transform 1 0 65632 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_576
timestamp 1698431365
transform 1 0 65856 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_579
timestamp 1698431365
transform 1 0 66192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_583
timestamp 1698431365
transform 1 0 66640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_587
timestamp 1698431365
transform 1 0 67088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_591
timestamp 1698431365
transform 1 0 67536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_597
timestamp 1698431365
transform 1 0 68208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_601
timestamp 1698431365
transform 1 0 68656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_610
timestamp 1698431365
transform 1 0 69664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_612
timestamp 1698431365
transform 1 0 69888 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_626
timestamp 1698431365
transform 1 0 71456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_648
timestamp 1698431365
transform 1 0 73920 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_664
timestamp 1698431365
transform 1 0 75712 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_681
timestamp 1698431365
transform 1 0 77616 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_717
timestamp 1698431365
transform 1 0 81648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_737
timestamp 1698431365
transform 1 0 83888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_739
timestamp 1698431365
transform 1 0 84112 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_749
timestamp 1698431365
transform 1 0 85232 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_753
timestamp 1698431365
transform 1 0 85680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_820
timestamp 1698431365
transform 1 0 93184 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_918
timestamp 1698431365
transform 1 0 104160 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_935
timestamp 1698431365
transform 1 0 106064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_961
timestamp 1698431365
transform 1 0 108976 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1012
timestamp 1698431365
transform 1 0 114688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1014
timestamp 1698431365
transform 1 0 114912 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1022
timestamp 1698431365
transform 1 0 115808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1026
timestamp 1698431365
transform 1 0 116256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1030
timestamp 1698431365
transform 1 0 116704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_1034
timestamp 1698431365
transform 1 0 117152 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_1066
timestamp 1698431365
transform 1 0 120736 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1082
timestamp 1698431365
transform 1 0 122528 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1084
timestamp 1698431365
transform 1 0 122752 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1087
timestamp 1698431365
transform 1 0 123088 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1151
timestamp 1698431365
transform 1 0 130256 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1157
timestamp 1698431365
transform 1 0 130928 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1221
timestamp 1698431365
transform 1 0 138096 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1227
timestamp 1698431365
transform 1 0 138768 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1291
timestamp 1698431365
transform 1 0 145936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1297
timestamp 1698431365
transform 1 0 146608 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1361
timestamp 1698431365
transform 1 0 153776 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_1367
timestamp 1698431365
transform 1 0 154448 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1399
timestamp 1698431365
transform 1 0 158032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1401
timestamp 1698431365
transform 1 0 158256 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_183
timestamp 1698431365
transform 1 0 21840 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_187
timestamp 1698431365
transform 1 0 22288 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_191
timestamp 1698431365
transform 1 0 22736 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_194
timestamp 1698431365
transform 1 0 23072 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_218
timestamp 1698431365
transform 1 0 25760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_223
timestamp 1698431365
transform 1 0 26320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_243
timestamp 1698431365
transform 1 0 28560 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_249
timestamp 1698431365
transform 1 0 29232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_253
timestamp 1698431365
transform 1 0 29680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_295
timestamp 1698431365
transform 1 0 34384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_316
timestamp 1698431365
transform 1 0 36736 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_366
timestamp 1698431365
transform 1 0 42336 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_370
timestamp 1698431365
transform 1 0 42784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_374
timestamp 1698431365
transform 1 0 43232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_392
timestamp 1698431365
transform 1 0 45248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_409
timestamp 1698431365
transform 1 0 47152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_411
timestamp 1698431365
transform 1 0 47376 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_443
timestamp 1698431365
transform 1 0 50960 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_449
timestamp 1698431365
transform 1 0 51632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_453
timestamp 1698431365
transform 1 0 52080 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_457
timestamp 1698431365
transform 1 0 52528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_461
timestamp 1698431365
transform 1 0 52976 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_465
timestamp 1698431365
transform 1 0 53424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_469
timestamp 1698431365
transform 1 0 53872 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_479
timestamp 1698431365
transform 1 0 54992 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_481
timestamp 1698431365
transform 1 0 55216 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_520
timestamp 1698431365
transform 1 0 59584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_522
timestamp 1698431365
transform 1 0 59808 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_557
timestamp 1698431365
transform 1 0 63728 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_559
timestamp 1698431365
transform 1 0 63952 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_562
timestamp 1698431365
transform 1 0 64288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_564
timestamp 1698431365
transform 1 0 64512 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_594
timestamp 1698431365
transform 1 0 67872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_598
timestamp 1698431365
transform 1 0 68320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_632
timestamp 1698431365
transform 1 0 72128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_688
timestamp 1698431365
transform 1 0 78400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_708
timestamp 1698431365
transform 1 0 80640 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_757
timestamp 1698431365
transform 1 0 86128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_761
timestamp 1698431365
transform 1 0 86576 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_772
timestamp 1698431365
transform 1 0 87808 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_908
timestamp 1698431365
transform 1 0 103040 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_962
timestamp 1698431365
transform 1 0 109088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_982
timestamp 1698431365
transform 1 0 111328 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_991
timestamp 1698431365
transform 1 0 112336 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1021
timestamp 1698431365
transform 1 0 115696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1025
timestamp 1698431365
transform 1 0 116144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_1029
timestamp 1698431365
transform 1 0 116592 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1045
timestamp 1698431365
transform 1 0 118384 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_1049
timestamp 1698431365
transform 1 0 118832 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1052
timestamp 1698431365
transform 1 0 119168 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1116
timestamp 1698431365
transform 1 0 126336 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1122
timestamp 1698431365
transform 1 0 127008 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1186
timestamp 1698431365
transform 1 0 134176 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1192
timestamp 1698431365
transform 1 0 134848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1256
timestamp 1698431365
transform 1 0 142016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1262
timestamp 1698431365
transform 1 0 142688 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1326
timestamp 1698431365
transform 1 0 149856 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1332
timestamp 1698431365
transform 1 0 150528 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1396
timestamp 1698431365
transform 1 0 157696 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_123
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_125
timestamp 1698431365
transform 1 0 15344 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_155
timestamp 1698431365
transform 1 0 18704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_183
timestamp 1698431365
transform 1 0 21840 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_187
timestamp 1698431365
transform 1 0 22288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_191
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_199
timestamp 1698431365
transform 1 0 23632 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_203
timestamp 1698431365
transform 1 0 24080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_211
timestamp 1698431365
transform 1 0 24976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_213
timestamp 1698431365
transform 1 0 25200 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_216
timestamp 1698431365
transform 1 0 25536 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_218
timestamp 1698431365
transform 1 0 25760 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_221
timestamp 1698431365
transform 1 0 26096 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_229
timestamp 1698431365
transform 1 0 26992 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_239
timestamp 1698431365
transform 1 0 28112 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_253
timestamp 1698431365
transform 1 0 29680 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_256
timestamp 1698431365
transform 1 0 30016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_340
timestamp 1698431365
transform 1 0 39424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_353
timestamp 1698431365
transform 1 0 40880 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_373
timestamp 1698431365
transform 1 0 43120 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_377
timestamp 1698431365
transform 1 0 43568 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_380
timestamp 1698431365
transform 1 0 43904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_391
timestamp 1698431365
transform 1 0 45136 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_395
timestamp 1698431365
transform 1 0 45584 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_399
timestamp 1698431365
transform 1 0 46032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_403
timestamp 1698431365
transform 1 0 46480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_405
timestamp 1698431365
transform 1 0 46704 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_408
timestamp 1698431365
transform 1 0 47040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_412
timestamp 1698431365
transform 1 0 47488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_416
timestamp 1698431365
transform 1 0 47936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_439
timestamp 1698431365
transform 1 0 50512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_443
timestamp 1698431365
transform 1 0 50960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_447
timestamp 1698431365
transform 1 0 51408 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_451
timestamp 1698431365
transform 1 0 51856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_473
timestamp 1698431365
transform 1 0 54320 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_524
timestamp 1698431365
transform 1 0 60032 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_531
timestamp 1698431365
transform 1 0 60816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_533
timestamp 1698431365
transform 1 0 61040 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_548
timestamp 1698431365
transform 1 0 62720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_552
timestamp 1698431365
transform 1 0 63168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_556
timestamp 1698431365
transform 1 0 63616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_560
timestamp 1698431365
transform 1 0 64064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_564
timestamp 1698431365
transform 1 0 64512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_574
timestamp 1698431365
transform 1 0 65632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_589
timestamp 1698431365
transform 1 0 67312 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_597
timestamp 1698431365
transform 1 0 68208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_601
timestamp 1698431365
transform 1 0 68656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_605
timestamp 1698431365
transform 1 0 69104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_609
timestamp 1698431365
transform 1 0 69552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_619
timestamp 1698431365
transform 1 0 70672 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_621
timestamp 1698431365
transform 1 0 70896 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_634
timestamp 1698431365
transform 1 0 72352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_641
timestamp 1698431365
transform 1 0 73136 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_643
timestamp 1698431365
transform 1 0 73360 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_650
timestamp 1698431365
transform 1 0 74144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_660
timestamp 1698431365
transform 1 0 75264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_662
timestamp 1698431365
transform 1 0 75488 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_681
timestamp 1698431365
transform 1 0 77616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_683
timestamp 1698431365
transform 1 0 77840 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_734
timestamp 1698431365
transform 1 0 83552 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_802
timestamp 1698431365
transform 1 0 91168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_804
timestamp 1698431365
transform 1 0 91392 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_807
timestamp 1698431365
transform 1 0 91728 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_826
timestamp 1698431365
transform 1 0 93856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_859
timestamp 1698431365
transform 1 0 97552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_863
timestamp 1698431365
transform 1 0 98000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_867
timestamp 1698431365
transform 1 0 98448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_871
timestamp 1698431365
transform 1 0 98896 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_877
timestamp 1698431365
transform 1 0 99568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_900
timestamp 1698431365
transform 1 0 102144 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_941
timestamp 1698431365
transform 1 0 106736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_973
timestamp 1698431365
transform 1 0 110320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_980
timestamp 1698431365
transform 1 0 111104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_987
timestamp 1698431365
transform 1 0 111888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_991
timestamp 1698431365
transform 1 0 112336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_995
timestamp 1698431365
transform 1 0 112784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_999
timestamp 1698431365
transform 1 0 113232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1003
timestamp 1698431365
transform 1 0 113680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1007
timestamp 1698431365
transform 1 0 114128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1011
timestamp 1698431365
transform 1 0 114576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1017
timestamp 1698431365
transform 1 0 115248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1081
timestamp 1698431365
transform 1 0 122416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1087
timestamp 1698431365
transform 1 0 123088 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1151
timestamp 1698431365
transform 1 0 130256 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1157
timestamp 1698431365
transform 1 0 130928 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1221
timestamp 1698431365
transform 1 0 138096 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1227
timestamp 1698431365
transform 1 0 138768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1291
timestamp 1698431365
transform 1 0 145936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1297
timestamp 1698431365
transform 1 0 146608 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1361
timestamp 1698431365
transform 1 0 153776 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_1367
timestamp 1698431365
transform 1 0 154448 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1399
timestamp 1698431365
transform 1 0 158032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_1401
timestamp 1698431365
transform 1 0 158256 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_148
timestamp 1698431365
transform 1 0 17920 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_151
timestamp 1698431365
transform 1 0 18256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_171
timestamp 1698431365
transform 1 0 20496 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_173
timestamp 1698431365
transform 1 0 20720 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_190
timestamp 1698431365
transform 1 0 22624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_194
timestamp 1698431365
transform 1 0 23072 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_198
timestamp 1698431365
transform 1 0 23520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_224
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_228
timestamp 1698431365
transform 1 0 26880 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_235
timestamp 1698431365
transform 1 0 27664 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_245
timestamp 1698431365
transform 1 0 28784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_255
timestamp 1698431365
transform 1 0 29904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_284
timestamp 1698431365
transform 1 0 33152 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_311
timestamp 1698431365
transform 1 0 36176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_313
timestamp 1698431365
transform 1 0 36400 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_328
timestamp 1698431365
transform 1 0 38080 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_332
timestamp 1698431365
transform 1 0 38528 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_335
timestamp 1698431365
transform 1 0 38864 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_339
timestamp 1698431365
transform 1 0 39312 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_342
timestamp 1698431365
transform 1 0 39648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_385
timestamp 1698431365
transform 1 0 44464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_406
timestamp 1698431365
transform 1 0 46816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_410
timestamp 1698431365
transform 1 0 47264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_414
timestamp 1698431365
transform 1 0 47712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_418
timestamp 1698431365
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_430
timestamp 1698431365
transform 1 0 49504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_434
timestamp 1698431365
transform 1 0 49952 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_441
timestamp 1698431365
transform 1 0 50736 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_471
timestamp 1698431365
transform 1 0 54096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_483
timestamp 1698431365
transform 1 0 55440 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_487
timestamp 1698431365
transform 1 0 55888 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_525
timestamp 1698431365
transform 1 0 60144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_533
timestamp 1698431365
transform 1 0 61040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_537
timestamp 1698431365
transform 1 0 61488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_541
timestamp 1698431365
transform 1 0 61936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_545
timestamp 1698431365
transform 1 0 62384 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_548
timestamp 1698431365
transform 1 0 62720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_552
timestamp 1698431365
transform 1 0 63168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_556
timestamp 1698431365
transform 1 0 63616 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_562
timestamp 1698431365
transform 1 0 64288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_564
timestamp 1698431365
transform 1 0 64512 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_573
timestamp 1698431365
transform 1 0 65520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_575
timestamp 1698431365
transform 1 0 65744 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_605
timestamp 1698431365
transform 1 0 69104 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_619
timestamp 1698431365
transform 1 0 70672 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_623
timestamp 1698431365
transform 1 0 71120 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_626
timestamp 1698431365
transform 1 0 71456 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_632
timestamp 1698431365
transform 1 0 72128 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_636
timestamp 1698431365
transform 1 0 72576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_640
timestamp 1698431365
transform 1 0 73024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_644
timestamp 1698431365
transform 1 0 73472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_648
timestamp 1698431365
transform 1 0 73920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_692
timestamp 1698431365
transform 1 0 78848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_694
timestamp 1698431365
transform 1 0 79072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_749
timestamp 1698431365
transform 1 0 85232 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_772
timestamp 1698431365
transform 1 0 87808 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_776
timestamp 1698431365
transform 1 0 88256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_780
timestamp 1698431365
transform 1 0 88704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_782
timestamp 1698431365
transform 1 0 88928 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_836
timestamp 1698431365
transform 1 0 94976 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_912
timestamp 1698431365
transform 1 0 103488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_914
timestamp 1698431365
transform 1 0 103712 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_926
timestamp 1698431365
transform 1 0 105056 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_960
timestamp 1698431365
transform 1 0 108864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_967
timestamp 1698431365
transform 1 0 109648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_971
timestamp 1698431365
transform 1 0 110096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_975
timestamp 1698431365
transform 1 0 110544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_979
timestamp 1698431365
transform 1 0 110992 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_982
timestamp 1698431365
transform 1 0 111328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_986
timestamp 1698431365
transform 1 0 111776 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_990
timestamp 1698431365
transform 1 0 112224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_994
timestamp 1698431365
transform 1 0 112672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_998
timestamp 1698431365
transform 1 0 113120 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_1002
timestamp 1698431365
transform 1 0 113568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_1006
timestamp 1698431365
transform 1 0 114016 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_1038
timestamp 1698431365
transform 1 0 117600 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1046
timestamp 1698431365
transform 1 0 118496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1052
timestamp 1698431365
transform 1 0 119168 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1116
timestamp 1698431365
transform 1 0 126336 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1122
timestamp 1698431365
transform 1 0 127008 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1186
timestamp 1698431365
transform 1 0 134176 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1192
timestamp 1698431365
transform 1 0 134848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1256
timestamp 1698431365
transform 1 0 142016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1262
timestamp 1698431365
transform 1 0 142688 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1326
timestamp 1698431365
transform 1 0 149856 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1332
timestamp 1698431365
transform 1 0 150528 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1396
timestamp 1698431365
transform 1 0 157696 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_155
timestamp 1698431365
transform 1 0 18704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_181
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_184
timestamp 1698431365
transform 1 0 21952 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_217
timestamp 1698431365
transform 1 0 25648 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_233
timestamp 1698431365
transform 1 0 27440 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_283
timestamp 1698431365
transform 1 0 33040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_285
timestamp 1698431365
transform 1 0 33264 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_323
timestamp 1698431365
transform 1 0 37520 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_332
timestamp 1698431365
transform 1 0 38528 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_336
timestamp 1698431365
transform 1 0 38976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_340
timestamp 1698431365
transform 1 0 39424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_344
timestamp 1698431365
transform 1 0 39872 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_346
timestamp 1698431365
transform 1 0 40096 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_349
timestamp 1698431365
transform 1 0 40432 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_382
timestamp 1698431365
transform 1 0 44128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_384
timestamp 1698431365
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_416
timestamp 1698431365
transform 1 0 47936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_436
timestamp 1698431365
transform 1 0 50176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_440
timestamp 1698431365
transform 1 0 50624 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_446
timestamp 1698431365
transform 1 0 51296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_450
timestamp 1698431365
transform 1 0 51744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_452
timestamp 1698431365
transform 1 0 51968 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_510
timestamp 1698431365
transform 1 0 58464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_514
timestamp 1698431365
transform 1 0 58912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_518
timestamp 1698431365
transform 1 0 59360 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_521
timestamp 1698431365
transform 1 0 59696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_535
timestamp 1698431365
transform 1 0 61264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_542
timestamp 1698431365
transform 1 0 62048 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_546
timestamp 1698431365
transform 1 0 62496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_550
timestamp 1698431365
transform 1 0 62944 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_585
timestamp 1698431365
transform 1 0 66864 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_589
timestamp 1698431365
transform 1 0 67312 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_592
timestamp 1698431365
transform 1 0 67648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_594
timestamp 1698431365
transform 1 0 67872 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_597
timestamp 1698431365
transform 1 0 68208 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_603
timestamp 1698431365
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_607
timestamp 1698431365
transform 1 0 69328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_609
timestamp 1698431365
transform 1 0 69552 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_639
timestamp 1698431365
transform 1 0 72912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_641
timestamp 1698431365
transform 1 0 73136 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_644
timestamp 1698431365
transform 1 0 73472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_648
timestamp 1698431365
transform 1 0 73920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_652
timestamp 1698431365
transform 1 0 74368 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_662
timestamp 1698431365
transform 1 0 75488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_664
timestamp 1698431365
transform 1 0 75712 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_671
timestamp 1698431365
transform 1 0 76496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_673
timestamp 1698431365
transform 1 0 76720 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_737
timestamp 1698431365
transform 1 0 83888 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_803
timestamp 1698431365
transform 1 0 91280 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_821
timestamp 1698431365
transform 1 0 93296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_825
timestamp 1698431365
transform 1 0 93744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_864
timestamp 1698431365
transform 1 0 98112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_868
timestamp 1698431365
transform 1 0 98560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_872
timestamp 1698431365
transform 1 0 99008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_874
timestamp 1698431365
transform 1 0 99232 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_877
timestamp 1698431365
transform 1 0 99568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_879
timestamp 1698431365
transform 1 0 99792 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_943
timestamp 1698431365
transform 1 0 106960 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_952
timestamp 1698431365
transform 1 0 107968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_956
timestamp 1698431365
transform 1 0 108416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_960
timestamp 1698431365
transform 1 0 108864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_964
timestamp 1698431365
transform 1 0 109312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_968
timestamp 1698431365
transform 1 0 109760 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_972
timestamp 1698431365
transform 1 0 110208 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_974
timestamp 1698431365
transform 1 0 110432 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_979
timestamp 1698431365
transform 1 0 110992 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_983
timestamp 1698431365
transform 1 0 111440 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_987
timestamp 1698431365
transform 1 0 111888 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_991
timestamp 1698431365
transform 1 0 112336 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_995
timestamp 1698431365
transform 1 0 112784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_999
timestamp 1698431365
transform 1 0 113232 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1017
timestamp 1698431365
transform 1 0 115248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1081
timestamp 1698431365
transform 1 0 122416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1087
timestamp 1698431365
transform 1 0 123088 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1151
timestamp 1698431365
transform 1 0 130256 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1157
timestamp 1698431365
transform 1 0 130928 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1221
timestamp 1698431365
transform 1 0 138096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1227
timestamp 1698431365
transform 1 0 138768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1291
timestamp 1698431365
transform 1 0 145936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1297
timestamp 1698431365
transform 1 0 146608 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1361
timestamp 1698431365
transform 1 0 153776 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_1367
timestamp 1698431365
transform 1 0 154448 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_1399
timestamp 1698431365
transform 1 0 158032 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_1401
timestamp 1698431365
transform 1 0 158256 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_158
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_162
timestamp 1698431365
transform 1 0 19488 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_165
timestamp 1698431365
transform 1 0 19824 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_172
timestamp 1698431365
transform 1 0 20608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_176
timestamp 1698431365
transform 1 0 21056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_180
timestamp 1698431365
transform 1 0 21504 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_196
timestamp 1698431365
transform 1 0 23296 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_204
timestamp 1698431365
transform 1 0 24192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_219
timestamp 1698431365
transform 1 0 25872 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_223
timestamp 1698431365
transform 1 0 26320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_261
timestamp 1698431365
transform 1 0 30576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_267
timestamp 1698431365
transform 1 0 31248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_269
timestamp 1698431365
transform 1 0 31472 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_272
timestamp 1698431365
transform 1 0 31808 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_305
timestamp 1698431365
transform 1 0 35504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_309
timestamp 1698431365
transform 1 0 35952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_313
timestamp 1698431365
transform 1 0 36400 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_317
timestamp 1698431365
transform 1 0 36848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_356
timestamp 1698431365
transform 1 0 41216 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_362
timestamp 1698431365
transform 1 0 41888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_366
timestamp 1698431365
transform 1 0 42336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_370
timestamp 1698431365
transform 1 0 42784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_372
timestamp 1698431365
transform 1 0 43008 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_375
timestamp 1698431365
transform 1 0 43344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_379
timestamp 1698431365
transform 1 0 43792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_383
timestamp 1698431365
transform 1 0 44240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_387
timestamp 1698431365
transform 1 0 44688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_391
timestamp 1698431365
transform 1 0 45136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_399
timestamp 1698431365
transform 1 0 46032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_403
timestamp 1698431365
transform 1 0 46480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_405
timestamp 1698431365
transform 1 0 46704 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_408
timestamp 1698431365
transform 1 0 47040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_412
timestamp 1698431365
transform 1 0 47488 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_426
timestamp 1698431365
transform 1 0 49056 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_429
timestamp 1698431365
transform 1 0 49392 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_433
timestamp 1698431365
transform 1 0 49840 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_437
timestamp 1698431365
transform 1 0 50288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_439
timestamp 1698431365
transform 1 0 50512 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_444
timestamp 1698431365
transform 1 0 51072 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_448
timestamp 1698431365
transform 1 0 51520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_478
timestamp 1698431365
transform 1 0 54880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_482
timestamp 1698431365
transform 1 0 55328 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_486
timestamp 1698431365
transform 1 0 55776 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_489
timestamp 1698431365
transform 1 0 56112 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_500
timestamp 1698431365
transform 1 0 57344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_504
timestamp 1698431365
transform 1 0 57792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_512
timestamp 1698431365
transform 1 0 58688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_551
timestamp 1698431365
transform 1 0 63056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_555
timestamp 1698431365
transform 1 0 63504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_559
timestamp 1698431365
transform 1 0 63952 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_570
timestamp 1698431365
transform 1 0 65184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_577
timestamp 1698431365
transform 1 0 65968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_581
timestamp 1698431365
transform 1 0 66416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_585
timestamp 1698431365
transform 1 0 66864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_589
timestamp 1698431365
transform 1 0 67312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_591
timestamp 1698431365
transform 1 0 67536 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_594
timestamp 1698431365
transform 1 0 67872 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_598
timestamp 1698431365
transform 1 0 68320 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_602
timestamp 1698431365
transform 1 0 68768 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_613
timestamp 1698431365
transform 1 0 70000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_615
timestamp 1698431365
transform 1 0 70224 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_618
timestamp 1698431365
transform 1 0 70560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_627
timestamp 1698431365
transform 1 0 71568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_629
timestamp 1698431365
transform 1 0 71792 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_637
timestamp 1698431365
transform 1 0 72688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_641
timestamp 1698431365
transform 1 0 73136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_643
timestamp 1698431365
transform 1 0 73360 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_646
timestamp 1698431365
transform 1 0 73696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_650
timestamp 1698431365
transform 1 0 74144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_698
timestamp 1698431365
transform 1 0 79520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_702
timestamp 1698431365
transform 1 0 79968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_704
timestamp 1698431365
transform 1 0 80192 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_707
timestamp 1698431365
transform 1 0 80528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_758
timestamp 1698431365
transform 1 0 86240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_762
timestamp 1698431365
transform 1 0 86688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_766
timestamp 1698431365
transform 1 0 87136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_772
timestamp 1698431365
transform 1 0 87808 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_776
timestamp 1698431365
transform 1 0 88256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_813
timestamp 1698431365
transform 1 0 92400 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_817
timestamp 1698431365
transform 1 0 92848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_821
timestamp 1698431365
transform 1 0 93296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_835
timestamp 1698431365
transform 1 0 94864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_839
timestamp 1698431365
transform 1 0 95312 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_903
timestamp 1698431365
transform 1 0 102480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_907
timestamp 1698431365
transform 1 0 102928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_909
timestamp 1698431365
transform 1 0 103152 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_938
timestamp 1698431365
transform 1 0 106400 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_942
timestamp 1698431365
transform 1 0 106848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_946
timestamp 1698431365
transform 1 0 107296 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_977
timestamp 1698431365
transform 1 0 110768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_979
timestamp 1698431365
transform 1 0 110992 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_986
timestamp 1698431365
transform 1 0 111776 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_990
timestamp 1698431365
transform 1 0 112224 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_1022
timestamp 1698431365
transform 1 0 115808 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_1038
timestamp 1698431365
transform 1 0 117600 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1046
timestamp 1698431365
transform 1 0 118496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1052
timestamp 1698431365
transform 1 0 119168 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1116
timestamp 1698431365
transform 1 0 126336 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1122
timestamp 1698431365
transform 1 0 127008 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1186
timestamp 1698431365
transform 1 0 134176 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1192
timestamp 1698431365
transform 1 0 134848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1256
timestamp 1698431365
transform 1 0 142016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1262
timestamp 1698431365
transform 1 0 142688 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1326
timestamp 1698431365
transform 1 0 149856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1332
timestamp 1698431365
transform 1 0 150528 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1396
timestamp 1698431365
transform 1 0 157696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_168
timestamp 1698431365
transform 1 0 20160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_209
timestamp 1698431365
transform 1 0 24752 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_215
timestamp 1698431365
transform 1 0 25424 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_231
timestamp 1698431365
transform 1 0 27216 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_251
timestamp 1698431365
transform 1 0 29456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_263
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_293
timestamp 1698431365
transform 1 0 34160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_297
timestamp 1698431365
transform 1 0 34608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_301
timestamp 1698431365
transform 1 0 35056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_305
timestamp 1698431365
transform 1 0 35504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_309
timestamp 1698431365
transform 1 0 35952 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_313
timestamp 1698431365
transform 1 0 36400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_321
timestamp 1698431365
transform 1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_325
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_329
timestamp 1698431365
transform 1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_333
timestamp 1698431365
transform 1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_337
timestamp 1698431365
transform 1 0 39088 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_341
timestamp 1698431365
transform 1 0 39536 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_345
timestamp 1698431365
transform 1 0 39984 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_353
timestamp 1698431365
transform 1 0 40880 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_357
timestamp 1698431365
transform 1 0 41328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_359
timestamp 1698431365
transform 1 0 41552 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_362
timestamp 1698431365
transform 1 0 41888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_366
timestamp 1698431365
transform 1 0 42336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_370
timestamp 1698431365
transform 1 0 42784 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_378
timestamp 1698431365
transform 1 0 43680 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_382
timestamp 1698431365
transform 1 0 44128 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_391
timestamp 1698431365
transform 1 0 45136 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_401
timestamp 1698431365
transform 1 0 46256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_409
timestamp 1698431365
transform 1 0 47152 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_419
timestamp 1698431365
transform 1 0 48272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_423
timestamp 1698431365
transform 1 0 48720 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_427
timestamp 1698431365
transform 1 0 49168 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_430
timestamp 1698431365
transform 1 0 49504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_434
timestamp 1698431365
transform 1 0 49952 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_450
timestamp 1698431365
transform 1 0 51744 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_454
timestamp 1698431365
transform 1 0 52192 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_465
timestamp 1698431365
transform 1 0 53424 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_469
timestamp 1698431365
transform 1 0 53872 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_472
timestamp 1698431365
transform 1 0 54208 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_476
timestamp 1698431365
transform 1 0 54656 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_492
timestamp 1698431365
transform 1 0 56448 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_498
timestamp 1698431365
transform 1 0 57120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_502
timestamp 1698431365
transform 1 0 57568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_506
timestamp 1698431365
transform 1 0 58016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_522
timestamp 1698431365
transform 1 0 59808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_524
timestamp 1698431365
transform 1 0 60032 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_527
timestamp 1698431365
transform 1 0 60368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_531
timestamp 1698431365
transform 1 0 60816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_543
timestamp 1698431365
transform 1 0 62160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_547
timestamp 1698431365
transform 1 0 62608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_551
timestamp 1698431365
transform 1 0 63056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_555
timestamp 1698431365
transform 1 0 63504 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_559
timestamp 1698431365
transform 1 0 63952 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_562
timestamp 1698431365
transform 1 0 64288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_566
timestamp 1698431365
transform 1 0 64736 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_586
timestamp 1698431365
transform 1 0 66976 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_594
timestamp 1698431365
transform 1 0 67872 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_597
timestamp 1698431365
transform 1 0 68208 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_601
timestamp 1698431365
transform 1 0 68656 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_631
timestamp 1698431365
transform 1 0 72016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_635
timestamp 1698431365
transform 1 0 72464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_637
timestamp 1698431365
transform 1 0 72688 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_640
timestamp 1698431365
transform 1 0 73024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_644
timestamp 1698431365
transform 1 0 73472 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_646
timestamp 1698431365
transform 1 0 73696 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_649
timestamp 1698431365
transform 1 0 74032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_653
timestamp 1698431365
transform 1 0 74480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_655
timestamp 1698431365
transform 1 0 74704 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_662
timestamp 1698431365
transform 1 0 75488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_664
timestamp 1698431365
transform 1 0 75712 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_667
timestamp 1698431365
transform 1 0 76048 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_671
timestamp 1698431365
transform 1 0 76496 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_728
timestamp 1698431365
transform 1 0 82880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_732
timestamp 1698431365
transform 1 0 83328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_734
timestamp 1698431365
transform 1 0 83552 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_747
timestamp 1698431365
transform 1 0 85008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_751
timestamp 1698431365
transform 1 0 85456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_755
timestamp 1698431365
transform 1 0 85904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_759
timestamp 1698431365
transform 1 0 86352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_795
timestamp 1698431365
transform 1 0 90384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_799
timestamp 1698431365
transform 1 0 90832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_803
timestamp 1698431365
transform 1 0 91280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_807
timestamp 1698431365
transform 1 0 91728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_811
timestamp 1698431365
transform 1 0 92176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_815
timestamp 1698431365
transform 1 0 92624 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_851
timestamp 1698431365
transform 1 0 96656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_855
timestamp 1698431365
transform 1 0 97104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_859
timestamp 1698431365
transform 1 0 97552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_863
timestamp 1698431365
transform 1 0 98000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_867
timestamp 1698431365
transform 1 0 98448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_977
timestamp 1698431365
transform 1 0 110768 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1009
timestamp 1698431365
transform 1 0 114352 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_1013
timestamp 1698431365
transform 1 0 114800 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1017
timestamp 1698431365
transform 1 0 115248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1081
timestamp 1698431365
transform 1 0 122416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1087
timestamp 1698431365
transform 1 0 123088 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1151
timestamp 1698431365
transform 1 0 130256 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1157
timestamp 1698431365
transform 1 0 130928 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1221
timestamp 1698431365
transform 1 0 138096 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1227
timestamp 1698431365
transform 1 0 138768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1291
timestamp 1698431365
transform 1 0 145936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1297
timestamp 1698431365
transform 1 0 146608 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1361
timestamp 1698431365
transform 1 0 153776 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_1367
timestamp 1698431365
transform 1 0 154448 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_1399
timestamp 1698431365
transform 1 0 158032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_1401
timestamp 1698431365
transform 1 0 158256 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_158
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_166
timestamp 1698431365
transform 1 0 19936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_168
timestamp 1698431365
transform 1 0 20160 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_179
timestamp 1698431365
transform 1 0 21392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_181
timestamp 1698431365
transform 1 0 21616 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_194
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_198
timestamp 1698431365
transform 1 0 23520 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_223
timestamp 1698431365
transform 1 0 26320 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_231
timestamp 1698431365
transform 1 0 27216 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_240
timestamp 1698431365
transform 1 0 28224 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_246
timestamp 1698431365
transform 1 0 28896 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_290
timestamp 1698431365
transform 1 0 33824 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_293
timestamp 1698431365
transform 1 0 34160 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_301
timestamp 1698431365
transform 1 0 35056 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_315
timestamp 1698431365
transform 1 0 36624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_317
timestamp 1698431365
transform 1 0 36848 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_331
timestamp 1698431365
transform 1 0 38416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_337
timestamp 1698431365
transform 1 0 39088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_341
timestamp 1698431365
transform 1 0 39536 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_381
timestamp 1698431365
transform 1 0 44016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_385
timestamp 1698431365
transform 1 0 44464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_389
timestamp 1698431365
transform 1 0 44912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_427
timestamp 1698431365
transform 1 0 49168 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_431
timestamp 1698431365
transform 1 0 49616 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_439
timestamp 1698431365
transform 1 0 50512 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_478
timestamp 1698431365
transform 1 0 54880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_482
timestamp 1698431365
transform 1 0 55328 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_496
timestamp 1698431365
transform 1 0 56896 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_505
timestamp 1698431365
transform 1 0 57904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_509
timestamp 1698431365
transform 1 0 58352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_513
timestamp 1698431365
transform 1 0 58800 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_517
timestamp 1698431365
transform 1 0 59248 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_520
timestamp 1698431365
transform 1 0 59584 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_524
timestamp 1698431365
transform 1 0 60032 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_549
timestamp 1698431365
transform 1 0 62832 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_559
timestamp 1698431365
transform 1 0 63952 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_591
timestamp 1698431365
transform 1 0 67536 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_603
timestamp 1698431365
transform 1 0 68880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_607
timestamp 1698431365
transform 1 0 69328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_611
timestamp 1698431365
transform 1 0 69776 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_615
timestamp 1698431365
transform 1 0 70224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_624
timestamp 1698431365
transform 1 0 71232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_628
timestamp 1698431365
transform 1 0 71680 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_632
timestamp 1698431365
transform 1 0 72128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_634
timestamp 1698431365
transform 1 0 72352 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_637
timestamp 1698431365
transform 1 0 72688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_639
timestamp 1698431365
transform 1 0 72912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_642
timestamp 1698431365
transform 1 0 73248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_646
timestamp 1698431365
transform 1 0 73696 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_649
timestamp 1698431365
transform 1 0 74032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_653
timestamp 1698431365
transform 1 0 74480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_686
timestamp 1698431365
transform 1 0 78176 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_690
timestamp 1698431365
transform 1 0 78624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_696
timestamp 1698431365
transform 1 0 79296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_731
timestamp 1698431365
transform 1 0 83216 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_735
timestamp 1698431365
transform 1 0 83664 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_765
timestamp 1698431365
transform 1 0 87024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_769
timestamp 1698431365
transform 1 0 87472 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_807
timestamp 1698431365
transform 1 0 91728 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_839
timestamp 1698431365
transform 1 0 95312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_877
timestamp 1698431365
transform 1 0 99568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_879
timestamp 1698431365
transform 1 0 99792 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_888
timestamp 1698431365
transform 1 0 100800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_906
timestamp 1698431365
transform 1 0 102816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_942
timestamp 1698431365
transform 1 0 106848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_946
timestamp 1698431365
transform 1 0 107296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_966
timestamp 1698431365
transform 1 0 109536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_970
timestamp 1698431365
transform 1 0 109984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_978
timestamp 1698431365
transform 1 0 110880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_982
timestamp 1698431365
transform 1 0 111328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1046
timestamp 1698431365
transform 1 0 118496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1052
timestamp 1698431365
transform 1 0 119168 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1116
timestamp 1698431365
transform 1 0 126336 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1122
timestamp 1698431365
transform 1 0 127008 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1186
timestamp 1698431365
transform 1 0 134176 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1192
timestamp 1698431365
transform 1 0 134848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1256
timestamp 1698431365
transform 1 0 142016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1262
timestamp 1698431365
transform 1 0 142688 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1326
timestamp 1698431365
transform 1 0 149856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1332
timestamp 1698431365
transform 1 0 150528 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1396
timestamp 1698431365
transform 1 0 157696 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_139
timestamp 1698431365
transform 1 0 16912 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_143
timestamp 1698431365
transform 1 0 17360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_145
timestamp 1698431365
transform 1 0 17584 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_179
timestamp 1698431365
transform 1 0 21392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_209
timestamp 1698431365
transform 1 0 24752 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_267
timestamp 1698431365
transform 1 0 31248 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_276
timestamp 1698431365
transform 1 0 32256 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_282
timestamp 1698431365
transform 1 0 32928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_284
timestamp 1698431365
transform 1 0 33152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_297
timestamp 1698431365
transform 1 0 34608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_301
timestamp 1698431365
transform 1 0 35056 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_303
timestamp 1698431365
transform 1 0 35280 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_367
timestamp 1698431365
transform 1 0 42448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_375
timestamp 1698431365
transform 1 0 43344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_379
timestamp 1698431365
transform 1 0 43792 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_383
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_403
timestamp 1698431365
transform 1 0 46480 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_435
timestamp 1698431365
transform 1 0 50064 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_443
timestamp 1698431365
transform 1 0 50960 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_447
timestamp 1698431365
transform 1 0 51408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_464
timestamp 1698431365
transform 1 0 53312 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_468
timestamp 1698431365
transform 1 0 53760 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_472
timestamp 1698431365
transform 1 0 54208 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_480
timestamp 1698431365
transform 1 0 55104 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_484
timestamp 1698431365
transform 1 0 55552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_486
timestamp 1698431365
transform 1 0 55776 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_503
timestamp 1698431365
transform 1 0 57680 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_519
timestamp 1698431365
transform 1 0 59472 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_523
timestamp 1698431365
transform 1 0 59920 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_527
timestamp 1698431365
transform 1 0 60368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_529
timestamp 1698431365
transform 1 0 60592 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_545
timestamp 1698431365
transform 1 0 62384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_549
timestamp 1698431365
transform 1 0 62832 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_553
timestamp 1698431365
transform 1 0 63280 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_580
timestamp 1698431365
transform 1 0 66304 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_588
timestamp 1698431365
transform 1 0 67200 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_592
timestamp 1698431365
transform 1 0 67648 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_594
timestamp 1698431365
transform 1 0 67872 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_626
timestamp 1698431365
transform 1 0 71456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_632
timestamp 1698431365
transform 1 0 72128 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_636
timestamp 1698431365
transform 1 0 72576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_638
timestamp 1698431365
transform 1 0 72800 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_647
timestamp 1698431365
transform 1 0 73808 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_653
timestamp 1698431365
transform 1 0 74480 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_667
timestamp 1698431365
transform 1 0 76048 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_671
timestamp 1698431365
transform 1 0 76496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_673
timestamp 1698431365
transform 1 0 76720 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_682
timestamp 1698431365
transform 1 0 77728 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_686
timestamp 1698431365
transform 1 0 78176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_690
timestamp 1698431365
transform 1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_694
timestamp 1698431365
transform 1 0 79072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_698
timestamp 1698431365
transform 1 0 79520 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_712
timestamp 1698431365
transform 1 0 81088 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_719
timestamp 1698431365
transform 1 0 81872 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_723
timestamp 1698431365
transform 1 0 82320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_727
timestamp 1698431365
transform 1 0 82768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_731
timestamp 1698431365
transform 1 0 83216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_737
timestamp 1698431365
transform 1 0 83888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_741
timestamp 1698431365
transform 1 0 84336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_745
timestamp 1698431365
transform 1 0 84784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_749
timestamp 1698431365
transform 1 0 85232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_753
timestamp 1698431365
transform 1 0 85680 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_757
timestamp 1698431365
transform 1 0 86128 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_804
timestamp 1698431365
transform 1 0 91392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_807
timestamp 1698431365
transform 1 0 91728 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_811
timestamp 1698431365
transform 1 0 92176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_815
timestamp 1698431365
transform 1 0 92624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_819
timestamp 1698431365
transform 1 0 93072 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_825
timestamp 1698431365
transform 1 0 93744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_829
timestamp 1698431365
transform 1 0 94192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_833
timestamp 1698431365
transform 1 0 94640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_837
timestamp 1698431365
transform 1 0 95088 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_841
timestamp 1698431365
transform 1 0 95536 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_872
timestamp 1698431365
transform 1 0 99008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_874
timestamp 1698431365
transform 1 0 99232 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_877
timestamp 1698431365
transform 1 0 99568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_881
timestamp 1698431365
transform 1 0 100016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_885
timestamp 1698431365
transform 1 0 100464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_887
timestamp 1698431365
transform 1 0 100688 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_890
timestamp 1698431365
transform 1 0 101024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_922
timestamp 1698431365
transform 1 0 104608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_926
timestamp 1698431365
transform 1 0 105056 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_930
timestamp 1698431365
transform 1 0 105504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_934
timestamp 1698431365
transform 1 0 105952 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_936
timestamp 1698431365
transform 1 0 106176 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_939
timestamp 1698431365
transform 1 0 106512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_947
timestamp 1698431365
transform 1 0 107408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_949
timestamp 1698431365
transform 1 0 107632 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_958
timestamp 1698431365
transform 1 0 108640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_962
timestamp 1698431365
transform 1 0 109088 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_970
timestamp 1698431365
transform 1 0 109984 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_975
timestamp 1698431365
transform 1 0 110544 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_983
timestamp 1698431365
transform 1 0 111440 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_987
timestamp 1698431365
transform 1 0 111888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_989
timestamp 1698431365
transform 1 0 112112 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_994
timestamp 1698431365
transform 1 0 112672 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1010
timestamp 1698431365
transform 1 0 114464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_1014
timestamp 1698431365
transform 1 0 114912 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1017
timestamp 1698431365
transform 1 0 115248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1081
timestamp 1698431365
transform 1 0 122416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1087
timestamp 1698431365
transform 1 0 123088 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1151
timestamp 1698431365
transform 1 0 130256 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1157
timestamp 1698431365
transform 1 0 130928 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1221
timestamp 1698431365
transform 1 0 138096 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1227
timestamp 1698431365
transform 1 0 138768 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1291
timestamp 1698431365
transform 1 0 145936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1297
timestamp 1698431365
transform 1 0 146608 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1361
timestamp 1698431365
transform 1 0 153776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_1367
timestamp 1698431365
transform 1 0 154448 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_1399
timestamp 1698431365
transform 1 0 158032 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_1401
timestamp 1698431365
transform 1 0 158256 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_158
timestamp 1698431365
transform 1 0 19040 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_161
timestamp 1698431365
transform 1 0 19376 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_183
timestamp 1698431365
transform 1 0 21840 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_191
timestamp 1698431365
transform 1 0 22736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_195
timestamp 1698431365
transform 1 0 23184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_197
timestamp 1698431365
transform 1 0 23408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_200
timestamp 1698431365
transform 1 0 23744 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698431365
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_220
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_222
timestamp 1698431365
transform 1 0 26208 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_231
timestamp 1698431365
transform 1 0 27216 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_235
timestamp 1698431365
transform 1 0 27664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_241
timestamp 1698431365
transform 1 0 28336 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_249
timestamp 1698431365
transform 1 0 29232 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_253
timestamp 1698431365
transform 1 0 29680 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_255
timestamp 1698431365
transform 1 0 29904 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_267
timestamp 1698431365
transform 1 0 31248 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_308
timestamp 1698431365
transform 1 0 35840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_312
timestamp 1698431365
transform 1 0 36288 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_320
timestamp 1698431365
transform 1 0 37184 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_324
timestamp 1698431365
transform 1 0 37632 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_338
timestamp 1698431365
transform 1 0 39200 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_381
timestamp 1698431365
transform 1 0 44016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_385
timestamp 1698431365
transform 1 0 44464 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_393
timestamp 1698431365
transform 1 0 45360 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_397
timestamp 1698431365
transform 1 0 45808 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_400
timestamp 1698431365
transform 1 0 46144 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_408
timestamp 1698431365
transform 1 0 47040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_418
timestamp 1698431365
transform 1 0 48160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_428
timestamp 1698431365
transform 1 0 49280 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_432
timestamp 1698431365
transform 1 0 49728 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_435
timestamp 1698431365
transform 1 0 50064 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_449
timestamp 1698431365
transform 1 0 51632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_453
timestamp 1698431365
transform 1 0 52080 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_457
timestamp 1698431365
transform 1 0 52528 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_487
timestamp 1698431365
transform 1 0 55888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_489
timestamp 1698431365
transform 1 0 56112 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_504
timestamp 1698431365
transform 1 0 57792 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_514
timestamp 1698431365
transform 1 0 58912 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_522
timestamp 1698431365
transform 1 0 59808 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_526
timestamp 1698431365
transform 1 0 60256 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_559
timestamp 1698431365
transform 1 0 63952 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_562
timestamp 1698431365
transform 1 0 64288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_566
timestamp 1698431365
transform 1 0 64736 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_574
timestamp 1698431365
transform 1 0 65632 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_632
timestamp 1698431365
transform 1 0 72128 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_662
timestamp 1698431365
transform 1 0 75488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_666
timestamp 1698431365
transform 1 0 75936 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_675
timestamp 1698431365
transform 1 0 76944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_679
timestamp 1698431365
transform 1 0 77392 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_683
timestamp 1698431365
transform 1 0 77840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_687
timestamp 1698431365
transform 1 0 78288 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_691
timestamp 1698431365
transform 1 0 78736 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_728
timestamp 1698431365
transform 1 0 82880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_732
timestamp 1698431365
transform 1 0 83328 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_766
timestamp 1698431365
transform 1 0 87136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_772
timestamp 1698431365
transform 1 0 87808 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_778
timestamp 1698431365
transform 1 0 88480 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_782
timestamp 1698431365
transform 1 0 88928 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_793
timestamp 1698431365
transform 1 0 90160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_797
timestamp 1698431365
transform 1 0 90608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_801
timestamp 1698431365
transform 1 0 91056 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_807
timestamp 1698431365
transform 1 0 91728 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_821
timestamp 1698431365
transform 1 0 93296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_833
timestamp 1698431365
transform 1 0 94640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_837
timestamp 1698431365
transform 1 0 95088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_839
timestamp 1698431365
transform 1 0 95312 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_842
timestamp 1698431365
transform 1 0 95648 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_868
timestamp 1698431365
transform 1 0 98560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_872
timestamp 1698431365
transform 1 0 99008 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_900
timestamp 1698431365
transform 1 0 102144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_904
timestamp 1698431365
transform 1 0 102592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_908
timestamp 1698431365
transform 1 0 103040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_912
timestamp 1698431365
transform 1 0 103488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_916
timestamp 1698431365
transform 1 0 103936 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_920
timestamp 1698431365
transform 1 0 104384 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_924
timestamp 1698431365
transform 1 0 104832 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_961
timestamp 1698431365
transform 1 0 108976 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_971
timestamp 1698431365
transform 1 0 110096 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_979
timestamp 1698431365
transform 1 0 110992 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_982
timestamp 1698431365
transform 1 0 111328 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_986
timestamp 1698431365
transform 1 0 111776 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_1023
timestamp 1698431365
transform 1 0 115920 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_1039
timestamp 1698431365
transform 1 0 117712 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_1047
timestamp 1698431365
transform 1 0 118608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_1049
timestamp 1698431365
transform 1 0 118832 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1052
timestamp 1698431365
transform 1 0 119168 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1116
timestamp 1698431365
transform 1 0 126336 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1122
timestamp 1698431365
transform 1 0 127008 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1186
timestamp 1698431365
transform 1 0 134176 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1192
timestamp 1698431365
transform 1 0 134848 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1256
timestamp 1698431365
transform 1 0 142016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1262
timestamp 1698431365
transform 1 0 142688 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1326
timestamp 1698431365
transform 1 0 149856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1332
timestamp 1698431365
transform 1 0 150528 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1396
timestamp 1698431365
transform 1 0 157696 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_205
timestamp 1698431365
transform 1 0 24304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_209
timestamp 1698431365
transform 1 0 24752 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_257
timestamp 1698431365
transform 1 0 30128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_301
timestamp 1698431365
transform 1 0 35056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_305
timestamp 1698431365
transform 1 0 35504 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_333
timestamp 1698431365
transform 1 0 38640 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_337
timestamp 1698431365
transform 1 0 39088 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_343
timestamp 1698431365
transform 1 0 39760 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_351
timestamp 1698431365
transform 1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_358
timestamp 1698431365
transform 1 0 41440 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_367
timestamp 1698431365
transform 1 0 42448 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_383
timestamp 1698431365
transform 1 0 44240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_399
timestamp 1698431365
transform 1 0 46032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_412
timestamp 1698431365
transform 1 0 47488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_414
timestamp 1698431365
transform 1 0 47712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_420
timestamp 1698431365
transform 1 0 48384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_422
timestamp 1698431365
transform 1 0 48608 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_446
timestamp 1698431365
transform 1 0 51296 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_454
timestamp 1698431365
transform 1 0 52192 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_461
timestamp 1698431365
transform 1 0 52976 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_477
timestamp 1698431365
transform 1 0 54768 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_517
timestamp 1698431365
transform 1 0 59248 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_521
timestamp 1698431365
transform 1 0 59696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_565
timestamp 1698431365
transform 1 0 64624 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_587
timestamp 1698431365
transform 1 0 67088 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_591
timestamp 1698431365
transform 1 0 67536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_597
timestamp 1698431365
transform 1 0 68208 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_599
timestamp 1698431365
transform 1 0 68432 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_642
timestamp 1698431365
transform 1 0 73248 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_648
timestamp 1698431365
transform 1 0 73920 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_652
timestamp 1698431365
transform 1 0 74368 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_660
timestamp 1698431365
transform 1 0 75264 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_664
timestamp 1698431365
transform 1 0 75712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_667
timestamp 1698431365
transform 1 0 76048 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_671
timestamp 1698431365
transform 1 0 76496 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_680
timestamp 1698431365
transform 1 0 77504 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_698
timestamp 1698431365
transform 1 0 79520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_732
timestamp 1698431365
transform 1 0 83328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_734
timestamp 1698431365
transform 1 0 83552 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_737
timestamp 1698431365
transform 1 0 83888 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_743
timestamp 1698431365
transform 1 0 84560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_757
timestamp 1698431365
transform 1 0 86128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_761
timestamp 1698431365
transform 1 0 86576 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_778
timestamp 1698431365
transform 1 0 88480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_782
timestamp 1698431365
transform 1 0 88928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_786
timestamp 1698431365
transform 1 0 89376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_790
timestamp 1698431365
transform 1 0 89824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_794
timestamp 1698431365
transform 1 0 90272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_800
timestamp 1698431365
transform 1 0 90944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_804
timestamp 1698431365
transform 1 0 91392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_807
timestamp 1698431365
transform 1 0 91728 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_813
timestamp 1698431365
transform 1 0 92400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_817
timestamp 1698431365
transform 1 0 92848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_821
timestamp 1698431365
transform 1 0 93296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_825
timestamp 1698431365
transform 1 0 93744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_827
timestamp 1698431365
transform 1 0 93968 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_858
timestamp 1698431365
transform 1 0 97440 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_867
timestamp 1698431365
transform 1 0 98448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_871
timestamp 1698431365
transform 1 0 98896 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_927
timestamp 1698431365
transform 1 0 105168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_943
timestamp 1698431365
transform 1 0 106960 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_955
timestamp 1698431365
transform 1 0 108304 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_959
timestamp 1698431365
transform 1 0 108752 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_992
timestamp 1698431365
transform 1 0 112448 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1008
timestamp 1698431365
transform 1 0 114240 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_1012
timestamp 1698431365
transform 1 0 114688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_1014
timestamp 1698431365
transform 1 0 114912 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1017
timestamp 1698431365
transform 1 0 115248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1081
timestamp 1698431365
transform 1 0 122416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1087
timestamp 1698431365
transform 1 0 123088 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1151
timestamp 1698431365
transform 1 0 130256 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1157
timestamp 1698431365
transform 1 0 130928 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1221
timestamp 1698431365
transform 1 0 138096 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1227
timestamp 1698431365
transform 1 0 138768 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1291
timestamp 1698431365
transform 1 0 145936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1297
timestamp 1698431365
transform 1 0 146608 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1361
timestamp 1698431365
transform 1 0 153776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_1367
timestamp 1698431365
transform 1 0 154448 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_1399
timestamp 1698431365
transform 1 0 158032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_1401
timestamp 1698431365
transform 1 0 158256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_174
timestamp 1698431365
transform 1 0 20832 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_216
timestamp 1698431365
transform 1 0 25536 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_222
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_230
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_234
timestamp 1698431365
transform 1 0 27552 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_242
timestamp 1698431365
transform 1 0 28448 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_244
timestamp 1698431365
transform 1 0 28672 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_247
timestamp 1698431365
transform 1 0 29008 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_251
timestamp 1698431365
transform 1 0 29456 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_253
timestamp 1698431365
transform 1 0 29680 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_262
timestamp 1698431365
transform 1 0 30688 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_270
timestamp 1698431365
transform 1 0 31584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_291
timestamp 1698431365
transform 1 0 33936 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_295
timestamp 1698431365
transform 1 0 34384 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_304
timestamp 1698431365
transform 1 0 35392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_308
timestamp 1698431365
transform 1 0 35840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_312
timestamp 1698431365
transform 1 0 36288 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_316
timestamp 1698431365
transform 1 0 36736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_356
timestamp 1698431365
transform 1 0 41216 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_358
timestamp 1698431365
transform 1 0 41440 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_380
timestamp 1698431365
transform 1 0 43904 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_388
timestamp 1698431365
transform 1 0 44800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_390
timestamp 1698431365
transform 1 0 45024 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_399
timestamp 1698431365
transform 1 0 46032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_403
timestamp 1698431365
transform 1 0 46480 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_407
timestamp 1698431365
transform 1 0 46928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_409
timestamp 1698431365
transform 1 0 47152 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_466
timestamp 1698431365
transform 1 0 53536 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_482
timestamp 1698431365
transform 1 0 55328 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_502
timestamp 1698431365
transform 1 0 57568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_506
timestamp 1698431365
transform 1 0 58016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_514
timestamp 1698431365
transform 1 0 58912 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_526
timestamp 1698431365
transform 1 0 60256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_599
timestamp 1698431365
transform 1 0 68432 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_603
timestamp 1698431365
transform 1 0 68880 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_616
timestamp 1698431365
transform 1 0 70336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_620
timestamp 1698431365
transform 1 0 70784 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_624
timestamp 1698431365
transform 1 0 71232 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_626
timestamp 1698431365
transform 1 0 71456 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_629
timestamp 1698431365
transform 1 0 71792 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_646
timestamp 1698431365
transform 1 0 73696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_656
timestamp 1698431365
transform 1 0 74816 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_660
timestamp 1698431365
transform 1 0 75264 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_670
timestamp 1698431365
transform 1 0 76384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_702
timestamp 1698431365
transform 1 0 79968 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_704
timestamp 1698431365
transform 1 0 80192 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_735
timestamp 1698431365
transform 1 0 83664 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_737
timestamp 1698431365
transform 1 0 83888 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_740
timestamp 1698431365
transform 1 0 84224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_744
timestamp 1698431365
transform 1 0 84672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_748
timestamp 1698431365
transform 1 0 85120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_752
timestamp 1698431365
transform 1 0 85568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_764
timestamp 1698431365
transform 1 0 86912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_768
timestamp 1698431365
transform 1 0 87360 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_802
timestamp 1698431365
transform 1 0 91168 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_812
timestamp 1698431365
transform 1 0 92288 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_821
timestamp 1698431365
transform 1 0 93296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_825
timestamp 1698431365
transform 1 0 93744 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_829
timestamp 1698431365
transform 1 0 94192 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_832
timestamp 1698431365
transform 1 0 94528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_836
timestamp 1698431365
transform 1 0 94976 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_876
timestamp 1698431365
transform 1 0 99456 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_886
timestamp 1698431365
transform 1 0 100576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_890
timestamp 1698431365
transform 1 0 101024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_900
timestamp 1698431365
transform 1 0 102144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_904
timestamp 1698431365
transform 1 0 102592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_908
timestamp 1698431365
transform 1 0 103040 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_912
timestamp 1698431365
transform 1 0 103488 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_928
timestamp 1698431365
transform 1 0 105280 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_940
timestamp 1698431365
transform 1 0 106624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_942
timestamp 1698431365
transform 1 0 106848 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_945
timestamp 1698431365
transform 1 0 107184 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_953
timestamp 1698431365
transform 1 0 108080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_957
timestamp 1698431365
transform 1 0 108528 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_968
timestamp 1698431365
transform 1 0 109760 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_976
timestamp 1698431365
transform 1 0 110656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_982
timestamp 1698431365
transform 1 0 111328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_984
timestamp 1698431365
transform 1 0 111552 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_993
timestamp 1698431365
transform 1 0 112560 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1009
timestamp 1698431365
transform 1 0 114352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_1017
timestamp 1698431365
transform 1 0 115248 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_1049
timestamp 1698431365
transform 1 0 118832 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1052
timestamp 1698431365
transform 1 0 119168 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1116
timestamp 1698431365
transform 1 0 126336 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1122
timestamp 1698431365
transform 1 0 127008 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1186
timestamp 1698431365
transform 1 0 134176 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1192
timestamp 1698431365
transform 1 0 134848 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1256
timestamp 1698431365
transform 1 0 142016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1262
timestamp 1698431365
transform 1 0 142688 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1326
timestamp 1698431365
transform 1 0 149856 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1332
timestamp 1698431365
transform 1 0 150528 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1396
timestamp 1698431365
transform 1 0 157696 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_185
timestamp 1698431365
transform 1 0 22064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_189
timestamp 1698431365
transform 1 0 22512 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_203
timestamp 1698431365
transform 1 0 24080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_207
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_211
timestamp 1698431365
transform 1 0 24976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_213
timestamp 1698431365
transform 1 0 25200 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_303
timestamp 1698431365
transform 1 0 35280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_329
timestamp 1698431365
transform 1 0 38192 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_333
timestamp 1698431365
transform 1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_335
timestamp 1698431365
transform 1 0 38864 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_379
timestamp 1698431365
transform 1 0 43792 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_383
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_439
timestamp 1698431365
transform 1 0 50512 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_468
timestamp 1698431365
transform 1 0 53760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_472
timestamp 1698431365
transform 1 0 54208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_474
timestamp 1698431365
transform 1 0 54432 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_484
timestamp 1698431365
transform 1 0 55552 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_490
timestamp 1698431365
transform 1 0 56224 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_506
timestamp 1698431365
transform 1 0 58016 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_519
timestamp 1698431365
transform 1 0 59472 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_523
timestamp 1698431365
transform 1 0 59920 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_527
timestamp 1698431365
transform 1 0 60368 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_538
timestamp 1698431365
transform 1 0 61600 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_589
timestamp 1698431365
transform 1 0 67312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_593
timestamp 1698431365
transform 1 0 67760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_597
timestamp 1698431365
transform 1 0 68208 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_649
timestamp 1698431365
transform 1 0 74032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_653
timestamp 1698431365
transform 1 0 74480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_717
timestamp 1698431365
transform 1 0 81648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_719
timestamp 1698431365
transform 1 0 81872 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_722
timestamp 1698431365
transform 1 0 82208 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_730
timestamp 1698431365
transform 1 0 83104 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_734
timestamp 1698431365
transform 1 0 83552 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_737
timestamp 1698431365
transform 1 0 83888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_745
timestamp 1698431365
transform 1 0 84784 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_748
timestamp 1698431365
transform 1 0 85120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_752
timestamp 1698431365
transform 1 0 85568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_756
timestamp 1698431365
transform 1 0 86016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_776
timestamp 1698431365
transform 1 0 88256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_780
timestamp 1698431365
transform 1 0 88704 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_796
timestamp 1698431365
transform 1 0 90496 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_807
timestamp 1698431365
transform 1 0 91728 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_811
timestamp 1698431365
transform 1 0 92176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_815
timestamp 1698431365
transform 1 0 92624 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_819
timestamp 1698431365
transform 1 0 93072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_821
timestamp 1698431365
transform 1 0 93296 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_824
timestamp 1698431365
transform 1 0 93632 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_828
timestamp 1698431365
transform 1 0 94080 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_831
timestamp 1698431365
transform 1 0 94416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_835
timestamp 1698431365
transform 1 0 94864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_837
timestamp 1698431365
transform 1 0 95088 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_840
timestamp 1698431365
transform 1 0 95424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_858
timestamp 1698431365
transform 1 0 97440 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_867
timestamp 1698431365
transform 1 0 98448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_871
timestamp 1698431365
transform 1 0 98896 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_877
timestamp 1698431365
transform 1 0 99568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_881
timestamp 1698431365
transform 1 0 100016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_885
timestamp 1698431365
transform 1 0 100464 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_917
timestamp 1698431365
transform 1 0 104048 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_927
timestamp 1698431365
transform 1 0 105168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_931
timestamp 1698431365
transform 1 0 105616 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_938
timestamp 1698431365
transform 1 0 106400 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_942
timestamp 1698431365
transform 1 0 106848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_944
timestamp 1698431365
transform 1 0 107072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_947
timestamp 1698431365
transform 1 0 107408 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_953
timestamp 1698431365
transform 1 0 108080 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_959
timestamp 1698431365
transform 1 0 108752 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_963
timestamp 1698431365
transform 1 0 109200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_967
timestamp 1698431365
transform 1 0 109648 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_983
timestamp 1698431365
transform 1 0 111440 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1001
timestamp 1698431365
transform 1 0 113456 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1009
timestamp 1698431365
transform 1 0 114352 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_1013
timestamp 1698431365
transform 1 0 114800 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1017
timestamp 1698431365
transform 1 0 115248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1081
timestamp 1698431365
transform 1 0 122416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1087
timestamp 1698431365
transform 1 0 123088 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1151
timestamp 1698431365
transform 1 0 130256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1157
timestamp 1698431365
transform 1 0 130928 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1221
timestamp 1698431365
transform 1 0 138096 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1227
timestamp 1698431365
transform 1 0 138768 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1291
timestamp 1698431365
transform 1 0 145936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1297
timestamp 1698431365
transform 1 0 146608 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1361
timestamp 1698431365
transform 1 0 153776 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_1367
timestamp 1698431365
transform 1 0 154448 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_1399
timestamp 1698431365
transform 1 0 158032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_1401
timestamp 1698431365
transform 1 0 158256 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_154
timestamp 1698431365
transform 1 0 18592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_156
timestamp 1698431365
transform 1 0 18816 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_186
timestamp 1698431365
transform 1 0 22176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_190
timestamp 1698431365
transform 1 0 22624 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_199
timestamp 1698431365
transform 1 0 23632 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698431365
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_231
timestamp 1698431365
transform 1 0 27216 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698431365
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_295
timestamp 1698431365
transform 1 0 34384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_297
timestamp 1698431365
transform 1 0 34608 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_334
timestamp 1698431365
transform 1 0 38752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_338
timestamp 1698431365
transform 1 0 39200 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_346
timestamp 1698431365
transform 1 0 40096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_361
timestamp 1698431365
transform 1 0 41776 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_369
timestamp 1698431365
transform 1 0 42672 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_385
timestamp 1698431365
transform 1 0 44464 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_417
timestamp 1698431365
transform 1 0 48048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_419
timestamp 1698431365
transform 1 0 48272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_426
timestamp 1698431365
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_428
timestamp 1698431365
transform 1 0 49280 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_455
timestamp 1698431365
transform 1 0 52304 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_466
timestamp 1698431365
transform 1 0 53536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_470
timestamp 1698431365
transform 1 0 53984 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_497
timestamp 1698431365
transform 1 0 57008 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_513
timestamp 1698431365
transform 1 0 58800 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_517
timestamp 1698431365
transform 1 0 59248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_536
timestamp 1698431365
transform 1 0 61376 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_552
timestamp 1698431365
transform 1 0 63168 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_566
timestamp 1698431365
transform 1 0 64736 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_596
timestamp 1698431365
transform 1 0 68096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_600
timestamp 1698431365
transform 1 0 68544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_618
timestamp 1698431365
transform 1 0 70560 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_626
timestamp 1698431365
transform 1 0 71456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_632
timestamp 1698431365
transform 1 0 72128 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_640
timestamp 1698431365
transform 1 0 73024 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_643
timestamp 1698431365
transform 1 0 73360 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_647
timestamp 1698431365
transform 1 0 73808 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_688
timestamp 1698431365
transform 1 0 78400 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_696
timestamp 1698431365
transform 1 0 79296 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_702
timestamp 1698431365
transform 1 0 79968 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_728
timestamp 1698431365
transform 1 0 82880 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_744
timestamp 1698431365
transform 1 0 84672 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_748
timestamp 1698431365
transform 1 0 85120 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_751
timestamp 1698431365
transform 1 0 85456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_769
timestamp 1698431365
transform 1 0 87472 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_772
timestamp 1698431365
transform 1 0 87808 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_788
timestamp 1698431365
transform 1 0 89600 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_822
timestamp 1698431365
transform 1 0 93408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_826
timestamp 1698431365
transform 1 0 93856 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_836
timestamp 1698431365
transform 1 0 94976 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_864
timestamp 1698431365
transform 1 0 98112 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_895
timestamp 1698431365
transform 1 0 101584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_899
timestamp 1698431365
transform 1 0 102032 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_907
timestamp 1698431365
transform 1 0 102928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_909
timestamp 1698431365
transform 1 0 103152 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_912
timestamp 1698431365
transform 1 0 103488 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_920
timestamp 1698431365
transform 1 0 104384 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_943
timestamp 1698431365
transform 1 0 106960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_947
timestamp 1698431365
transform 1 0 107408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_975
timestamp 1698431365
transform 1 0 110544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_977
timestamp 1698431365
transform 1 0 110768 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_982
timestamp 1698431365
transform 1 0 111328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_986
timestamp 1698431365
transform 1 0 111776 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_1003
timestamp 1698431365
transform 1 0 113680 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_1007
timestamp 1698431365
transform 1 0 114128 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_1039
timestamp 1698431365
transform 1 0 117712 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_1047
timestamp 1698431365
transform 1 0 118608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_1049
timestamp 1698431365
transform 1 0 118832 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1052
timestamp 1698431365
transform 1 0 119168 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1116
timestamp 1698431365
transform 1 0 126336 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1122
timestamp 1698431365
transform 1 0 127008 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1186
timestamp 1698431365
transform 1 0 134176 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1192
timestamp 1698431365
transform 1 0 134848 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1256
timestamp 1698431365
transform 1 0 142016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1262
timestamp 1698431365
transform 1 0 142688 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1326
timestamp 1698431365
transform 1 0 149856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1332
timestamp 1698431365
transform 1 0 150528 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1396
timestamp 1698431365
transform 1 0 157696 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_193
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_205
timestamp 1698431365
transform 1 0 24304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_209
timestamp 1698431365
transform 1 0 24752 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_213
timestamp 1698431365
transform 1 0 25200 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_221
timestamp 1698431365
transform 1 0 26096 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_229
timestamp 1698431365
transform 1 0 26992 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_253
timestamp 1698431365
transform 1 0 29680 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_257
timestamp 1698431365
transform 1 0 30128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_259
timestamp 1698431365
transform 1 0 30352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698431365
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_330
timestamp 1698431365
transform 1 0 38304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_334
timestamp 1698431365
transform 1 0 38752 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_350
timestamp 1698431365
transform 1 0 40544 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_371
timestamp 1698431365
transform 1 0 42896 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_379
timestamp 1698431365
transform 1 0 43792 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_389
timestamp 1698431365
transform 1 0 44912 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_403
timestamp 1698431365
transform 1 0 46480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_405
timestamp 1698431365
transform 1 0 46704 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_437
timestamp 1698431365
transform 1 0 50288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_465
timestamp 1698431365
transform 1 0 53424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_469
timestamp 1698431365
transform 1 0 53872 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_482
timestamp 1698431365
transform 1 0 55328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_502
timestamp 1698431365
transform 1 0 57568 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_506
timestamp 1698431365
transform 1 0 58016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_510
timestamp 1698431365
transform 1 0 58464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_539
timestamp 1698431365
transform 1 0 61712 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_547
timestamp 1698431365
transform 1 0 62608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_551
timestamp 1698431365
transform 1 0 63056 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_589
timestamp 1698431365
transform 1 0 67312 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_593
timestamp 1698431365
transform 1 0 67760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_597
timestamp 1698431365
transform 1 0 68208 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_629
timestamp 1698431365
transform 1 0 71792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_661
timestamp 1698431365
transform 1 0 75376 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_667
timestamp 1698431365
transform 1 0 76048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_669
timestamp 1698431365
transform 1 0 76272 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_694
timestamp 1698431365
transform 1 0 79072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_698
timestamp 1698431365
transform 1 0 79520 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_718
timestamp 1698431365
transform 1 0 81760 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_734
timestamp 1698431365
transform 1 0 83552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_737
timestamp 1698431365
transform 1 0 83888 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_745
timestamp 1698431365
transform 1 0 84784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_747
timestamp 1698431365
transform 1 0 85008 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_778
timestamp 1698431365
transform 1 0 88480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_782
timestamp 1698431365
transform 1 0 88928 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_798
timestamp 1698431365
transform 1 0 90720 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_802
timestamp 1698431365
transform 1 0 91168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_823
timestamp 1698431365
transform 1 0 93520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_827
timestamp 1698431365
transform 1 0 93968 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_835
timestamp 1698431365
transform 1 0 94864 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_839
timestamp 1698431365
transform 1 0 95312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_871
timestamp 1698431365
transform 1 0 98896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_877
timestamp 1698431365
transform 1 0 99568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_909
timestamp 1698431365
transform 1 0 103152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_942
timestamp 1698431365
transform 1 0 106848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_944
timestamp 1698431365
transform 1 0 107072 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_947
timestamp 1698431365
transform 1 0 107408 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_951
timestamp 1698431365
transform 1 0 107856 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_984
timestamp 1698431365
transform 1 0 111552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1017
timestamp 1698431365
transform 1 0 115248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1081
timestamp 1698431365
transform 1 0 122416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1087
timestamp 1698431365
transform 1 0 123088 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1151
timestamp 1698431365
transform 1 0 130256 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1157
timestamp 1698431365
transform 1 0 130928 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1221
timestamp 1698431365
transform 1 0 138096 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1227
timestamp 1698431365
transform 1 0 138768 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1291
timestamp 1698431365
transform 1 0 145936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1297
timestamp 1698431365
transform 1 0 146608 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1361
timestamp 1698431365
transform 1 0 153776 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_1367
timestamp 1698431365
transform 1 0 154448 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_1399
timestamp 1698431365
transform 1 0 158032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_1401
timestamp 1698431365
transform 1 0 158256 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_174
timestamp 1698431365
transform 1 0 20832 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_216
timestamp 1698431365
transform 1 0 25536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_218
timestamp 1698431365
transform 1 0 25760 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_254
timestamp 1698431365
transform 1 0 29792 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_258
timestamp 1698431365
transform 1 0 30240 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_266
timestamp 1698431365
transform 1 0 31136 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_273
timestamp 1698431365
transform 1 0 31920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698431365
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_288
timestamp 1698431365
transform 1 0 33600 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_297
timestamp 1698431365
transform 1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_301
timestamp 1698431365
transform 1 0 35056 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_309
timestamp 1698431365
transform 1 0 35952 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_313
timestamp 1698431365
transform 1 0 36400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_317
timestamp 1698431365
transform 1 0 36848 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_356
timestamp 1698431365
transform 1 0 41216 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_365
timestamp 1698431365
transform 1 0 42224 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_369
timestamp 1698431365
transform 1 0 42672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_371
timestamp 1698431365
transform 1 0 42896 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_374
timestamp 1698431365
transform 1 0 43232 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_383
timestamp 1698431365
transform 1 0 44240 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_399
timestamp 1698431365
transform 1 0 46032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_417
timestamp 1698431365
transform 1 0 48048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_419
timestamp 1698431365
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_426
timestamp 1698431365
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_430
timestamp 1698431365
transform 1 0 49504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_432
timestamp 1698431365
transform 1 0 49728 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_435
timestamp 1698431365
transform 1 0 50064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_447
timestamp 1698431365
transform 1 0 51408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_464
timestamp 1698431365
transform 1 0 53312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_474
timestamp 1698431365
transform 1 0 54432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_476
timestamp 1698431365
transform 1 0 54656 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_500
timestamp 1698431365
transform 1 0 57344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_508
timestamp 1698431365
transform 1 0 58240 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_512
timestamp 1698431365
transform 1 0 58688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_514
timestamp 1698431365
transform 1 0 58912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_533
timestamp 1698431365
transform 1 0 61040 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_549
timestamp 1698431365
transform 1 0 62832 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_557
timestamp 1698431365
transform 1 0 63728 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_559
timestamp 1698431365
transform 1 0 63952 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_591
timestamp 1698431365
transform 1 0 67536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_595
timestamp 1698431365
transform 1 0 67984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_599
timestamp 1698431365
transform 1 0 68432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_601
timestamp 1698431365
transform 1 0 68656 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_610
timestamp 1698431365
transform 1 0 69664 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_626
timestamp 1698431365
transform 1 0 71456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_632
timestamp 1698431365
transform 1 0 72128 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_640
timestamp 1698431365
transform 1 0 73024 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_644
timestamp 1698431365
transform 1 0 73472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_654
timestamp 1698431365
transform 1 0 74592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_659
timestamp 1698431365
transform 1 0 75152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_663
timestamp 1698431365
transform 1 0 75600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_667
timestamp 1698431365
transform 1 0 76048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_669
timestamp 1698431365
transform 1 0 76272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_702
timestamp 1698431365
transform 1 0 79968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_706
timestamp 1698431365
transform 1 0 80416 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_714
timestamp 1698431365
transform 1 0 81312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_724
timestamp 1698431365
transform 1 0 82432 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_768
timestamp 1698431365
transform 1 0 87360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_780
timestamp 1698431365
transform 1 0 88704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_788
timestamp 1698431365
transform 1 0 89600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_792
timestamp 1698431365
transform 1 0 90048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_832
timestamp 1698431365
transform 1 0 94528 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_842
timestamp 1698431365
transform 1 0 95648 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_868
timestamp 1698431365
transform 1 0 98560 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_900
timestamp 1698431365
transform 1 0 102144 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_912
timestamp 1698431365
transform 1 0 103488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_914
timestamp 1698431365
transform 1 0 103712 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_923
timestamp 1698431365
transform 1 0 104720 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_963
timestamp 1698431365
transform 1 0 109200 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_979
timestamp 1698431365
transform 1 0 110992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_982
timestamp 1698431365
transform 1 0 111328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1046
timestamp 1698431365
transform 1 0 118496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1052
timestamp 1698431365
transform 1 0 119168 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1116
timestamp 1698431365
transform 1 0 126336 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1122
timestamp 1698431365
transform 1 0 127008 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1186
timestamp 1698431365
transform 1 0 134176 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1192
timestamp 1698431365
transform 1 0 134848 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1256
timestamp 1698431365
transform 1 0 142016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1262
timestamp 1698431365
transform 1 0 142688 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1326
timestamp 1698431365
transform 1 0 149856 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1332
timestamp 1698431365
transform 1 0 150528 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1396
timestamp 1698431365
transform 1 0 157696 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_193
timestamp 1698431365
transform 1 0 22960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_205
timestamp 1698431365
transform 1 0 24304 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_221
timestamp 1698431365
transform 1 0 26096 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_229
timestamp 1698431365
transform 1 0 26992 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_233
timestamp 1698431365
transform 1 0 27440 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_252
timestamp 1698431365
transform 1 0 29568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_256
timestamp 1698431365
transform 1 0 30016 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_272
timestamp 1698431365
transform 1 0 31808 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_276
timestamp 1698431365
transform 1 0 32256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_346
timestamp 1698431365
transform 1 0 40096 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_350
timestamp 1698431365
transform 1 0 40544 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_358
timestamp 1698431365
transform 1 0 41440 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_362
timestamp 1698431365
transform 1 0 41888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_380
timestamp 1698431365
transform 1 0 43904 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_384
timestamp 1698431365
transform 1 0 44352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_451
timestamp 1698431365
transform 1 0 51856 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_513
timestamp 1698431365
transform 1 0 58800 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_517
timestamp 1698431365
transform 1 0 59248 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_535
timestamp 1698431365
transform 1 0 61264 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_567
timestamp 1698431365
transform 1 0 64848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_571
timestamp 1698431365
transform 1 0 65296 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_587
timestamp 1698431365
transform 1 0 67088 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_626
timestamp 1698431365
transform 1 0 71456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_630
timestamp 1698431365
transform 1 0 71904 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_646
timestamp 1698431365
transform 1 0 73696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_650
timestamp 1698431365
transform 1 0 74144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_660
timestamp 1698431365
transform 1 0 75264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_662
timestamp 1698431365
transform 1 0 75488 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_667
timestamp 1698431365
transform 1 0 76048 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_683
timestamp 1698431365
transform 1 0 77840 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_691
timestamp 1698431365
transform 1 0 78736 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_696
timestamp 1698431365
transform 1 0 79296 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_704
timestamp 1698431365
transform 1 0 80192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_737
timestamp 1698431365
transform 1 0 83888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_741
timestamp 1698431365
transform 1 0 84336 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_781
timestamp 1698431365
transform 1 0 88816 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_789
timestamp 1698431365
transform 1 0 89712 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_793
timestamp 1698431365
transform 1 0 90160 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_804
timestamp 1698431365
transform 1 0 91392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_815
timestamp 1698431365
transform 1 0 92624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_847
timestamp 1698431365
transform 1 0 96208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_851
timestamp 1698431365
transform 1 0 96656 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_867
timestamp 1698431365
transform 1 0 98448 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_927
timestamp 1698431365
transform 1 0 105168 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_943
timestamp 1698431365
transform 1 0 106960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_947
timestamp 1698431365
transform 1 0 107408 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1011
timestamp 1698431365
transform 1 0 114576 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1017
timestamp 1698431365
transform 1 0 115248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1081
timestamp 1698431365
transform 1 0 122416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1087
timestamp 1698431365
transform 1 0 123088 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1151
timestamp 1698431365
transform 1 0 130256 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1157
timestamp 1698431365
transform 1 0 130928 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1221
timestamp 1698431365
transform 1 0 138096 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1227
timestamp 1698431365
transform 1 0 138768 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1291
timestamp 1698431365
transform 1 0 145936 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1297
timestamp 1698431365
transform 1 0 146608 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1361
timestamp 1698431365
transform 1 0 153776 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_1367
timestamp 1698431365
transform 1 0 154448 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_1399
timestamp 1698431365
transform 1 0 158032 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_1401
timestamp 1698431365
transform 1 0 158256 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_174
timestamp 1698431365
transform 1 0 20832 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_178
timestamp 1698431365
transform 1 0 21280 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_180
timestamp 1698431365
transform 1 0 21504 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_217
timestamp 1698431365
transform 1 0 25648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_221
timestamp 1698431365
transform 1 0 26096 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_229
timestamp 1698431365
transform 1 0 26992 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_233
timestamp 1698431365
transform 1 0 27440 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_239
timestamp 1698431365
transform 1 0 28112 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_271
timestamp 1698431365
transform 1 0 31696 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_284
timestamp 1698431365
transform 1 0 33152 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_295
timestamp 1698431365
transform 1 0 34384 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_327
timestamp 1698431365
transform 1 0 37968 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_335
timestamp 1698431365
transform 1 0 38864 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_343
timestamp 1698431365
transform 1 0 39760 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_347
timestamp 1698431365
transform 1 0 40208 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_370
timestamp 1698431365
transform 1 0 42784 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_374
timestamp 1698431365
transform 1 0 43232 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_384
timestamp 1698431365
transform 1 0 44352 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_388
timestamp 1698431365
transform 1 0 44800 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_428
timestamp 1698431365
transform 1 0 49280 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_450
timestamp 1698431365
transform 1 0 51744 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_454
timestamp 1698431365
transform 1 0 52192 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_471
timestamp 1698431365
transform 1 0 54096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_502
timestamp 1698431365
transform 1 0 57568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_506
timestamp 1698431365
transform 1 0 58016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_517
timestamp 1698431365
transform 1 0 59248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_521
timestamp 1698431365
transform 1 0 59696 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_555
timestamp 1698431365
transform 1 0 63504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_557
timestamp 1698431365
transform 1 0 63728 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_568
timestamp 1698431365
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_570
timestamp 1698431365
transform 1 0 65184 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_577
timestamp 1698431365
transform 1 0 65968 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_609
timestamp 1698431365
transform 1 0 69552 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_625
timestamp 1698431365
transform 1 0 71344 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_629
timestamp 1698431365
transform 1 0 71792 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_632
timestamp 1698431365
transform 1 0 72128 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_671
timestamp 1698431365
transform 1 0 76496 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_687
timestamp 1698431365
transform 1 0 78288 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_696
timestamp 1698431365
transform 1 0 79296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_736
timestamp 1698431365
transform 1 0 83776 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_740
timestamp 1698431365
transform 1 0 84224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_744
timestamp 1698431365
transform 1 0 84672 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_752
timestamp 1698431365
transform 1 0 85568 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_756
timestamp 1698431365
transform 1 0 86016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_766
timestamp 1698431365
transform 1 0 87136 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_772
timestamp 1698431365
transform 1 0 87808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_780
timestamp 1698431365
transform 1 0 88704 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_784
timestamp 1698431365
transform 1 0 89152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_786
timestamp 1698431365
transform 1 0 89376 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_825
timestamp 1698431365
transform 1 0 93744 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_833
timestamp 1698431365
transform 1 0 94640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_837
timestamp 1698431365
transform 1 0 95088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_839
timestamp 1698431365
transform 1 0 95312 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_842
timestamp 1698431365
transform 1 0 95648 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_906
timestamp 1698431365
transform 1 0 102816 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_912
timestamp 1698431365
transform 1 0 103488 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_976
timestamp 1698431365
transform 1 0 110656 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_982
timestamp 1698431365
transform 1 0 111328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1046
timestamp 1698431365
transform 1 0 118496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1052
timestamp 1698431365
transform 1 0 119168 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1116
timestamp 1698431365
transform 1 0 126336 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1122
timestamp 1698431365
transform 1 0 127008 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1186
timestamp 1698431365
transform 1 0 134176 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1192
timestamp 1698431365
transform 1 0 134848 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1256
timestamp 1698431365
transform 1 0 142016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1262
timestamp 1698431365
transform 1 0 142688 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1326
timestamp 1698431365
transform 1 0 149856 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1332
timestamp 1698431365
transform 1 0 150528 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1396
timestamp 1698431365
transform 1 0 157696 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_209
timestamp 1698431365
transform 1 0 24752 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_225
timestamp 1698431365
transform 1 0 26544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_227
timestamp 1698431365
transform 1 0 26768 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_263
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_293
timestamp 1698431365
transform 1 0 34160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_297
timestamp 1698431365
transform 1 0 34608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_307
timestamp 1698431365
transform 1 0 35728 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_333
timestamp 1698431365
transform 1 0 38640 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_337
timestamp 1698431365
transform 1 0 39088 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_346
timestamp 1698431365
transform 1 0 40096 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_350
timestamp 1698431365
transform 1 0 40544 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_366
timestamp 1698431365
transform 1 0 42336 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_368
timestamp 1698431365
transform 1 0 42560 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_375
timestamp 1698431365
transform 1 0 43344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_379
timestamp 1698431365
transform 1 0 43792 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_383
timestamp 1698431365
transform 1 0 44240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_391
timestamp 1698431365
transform 1 0 45136 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_416
timestamp 1698431365
transform 1 0 47936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_420
timestamp 1698431365
transform 1 0 48384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_424
timestamp 1698431365
transform 1 0 48832 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_432
timestamp 1698431365
transform 1 0 49728 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_434
timestamp 1698431365
transform 1 0 49952 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_461
timestamp 1698431365
transform 1 0 52976 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_465
timestamp 1698431365
transform 1 0 53424 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_509
timestamp 1698431365
transform 1 0 58352 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_513
timestamp 1698431365
transform 1 0 58800 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_519
timestamp 1698431365
transform 1 0 59472 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_523
timestamp 1698431365
transform 1 0 59920 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_527
timestamp 1698431365
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_536
timestamp 1698431365
transform 1 0 61376 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_552
timestamp 1698431365
transform 1 0 63168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_560
timestamp 1698431365
transform 1 0 64064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_562
timestamp 1698431365
transform 1 0 64288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_597
timestamp 1698431365
transform 1 0 68208 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_599
timestamp 1698431365
transform 1 0 68432 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_609
timestamp 1698431365
transform 1 0 69552 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_625
timestamp 1698431365
transform 1 0 71344 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_633
timestamp 1698431365
transform 1 0 72240 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_637
timestamp 1698431365
transform 1 0 72688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_647
timestamp 1698431365
transform 1 0 73808 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_661
timestamp 1698431365
transform 1 0 75376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_667
timestamp 1698431365
transform 1 0 76048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_669
timestamp 1698431365
transform 1 0 76272 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_676
timestamp 1698431365
transform 1 0 77056 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_684
timestamp 1698431365
transform 1 0 77952 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_737
timestamp 1698431365
transform 1 0 83888 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_753
timestamp 1698431365
transform 1 0 85680 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_757
timestamp 1698431365
transform 1 0 86128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_759
timestamp 1698431365
transform 1 0 86352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_766
timestamp 1698431365
transform 1 0 87136 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_798
timestamp 1698431365
transform 1 0 90720 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_802
timestamp 1698431365
transform 1 0 91168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_804
timestamp 1698431365
transform 1 0 91392 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_807
timestamp 1698431365
transform 1 0 91728 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_817
timestamp 1698431365
transform 1 0 92848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_821
timestamp 1698431365
transform 1 0 93296 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_853
timestamp 1698431365
transform 1 0 96880 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_869
timestamp 1698431365
transform 1 0 98672 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_873
timestamp 1698431365
transform 1 0 99120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_877
timestamp 1698431365
transform 1 0 99568 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_941
timestamp 1698431365
transform 1 0 106736 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_947
timestamp 1698431365
transform 1 0 107408 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1011
timestamp 1698431365
transform 1 0 114576 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1017
timestamp 1698431365
transform 1 0 115248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1081
timestamp 1698431365
transform 1 0 122416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1087
timestamp 1698431365
transform 1 0 123088 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1151
timestamp 1698431365
transform 1 0 130256 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1157
timestamp 1698431365
transform 1 0 130928 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1221
timestamp 1698431365
transform 1 0 138096 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1227
timestamp 1698431365
transform 1 0 138768 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1291
timestamp 1698431365
transform 1 0 145936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1297
timestamp 1698431365
transform 1 0 146608 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1361
timestamp 1698431365
transform 1 0 153776 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_1367
timestamp 1698431365
transform 1 0 154448 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_1399
timestamp 1698431365
transform 1 0 158032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_1401
timestamp 1698431365
transform 1 0 158256 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_174
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_190
timestamp 1698431365
transform 1 0 22624 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_194
timestamp 1698431365
transform 1 0 23072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_228
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_258
timestamp 1698431365
transform 1 0 30240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_262
timestamp 1698431365
transform 1 0 30688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_294
timestamp 1698431365
transform 1 0 34272 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_296
timestamp 1698431365
transform 1 0 34496 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_325
timestamp 1698431365
transform 1 0 37744 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_333
timestamp 1698431365
transform 1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_335
timestamp 1698431365
transform 1 0 38864 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_338
timestamp 1698431365
transform 1 0 39200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_368
timestamp 1698431365
transform 1 0 42560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_370
timestamp 1698431365
transform 1 0 42784 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_388
timestamp 1698431365
transform 1 0 44800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_392
timestamp 1698431365
transform 1 0 45248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_400
timestamp 1698431365
transform 1 0 46144 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_409
timestamp 1698431365
transform 1 0 47152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_417
timestamp 1698431365
transform 1 0 48048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_419
timestamp 1698431365
transform 1 0 48272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_424
timestamp 1698431365
transform 1 0 48832 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_431
timestamp 1698431365
transform 1 0 49616 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_435
timestamp 1698431365
transform 1 0 50064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_447
timestamp 1698431365
transform 1 0 51408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_451
timestamp 1698431365
transform 1 0 51856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_461
timestamp 1698431365
transform 1 0 52976 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_477
timestamp 1698431365
transform 1 0 54768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_513
timestamp 1698431365
transform 1 0 58800 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_522
timestamp 1698431365
transform 1 0 59808 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_538
timestamp 1698431365
transform 1 0 61600 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_542
timestamp 1698431365
transform 1 0 62048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_544
timestamp 1698431365
transform 1 0 62272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_547
timestamp 1698431365
transform 1 0 62608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_551
timestamp 1698431365
transform 1 0 63056 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_559
timestamp 1698431365
transform 1 0 63952 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_568
timestamp 1698431365
transform 1 0 64960 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_584
timestamp 1698431365
transform 1 0 66752 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_588
timestamp 1698431365
transform 1 0 67200 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_626
timestamp 1698431365
transform 1 0 71456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_632
timestamp 1698431365
transform 1 0 72128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_667
timestamp 1698431365
transform 1 0 76048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_669
timestamp 1698431365
transform 1 0 76272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_676
timestamp 1698431365
transform 1 0 77056 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_684
timestamp 1698431365
transform 1 0 77952 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_693
timestamp 1698431365
transform 1 0 78960 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_697
timestamp 1698431365
transform 1 0 79408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_699
timestamp 1698431365
transform 1 0 79632 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_702
timestamp 1698431365
transform 1 0 79968 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_706
timestamp 1698431365
transform 1 0 80416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_744
timestamp 1698431365
transform 1 0 84672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_748
timestamp 1698431365
transform 1 0 85120 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_764
timestamp 1698431365
transform 1 0 86912 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_768
timestamp 1698431365
transform 1 0 87360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_772
timestamp 1698431365
transform 1 0 87808 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_836
timestamp 1698431365
transform 1 0 94976 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_842
timestamp 1698431365
transform 1 0 95648 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_906
timestamp 1698431365
transform 1 0 102816 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_912
timestamp 1698431365
transform 1 0 103488 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_944
timestamp 1698431365
transform 1 0 107072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_947
timestamp 1698431365
transform 1 0 107408 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_979
timestamp 1698431365
transform 1 0 110992 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_982
timestamp 1698431365
transform 1 0 111328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1046
timestamp 1698431365
transform 1 0 118496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1052
timestamp 1698431365
transform 1 0 119168 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1116
timestamp 1698431365
transform 1 0 126336 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1122
timestamp 1698431365
transform 1 0 127008 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1186
timestamp 1698431365
transform 1 0 134176 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1192
timestamp 1698431365
transform 1 0 134848 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1256
timestamp 1698431365
transform 1 0 142016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1262
timestamp 1698431365
transform 1 0 142688 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1326
timestamp 1698431365
transform 1 0 149856 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1332
timestamp 1698431365
transform 1 0 150528 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1396
timestamp 1698431365
transform 1 0 157696 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_193
timestamp 1698431365
transform 1 0 22960 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_195
timestamp 1698431365
transform 1 0 23184 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_226
timestamp 1698431365
transform 1 0 26656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_230
timestamp 1698431365
transform 1 0 27104 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698431365
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698431365
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_275
timestamp 1698431365
transform 1 0 32144 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_283
timestamp 1698431365
transform 1 0 33040 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_287
timestamp 1698431365
transform 1 0 33488 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_319
timestamp 1698431365
transform 1 0 37072 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_352
timestamp 1698431365
transform 1 0 40768 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_361
timestamp 1698431365
transform 1 0 41776 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_369
timestamp 1698431365
transform 1 0 42672 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_373
timestamp 1698431365
transform 1 0 43120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_382
timestamp 1698431365
transform 1 0 44128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_395
timestamp 1698431365
transform 1 0 45584 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_404
timestamp 1698431365
transform 1 0 46592 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_408
timestamp 1698431365
transform 1 0 47040 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_419
timestamp 1698431365
transform 1 0 48272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_431
timestamp 1698431365
transform 1 0 49616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_433
timestamp 1698431365
transform 1 0 49840 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_444
timestamp 1698431365
transform 1 0 51072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_448
timestamp 1698431365
transform 1 0 51520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_452
timestamp 1698431365
transform 1 0 51968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_459
timestamp 1698431365
transform 1 0 52752 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_523
timestamp 1698431365
transform 1 0 59920 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_527
timestamp 1698431365
transform 1 0 60368 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_545
timestamp 1698431365
transform 1 0 62384 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_575
timestamp 1698431365
transform 1 0 65744 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_591
timestamp 1698431365
transform 1 0 67536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_597
timestamp 1698431365
transform 1 0 68208 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_601
timestamp 1698431365
transform 1 0 68656 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_625
timestamp 1698431365
transform 1 0 71344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_629
timestamp 1698431365
transform 1 0 71792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_633
timestamp 1698431365
transform 1 0 72240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_659
timestamp 1698431365
transform 1 0 75152 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_663
timestamp 1698431365
transform 1 0 75600 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_667
timestamp 1698431365
transform 1 0 76048 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_675
timestamp 1698431365
transform 1 0 76944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_677
timestamp 1698431365
transform 1 0 77168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_708
timestamp 1698431365
transform 1 0 80640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_712
timestamp 1698431365
transform 1 0 81088 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_728
timestamp 1698431365
transform 1 0 82880 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_732
timestamp 1698431365
transform 1 0 83328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_734
timestamp 1698431365
transform 1 0 83552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_737
timestamp 1698431365
transform 1 0 83888 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_753
timestamp 1698431365
transform 1 0 85680 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_761
timestamp 1698431365
transform 1 0 86576 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_765
timestamp 1698431365
transform 1 0 87024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_777
timestamp 1698431365
transform 1 0 88368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_792
timestamp 1698431365
transform 1 0 90048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_796
timestamp 1698431365
transform 1 0 90496 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_804
timestamp 1698431365
transform 1 0 91392 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_807
timestamp 1698431365
transform 1 0 91728 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_871
timestamp 1698431365
transform 1 0 98896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_877
timestamp 1698431365
transform 1 0 99568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_881
timestamp 1698431365
transform 1 0 100016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_883
timestamp 1698431365
transform 1 0 100240 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_895
timestamp 1698431365
transform 1 0 101584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_899
timestamp 1698431365
transform 1 0 102032 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_915
timestamp 1698431365
transform 1 0 103824 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_923
timestamp 1698431365
transform 1 0 104720 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_927
timestamp 1698431365
transform 1 0 105168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_929
timestamp 1698431365
transform 1 0 105392 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_932
timestamp 1698431365
transform 1 0 105728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_956
timestamp 1698431365
transform 1 0 108416 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_960
timestamp 1698431365
transform 1 0 108864 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_992
timestamp 1698431365
transform 1 0 112448 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1008
timestamp 1698431365
transform 1 0 114240 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_1012
timestamp 1698431365
transform 1 0 114688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_1014
timestamp 1698431365
transform 1 0 114912 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1017
timestamp 1698431365
transform 1 0 115248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1081
timestamp 1698431365
transform 1 0 122416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1087
timestamp 1698431365
transform 1 0 123088 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1151
timestamp 1698431365
transform 1 0 130256 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1157
timestamp 1698431365
transform 1 0 130928 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1221
timestamp 1698431365
transform 1 0 138096 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1227
timestamp 1698431365
transform 1 0 138768 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1291
timestamp 1698431365
transform 1 0 145936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1297
timestamp 1698431365
transform 1 0 146608 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1361
timestamp 1698431365
transform 1 0 153776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_1367
timestamp 1698431365
transform 1 0 154448 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_1399
timestamp 1698431365
transform 1 0 158032 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_1401
timestamp 1698431365
transform 1 0 158256 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698431365
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_174
timestamp 1698431365
transform 1 0 20832 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_190
timestamp 1698431365
transform 1 0 22624 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_198
timestamp 1698431365
transform 1 0 23520 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_202
timestamp 1698431365
transform 1 0 23968 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_222
timestamp 1698431365
transform 1 0 26208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_228
timestamp 1698431365
transform 1 0 26880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_232
timestamp 1698431365
transform 1 0 27328 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_248
timestamp 1698431365
transform 1 0 29120 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_302
timestamp 1698431365
transform 1 0 35168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_318
timestamp 1698431365
transform 1 0 36960 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_326
timestamp 1698431365
transform 1 0 37856 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_365
timestamp 1698431365
transform 1 0 42224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_379
timestamp 1698431365
transform 1 0 43792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_381
timestamp 1698431365
transform 1 0 44016 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_396
timestamp 1698431365
transform 1 0 45696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_400
timestamp 1698431365
transform 1 0 46144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_404
timestamp 1698431365
transform 1 0 46592 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_412
timestamp 1698431365
transform 1 0 47488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_414
timestamp 1698431365
transform 1 0 47712 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_446
timestamp 1698431365
transform 1 0 51296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_448
timestamp 1698431365
transform 1 0 51520 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_455
timestamp 1698431365
transform 1 0 52304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_457
timestamp 1698431365
transform 1 0 52528 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_478
timestamp 1698431365
transform 1 0 54880 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_482
timestamp 1698431365
transform 1 0 55328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_484
timestamp 1698431365
transform 1 0 55552 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_494
timestamp 1698431365
transform 1 0 56672 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_535
timestamp 1698431365
transform 1 0 61264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_539
timestamp 1698431365
transform 1 0 61712 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_543
timestamp 1698431365
transform 1 0 62160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_570
timestamp 1698431365
transform 1 0 65184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_574
timestamp 1698431365
transform 1 0 65632 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_582
timestamp 1698431365
transform 1 0 66528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_584
timestamp 1698431365
transform 1 0 66752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_621
timestamp 1698431365
transform 1 0 70896 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_625
timestamp 1698431365
transform 1 0 71344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_627
timestamp 1698431365
transform 1 0 71568 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_667
timestamp 1698431365
transform 1 0 76048 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_671
timestamp 1698431365
transform 1 0 76496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_673
timestamp 1698431365
transform 1 0 76720 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_684
timestamp 1698431365
transform 1 0 77952 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_702
timestamp 1698431365
transform 1 0 79968 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_734
timestamp 1698431365
transform 1 0 83552 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_750
timestamp 1698431365
transform 1 0 85344 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_754
timestamp 1698431365
transform 1 0 85792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_756
timestamp 1698431365
transform 1 0 86016 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_767
timestamp 1698431365
transform 1 0 87248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_769
timestamp 1698431365
transform 1 0 87472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_772
timestamp 1698431365
transform 1 0 87808 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_836
timestamp 1698431365
transform 1 0 94976 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_842
timestamp 1698431365
transform 1 0 95648 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_906
timestamp 1698431365
transform 1 0 102816 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_912
timestamp 1698431365
transform 1 0 103488 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_920
timestamp 1698431365
transform 1 0 104384 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_941
timestamp 1698431365
transform 1 0 106736 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_945
timestamp 1698431365
transform 1 0 107184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_949
timestamp 1698431365
transform 1 0 107632 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_965
timestamp 1698431365
transform 1 0 109424 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_973
timestamp 1698431365
transform 1 0 110320 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_977
timestamp 1698431365
transform 1 0 110768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_979
timestamp 1698431365
transform 1 0 110992 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_982
timestamp 1698431365
transform 1 0 111328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1046
timestamp 1698431365
transform 1 0 118496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1052
timestamp 1698431365
transform 1 0 119168 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1116
timestamp 1698431365
transform 1 0 126336 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1122
timestamp 1698431365
transform 1 0 127008 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1186
timestamp 1698431365
transform 1 0 134176 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1192
timestamp 1698431365
transform 1 0 134848 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1256
timestamp 1698431365
transform 1 0 142016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1262
timestamp 1698431365
transform 1 0 142688 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1326
timestamp 1698431365
transform 1 0 149856 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1332
timestamp 1698431365
transform 1 0 150528 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1396
timestamp 1698431365
transform 1 0 157696 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_209
timestamp 1698431365
transform 1 0 24752 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_217
timestamp 1698431365
transform 1 0 25648 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_221
timestamp 1698431365
transform 1 0 26096 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_224
timestamp 1698431365
transform 1 0 26432 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_240
timestamp 1698431365
transform 1 0 28224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_259
timestamp 1698431365
transform 1 0 30352 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_261
timestamp 1698431365
transform 1 0 30576 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_274
timestamp 1698431365
transform 1 0 32032 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_290
timestamp 1698431365
transform 1 0 33824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_292
timestamp 1698431365
transform 1 0 34048 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_333
timestamp 1698431365
transform 1 0 38640 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_357
timestamp 1698431365
transform 1 0 41328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_373
timestamp 1698431365
transform 1 0 43120 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_381
timestamp 1698431365
transform 1 0 44016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_389
timestamp 1698431365
transform 1 0 44912 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_392
timestamp 1698431365
transform 1 0 45248 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_402
timestamp 1698431365
transform 1 0 46368 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_410
timestamp 1698431365
transform 1 0 47264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_452
timestamp 1698431365
transform 1 0 51968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_454
timestamp 1698431365
transform 1 0 52192 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_465
timestamp 1698431365
transform 1 0 53424 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_469
timestamp 1698431365
transform 1 0 53872 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_471
timestamp 1698431365
transform 1 0 54096 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_515
timestamp 1698431365
transform 1 0 59024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_527
timestamp 1698431365
transform 1 0 60368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_543
timestamp 1698431365
transform 1 0 62160 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_547
timestamp 1698431365
transform 1 0 62608 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_550
timestamp 1698431365
transform 1 0 62944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_554
timestamp 1698431365
transform 1 0 63392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_597
timestamp 1698431365
transform 1 0 68208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_619
timestamp 1698431365
transform 1 0 70672 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_623
timestamp 1698431365
transform 1 0 71120 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_635
timestamp 1698431365
transform 1 0 72464 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_654
timestamp 1698431365
transform 1 0 74592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_656
timestamp 1698431365
transform 1 0 74816 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_697
timestamp 1698431365
transform 1 0 79408 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_701
timestamp 1698431365
transform 1 0 79856 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_733
timestamp 1698431365
transform 1 0 83440 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_737
timestamp 1698431365
transform 1 0 83888 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_801
timestamp 1698431365
transform 1 0 91056 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_807
timestamp 1698431365
transform 1 0 91728 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_871
timestamp 1698431365
transform 1 0 98896 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_877
timestamp 1698431365
transform 1 0 99568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_909
timestamp 1698431365
transform 1 0 103152 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_925
timestamp 1698431365
transform 1 0 104944 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_929
timestamp 1698431365
transform 1 0 105392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_931
timestamp 1698431365
transform 1 0 105616 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_934
timestamp 1698431365
transform 1 0 105952 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_942
timestamp 1698431365
transform 1 0 106848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_944
timestamp 1698431365
transform 1 0 107072 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_947
timestamp 1698431365
transform 1 0 107408 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1011
timestamp 1698431365
transform 1 0 114576 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1017
timestamp 1698431365
transform 1 0 115248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1081
timestamp 1698431365
transform 1 0 122416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1087
timestamp 1698431365
transform 1 0 123088 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1151
timestamp 1698431365
transform 1 0 130256 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1157
timestamp 1698431365
transform 1 0 130928 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1221
timestamp 1698431365
transform 1 0 138096 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1227
timestamp 1698431365
transform 1 0 138768 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1291
timestamp 1698431365
transform 1 0 145936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1297
timestamp 1698431365
transform 1 0 146608 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1361
timestamp 1698431365
transform 1 0 153776 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_1367
timestamp 1698431365
transform 1 0 154448 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_1399
timestamp 1698431365
transform 1 0 158032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_1401
timestamp 1698431365
transform 1 0 158256 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_224
timestamp 1698431365
transform 1 0 26432 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_255
timestamp 1698431365
transform 1 0 29904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_259
timestamp 1698431365
transform 1 0 30352 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_266
timestamp 1698431365
transform 1 0 31136 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_274
timestamp 1698431365
transform 1 0 32032 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_278
timestamp 1698431365
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_295
timestamp 1698431365
transform 1 0 34384 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_327
timestamp 1698431365
transform 1 0 37968 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_343
timestamp 1698431365
transform 1 0 39760 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_368
timestamp 1698431365
transform 1 0 42560 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_376
timestamp 1698431365
transform 1 0 43456 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_380
timestamp 1698431365
transform 1 0 43904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_394
timestamp 1698431365
transform 1 0 45472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_398
timestamp 1698431365
transform 1 0 45920 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_414
timestamp 1698431365
transform 1 0 47712 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_418
timestamp 1698431365
transform 1 0 48160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_447
timestamp 1698431365
transform 1 0 51408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_451
timestamp 1698431365
transform 1 0 51856 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_459
timestamp 1698431365
transform 1 0 52752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_461
timestamp 1698431365
transform 1 0 52976 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_466
timestamp 1698431365
transform 1 0 53536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_468
timestamp 1698431365
transform 1 0 53760 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_475
timestamp 1698431365
transform 1 0 54544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_479
timestamp 1698431365
transform 1 0 54992 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_511
timestamp 1698431365
transform 1 0 58576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_515
timestamp 1698431365
transform 1 0 59024 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_525
timestamp 1698431365
transform 1 0 60144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_527
timestamp 1698431365
transform 1 0 60368 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_548
timestamp 1698431365
transform 1 0 62720 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_552
timestamp 1698431365
transform 1 0 63168 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_581
timestamp 1698431365
transform 1 0 66416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_583
timestamp 1698431365
transform 1 0 66640 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_617
timestamp 1698431365
transform 1 0 70448 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_628
timestamp 1698431365
transform 1 0 71680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_653
timestamp 1698431365
transform 1 0 74480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_657
timestamp 1698431365
transform 1 0 74928 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_673
timestamp 1698431365
transform 1 0 76720 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_677
timestamp 1698431365
transform 1 0 77168 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_688
timestamp 1698431365
transform 1 0 78400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_692
timestamp 1698431365
transform 1 0 78848 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_702
timestamp 1698431365
transform 1 0 79968 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_766
timestamp 1698431365
transform 1 0 87136 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_772
timestamp 1698431365
transform 1 0 87808 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_836
timestamp 1698431365
transform 1 0 94976 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_842
timestamp 1698431365
transform 1 0 95648 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_906
timestamp 1698431365
transform 1 0 102816 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_912
timestamp 1698431365
transform 1 0 103488 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_976
timestamp 1698431365
transform 1 0 110656 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_982
timestamp 1698431365
transform 1 0 111328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1046
timestamp 1698431365
transform 1 0 118496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1052
timestamp 1698431365
transform 1 0 119168 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1116
timestamp 1698431365
transform 1 0 126336 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1122
timestamp 1698431365
transform 1 0 127008 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1186
timestamp 1698431365
transform 1 0 134176 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1192
timestamp 1698431365
transform 1 0 134848 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1256
timestamp 1698431365
transform 1 0 142016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1262
timestamp 1698431365
transform 1 0 142688 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1326
timestamp 1698431365
transform 1 0 149856 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1332
timestamp 1698431365
transform 1 0 150528 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1396
timestamp 1698431365
transform 1 0 157696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_251
timestamp 1698431365
transform 1 0 29456 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_281
timestamp 1698431365
transform 1 0 32816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_285
timestamp 1698431365
transform 1 0 33264 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_301
timestamp 1698431365
transform 1 0 35056 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_309
timestamp 1698431365
transform 1 0 35952 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_313
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_381
timestamp 1698431365
transform 1 0 44016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_393
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_409
timestamp 1698431365
transform 1 0 47152 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_417
timestamp 1698431365
transform 1 0 48048 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_421
timestamp 1698431365
transform 1 0 48496 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_441
timestamp 1698431365
transform 1 0 50736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_445
timestamp 1698431365
transform 1 0 51184 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_453
timestamp 1698431365
transform 1 0 52080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_459
timestamp 1698431365
transform 1 0 52752 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_507
timestamp 1698431365
transform 1 0 58128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_523
timestamp 1698431365
transform 1 0 59920 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_527
timestamp 1698431365
transform 1 0 60368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_531
timestamp 1698431365
transform 1 0 60816 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_579
timestamp 1698431365
transform 1 0 66192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_583
timestamp 1698431365
transform 1 0 66640 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_591
timestamp 1698431365
transform 1 0 67536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_597
timestamp 1698431365
transform 1 0 68208 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_601
timestamp 1698431365
transform 1 0 68656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_609
timestamp 1698431365
transform 1 0 69552 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_619
timestamp 1698431365
transform 1 0 70672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_623
timestamp 1698431365
transform 1 0 71120 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_631
timestamp 1698431365
transform 1 0 72016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_641
timestamp 1698431365
transform 1 0 73136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_645
timestamp 1698431365
transform 1 0 73584 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_661
timestamp 1698431365
transform 1 0 75376 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_667
timestamp 1698431365
transform 1 0 76048 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_731
timestamp 1698431365
transform 1 0 83216 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_737
timestamp 1698431365
transform 1 0 83888 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_801
timestamp 1698431365
transform 1 0 91056 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_807
timestamp 1698431365
transform 1 0 91728 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_871
timestamp 1698431365
transform 1 0 98896 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_877
timestamp 1698431365
transform 1 0 99568 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_941
timestamp 1698431365
transform 1 0 106736 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_947
timestamp 1698431365
transform 1 0 107408 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1011
timestamp 1698431365
transform 1 0 114576 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1017
timestamp 1698431365
transform 1 0 115248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1081
timestamp 1698431365
transform 1 0 122416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1087
timestamp 1698431365
transform 1 0 123088 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1151
timestamp 1698431365
transform 1 0 130256 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1157
timestamp 1698431365
transform 1 0 130928 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1221
timestamp 1698431365
transform 1 0 138096 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1227
timestamp 1698431365
transform 1 0 138768 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1291
timestamp 1698431365
transform 1 0 145936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1297
timestamp 1698431365
transform 1 0 146608 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1361
timestamp 1698431365
transform 1 0 153776 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_1367
timestamp 1698431365
transform 1 0 154448 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_1399
timestamp 1698431365
transform 1 0 158032 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_1401
timestamp 1698431365
transform 1 0 158256 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_368
timestamp 1698431365
transform 1 0 42560 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_372
timestamp 1698431365
transform 1 0 43008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_374
timestamp 1698431365
transform 1 0 43232 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_408
timestamp 1698431365
transform 1 0 47040 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_412
timestamp 1698431365
transform 1 0 47488 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_428
timestamp 1698431365
transform 1 0 49280 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_436
timestamp 1698431365
transform 1 0 50176 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_440
timestamp 1698431365
transform 1 0 50624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_471
timestamp 1698431365
transform 1 0 54096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_477
timestamp 1698431365
transform 1 0 54768 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_500
timestamp 1698431365
transform 1 0 57344 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_516
timestamp 1698431365
transform 1 0 59136 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_522
timestamp 1698431365
transform 1 0 59808 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_554
timestamp 1698431365
transform 1 0 63392 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_558
timestamp 1698431365
transform 1 0 63840 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_562
timestamp 1698431365
transform 1 0 64288 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_572
timestamp 1698431365
transform 1 0 65408 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_604
timestamp 1698431365
transform 1 0 68992 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_620
timestamp 1698431365
transform 1 0 70784 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_628
timestamp 1698431365
transform 1 0 71680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_632
timestamp 1698431365
transform 1 0 72128 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_696
timestamp 1698431365
transform 1 0 79296 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_702
timestamp 1698431365
transform 1 0 79968 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_766
timestamp 1698431365
transform 1 0 87136 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_772
timestamp 1698431365
transform 1 0 87808 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_836
timestamp 1698431365
transform 1 0 94976 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_842
timestamp 1698431365
transform 1 0 95648 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_906
timestamp 1698431365
transform 1 0 102816 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_912
timestamp 1698431365
transform 1 0 103488 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_976
timestamp 1698431365
transform 1 0 110656 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_982
timestamp 1698431365
transform 1 0 111328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1046
timestamp 1698431365
transform 1 0 118496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1052
timestamp 1698431365
transform 1 0 119168 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1116
timestamp 1698431365
transform 1 0 126336 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1122
timestamp 1698431365
transform 1 0 127008 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1186
timestamp 1698431365
transform 1 0 134176 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1192
timestamp 1698431365
transform 1 0 134848 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1256
timestamp 1698431365
transform 1 0 142016 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1262
timestamp 1698431365
transform 1 0 142688 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1326
timestamp 1698431365
transform 1 0 149856 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1332
timestamp 1698431365
transform 1 0 150528 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1396
timestamp 1698431365
transform 1 0 157696 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698431365
transform 1 0 44016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_395
timestamp 1698431365
transform 1 0 45584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_461
timestamp 1698431365
transform 1 0 52976 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_469
timestamp 1698431365
transform 1 0 53872 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_473
timestamp 1698431365
transform 1 0 54320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_475
timestamp 1698431365
transform 1 0 54544 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_492
timestamp 1698431365
transform 1 0 56448 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_524
timestamp 1698431365
transform 1 0 60032 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_535
timestamp 1698431365
transform 1 0 61264 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_567
timestamp 1698431365
transform 1 0 64848 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_583
timestamp 1698431365
transform 1 0 66640 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_591
timestamp 1698431365
transform 1 0 67536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_597
timestamp 1698431365
transform 1 0 68208 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_661
timestamp 1698431365
transform 1 0 75376 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_667
timestamp 1698431365
transform 1 0 76048 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_731
timestamp 1698431365
transform 1 0 83216 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_737
timestamp 1698431365
transform 1 0 83888 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_801
timestamp 1698431365
transform 1 0 91056 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_807
timestamp 1698431365
transform 1 0 91728 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_871
timestamp 1698431365
transform 1 0 98896 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_877
timestamp 1698431365
transform 1 0 99568 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_941
timestamp 1698431365
transform 1 0 106736 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_947
timestamp 1698431365
transform 1 0 107408 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1011
timestamp 1698431365
transform 1 0 114576 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1017
timestamp 1698431365
transform 1 0 115248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1081
timestamp 1698431365
transform 1 0 122416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1087
timestamp 1698431365
transform 1 0 123088 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1151
timestamp 1698431365
transform 1 0 130256 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1157
timestamp 1698431365
transform 1 0 130928 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1221
timestamp 1698431365
transform 1 0 138096 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1227
timestamp 1698431365
transform 1 0 138768 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1291
timestamp 1698431365
transform 1 0 145936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1297
timestamp 1698431365
transform 1 0 146608 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1361
timestamp 1698431365
transform 1 0 153776 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_1367
timestamp 1698431365
transform 1 0 154448 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_1399
timestamp 1698431365
transform 1 0 158032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_1401
timestamp 1698431365
transform 1 0 158256 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698431365
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_416
timestamp 1698431365
transform 1 0 47936 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698431365
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_556
timestamp 1698431365
transform 1 0 63616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_562
timestamp 1698431365
transform 1 0 64288 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_626
timestamp 1698431365
transform 1 0 71456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_632
timestamp 1698431365
transform 1 0 72128 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_696
timestamp 1698431365
transform 1 0 79296 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_702
timestamp 1698431365
transform 1 0 79968 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_766
timestamp 1698431365
transform 1 0 87136 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_772
timestamp 1698431365
transform 1 0 87808 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_836
timestamp 1698431365
transform 1 0 94976 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_842
timestamp 1698431365
transform 1 0 95648 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_906
timestamp 1698431365
transform 1 0 102816 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_912
timestamp 1698431365
transform 1 0 103488 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_976
timestamp 1698431365
transform 1 0 110656 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_982
timestamp 1698431365
transform 1 0 111328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1046
timestamp 1698431365
transform 1 0 118496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1052
timestamp 1698431365
transform 1 0 119168 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1116
timestamp 1698431365
transform 1 0 126336 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1122
timestamp 1698431365
transform 1 0 127008 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1186
timestamp 1698431365
transform 1 0 134176 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1192
timestamp 1698431365
transform 1 0 134848 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1256
timestamp 1698431365
transform 1 0 142016 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1262
timestamp 1698431365
transform 1 0 142688 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1326
timestamp 1698431365
transform 1 0 149856 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1332
timestamp 1698431365
transform 1 0 150528 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1396
timestamp 1698431365
transform 1 0 157696 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_381
timestamp 1698431365
transform 1 0 44016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1698431365
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_521
timestamp 1698431365
transform 1 0 59696 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_527
timestamp 1698431365
transform 1 0 60368 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_591
timestamp 1698431365
transform 1 0 67536 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_597
timestamp 1698431365
transform 1 0 68208 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_661
timestamp 1698431365
transform 1 0 75376 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_667
timestamp 1698431365
transform 1 0 76048 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_731
timestamp 1698431365
transform 1 0 83216 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_737
timestamp 1698431365
transform 1 0 83888 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_801
timestamp 1698431365
transform 1 0 91056 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_807
timestamp 1698431365
transform 1 0 91728 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_871
timestamp 1698431365
transform 1 0 98896 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_877
timestamp 1698431365
transform 1 0 99568 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_941
timestamp 1698431365
transform 1 0 106736 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_947
timestamp 1698431365
transform 1 0 107408 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1011
timestamp 1698431365
transform 1 0 114576 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1017
timestamp 1698431365
transform 1 0 115248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1081
timestamp 1698431365
transform 1 0 122416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1087
timestamp 1698431365
transform 1 0 123088 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1151
timestamp 1698431365
transform 1 0 130256 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1157
timestamp 1698431365
transform 1 0 130928 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1221
timestamp 1698431365
transform 1 0 138096 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1227
timestamp 1698431365
transform 1 0 138768 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1291
timestamp 1698431365
transform 1 0 145936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1297
timestamp 1698431365
transform 1 0 146608 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1361
timestamp 1698431365
transform 1 0 153776 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_1367
timestamp 1698431365
transform 1 0 154448 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_1399
timestamp 1698431365
transform 1 0 158032 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_1401
timestamp 1698431365
transform 1 0 158256 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_416
timestamp 1698431365
transform 1 0 47936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698431365
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_556
timestamp 1698431365
transform 1 0 63616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_562
timestamp 1698431365
transform 1 0 64288 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_626
timestamp 1698431365
transform 1 0 71456 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_632
timestamp 1698431365
transform 1 0 72128 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_696
timestamp 1698431365
transform 1 0 79296 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_702
timestamp 1698431365
transform 1 0 79968 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_766
timestamp 1698431365
transform 1 0 87136 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_772
timestamp 1698431365
transform 1 0 87808 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_836
timestamp 1698431365
transform 1 0 94976 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_842
timestamp 1698431365
transform 1 0 95648 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_906
timestamp 1698431365
transform 1 0 102816 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_912
timestamp 1698431365
transform 1 0 103488 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_976
timestamp 1698431365
transform 1 0 110656 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_982
timestamp 1698431365
transform 1 0 111328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1046
timestamp 1698431365
transform 1 0 118496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1052
timestamp 1698431365
transform 1 0 119168 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1116
timestamp 1698431365
transform 1 0 126336 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1122
timestamp 1698431365
transform 1 0 127008 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1186
timestamp 1698431365
transform 1 0 134176 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1192
timestamp 1698431365
transform 1 0 134848 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1256
timestamp 1698431365
transform 1 0 142016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1262
timestamp 1698431365
transform 1 0 142688 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1326
timestamp 1698431365
transform 1 0 149856 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1332
timestamp 1698431365
transform 1 0 150528 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1396
timestamp 1698431365
transform 1 0 157696 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_451
timestamp 1698431365
transform 1 0 51856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_521
timestamp 1698431365
transform 1 0 59696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_527
timestamp 1698431365
transform 1 0 60368 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_591
timestamp 1698431365
transform 1 0 67536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_597
timestamp 1698431365
transform 1 0 68208 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_661
timestamp 1698431365
transform 1 0 75376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_667
timestamp 1698431365
transform 1 0 76048 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_731
timestamp 1698431365
transform 1 0 83216 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_737
timestamp 1698431365
transform 1 0 83888 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_801
timestamp 1698431365
transform 1 0 91056 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_807
timestamp 1698431365
transform 1 0 91728 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_871
timestamp 1698431365
transform 1 0 98896 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_877
timestamp 1698431365
transform 1 0 99568 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_941
timestamp 1698431365
transform 1 0 106736 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_947
timestamp 1698431365
transform 1 0 107408 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1011
timestamp 1698431365
transform 1 0 114576 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1017
timestamp 1698431365
transform 1 0 115248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1081
timestamp 1698431365
transform 1 0 122416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1087
timestamp 1698431365
transform 1 0 123088 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1151
timestamp 1698431365
transform 1 0 130256 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1157
timestamp 1698431365
transform 1 0 130928 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1221
timestamp 1698431365
transform 1 0 138096 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1227
timestamp 1698431365
transform 1 0 138768 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1291
timestamp 1698431365
transform 1 0 145936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1297
timestamp 1698431365
transform 1 0 146608 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1361
timestamp 1698431365
transform 1 0 153776 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_1367
timestamp 1698431365
transform 1 0 154448 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_1399
timestamp 1698431365
transform 1 0 158032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_1401
timestamp 1698431365
transform 1 0 158256 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1698431365
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_556
timestamp 1698431365
transform 1 0 63616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_562
timestamp 1698431365
transform 1 0 64288 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_626
timestamp 1698431365
transform 1 0 71456 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_632
timestamp 1698431365
transform 1 0 72128 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_696
timestamp 1698431365
transform 1 0 79296 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_702
timestamp 1698431365
transform 1 0 79968 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_766
timestamp 1698431365
transform 1 0 87136 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_772
timestamp 1698431365
transform 1 0 87808 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_836
timestamp 1698431365
transform 1 0 94976 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_842
timestamp 1698431365
transform 1 0 95648 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_906
timestamp 1698431365
transform 1 0 102816 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_912
timestamp 1698431365
transform 1 0 103488 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_976
timestamp 1698431365
transform 1 0 110656 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_982
timestamp 1698431365
transform 1 0 111328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1046
timestamp 1698431365
transform 1 0 118496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1052
timestamp 1698431365
transform 1 0 119168 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1116
timestamp 1698431365
transform 1 0 126336 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1122
timestamp 1698431365
transform 1 0 127008 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1186
timestamp 1698431365
transform 1 0 134176 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1192
timestamp 1698431365
transform 1 0 134848 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1256
timestamp 1698431365
transform 1 0 142016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1262
timestamp 1698431365
transform 1 0 142688 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1326
timestamp 1698431365
transform 1 0 149856 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1332
timestamp 1698431365
transform 1 0 150528 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1396
timestamp 1698431365
transform 1 0 157696 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_451
timestamp 1698431365
transform 1 0 51856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_521
timestamp 1698431365
transform 1 0 59696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_527
timestamp 1698431365
transform 1 0 60368 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_591
timestamp 1698431365
transform 1 0 67536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_597
timestamp 1698431365
transform 1 0 68208 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_661
timestamp 1698431365
transform 1 0 75376 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_667
timestamp 1698431365
transform 1 0 76048 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_731
timestamp 1698431365
transform 1 0 83216 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_737
timestamp 1698431365
transform 1 0 83888 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_801
timestamp 1698431365
transform 1 0 91056 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_807
timestamp 1698431365
transform 1 0 91728 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_871
timestamp 1698431365
transform 1 0 98896 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_877
timestamp 1698431365
transform 1 0 99568 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_941
timestamp 1698431365
transform 1 0 106736 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_947
timestamp 1698431365
transform 1 0 107408 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1011
timestamp 1698431365
transform 1 0 114576 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1017
timestamp 1698431365
transform 1 0 115248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1081
timestamp 1698431365
transform 1 0 122416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1087
timestamp 1698431365
transform 1 0 123088 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1151
timestamp 1698431365
transform 1 0 130256 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1157
timestamp 1698431365
transform 1 0 130928 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1221
timestamp 1698431365
transform 1 0 138096 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1227
timestamp 1698431365
transform 1 0 138768 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1291
timestamp 1698431365
transform 1 0 145936 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1297
timestamp 1698431365
transform 1 0 146608 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1361
timestamp 1698431365
transform 1 0 153776 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_1367
timestamp 1698431365
transform 1 0 154448 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_1399
timestamp 1698431365
transform 1 0 158032 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_1401
timestamp 1698431365
transform 1 0 158256 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698431365
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698431365
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_556
timestamp 1698431365
transform 1 0 63616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_562
timestamp 1698431365
transform 1 0 64288 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_626
timestamp 1698431365
transform 1 0 71456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_632
timestamp 1698431365
transform 1 0 72128 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_696
timestamp 1698431365
transform 1 0 79296 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_702
timestamp 1698431365
transform 1 0 79968 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_766
timestamp 1698431365
transform 1 0 87136 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_772
timestamp 1698431365
transform 1 0 87808 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_836
timestamp 1698431365
transform 1 0 94976 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_842
timestamp 1698431365
transform 1 0 95648 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_906
timestamp 1698431365
transform 1 0 102816 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_912
timestamp 1698431365
transform 1 0 103488 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_976
timestamp 1698431365
transform 1 0 110656 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_982
timestamp 1698431365
transform 1 0 111328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1046
timestamp 1698431365
transform 1 0 118496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1052
timestamp 1698431365
transform 1 0 119168 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1116
timestamp 1698431365
transform 1 0 126336 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1122
timestamp 1698431365
transform 1 0 127008 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1186
timestamp 1698431365
transform 1 0 134176 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1192
timestamp 1698431365
transform 1 0 134848 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1256
timestamp 1698431365
transform 1 0 142016 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1262
timestamp 1698431365
transform 1 0 142688 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1326
timestamp 1698431365
transform 1 0 149856 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1332
timestamp 1698431365
transform 1 0 150528 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1396
timestamp 1698431365
transform 1 0 157696 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_381
timestamp 1698431365
transform 1 0 44016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_451
timestamp 1698431365
transform 1 0 51856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_521
timestamp 1698431365
transform 1 0 59696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_527
timestamp 1698431365
transform 1 0 60368 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_591
timestamp 1698431365
transform 1 0 67536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_597
timestamp 1698431365
transform 1 0 68208 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_661
timestamp 1698431365
transform 1 0 75376 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_667
timestamp 1698431365
transform 1 0 76048 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_731
timestamp 1698431365
transform 1 0 83216 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_737
timestamp 1698431365
transform 1 0 83888 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_801
timestamp 1698431365
transform 1 0 91056 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_807
timestamp 1698431365
transform 1 0 91728 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_871
timestamp 1698431365
transform 1 0 98896 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_877
timestamp 1698431365
transform 1 0 99568 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_941
timestamp 1698431365
transform 1 0 106736 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_947
timestamp 1698431365
transform 1 0 107408 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1011
timestamp 1698431365
transform 1 0 114576 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1017
timestamp 1698431365
transform 1 0 115248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1081
timestamp 1698431365
transform 1 0 122416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1087
timestamp 1698431365
transform 1 0 123088 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1151
timestamp 1698431365
transform 1 0 130256 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1157
timestamp 1698431365
transform 1 0 130928 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1221
timestamp 1698431365
transform 1 0 138096 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1227
timestamp 1698431365
transform 1 0 138768 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1291
timestamp 1698431365
transform 1 0 145936 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1297
timestamp 1698431365
transform 1 0 146608 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1361
timestamp 1698431365
transform 1 0 153776 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_1367
timestamp 1698431365
transform 1 0 154448 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_1399
timestamp 1698431365
transform 1 0 158032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_1401
timestamp 1698431365
transform 1 0 158256 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698431365
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698431365
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_556
timestamp 1698431365
transform 1 0 63616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_562
timestamp 1698431365
transform 1 0 64288 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_626
timestamp 1698431365
transform 1 0 71456 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_632
timestamp 1698431365
transform 1 0 72128 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_696
timestamp 1698431365
transform 1 0 79296 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_702
timestamp 1698431365
transform 1 0 79968 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_766
timestamp 1698431365
transform 1 0 87136 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_772
timestamp 1698431365
transform 1 0 87808 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_836
timestamp 1698431365
transform 1 0 94976 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_842
timestamp 1698431365
transform 1 0 95648 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_906
timestamp 1698431365
transform 1 0 102816 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_912
timestamp 1698431365
transform 1 0 103488 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_976
timestamp 1698431365
transform 1 0 110656 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_982
timestamp 1698431365
transform 1 0 111328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1046
timestamp 1698431365
transform 1 0 118496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1052
timestamp 1698431365
transform 1 0 119168 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1116
timestamp 1698431365
transform 1 0 126336 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1122
timestamp 1698431365
transform 1 0 127008 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1186
timestamp 1698431365
transform 1 0 134176 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1192
timestamp 1698431365
transform 1 0 134848 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1256
timestamp 1698431365
transform 1 0 142016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1262
timestamp 1698431365
transform 1 0 142688 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1326
timestamp 1698431365
transform 1 0 149856 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1332
timestamp 1698431365
transform 1 0 150528 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1396
timestamp 1698431365
transform 1 0 157696 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_381
timestamp 1698431365
transform 1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698431365
transform 1 0 51856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_521
timestamp 1698431365
transform 1 0 59696 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_527
timestamp 1698431365
transform 1 0 60368 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_591
timestamp 1698431365
transform 1 0 67536 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_597
timestamp 1698431365
transform 1 0 68208 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_661
timestamp 1698431365
transform 1 0 75376 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_667
timestamp 1698431365
transform 1 0 76048 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_731
timestamp 1698431365
transform 1 0 83216 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_737
timestamp 1698431365
transform 1 0 83888 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_801
timestamp 1698431365
transform 1 0 91056 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_807
timestamp 1698431365
transform 1 0 91728 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_871
timestamp 1698431365
transform 1 0 98896 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_877
timestamp 1698431365
transform 1 0 99568 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_941
timestamp 1698431365
transform 1 0 106736 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_947
timestamp 1698431365
transform 1 0 107408 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1011
timestamp 1698431365
transform 1 0 114576 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1017
timestamp 1698431365
transform 1 0 115248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1081
timestamp 1698431365
transform 1 0 122416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1087
timestamp 1698431365
transform 1 0 123088 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1151
timestamp 1698431365
transform 1 0 130256 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1157
timestamp 1698431365
transform 1 0 130928 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1221
timestamp 1698431365
transform 1 0 138096 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1227
timestamp 1698431365
transform 1 0 138768 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1291
timestamp 1698431365
transform 1 0 145936 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1297
timestamp 1698431365
transform 1 0 146608 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1361
timestamp 1698431365
transform 1 0 153776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_1367
timestamp 1698431365
transform 1 0 154448 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_1399
timestamp 1698431365
transform 1 0 158032 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_1401
timestamp 1698431365
transform 1 0 158256 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_416
timestamp 1698431365
transform 1 0 47936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698431365
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_556
timestamp 1698431365
transform 1 0 63616 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_562
timestamp 1698431365
transform 1 0 64288 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_626
timestamp 1698431365
transform 1 0 71456 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_632
timestamp 1698431365
transform 1 0 72128 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_696
timestamp 1698431365
transform 1 0 79296 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_702
timestamp 1698431365
transform 1 0 79968 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_766
timestamp 1698431365
transform 1 0 87136 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_772
timestamp 1698431365
transform 1 0 87808 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_836
timestamp 1698431365
transform 1 0 94976 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_842
timestamp 1698431365
transform 1 0 95648 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_906
timestamp 1698431365
transform 1 0 102816 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_912
timestamp 1698431365
transform 1 0 103488 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_976
timestamp 1698431365
transform 1 0 110656 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_982
timestamp 1698431365
transform 1 0 111328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1046
timestamp 1698431365
transform 1 0 118496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1052
timestamp 1698431365
transform 1 0 119168 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1116
timestamp 1698431365
transform 1 0 126336 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1122
timestamp 1698431365
transform 1 0 127008 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1186
timestamp 1698431365
transform 1 0 134176 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1192
timestamp 1698431365
transform 1 0 134848 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1256
timestamp 1698431365
transform 1 0 142016 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1262
timestamp 1698431365
transform 1 0 142688 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1326
timestamp 1698431365
transform 1 0 149856 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1332
timestamp 1698431365
transform 1 0 150528 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1396
timestamp 1698431365
transform 1 0 157696 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698431365
transform 1 0 44016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_451
timestamp 1698431365
transform 1 0 51856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_521
timestamp 1698431365
transform 1 0 59696 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_527
timestamp 1698431365
transform 1 0 60368 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_591
timestamp 1698431365
transform 1 0 67536 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_597
timestamp 1698431365
transform 1 0 68208 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_661
timestamp 1698431365
transform 1 0 75376 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_667
timestamp 1698431365
transform 1 0 76048 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_731
timestamp 1698431365
transform 1 0 83216 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_737
timestamp 1698431365
transform 1 0 83888 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_801
timestamp 1698431365
transform 1 0 91056 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_807
timestamp 1698431365
transform 1 0 91728 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_871
timestamp 1698431365
transform 1 0 98896 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_877
timestamp 1698431365
transform 1 0 99568 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_941
timestamp 1698431365
transform 1 0 106736 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_947
timestamp 1698431365
transform 1 0 107408 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1011
timestamp 1698431365
transform 1 0 114576 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1017
timestamp 1698431365
transform 1 0 115248 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1081
timestamp 1698431365
transform 1 0 122416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1087
timestamp 1698431365
transform 1 0 123088 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1151
timestamp 1698431365
transform 1 0 130256 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1157
timestamp 1698431365
transform 1 0 130928 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1221
timestamp 1698431365
transform 1 0 138096 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1227
timestamp 1698431365
transform 1 0 138768 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1291
timestamp 1698431365
transform 1 0 145936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1297
timestamp 1698431365
transform 1 0 146608 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1361
timestamp 1698431365
transform 1 0 153776 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_1367
timestamp 1698431365
transform 1 0 154448 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_1399
timestamp 1698431365
transform 1 0 158032 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_1401
timestamp 1698431365
transform 1 0 158256 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698431365
transform 1 0 55776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_556
timestamp 1698431365
transform 1 0 63616 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_562
timestamp 1698431365
transform 1 0 64288 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_626
timestamp 1698431365
transform 1 0 71456 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_632
timestamp 1698431365
transform 1 0 72128 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_696
timestamp 1698431365
transform 1 0 79296 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_702
timestamp 1698431365
transform 1 0 79968 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_766
timestamp 1698431365
transform 1 0 87136 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_772
timestamp 1698431365
transform 1 0 87808 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_836
timestamp 1698431365
transform 1 0 94976 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_842
timestamp 1698431365
transform 1 0 95648 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_906
timestamp 1698431365
transform 1 0 102816 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_912
timestamp 1698431365
transform 1 0 103488 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_976
timestamp 1698431365
transform 1 0 110656 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_982
timestamp 1698431365
transform 1 0 111328 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1046
timestamp 1698431365
transform 1 0 118496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1052
timestamp 1698431365
transform 1 0 119168 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1116
timestamp 1698431365
transform 1 0 126336 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1122
timestamp 1698431365
transform 1 0 127008 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1186
timestamp 1698431365
transform 1 0 134176 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1192
timestamp 1698431365
transform 1 0 134848 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1256
timestamp 1698431365
transform 1 0 142016 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1262
timestamp 1698431365
transform 1 0 142688 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1326
timestamp 1698431365
transform 1 0 149856 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1332
timestamp 1698431365
transform 1 0 150528 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1396
timestamp 1698431365
transform 1 0 157696 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698431365
transform 1 0 51856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_521
timestamp 1698431365
transform 1 0 59696 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_527
timestamp 1698431365
transform 1 0 60368 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_591
timestamp 1698431365
transform 1 0 67536 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_597
timestamp 1698431365
transform 1 0 68208 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_661
timestamp 1698431365
transform 1 0 75376 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_667
timestamp 1698431365
transform 1 0 76048 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_731
timestamp 1698431365
transform 1 0 83216 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_737
timestamp 1698431365
transform 1 0 83888 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_801
timestamp 1698431365
transform 1 0 91056 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_807
timestamp 1698431365
transform 1 0 91728 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_871
timestamp 1698431365
transform 1 0 98896 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_877
timestamp 1698431365
transform 1 0 99568 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_941
timestamp 1698431365
transform 1 0 106736 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_947
timestamp 1698431365
transform 1 0 107408 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1011
timestamp 1698431365
transform 1 0 114576 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1017
timestamp 1698431365
transform 1 0 115248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1081
timestamp 1698431365
transform 1 0 122416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1087
timestamp 1698431365
transform 1 0 123088 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1151
timestamp 1698431365
transform 1 0 130256 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1157
timestamp 1698431365
transform 1 0 130928 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1221
timestamp 1698431365
transform 1 0 138096 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1227
timestamp 1698431365
transform 1 0 138768 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1291
timestamp 1698431365
transform 1 0 145936 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1297
timestamp 1698431365
transform 1 0 146608 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1361
timestamp 1698431365
transform 1 0 153776 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_1367
timestamp 1698431365
transform 1 0 154448 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_1399
timestamp 1698431365
transform 1 0 158032 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_1401
timestamp 1698431365
transform 1 0 158256 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_346
timestamp 1698431365
transform 1 0 40096 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_416
timestamp 1698431365
transform 1 0 47936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_486
timestamp 1698431365
transform 1 0 55776 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_556
timestamp 1698431365
transform 1 0 63616 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_562
timestamp 1698431365
transform 1 0 64288 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_626
timestamp 1698431365
transform 1 0 71456 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_632
timestamp 1698431365
transform 1 0 72128 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_696
timestamp 1698431365
transform 1 0 79296 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_702
timestamp 1698431365
transform 1 0 79968 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_766
timestamp 1698431365
transform 1 0 87136 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_772
timestamp 1698431365
transform 1 0 87808 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_836
timestamp 1698431365
transform 1 0 94976 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_842
timestamp 1698431365
transform 1 0 95648 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_906
timestamp 1698431365
transform 1 0 102816 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_912
timestamp 1698431365
transform 1 0 103488 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_976
timestamp 1698431365
transform 1 0 110656 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_982
timestamp 1698431365
transform 1 0 111328 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1046
timestamp 1698431365
transform 1 0 118496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1052
timestamp 1698431365
transform 1 0 119168 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1116
timestamp 1698431365
transform 1 0 126336 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1122
timestamp 1698431365
transform 1 0 127008 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1186
timestamp 1698431365
transform 1 0 134176 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1192
timestamp 1698431365
transform 1 0 134848 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1256
timestamp 1698431365
transform 1 0 142016 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1262
timestamp 1698431365
transform 1 0 142688 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1326
timestamp 1698431365
transform 1 0 149856 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1332
timestamp 1698431365
transform 1 0 150528 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1396
timestamp 1698431365
transform 1 0 157696 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698431365
transform 1 0 20496 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698431365
transform 1 0 51856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_521
timestamp 1698431365
transform 1 0 59696 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_527
timestamp 1698431365
transform 1 0 60368 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_591
timestamp 1698431365
transform 1 0 67536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_597
timestamp 1698431365
transform 1 0 68208 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_661
timestamp 1698431365
transform 1 0 75376 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_667
timestamp 1698431365
transform 1 0 76048 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_731
timestamp 1698431365
transform 1 0 83216 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_737
timestamp 1698431365
transform 1 0 83888 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_801
timestamp 1698431365
transform 1 0 91056 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_807
timestamp 1698431365
transform 1 0 91728 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_871
timestamp 1698431365
transform 1 0 98896 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_877
timestamp 1698431365
transform 1 0 99568 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_941
timestamp 1698431365
transform 1 0 106736 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_947
timestamp 1698431365
transform 1 0 107408 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1011
timestamp 1698431365
transform 1 0 114576 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1017
timestamp 1698431365
transform 1 0 115248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1081
timestamp 1698431365
transform 1 0 122416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1087
timestamp 1698431365
transform 1 0 123088 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1151
timestamp 1698431365
transform 1 0 130256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1157
timestamp 1698431365
transform 1 0 130928 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1221
timestamp 1698431365
transform 1 0 138096 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1227
timestamp 1698431365
transform 1 0 138768 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1291
timestamp 1698431365
transform 1 0 145936 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1297
timestamp 1698431365
transform 1 0 146608 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1361
timestamp 1698431365
transform 1 0 153776 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_1367
timestamp 1698431365
transform 1 0 154448 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_1399
timestamp 1698431365
transform 1 0 158032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_1401
timestamp 1698431365
transform 1 0 158256 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_276
timestamp 1698431365
transform 1 0 32256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_346
timestamp 1698431365
transform 1 0 40096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_416
timestamp 1698431365
transform 1 0 47936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_486
timestamp 1698431365
transform 1 0 55776 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_556
timestamp 1698431365
transform 1 0 63616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_562
timestamp 1698431365
transform 1 0 64288 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_626
timestamp 1698431365
transform 1 0 71456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_632
timestamp 1698431365
transform 1 0 72128 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_696
timestamp 1698431365
transform 1 0 79296 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_702
timestamp 1698431365
transform 1 0 79968 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_766
timestamp 1698431365
transform 1 0 87136 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_772
timestamp 1698431365
transform 1 0 87808 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_836
timestamp 1698431365
transform 1 0 94976 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_842
timestamp 1698431365
transform 1 0 95648 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_906
timestamp 1698431365
transform 1 0 102816 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_912
timestamp 1698431365
transform 1 0 103488 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_976
timestamp 1698431365
transform 1 0 110656 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_982
timestamp 1698431365
transform 1 0 111328 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1046
timestamp 1698431365
transform 1 0 118496 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1052
timestamp 1698431365
transform 1 0 119168 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1116
timestamp 1698431365
transform 1 0 126336 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1122
timestamp 1698431365
transform 1 0 127008 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1186
timestamp 1698431365
transform 1 0 134176 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1192
timestamp 1698431365
transform 1 0 134848 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1256
timestamp 1698431365
transform 1 0 142016 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1262
timestamp 1698431365
transform 1 0 142688 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1326
timestamp 1698431365
transform 1 0 149856 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1332
timestamp 1698431365
transform 1 0 150528 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1396
timestamp 1698431365
transform 1 0 157696 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_311
timestamp 1698431365
transform 1 0 36176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_381
timestamp 1698431365
transform 1 0 44016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_451
timestamp 1698431365
transform 1 0 51856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_521
timestamp 1698431365
transform 1 0 59696 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_527
timestamp 1698431365
transform 1 0 60368 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_591
timestamp 1698431365
transform 1 0 67536 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_597
timestamp 1698431365
transform 1 0 68208 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_661
timestamp 1698431365
transform 1 0 75376 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_667
timestamp 1698431365
transform 1 0 76048 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_731
timestamp 1698431365
transform 1 0 83216 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_737
timestamp 1698431365
transform 1 0 83888 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_801
timestamp 1698431365
transform 1 0 91056 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_807
timestamp 1698431365
transform 1 0 91728 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_871
timestamp 1698431365
transform 1 0 98896 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_877
timestamp 1698431365
transform 1 0 99568 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_941
timestamp 1698431365
transform 1 0 106736 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_947
timestamp 1698431365
transform 1 0 107408 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1011
timestamp 1698431365
transform 1 0 114576 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1017
timestamp 1698431365
transform 1 0 115248 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1081
timestamp 1698431365
transform 1 0 122416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1087
timestamp 1698431365
transform 1 0 123088 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1151
timestamp 1698431365
transform 1 0 130256 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1157
timestamp 1698431365
transform 1 0 130928 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1221
timestamp 1698431365
transform 1 0 138096 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1227
timestamp 1698431365
transform 1 0 138768 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1291
timestamp 1698431365
transform 1 0 145936 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1297
timestamp 1698431365
transform 1 0 146608 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1361
timestamp 1698431365
transform 1 0 153776 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_1367
timestamp 1698431365
transform 1 0 154448 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_1399
timestamp 1698431365
transform 1 0 158032 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_1401
timestamp 1698431365
transform 1 0 158256 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_276
timestamp 1698431365
transform 1 0 32256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_346
timestamp 1698431365
transform 1 0 40096 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_416
timestamp 1698431365
transform 1 0 47936 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_486
timestamp 1698431365
transform 1 0 55776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_556
timestamp 1698431365
transform 1 0 63616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_562
timestamp 1698431365
transform 1 0 64288 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_626
timestamp 1698431365
transform 1 0 71456 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_632
timestamp 1698431365
transform 1 0 72128 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_696
timestamp 1698431365
transform 1 0 79296 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_702
timestamp 1698431365
transform 1 0 79968 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_766
timestamp 1698431365
transform 1 0 87136 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_772
timestamp 1698431365
transform 1 0 87808 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_836
timestamp 1698431365
transform 1 0 94976 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_842
timestamp 1698431365
transform 1 0 95648 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_906
timestamp 1698431365
transform 1 0 102816 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_912
timestamp 1698431365
transform 1 0 103488 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_976
timestamp 1698431365
transform 1 0 110656 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_982
timestamp 1698431365
transform 1 0 111328 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1046
timestamp 1698431365
transform 1 0 118496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1052
timestamp 1698431365
transform 1 0 119168 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1116
timestamp 1698431365
transform 1 0 126336 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1122
timestamp 1698431365
transform 1 0 127008 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1186
timestamp 1698431365
transform 1 0 134176 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1192
timestamp 1698431365
transform 1 0 134848 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1256
timestamp 1698431365
transform 1 0 142016 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1262
timestamp 1698431365
transform 1 0 142688 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1326
timestamp 1698431365
transform 1 0 149856 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1332
timestamp 1698431365
transform 1 0 150528 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1396
timestamp 1698431365
transform 1 0 157696 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_101
timestamp 1698431365
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_241
timestamp 1698431365
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_311
timestamp 1698431365
transform 1 0 36176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_381
timestamp 1698431365
transform 1 0 44016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698431365
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_521
timestamp 1698431365
transform 1 0 59696 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_527
timestamp 1698431365
transform 1 0 60368 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_591
timestamp 1698431365
transform 1 0 67536 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_597
timestamp 1698431365
transform 1 0 68208 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_661
timestamp 1698431365
transform 1 0 75376 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_667
timestamp 1698431365
transform 1 0 76048 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_731
timestamp 1698431365
transform 1 0 83216 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_737
timestamp 1698431365
transform 1 0 83888 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_801
timestamp 1698431365
transform 1 0 91056 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_807
timestamp 1698431365
transform 1 0 91728 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_871
timestamp 1698431365
transform 1 0 98896 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_877
timestamp 1698431365
transform 1 0 99568 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_941
timestamp 1698431365
transform 1 0 106736 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_947
timestamp 1698431365
transform 1 0 107408 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1011
timestamp 1698431365
transform 1 0 114576 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1017
timestamp 1698431365
transform 1 0 115248 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1081
timestamp 1698431365
transform 1 0 122416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1087
timestamp 1698431365
transform 1 0 123088 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1151
timestamp 1698431365
transform 1 0 130256 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1157
timestamp 1698431365
transform 1 0 130928 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1221
timestamp 1698431365
transform 1 0 138096 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1227
timestamp 1698431365
transform 1 0 138768 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1291
timestamp 1698431365
transform 1 0 145936 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1297
timestamp 1698431365
transform 1 0 146608 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1361
timestamp 1698431365
transform 1 0 153776 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_1367
timestamp 1698431365
transform 1 0 154448 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1399
timestamp 1698431365
transform 1 0 158032 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1401
timestamp 1698431365
transform 1 0 158256 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_66
timestamp 1698431365
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_136
timestamp 1698431365
transform 1 0 16576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_206
timestamp 1698431365
transform 1 0 24416 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_276
timestamp 1698431365
transform 1 0 32256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_346
timestamp 1698431365
transform 1 0 40096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_416
timestamp 1698431365
transform 1 0 47936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_422
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_486
timestamp 1698431365
transform 1 0 55776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_556
timestamp 1698431365
transform 1 0 63616 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_562
timestamp 1698431365
transform 1 0 64288 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_626
timestamp 1698431365
transform 1 0 71456 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_632
timestamp 1698431365
transform 1 0 72128 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_696
timestamp 1698431365
transform 1 0 79296 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_702
timestamp 1698431365
transform 1 0 79968 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_766
timestamp 1698431365
transform 1 0 87136 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_772
timestamp 1698431365
transform 1 0 87808 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_836
timestamp 1698431365
transform 1 0 94976 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_842
timestamp 1698431365
transform 1 0 95648 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_906
timestamp 1698431365
transform 1 0 102816 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_912
timestamp 1698431365
transform 1 0 103488 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_976
timestamp 1698431365
transform 1 0 110656 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_982
timestamp 1698431365
transform 1 0 111328 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1046
timestamp 1698431365
transform 1 0 118496 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1052
timestamp 1698431365
transform 1 0 119168 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1116
timestamp 1698431365
transform 1 0 126336 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1122
timestamp 1698431365
transform 1 0 127008 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1186
timestamp 1698431365
transform 1 0 134176 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1192
timestamp 1698431365
transform 1 0 134848 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1256
timestamp 1698431365
transform 1 0 142016 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1262
timestamp 1698431365
transform 1 0 142688 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1326
timestamp 1698431365
transform 1 0 149856 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1332
timestamp 1698431365
transform 1 0 150528 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1396
timestamp 1698431365
transform 1 0 157696 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_101
timestamp 1698431365
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_241
timestamp 1698431365
transform 1 0 28336 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_311
timestamp 1698431365
transform 1 0 36176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_381
timestamp 1698431365
transform 1 0 44016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_451
timestamp 1698431365
transform 1 0 51856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_521
timestamp 1698431365
transform 1 0 59696 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_527
timestamp 1698431365
transform 1 0 60368 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_591
timestamp 1698431365
transform 1 0 67536 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_597
timestamp 1698431365
transform 1 0 68208 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_661
timestamp 1698431365
transform 1 0 75376 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_667
timestamp 1698431365
transform 1 0 76048 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_731
timestamp 1698431365
transform 1 0 83216 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_737
timestamp 1698431365
transform 1 0 83888 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_801
timestamp 1698431365
transform 1 0 91056 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_807
timestamp 1698431365
transform 1 0 91728 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_871
timestamp 1698431365
transform 1 0 98896 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_877
timestamp 1698431365
transform 1 0 99568 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_941
timestamp 1698431365
transform 1 0 106736 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_947
timestamp 1698431365
transform 1 0 107408 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1011
timestamp 1698431365
transform 1 0 114576 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1017
timestamp 1698431365
transform 1 0 115248 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1081
timestamp 1698431365
transform 1 0 122416 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1087
timestamp 1698431365
transform 1 0 123088 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1151
timestamp 1698431365
transform 1 0 130256 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1157
timestamp 1698431365
transform 1 0 130928 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1221
timestamp 1698431365
transform 1 0 138096 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1227
timestamp 1698431365
transform 1 0 138768 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1291
timestamp 1698431365
transform 1 0 145936 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1297
timestamp 1698431365
transform 1 0 146608 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1361
timestamp 1698431365
transform 1 0 153776 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_1367
timestamp 1698431365
transform 1 0 154448 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_1399
timestamp 1698431365
transform 1 0 158032 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_1401
timestamp 1698431365
transform 1 0 158256 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_66
timestamp 1698431365
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698431365
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_206
timestamp 1698431365
transform 1 0 24416 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_276
timestamp 1698431365
transform 1 0 32256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_346
timestamp 1698431365
transform 1 0 40096 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_416
timestamp 1698431365
transform 1 0 47936 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_486
timestamp 1698431365
transform 1 0 55776 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_556
timestamp 1698431365
transform 1 0 63616 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_562
timestamp 1698431365
transform 1 0 64288 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_626
timestamp 1698431365
transform 1 0 71456 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_632
timestamp 1698431365
transform 1 0 72128 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_696
timestamp 1698431365
transform 1 0 79296 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_702
timestamp 1698431365
transform 1 0 79968 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_766
timestamp 1698431365
transform 1 0 87136 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_772
timestamp 1698431365
transform 1 0 87808 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_836
timestamp 1698431365
transform 1 0 94976 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_842
timestamp 1698431365
transform 1 0 95648 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_906
timestamp 1698431365
transform 1 0 102816 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_912
timestamp 1698431365
transform 1 0 103488 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_976
timestamp 1698431365
transform 1 0 110656 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_982
timestamp 1698431365
transform 1 0 111328 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1046
timestamp 1698431365
transform 1 0 118496 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1052
timestamp 1698431365
transform 1 0 119168 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1116
timestamp 1698431365
transform 1 0 126336 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1122
timestamp 1698431365
transform 1 0 127008 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1186
timestamp 1698431365
transform 1 0 134176 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1192
timestamp 1698431365
transform 1 0 134848 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1256
timestamp 1698431365
transform 1 0 142016 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1262
timestamp 1698431365
transform 1 0 142688 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1326
timestamp 1698431365
transform 1 0 149856 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1332
timestamp 1698431365
transform 1 0 150528 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1396
timestamp 1698431365
transform 1 0 157696 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_171
timestamp 1698431365
transform 1 0 20496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_241
timestamp 1698431365
transform 1 0 28336 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_311
timestamp 1698431365
transform 1 0 36176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_381
timestamp 1698431365
transform 1 0 44016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_451
timestamp 1698431365
transform 1 0 51856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_521
timestamp 1698431365
transform 1 0 59696 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_527
timestamp 1698431365
transform 1 0 60368 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_591
timestamp 1698431365
transform 1 0 67536 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_597
timestamp 1698431365
transform 1 0 68208 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_661
timestamp 1698431365
transform 1 0 75376 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_667
timestamp 1698431365
transform 1 0 76048 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_731
timestamp 1698431365
transform 1 0 83216 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_737
timestamp 1698431365
transform 1 0 83888 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_801
timestamp 1698431365
transform 1 0 91056 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_807
timestamp 1698431365
transform 1 0 91728 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_871
timestamp 1698431365
transform 1 0 98896 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_877
timestamp 1698431365
transform 1 0 99568 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_941
timestamp 1698431365
transform 1 0 106736 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_947
timestamp 1698431365
transform 1 0 107408 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1011
timestamp 1698431365
transform 1 0 114576 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1017
timestamp 1698431365
transform 1 0 115248 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1081
timestamp 1698431365
transform 1 0 122416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1087
timestamp 1698431365
transform 1 0 123088 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1151
timestamp 1698431365
transform 1 0 130256 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1157
timestamp 1698431365
transform 1 0 130928 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1221
timestamp 1698431365
transform 1 0 138096 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1227
timestamp 1698431365
transform 1 0 138768 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1291
timestamp 1698431365
transform 1 0 145936 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1297
timestamp 1698431365
transform 1 0 146608 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1361
timestamp 1698431365
transform 1 0 153776 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_1367
timestamp 1698431365
transform 1 0 154448 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_1399
timestamp 1698431365
transform 1 0 158032 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_1401
timestamp 1698431365
transform 1 0 158256 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1698431365
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_276
timestamp 1698431365
transform 1 0 32256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_346
timestamp 1698431365
transform 1 0 40096 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_416
timestamp 1698431365
transform 1 0 47936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_422
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_486
timestamp 1698431365
transform 1 0 55776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_556
timestamp 1698431365
transform 1 0 63616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_562
timestamp 1698431365
transform 1 0 64288 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_626
timestamp 1698431365
transform 1 0 71456 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_632
timestamp 1698431365
transform 1 0 72128 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_696
timestamp 1698431365
transform 1 0 79296 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_702
timestamp 1698431365
transform 1 0 79968 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_766
timestamp 1698431365
transform 1 0 87136 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_772
timestamp 1698431365
transform 1 0 87808 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_836
timestamp 1698431365
transform 1 0 94976 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_842
timestamp 1698431365
transform 1 0 95648 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_906
timestamp 1698431365
transform 1 0 102816 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_912
timestamp 1698431365
transform 1 0 103488 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_976
timestamp 1698431365
transform 1 0 110656 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_982
timestamp 1698431365
transform 1 0 111328 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1046
timestamp 1698431365
transform 1 0 118496 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1052
timestamp 1698431365
transform 1 0 119168 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1116
timestamp 1698431365
transform 1 0 126336 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1122
timestamp 1698431365
transform 1 0 127008 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1186
timestamp 1698431365
transform 1 0 134176 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1192
timestamp 1698431365
transform 1 0 134848 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1256
timestamp 1698431365
transform 1 0 142016 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1262
timestamp 1698431365
transform 1 0 142688 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1326
timestamp 1698431365
transform 1 0 149856 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1332
timestamp 1698431365
transform 1 0 150528 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1396
timestamp 1698431365
transform 1 0 157696 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_171
timestamp 1698431365
transform 1 0 20496 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_241
timestamp 1698431365
transform 1 0 28336 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_311
timestamp 1698431365
transform 1 0 36176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_381
timestamp 1698431365
transform 1 0 44016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_451
timestamp 1698431365
transform 1 0 51856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_521
timestamp 1698431365
transform 1 0 59696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_527
timestamp 1698431365
transform 1 0 60368 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_591
timestamp 1698431365
transform 1 0 67536 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_597
timestamp 1698431365
transform 1 0 68208 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_661
timestamp 1698431365
transform 1 0 75376 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_667
timestamp 1698431365
transform 1 0 76048 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_731
timestamp 1698431365
transform 1 0 83216 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_737
timestamp 1698431365
transform 1 0 83888 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_801
timestamp 1698431365
transform 1 0 91056 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_807
timestamp 1698431365
transform 1 0 91728 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_871
timestamp 1698431365
transform 1 0 98896 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_877
timestamp 1698431365
transform 1 0 99568 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_941
timestamp 1698431365
transform 1 0 106736 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_947
timestamp 1698431365
transform 1 0 107408 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1011
timestamp 1698431365
transform 1 0 114576 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1017
timestamp 1698431365
transform 1 0 115248 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1081
timestamp 1698431365
transform 1 0 122416 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1087
timestamp 1698431365
transform 1 0 123088 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1151
timestamp 1698431365
transform 1 0 130256 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1157
timestamp 1698431365
transform 1 0 130928 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1221
timestamp 1698431365
transform 1 0 138096 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1227
timestamp 1698431365
transform 1 0 138768 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1291
timestamp 1698431365
transform 1 0 145936 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1297
timestamp 1698431365
transform 1 0 146608 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1361
timestamp 1698431365
transform 1 0 153776 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_1367
timestamp 1698431365
transform 1 0 154448 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_1399
timestamp 1698431365
transform 1 0 158032 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_1401
timestamp 1698431365
transform 1 0 158256 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1698431365
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_136
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698431365
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_276
timestamp 1698431365
transform 1 0 32256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_346
timestamp 1698431365
transform 1 0 40096 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_416
timestamp 1698431365
transform 1 0 47936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_422
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_486
timestamp 1698431365
transform 1 0 55776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_556
timestamp 1698431365
transform 1 0 63616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_562
timestamp 1698431365
transform 1 0 64288 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_626
timestamp 1698431365
transform 1 0 71456 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_632
timestamp 1698431365
transform 1 0 72128 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_696
timestamp 1698431365
transform 1 0 79296 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_702
timestamp 1698431365
transform 1 0 79968 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_766
timestamp 1698431365
transform 1 0 87136 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_772
timestamp 1698431365
transform 1 0 87808 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_836
timestamp 1698431365
transform 1 0 94976 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_842
timestamp 1698431365
transform 1 0 95648 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_906
timestamp 1698431365
transform 1 0 102816 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_912
timestamp 1698431365
transform 1 0 103488 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_976
timestamp 1698431365
transform 1 0 110656 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_982
timestamp 1698431365
transform 1 0 111328 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1046
timestamp 1698431365
transform 1 0 118496 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1052
timestamp 1698431365
transform 1 0 119168 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1116
timestamp 1698431365
transform 1 0 126336 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1122
timestamp 1698431365
transform 1 0 127008 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1186
timestamp 1698431365
transform 1 0 134176 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1192
timestamp 1698431365
transform 1 0 134848 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1256
timestamp 1698431365
transform 1 0 142016 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1262
timestamp 1698431365
transform 1 0 142688 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1326
timestamp 1698431365
transform 1 0 149856 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1332
timestamp 1698431365
transform 1 0 150528 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1396
timestamp 1698431365
transform 1 0 157696 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_171
timestamp 1698431365
transform 1 0 20496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_241
timestamp 1698431365
transform 1 0 28336 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_311
timestamp 1698431365
transform 1 0 36176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_381
timestamp 1698431365
transform 1 0 44016 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_451
timestamp 1698431365
transform 1 0 51856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_521
timestamp 1698431365
transform 1 0 59696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_527
timestamp 1698431365
transform 1 0 60368 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_591
timestamp 1698431365
transform 1 0 67536 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_597
timestamp 1698431365
transform 1 0 68208 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_661
timestamp 1698431365
transform 1 0 75376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_667
timestamp 1698431365
transform 1 0 76048 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_731
timestamp 1698431365
transform 1 0 83216 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_737
timestamp 1698431365
transform 1 0 83888 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_801
timestamp 1698431365
transform 1 0 91056 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_807
timestamp 1698431365
transform 1 0 91728 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_871
timestamp 1698431365
transform 1 0 98896 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_877
timestamp 1698431365
transform 1 0 99568 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_941
timestamp 1698431365
transform 1 0 106736 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_947
timestamp 1698431365
transform 1 0 107408 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1011
timestamp 1698431365
transform 1 0 114576 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1017
timestamp 1698431365
transform 1 0 115248 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1081
timestamp 1698431365
transform 1 0 122416 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1087
timestamp 1698431365
transform 1 0 123088 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1151
timestamp 1698431365
transform 1 0 130256 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1157
timestamp 1698431365
transform 1 0 130928 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1221
timestamp 1698431365
transform 1 0 138096 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1227
timestamp 1698431365
transform 1 0 138768 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1291
timestamp 1698431365
transform 1 0 145936 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1297
timestamp 1698431365
transform 1 0 146608 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1361
timestamp 1698431365
transform 1 0 153776 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_1367
timestamp 1698431365
transform 1 0 154448 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_1399
timestamp 1698431365
transform 1 0 158032 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_1401
timestamp 1698431365
transform 1 0 158256 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_136
timestamp 1698431365
transform 1 0 16576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_276
timestamp 1698431365
transform 1 0 32256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_346
timestamp 1698431365
transform 1 0 40096 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_416
timestamp 1698431365
transform 1 0 47936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_486
timestamp 1698431365
transform 1 0 55776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_556
timestamp 1698431365
transform 1 0 63616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_562
timestamp 1698431365
transform 1 0 64288 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_626
timestamp 1698431365
transform 1 0 71456 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_632
timestamp 1698431365
transform 1 0 72128 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_696
timestamp 1698431365
transform 1 0 79296 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_702
timestamp 1698431365
transform 1 0 79968 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_766
timestamp 1698431365
transform 1 0 87136 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_772
timestamp 1698431365
transform 1 0 87808 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_836
timestamp 1698431365
transform 1 0 94976 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_842
timestamp 1698431365
transform 1 0 95648 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_906
timestamp 1698431365
transform 1 0 102816 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_912
timestamp 1698431365
transform 1 0 103488 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_976
timestamp 1698431365
transform 1 0 110656 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_982
timestamp 1698431365
transform 1 0 111328 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1046
timestamp 1698431365
transform 1 0 118496 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1052
timestamp 1698431365
transform 1 0 119168 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1116
timestamp 1698431365
transform 1 0 126336 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1122
timestamp 1698431365
transform 1 0 127008 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1186
timestamp 1698431365
transform 1 0 134176 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1192
timestamp 1698431365
transform 1 0 134848 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1256
timestamp 1698431365
transform 1 0 142016 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1262
timestamp 1698431365
transform 1 0 142688 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1326
timestamp 1698431365
transform 1 0 149856 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1332
timestamp 1698431365
transform 1 0 150528 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1396
timestamp 1698431365
transform 1 0 157696 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_171
timestamp 1698431365
transform 1 0 20496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_241
timestamp 1698431365
transform 1 0 28336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698431365
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_381
timestamp 1698431365
transform 1 0 44016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698431365
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_521
timestamp 1698431365
transform 1 0 59696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_527
timestamp 1698431365
transform 1 0 60368 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_591
timestamp 1698431365
transform 1 0 67536 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_597
timestamp 1698431365
transform 1 0 68208 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_661
timestamp 1698431365
transform 1 0 75376 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_667
timestamp 1698431365
transform 1 0 76048 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_731
timestamp 1698431365
transform 1 0 83216 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_737
timestamp 1698431365
transform 1 0 83888 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_801
timestamp 1698431365
transform 1 0 91056 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_807
timestamp 1698431365
transform 1 0 91728 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_871
timestamp 1698431365
transform 1 0 98896 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_877
timestamp 1698431365
transform 1 0 99568 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_941
timestamp 1698431365
transform 1 0 106736 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_947
timestamp 1698431365
transform 1 0 107408 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1011
timestamp 1698431365
transform 1 0 114576 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1017
timestamp 1698431365
transform 1 0 115248 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1081
timestamp 1698431365
transform 1 0 122416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1087
timestamp 1698431365
transform 1 0 123088 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1151
timestamp 1698431365
transform 1 0 130256 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1157
timestamp 1698431365
transform 1 0 130928 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1221
timestamp 1698431365
transform 1 0 138096 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1227
timestamp 1698431365
transform 1 0 138768 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1291
timestamp 1698431365
transform 1 0 145936 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1297
timestamp 1698431365
transform 1 0 146608 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1361
timestamp 1698431365
transform 1 0 153776 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_1367
timestamp 1698431365
transform 1 0 154448 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1399
timestamp 1698431365
transform 1 0 158032 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_1401
timestamp 1698431365
transform 1 0 158256 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698431365
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_206
timestamp 1698431365
transform 1 0 24416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_276
timestamp 1698431365
transform 1 0 32256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_346
timestamp 1698431365
transform 1 0 40096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_416
timestamp 1698431365
transform 1 0 47936 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_556
timestamp 1698431365
transform 1 0 63616 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_562
timestamp 1698431365
transform 1 0 64288 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_626
timestamp 1698431365
transform 1 0 71456 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_632
timestamp 1698431365
transform 1 0 72128 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_696
timestamp 1698431365
transform 1 0 79296 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_702
timestamp 1698431365
transform 1 0 79968 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_766
timestamp 1698431365
transform 1 0 87136 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_772
timestamp 1698431365
transform 1 0 87808 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_836
timestamp 1698431365
transform 1 0 94976 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_842
timestamp 1698431365
transform 1 0 95648 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_906
timestamp 1698431365
transform 1 0 102816 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_912
timestamp 1698431365
transform 1 0 103488 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_976
timestamp 1698431365
transform 1 0 110656 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_982
timestamp 1698431365
transform 1 0 111328 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1014
timestamp 1698431365
transform 1 0 114912 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1018
timestamp 1698431365
transform 1 0 115360 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1026
timestamp 1698431365
transform 1 0 116256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_1030
timestamp 1698431365
transform 1 0 116704 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1046
timestamp 1698431365
transform 1 0 118496 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1052
timestamp 1698431365
transform 1 0 119168 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1116
timestamp 1698431365
transform 1 0 126336 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1122
timestamp 1698431365
transform 1 0 127008 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1186
timestamp 1698431365
transform 1 0 134176 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1192
timestamp 1698431365
transform 1 0 134848 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1256
timestamp 1698431365
transform 1 0 142016 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1262
timestamp 1698431365
transform 1 0 142688 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1326
timestamp 1698431365
transform 1 0 149856 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1332
timestamp 1698431365
transform 1 0 150528 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1396
timestamp 1698431365
transform 1 0 157696 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_171
timestamp 1698431365
transform 1 0 20496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_209
timestamp 1698431365
transform 1 0 24752 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_225
timestamp 1698431365
transform 1 0 26544 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_233
timestamp 1698431365
transform 1 0 27440 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_244
timestamp 1698431365
transform 1 0 28672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_251
timestamp 1698431365
transform 1 0 29456 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_381
timestamp 1698431365
transform 1 0 44016 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_419
timestamp 1698431365
transform 1 0 48272 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_427
timestamp 1698431365
transform 1 0 49168 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_437
timestamp 1698431365
transform 1 0 50288 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_453
timestamp 1698431365
transform 1 0 52080 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_473
timestamp 1698431365
transform 1 0 54320 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_477
timestamp 1698431365
transform 1 0 54768 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_481
timestamp 1698431365
transform 1 0 55216 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_513
timestamp 1698431365
transform 1 0 58800 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_521
timestamp 1698431365
transform 1 0 59696 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_537
timestamp 1698431365
transform 1 0 61488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_541
timestamp 1698431365
transform 1 0 61936 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_545
timestamp 1698431365
transform 1 0 62384 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_577
timestamp 1698431365
transform 1 0 65968 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_583
timestamp 1698431365
transform 1 0 66640 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_591
timestamp 1698431365
transform 1 0 67536 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_597
timestamp 1698431365
transform 1 0 68208 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_605
timestamp 1698431365
transform 1 0 69104 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_609
timestamp 1698431365
transform 1 0 69552 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_624
timestamp 1698431365
transform 1 0 71232 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_628
timestamp 1698431365
transform 1 0 71680 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_660
timestamp 1698431365
transform 1 0 75264 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_664
timestamp 1698431365
transform 1 0 75712 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_667
timestamp 1698431365
transform 1 0 76048 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_675
timestamp 1698431365
transform 1 0 76944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_679
timestamp 1698431365
transform 1 0 77392 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_685
timestamp 1698431365
transform 1 0 78064 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_701
timestamp 1698431365
transform 1 0 79856 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_709
timestamp 1698431365
transform 1 0 80752 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_711
timestamp 1698431365
transform 1 0 80976 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_720
timestamp 1698431365
transform 1 0 81984 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_728
timestamp 1698431365
transform 1 0 82880 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_732
timestamp 1698431365
transform 1 0 83328 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_734
timestamp 1698431365
transform 1 0 83552 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_737
timestamp 1698431365
transform 1 0 83888 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_769
timestamp 1698431365
transform 1 0 87472 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_777
timestamp 1698431365
transform 1 0 88368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_781
timestamp 1698431365
transform 1 0 88816 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_787
timestamp 1698431365
transform 1 0 89488 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_803
timestamp 1698431365
transform 1 0 91280 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_807
timestamp 1698431365
transform 1 0 91728 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_811
timestamp 1698431365
transform 1 0 92176 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_813
timestamp 1698431365
transform 1 0 92400 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_822
timestamp 1698431365
transform 1 0 93408 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_838
timestamp 1698431365
transform 1 0 95200 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_846
timestamp 1698431365
transform 1 0 96096 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_850
timestamp 1698431365
transform 1 0 96544 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_852
timestamp 1698431365
transform 1 0 96768 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_855
timestamp 1698431365
transform 1 0 97104 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_871
timestamp 1698431365
transform 1 0 98896 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_877
timestamp 1698431365
transform 1 0 99568 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_885
timestamp 1698431365
transform 1 0 100464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_889
timestamp 1698431365
transform 1 0 100912 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_905
timestamp 1698431365
transform 1 0 102704 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_913
timestamp 1698431365
transform 1 0 103600 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_915
timestamp 1698431365
transform 1 0 103824 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_924
timestamp 1698431365
transform 1 0 104832 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_940
timestamp 1698431365
transform 1 0 106624 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_944
timestamp 1698431365
transform 1 0 107072 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_947
timestamp 1698431365
transform 1 0 107408 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_957
timestamp 1698431365
transform 1 0 108528 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_991
timestamp 1698431365
transform 1 0 112336 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1007
timestamp 1698431365
transform 1 0 114128 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1017
timestamp 1698431365
transform 1 0 115248 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1019
timestamp 1698431365
transform 1 0 115472 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1030
timestamp 1698431365
transform 1 0 116704 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1046
timestamp 1698431365
transform 1 0 118496 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1054
timestamp 1698431365
transform 1 0 119392 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1056
timestamp 1698431365
transform 1 0 119616 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1059
timestamp 1698431365
transform 1 0 119952 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1075
timestamp 1698431365
transform 1 0 121744 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1083
timestamp 1698431365
transform 1 0 122640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1087
timestamp 1698431365
transform 1 0 123088 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1093
timestamp 1698431365
transform 1 0 123760 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1109
timestamp 1698431365
transform 1 0 125552 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1117
timestamp 1698431365
transform 1 0 126448 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1119
timestamp 1698431365
transform 1 0 126672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1128
timestamp 1698431365
transform 1 0 127680 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1144
timestamp 1698431365
transform 1 0 129472 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1152
timestamp 1698431365
transform 1 0 130368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1154
timestamp 1698431365
transform 1 0 130592 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1157
timestamp 1698431365
transform 1 0 130928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_1161
timestamp 1698431365
transform 1 0 131376 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1195
timestamp 1698431365
transform 1 0 135184 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1211
timestamp 1698431365
transform 1 0 136976 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1219
timestamp 1698431365
transform 1 0 137872 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1233
timestamp 1698431365
transform 1 0 139440 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1249
timestamp 1698431365
transform 1 0 141232 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1257
timestamp 1698431365
transform 1 0 142128 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_1263
timestamp 1698431365
transform 1 0 142800 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1297
timestamp 1698431365
transform 1 0 146608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_1301
timestamp 1698431365
transform 1 0 147056 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1333
timestamp 1698431365
transform 1 0 150640 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1349
timestamp 1698431365
transform 1 0 152432 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1357
timestamp 1698431365
transform 1 0 153328 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1361
timestamp 1698431365
transform 1 0 153776 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_1367
timestamp 1698431365
transform 1 0 154448 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1399
timestamp 1698431365
transform 1 0 158032 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1401
timestamp 1698431365
transform 1 0 158256 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_18
timestamp 1698431365
transform 1 0 3360 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_26
timestamp 1698431365
transform 1 0 4256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_30
timestamp 1698431365
transform 1 0 4704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_36
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_38
timestamp 1698431365
transform 1 0 5600 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_45
timestamp 1698431365
transform 1 0 6384 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_61
timestamp 1698431365
transform 1 0 8176 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_65
timestamp 1698431365
transform 1 0 8624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_67
timestamp 1698431365
transform 1 0 8848 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_104
timestamp 1698431365
transform 1 0 12992 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_106
timestamp 1698431365
transform 1 0 13216 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_111
timestamp 1698431365
transform 1 0 13776 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_127
timestamp 1698431365
transform 1 0 15568 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_135
timestamp 1698431365
transform 1 0 16464 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_140
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_167
timestamp 1698431365
transform 1 0 20048 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_169
timestamp 1698431365
transform 1 0 20272 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_172
timestamp 1698431365
transform 1 0 20608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_176
timestamp 1698431365
transform 1 0 21056 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_192
timestamp 1698431365
transform 1 0 22848 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_200
timestamp 1698431365
transform 1 0 23744 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_206
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_208
timestamp 1698431365
transform 1 0 24640 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_213
timestamp 1698431365
transform 1 0 25200 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_229
timestamp 1698431365
transform 1 0 26992 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_237
timestamp 1698431365
transform 1 0 27888 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_240
timestamp 1698431365
transform 1 0 28224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_242
timestamp 1698431365
transform 1 0 28448 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_269
timestamp 1698431365
transform 1 0 31472 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_271
timestamp 1698431365
transform 1 0 31696 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_274
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_308
timestamp 1698431365
transform 1 0 35840 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_310
timestamp 1698431365
transform 1 0 36064 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_315
timestamp 1698431365
transform 1 0 36624 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_331
timestamp 1698431365
transform 1 0 38416 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_339
timestamp 1698431365
transform 1 0 39312 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_342
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_344
timestamp 1698431365
transform 1 0 39872 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_371
timestamp 1698431365
transform 1 0 42896 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_373
timestamp 1698431365
transform 1 0 43120 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_376
timestamp 1698431365
transform 1 0 43456 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_380
timestamp 1698431365
transform 1 0 43904 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_396
timestamp 1698431365
transform 1 0 45696 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_404
timestamp 1698431365
transform 1 0 46592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_410
timestamp 1698431365
transform 1 0 47264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_412
timestamp 1698431365
transform 1 0 47488 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_417
timestamp 1698431365
transform 1 0 48048 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_433
timestamp 1698431365
transform 1 0 49840 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_441
timestamp 1698431365
transform 1 0 50736 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_444
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_446
timestamp 1698431365
transform 1 0 51296 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_473
timestamp 1698431365
transform 1 0 54320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_475
timestamp 1698431365
transform 1 0 54544 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_478
timestamp 1698431365
transform 1 0 54880 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_480
timestamp 1698431365
transform 1 0 55104 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_489
timestamp 1698431365
transform 1 0 56112 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_505
timestamp 1698431365
transform 1 0 57904 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_509
timestamp 1698431365
transform 1 0 58352 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_512
timestamp 1698431365
transform 1 0 58688 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_514
timestamp 1698431365
transform 1 0 58912 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_541
timestamp 1698431365
transform 1 0 61936 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_543
timestamp 1698431365
transform 1 0 62160 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_546
timestamp 1698431365
transform 1 0 62496 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_548
timestamp 1698431365
transform 1 0 62720 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_575
timestamp 1698431365
transform 1 0 65744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_577
timestamp 1698431365
transform 1 0 65968 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_580
timestamp 1698431365
transform 1 0 66304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_582
timestamp 1698431365
transform 1 0 66528 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_589
timestamp 1698431365
transform 1 0 67312 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_605
timestamp 1698431365
transform 1 0 69104 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_609
timestamp 1698431365
transform 1 0 69552 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_611
timestamp 1698431365
transform 1 0 69776 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_614
timestamp 1698431365
transform 1 0 70112 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_616
timestamp 1698431365
transform 1 0 70336 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_643
timestamp 1698431365
transform 1 0 73360 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_645
timestamp 1698431365
transform 1 0 73584 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_648
timestamp 1698431365
transform 1 0 73920 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_650
timestamp 1698431365
transform 1 0 74144 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_677
timestamp 1698431365
transform 1 0 77168 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_679
timestamp 1698431365
transform 1 0 77392 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_682
timestamp 1698431365
transform 1 0 77728 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_684
timestamp 1698431365
transform 1 0 77952 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_691
timestamp 1698431365
transform 1 0 78736 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_707
timestamp 1698431365
transform 1 0 80528 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_711
timestamp 1698431365
transform 1 0 80976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_713
timestamp 1698431365
transform 1 0 81200 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_716
timestamp 1698431365
transform 1 0 81536 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_718
timestamp 1698431365
transform 1 0 81760 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_745
timestamp 1698431365
transform 1 0 84784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_747
timestamp 1698431365
transform 1 0 85008 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_750
timestamp 1698431365
transform 1 0 85344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_752
timestamp 1698431365
transform 1 0 85568 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_779
timestamp 1698431365
transform 1 0 88592 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_781
timestamp 1698431365
transform 1 0 88816 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_784
timestamp 1698431365
transform 1 0 89152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_786
timestamp 1698431365
transform 1 0 89376 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_793
timestamp 1698431365
transform 1 0 90160 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_809
timestamp 1698431365
transform 1 0 91952 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_813
timestamp 1698431365
transform 1 0 92400 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_815
timestamp 1698431365
transform 1 0 92624 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_818
timestamp 1698431365
transform 1 0 92960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_820
timestamp 1698431365
transform 1 0 93184 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_847
timestamp 1698431365
transform 1 0 96208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_849
timestamp 1698431365
transform 1 0 96432 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_852
timestamp 1698431365
transform 1 0 96768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_854
timestamp 1698431365
transform 1 0 96992 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_881
timestamp 1698431365
transform 1 0 100016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_883
timestamp 1698431365
transform 1 0 100240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_886
timestamp 1698431365
transform 1 0 100576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_888
timestamp 1698431365
transform 1 0 100800 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_895
timestamp 1698431365
transform 1 0 101584 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_911
timestamp 1698431365
transform 1 0 103376 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_915
timestamp 1698431365
transform 1 0 103824 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_917
timestamp 1698431365
transform 1 0 104048 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_920
timestamp 1698431365
transform 1 0 104384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_922
timestamp 1698431365
transform 1 0 104608 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_949
timestamp 1698431365
transform 1 0 107632 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_951
timestamp 1698431365
transform 1 0 107856 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_954
timestamp 1698431365
transform 1 0 108192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_956
timestamp 1698431365
transform 1 0 108416 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_983
timestamp 1698431365
transform 1 0 111440 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_985
timestamp 1698431365
transform 1 0 111664 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_988
timestamp 1698431365
transform 1 0 112000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_990
timestamp 1698431365
transform 1 0 112224 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_997
timestamp 1698431365
transform 1 0 113008 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1013
timestamp 1698431365
transform 1 0 114800 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1017
timestamp 1698431365
transform 1 0 115248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1019
timestamp 1698431365
transform 1 0 115472 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1022
timestamp 1698431365
transform 1 0 115808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1024
timestamp 1698431365
transform 1 0 116032 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1051
timestamp 1698431365
transform 1 0 119056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1053
timestamp 1698431365
transform 1 0 119280 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1056
timestamp 1698431365
transform 1 0 119616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1058
timestamp 1698431365
transform 1 0 119840 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1085
timestamp 1698431365
transform 1 0 122864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1087
timestamp 1698431365
transform 1 0 123088 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1090
timestamp 1698431365
transform 1 0 123424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1092
timestamp 1698431365
transform 1 0 123648 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1099
timestamp 1698431365
transform 1 0 124432 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1115
timestamp 1698431365
transform 1 0 126224 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1119
timestamp 1698431365
transform 1 0 126672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1121
timestamp 1698431365
transform 1 0 126896 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1124
timestamp 1698431365
transform 1 0 127232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1126
timestamp 1698431365
transform 1 0 127456 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1153
timestamp 1698431365
transform 1 0 130480 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1155
timestamp 1698431365
transform 1 0 130704 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1158
timestamp 1698431365
transform 1 0 131040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1160
timestamp 1698431365
transform 1 0 131264 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1187
timestamp 1698431365
transform 1 0 134288 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1189
timestamp 1698431365
transform 1 0 134512 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1192
timestamp 1698431365
transform 1 0 134848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1194
timestamp 1698431365
transform 1 0 135072 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1203
timestamp 1698431365
transform 1 0 136080 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1219
timestamp 1698431365
transform 1 0 137872 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1223
timestamp 1698431365
transform 1 0 138320 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1226
timestamp 1698431365
transform 1 0 138656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1228
timestamp 1698431365
transform 1 0 138880 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1255
timestamp 1698431365
transform 1 0 141904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1257
timestamp 1698431365
transform 1 0 142128 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1260
timestamp 1698431365
transform 1 0 142464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1262
timestamp 1698431365
transform 1 0 142688 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1289
timestamp 1698431365
transform 1 0 145712 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1291
timestamp 1698431365
transform 1 0 145936 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1294
timestamp 1698431365
transform 1 0 146272 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1296
timestamp 1698431365
transform 1 0 146496 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1305
timestamp 1698431365
transform 1 0 147504 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1321
timestamp 1698431365
transform 1 0 149296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1323
timestamp 1698431365
transform 1 0 149520 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1328
timestamp 1698431365
transform 1 0 150080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1330
timestamp 1698431365
transform 1 0 150304 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1357
timestamp 1698431365
transform 1 0 153328 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1359
timestamp 1698431365
transform 1 0 153552 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1362
timestamp 1698431365
transform 1 0 153888 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1364
timestamp 1698431365
transform 1 0 154112 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1391
timestamp 1698431365
transform 1 0 157136 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1393
timestamp 1698431365
transform 1 0 157360 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1396
timestamp 1698431365
transform 1 0 157696 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1400
timestamp 1698431365
transform 1 0 158144 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 95200 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform 1 0 46032 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 71232 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform -1 0 58912 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform -1 0 81760 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform -1 0 117040 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform -1 0 105728 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform -1 0 75712 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform -1 0 64064 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform -1 0 111104 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform 1 0 107408 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform -1 0 86352 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform -1 0 102368 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform -1 0 105392 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform -1 0 123872 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform 1 0 101360 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform 1 0 58352 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform -1 0 91056 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform -1 0 24864 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform 1 0 119168 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform -1 0 48160 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform -1 0 23968 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform -1 0 71904 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform 1 0 41664 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold26
timestamp 1698431365
transform -1 0 75824 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform -1 0 32704 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform -1 0 29904 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform 1 0 98784 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold30
timestamp 1698431365
transform 1 0 115248 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform 1 0 108640 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform 1 0 124992 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform 1 0 80080 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold34
timestamp 1698431365
transform 1 0 61264 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform -1 0 31472 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold36
timestamp 1698431365
transform -1 0 78736 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold37
timestamp 1698431365
transform -1 0 91504 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold38
timestamp 1698431365
transform -1 0 132384 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold39
timestamp 1698431365
transform -1 0 102368 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold40
timestamp 1698431365
transform 1 0 91728 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold41
timestamp 1698431365
transform -1 0 54992 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold42
timestamp 1698431365
transform 1 0 67648 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold43
timestamp 1698431365
transform 1 0 57008 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold44
timestamp 1698431365
transform 1 0 133616 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold45
timestamp 1698431365
transform -1 0 36624 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold46
timestamp 1698431365
transform 1 0 53648 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold47
timestamp 1698431365
transform -1 0 36512 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold48
timestamp 1698431365
transform -1 0 34720 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold49
timestamp 1698431365
transform 1 0 17920 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold50 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38416 0 1 9408
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold51
timestamp 1698431365
transform -1 0 27888 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold52
timestamp 1698431365
transform 1 0 137536 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold53
timestamp 1698431365
transform 1 0 49504 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold54
timestamp 1698431365
transform -1 0 32704 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold55
timestamp 1698431365
transform -1 0 144592 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold56
timestamp 1698431365
transform 1 0 149296 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold57
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold58
timestamp 1698431365
transform -1 0 149520 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold59
timestamp 1698431365
transform 1 0 45920 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold60
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold61
timestamp 1698431365
transform 1 0 41216 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold62
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold63
timestamp 1698431365
transform -1 0 122752 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  hold64
timestamp 1698431365
transform -1 0 111104 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  hold65
timestamp 1698431365
transform -1 0 69552 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold66
timestamp 1698431365
transform 1 0 115808 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold67
timestamp 1698431365
transform 1 0 143920 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold68
timestamp 1698431365
transform -1 0 141792 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold69
timestamp 1698431365
transform 1 0 104048 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold70
timestamp 1698431365
transform -1 0 56224 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold71
timestamp 1698431365
transform 1 0 95984 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold72
timestamp 1698431365
transform -1 0 94640 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold73
timestamp 1698431365
transform -1 0 48720 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold74
timestamp 1698431365
transform 1 0 69104 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold75
timestamp 1698431365
transform -1 0 27888 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold76
timestamp 1698431365
transform -1 0 82768 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold77
timestamp 1698431365
transform -1 0 93408 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold78
timestamp 1698431365
transform 1 0 86352 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold79
timestamp 1698431365
transform -1 0 44464 0 1 7840
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold80
timestamp 1698431365
transform 1 0 46256 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold81
timestamp 1698431365
transform -1 0 64064 0 -1 7840
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold82
timestamp 1698431365
transform -1 0 60144 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold83
timestamp 1698431365
transform 1 0 99792 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold84
timestamp 1698431365
transform -1 0 110656 0 1 7840
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold86
timestamp 1698431365
transform -1 0 71008 0 1 7840
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold87
timestamp 1698431365
transform 1 0 76720 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold88
timestamp 1698431365
transform 1 0 29568 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold89
timestamp 1698431365
transform 1 0 112000 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold90
timestamp 1698431365
transform -1 0 39648 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold91
timestamp 1698431365
transform 1 0 61264 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold92
timestamp 1698431365
transform 1 0 114576 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold93
timestamp 1698431365
transform -1 0 72352 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold94
timestamp 1698431365
transform -1 0 82768 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold95
timestamp 1698431365
transform -1 0 125888 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold96
timestamp 1698431365
transform -1 0 60144 0 1 7840
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold97
timestamp 1698431365
transform -1 0 108528 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold98
timestamp 1698431365
transform -1 0 61264 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold99
timestamp 1698431365
transform -1 0 90608 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold100
timestamp 1698431365
transform 1 0 91280 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold101
timestamp 1698431365
transform -1 0 79744 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold102
timestamp 1698431365
transform -1 0 130592 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold103
timestamp 1698431365
transform -1 0 120624 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold104
timestamp 1698431365
transform 1 0 95984 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold105
timestamp 1698431365
transform -1 0 114128 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold106
timestamp 1698431365
transform -1 0 128688 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold107
timestamp 1698431365
transform 1 0 73024 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold108
timestamp 1698431365
transform 1 0 118160 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold109
timestamp 1698431365
transform 1 0 98560 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold110
timestamp 1698431365
transform -1 0 107184 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform -1 0 124432 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2
timestamp 1698431365
transform 1 0 135184 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform 1 0 146608 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input4
timestamp 1698431365
transform 1 0 55216 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform 1 0 66640 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 78064 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698431365
transform 1 0 89488 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input8
timestamp 1698431365
transform 1 0 100912 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform -1 0 113008 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input10
timestamp 1698431365
transform 1 0 5712 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform 1 0 10640 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input12
timestamp 1698431365
transform -1 0 19264 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input13
timestamp 1698431365
transform 1 0 64288 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input14
timestamp 1698431365
transform -1 0 67984 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input15
timestamp 1698431365
transform 1 0 71008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input16
timestamp 1698431365
transform -1 0 76944 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input17
timestamp 1698431365
transform -1 0 82208 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input18
timestamp 1698431365
transform -1 0 86912 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 86016 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input20
timestamp 1698431365
transform 1 0 94080 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input21
timestamp 1698431365
transform -1 0 101248 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input22
timestamp 1698431365
transform -1 0 102144 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input23
timestamp 1698431365
transform -1 0 22064 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 108864 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input25
timestamp 1698431365
transform -1 0 115584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input26
timestamp 1698431365
transform -1 0 119392 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input27
timestamp 1698431365
transform 1 0 117600 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 120736 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 123872 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 127792 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 133056 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 135296 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 143360 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input34
timestamp 1698431365
transform -1 0 26992 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform -1 0 145264 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform -1 0 148400 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 24192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input39
timestamp 1698431365
transform -1 0 43456 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input40
timestamp 1698431365
transform -1 0 42784 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input41
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input42
timestamp 1698431365
transform 1 0 54992 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input43
timestamp 1698431365
transform -1 0 58464 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform 1 0 13328 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform 1 0 16352 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform -1 0 63168 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform -1 0 69104 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform 1 0 72128 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform -1 0 73696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform 1 0 79296 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698431365
transform 1 0 83888 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1698431365
transform -1 0 89824 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1698431365
transform -1 0 97440 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1698431365
transform -1 0 107856 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform 1 0 101696 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1698431365
transform 1 0 22400 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1698431365
transform 1 0 104384 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1698431365
transform 1 0 108976 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1698431365
transform -1 0 115360 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1698431365
transform -1 0 123200 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1698431365
transform -1 0 121632 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1698431365
transform -1 0 127008 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1698431365
transform -1 0 129360 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1698431365
transform -1 0 134624 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input65
timestamp 1698431365
transform -1 0 138432 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input66
timestamp 1698431365
transform -1 0 142240 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input67
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input68
timestamp 1698431365
transform -1 0 146048 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input69
timestamp 1698431365
transform -1 0 150192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input70
timestamp 1698431365
transform -1 0 28896 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input71
timestamp 1698431365
transform -1 0 43232 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input72
timestamp 1698431365
transform -1 0 47936 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input73
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1698431365
transform 1 0 53424 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1698431365
transform 1 0 55552 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1698431365
transform -1 0 62272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input77
timestamp 1698431365
transform -1 0 18144 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1698431365
transform 1 0 22624 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input79
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input80
timestamp 1698431365
transform 1 0 34720 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input81
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input82
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output83 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 127568 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output84
timestamp 1698431365
transform 1 0 138992 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output85
timestamp 1698431365
transform 1 0 150416 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output86
timestamp 1698431365
transform -1 0 61936 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output87
timestamp 1698431365
transform 1 0 70448 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output88
timestamp 1698431365
transform 1 0 81872 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output89
timestamp 1698431365
transform 1 0 93296 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output90
timestamp 1698431365
transform 1 0 104720 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output91
timestamp 1698431365
transform 1 0 116144 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output92
timestamp 1698431365
transform -1 0 20048 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output93
timestamp 1698431365
transform 1 0 131376 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output94
timestamp 1698431365
transform 1 0 142800 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output95
timestamp 1698431365
transform 1 0 154224 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output96
timestamp 1698431365
transform 1 0 28560 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output97
timestamp 1698431365
transform -1 0 42896 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output98
timestamp 1698431365
transform 1 0 51408 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output99
timestamp 1698431365
transform 1 0 62832 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output100
timestamp 1698431365
transform -1 0 77168 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output101
timestamp 1698431365
transform -1 0 88592 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output102
timestamp 1698431365
transform 1 0 97104 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output103
timestamp 1698431365
transform 1 0 108528 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output104
timestamp 1698431365
transform 1 0 119952 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output105
timestamp 1698431365
transform -1 0 15904 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output106
timestamp 1698431365
transform -1 0 23520 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output107
timestamp 1698431365
transform -1 0 66080 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output108
timestamp 1698431365
transform -1 0 73024 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output109
timestamp 1698431365
transform -1 0 76720 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output110
timestamp 1698431365
transform 1 0 77840 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output111
timestamp 1698431365
transform 1 0 81872 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output112
timestamp 1698431365
transform 1 0 85904 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output113
timestamp 1698431365
transform -1 0 92736 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output114
timestamp 1698431365
transform -1 0 98560 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output115
timestamp 1698431365
transform -1 0 100352 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output116
timestamp 1698431365
transform -1 0 104160 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output117
timestamp 1698431365
transform -1 0 28000 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output118
timestamp 1698431365
transform 1 0 106064 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output119
timestamp 1698431365
transform 1 0 108864 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output120
timestamp 1698431365
transform 1 0 115808 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output121
timestamp 1698431365
transform 1 0 119616 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output122
timestamp 1698431365
transform 1 0 123424 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output123
timestamp 1698431365
transform 1 0 127232 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output124
timestamp 1698431365
transform 1 0 131040 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output125
timestamp 1698431365
transform 1 0 134848 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output126
timestamp 1698431365
transform 1 0 138656 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output127
timestamp 1698431365
transform 1 0 142464 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output128
timestamp 1698431365
transform -1 0 31808 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output129
timestamp 1698431365
transform 1 0 146384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output130
timestamp 1698431365
transform 1 0 150416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output131
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output132
timestamp 1698431365
transform 1 0 43456 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output133
timestamp 1698431365
transform -1 0 47040 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output134
timestamp 1698431365
transform 1 0 47936 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output135
timestamp 1698431365
transform 1 0 51744 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output136
timestamp 1698431365
transform -1 0 61600 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output137
timestamp 1698431365
transform -1 0 63840 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 158592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 158592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 158592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 158592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 158592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 158592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 158592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 158592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 158592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 158592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 158592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 158592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 158592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 158592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 158592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 158592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 158592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 158592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 158592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 158592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 158592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 158592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 158592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 158592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 158592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 158592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 158592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 158592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 158592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 158592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 158592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 158592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 158592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 158592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 158592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 158592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 158592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 158592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 158592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 158592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 158592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 158592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 158592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 158592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 158592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 158592 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 158592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 158592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 158592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 158592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 158592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 158592 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 158592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 158592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 158592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 158592 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 158592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 158592 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 158592 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 158592 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 158592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 158592 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 158592 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 158592 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 158592 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 158592 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 158592 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 158592 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_150
timestamp 1698431365
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_151
timestamp 1698431365
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_152
timestamp 1698431365
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_153
timestamp 1698431365
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_154
timestamp 1698431365
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_155
timestamp 1698431365
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_156
timestamp 1698431365
transform 1 0 81312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_157
timestamp 1698431365
transform 1 0 85120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_158
timestamp 1698431365
transform 1 0 88928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_159
timestamp 1698431365
transform 1 0 92736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_160
timestamp 1698431365
transform 1 0 96544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_161
timestamp 1698431365
transform 1 0 100352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_162
timestamp 1698431365
transform 1 0 104160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_163
timestamp 1698431365
transform 1 0 107968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_164
timestamp 1698431365
transform 1 0 111776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_165
timestamp 1698431365
transform 1 0 115584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_166
timestamp 1698431365
transform 1 0 119392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_167
timestamp 1698431365
transform 1 0 123200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_168
timestamp 1698431365
transform 1 0 127008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_169
timestamp 1698431365
transform 1 0 130816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_170
timestamp 1698431365
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_171
timestamp 1698431365
transform 1 0 138432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_172
timestamp 1698431365
transform 1 0 142240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_173
timestamp 1698431365
transform 1 0 146048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_174
timestamp 1698431365
transform 1 0 149856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_175
timestamp 1698431365
transform 1 0 153664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_176
timestamp 1698431365
transform 1 0 157472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_177
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_178
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_179
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_180
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_181
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_182
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_183
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_184
timestamp 1698431365
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_185
timestamp 1698431365
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_186
timestamp 1698431365
transform 1 0 79744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_187
timestamp 1698431365
transform 1 0 87584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_188
timestamp 1698431365
transform 1 0 95424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_189
timestamp 1698431365
transform 1 0 103264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_190
timestamp 1698431365
transform 1 0 111104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_191
timestamp 1698431365
transform 1 0 118944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_192
timestamp 1698431365
transform 1 0 126784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_193
timestamp 1698431365
transform 1 0 134624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_194
timestamp 1698431365
transform 1 0 142464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_195
timestamp 1698431365
transform 1 0 150304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_196
timestamp 1698431365
transform 1 0 158144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_197
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_198
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_199
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_200
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_201
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_202
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_203
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_204
timestamp 1698431365
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_205
timestamp 1698431365
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_206
timestamp 1698431365
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_207
timestamp 1698431365
transform 1 0 83664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_208
timestamp 1698431365
transform 1 0 91504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_209
timestamp 1698431365
transform 1 0 99344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_210
timestamp 1698431365
transform 1 0 107184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_211
timestamp 1698431365
transform 1 0 115024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_212
timestamp 1698431365
transform 1 0 122864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_213
timestamp 1698431365
transform 1 0 130704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_214
timestamp 1698431365
transform 1 0 138544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_215
timestamp 1698431365
transform 1 0 146384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_216
timestamp 1698431365
transform 1 0 154224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_217
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_218
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_219
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_220
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_221
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_222
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_223
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_224
timestamp 1698431365
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_225
timestamp 1698431365
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_226
timestamp 1698431365
transform 1 0 79744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_227
timestamp 1698431365
transform 1 0 87584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_228
timestamp 1698431365
transform 1 0 95424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_229
timestamp 1698431365
transform 1 0 103264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_230
timestamp 1698431365
transform 1 0 111104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_231
timestamp 1698431365
transform 1 0 118944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_232
timestamp 1698431365
transform 1 0 126784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_233
timestamp 1698431365
transform 1 0 134624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_234
timestamp 1698431365
transform 1 0 142464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_235
timestamp 1698431365
transform 1 0 150304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_236
timestamp 1698431365
transform 1 0 158144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_237
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_238
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_239
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_240
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_241
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_242
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_243
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_244
timestamp 1698431365
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_245
timestamp 1698431365
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_246
timestamp 1698431365
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_247
timestamp 1698431365
transform 1 0 83664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_248
timestamp 1698431365
transform 1 0 91504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_249
timestamp 1698431365
transform 1 0 99344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_250
timestamp 1698431365
transform 1 0 107184 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_251
timestamp 1698431365
transform 1 0 115024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_252
timestamp 1698431365
transform 1 0 122864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_253
timestamp 1698431365
transform 1 0 130704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_254
timestamp 1698431365
transform 1 0 138544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_255
timestamp 1698431365
transform 1 0 146384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_256
timestamp 1698431365
transform 1 0 154224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_257
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_258
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_259
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_260
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_261
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_262
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_263
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_264
timestamp 1698431365
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_265
timestamp 1698431365
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_266
timestamp 1698431365
transform 1 0 79744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_267
timestamp 1698431365
transform 1 0 87584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_268
timestamp 1698431365
transform 1 0 95424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_269
timestamp 1698431365
transform 1 0 103264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_270
timestamp 1698431365
transform 1 0 111104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_271
timestamp 1698431365
transform 1 0 118944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_272
timestamp 1698431365
transform 1 0 126784 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_273
timestamp 1698431365
transform 1 0 134624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_274
timestamp 1698431365
transform 1 0 142464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_275
timestamp 1698431365
transform 1 0 150304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_276
timestamp 1698431365
transform 1 0 158144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_277
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_278
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_279
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_280
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_281
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_282
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_283
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_284
timestamp 1698431365
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_285
timestamp 1698431365
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_286
timestamp 1698431365
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_287
timestamp 1698431365
transform 1 0 83664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_288
timestamp 1698431365
transform 1 0 91504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_289
timestamp 1698431365
transform 1 0 99344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_290
timestamp 1698431365
transform 1 0 107184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_291
timestamp 1698431365
transform 1 0 115024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_292
timestamp 1698431365
transform 1 0 122864 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_293
timestamp 1698431365
transform 1 0 130704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_294
timestamp 1698431365
transform 1 0 138544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_295
timestamp 1698431365
transform 1 0 146384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_296
timestamp 1698431365
transform 1 0 154224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_297
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_298
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_299
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_300
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_301
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_302
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_303
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_304
timestamp 1698431365
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_305
timestamp 1698431365
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_306
timestamp 1698431365
transform 1 0 79744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_307
timestamp 1698431365
transform 1 0 87584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_308
timestamp 1698431365
transform 1 0 95424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_309
timestamp 1698431365
transform 1 0 103264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_310
timestamp 1698431365
transform 1 0 111104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_311
timestamp 1698431365
transform 1 0 118944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_312
timestamp 1698431365
transform 1 0 126784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_313
timestamp 1698431365
transform 1 0 134624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_314
timestamp 1698431365
transform 1 0 142464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_315
timestamp 1698431365
transform 1 0 150304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_316
timestamp 1698431365
transform 1 0 158144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_317
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_318
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_319
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_320
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_321
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_322
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_323
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_324
timestamp 1698431365
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_325
timestamp 1698431365
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_326
timestamp 1698431365
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_327
timestamp 1698431365
transform 1 0 83664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_328
timestamp 1698431365
transform 1 0 91504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_329
timestamp 1698431365
transform 1 0 99344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_330
timestamp 1698431365
transform 1 0 107184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_331
timestamp 1698431365
transform 1 0 115024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_332
timestamp 1698431365
transform 1 0 122864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_333
timestamp 1698431365
transform 1 0 130704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_334
timestamp 1698431365
transform 1 0 138544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_335
timestamp 1698431365
transform 1 0 146384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_336
timestamp 1698431365
transform 1 0 154224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_337
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_338
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_339
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_340
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_341
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_342
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_343
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_344
timestamp 1698431365
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_345
timestamp 1698431365
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_346
timestamp 1698431365
transform 1 0 79744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_347
timestamp 1698431365
transform 1 0 87584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_348
timestamp 1698431365
transform 1 0 95424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_349
timestamp 1698431365
transform 1 0 103264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_350
timestamp 1698431365
transform 1 0 111104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_351
timestamp 1698431365
transform 1 0 118944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_352
timestamp 1698431365
transform 1 0 126784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_353
timestamp 1698431365
transform 1 0 134624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_354
timestamp 1698431365
transform 1 0 142464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_355
timestamp 1698431365
transform 1 0 150304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_356
timestamp 1698431365
transform 1 0 158144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_357
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_358
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_359
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_360
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_361
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_362
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_363
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_364
timestamp 1698431365
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_365
timestamp 1698431365
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_366
timestamp 1698431365
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_367
timestamp 1698431365
transform 1 0 83664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_368
timestamp 1698431365
transform 1 0 91504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_369
timestamp 1698431365
transform 1 0 99344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_370
timestamp 1698431365
transform 1 0 107184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_371
timestamp 1698431365
transform 1 0 115024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_372
timestamp 1698431365
transform 1 0 122864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_373
timestamp 1698431365
transform 1 0 130704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_374
timestamp 1698431365
transform 1 0 138544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_375
timestamp 1698431365
transform 1 0 146384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_376
timestamp 1698431365
transform 1 0 154224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_377
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_378
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_379
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_380
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_381
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_382
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_383
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_384
timestamp 1698431365
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_385
timestamp 1698431365
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_386
timestamp 1698431365
transform 1 0 79744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_387
timestamp 1698431365
transform 1 0 87584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_388
timestamp 1698431365
transform 1 0 95424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_389
timestamp 1698431365
transform 1 0 103264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_390
timestamp 1698431365
transform 1 0 111104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_391
timestamp 1698431365
transform 1 0 118944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_392
timestamp 1698431365
transform 1 0 126784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_393
timestamp 1698431365
transform 1 0 134624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_394
timestamp 1698431365
transform 1 0 142464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_395
timestamp 1698431365
transform 1 0 150304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_396
timestamp 1698431365
transform 1 0 158144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_397
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_398
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_399
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_400
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_401
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_402
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_403
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_404
timestamp 1698431365
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_405
timestamp 1698431365
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_406
timestamp 1698431365
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_407
timestamp 1698431365
transform 1 0 83664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_408
timestamp 1698431365
transform 1 0 91504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_409
timestamp 1698431365
transform 1 0 99344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_410
timestamp 1698431365
transform 1 0 107184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_411
timestamp 1698431365
transform 1 0 115024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_412
timestamp 1698431365
transform 1 0 122864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_413
timestamp 1698431365
transform 1 0 130704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_414
timestamp 1698431365
transform 1 0 138544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_415
timestamp 1698431365
transform 1 0 146384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_416
timestamp 1698431365
transform 1 0 154224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_417
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_418
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_419
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_420
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_421
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_422
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_423
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_424
timestamp 1698431365
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_425
timestamp 1698431365
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_426
timestamp 1698431365
transform 1 0 79744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_427
timestamp 1698431365
transform 1 0 87584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_428
timestamp 1698431365
transform 1 0 95424 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_429
timestamp 1698431365
transform 1 0 103264 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_430
timestamp 1698431365
transform 1 0 111104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_431
timestamp 1698431365
transform 1 0 118944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_432
timestamp 1698431365
transform 1 0 126784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_433
timestamp 1698431365
transform 1 0 134624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_434
timestamp 1698431365
transform 1 0 142464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_435
timestamp 1698431365
transform 1 0 150304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_436
timestamp 1698431365
transform 1 0 158144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_437
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_438
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_439
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_440
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_441
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_442
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_443
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_444
timestamp 1698431365
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_445
timestamp 1698431365
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_446
timestamp 1698431365
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_447
timestamp 1698431365
transform 1 0 83664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_448
timestamp 1698431365
transform 1 0 91504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_449
timestamp 1698431365
transform 1 0 99344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_450
timestamp 1698431365
transform 1 0 107184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_451
timestamp 1698431365
transform 1 0 115024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_452
timestamp 1698431365
transform 1 0 122864 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_453
timestamp 1698431365
transform 1 0 130704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_454
timestamp 1698431365
transform 1 0 138544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_455
timestamp 1698431365
transform 1 0 146384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_456
timestamp 1698431365
transform 1 0 154224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_457
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_458
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_459
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_460
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_461
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_462
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_463
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_464
timestamp 1698431365
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_465
timestamp 1698431365
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_466
timestamp 1698431365
transform 1 0 79744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_467
timestamp 1698431365
transform 1 0 87584 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_468
timestamp 1698431365
transform 1 0 95424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_469
timestamp 1698431365
transform 1 0 103264 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_470
timestamp 1698431365
transform 1 0 111104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_471
timestamp 1698431365
transform 1 0 118944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_472
timestamp 1698431365
transform 1 0 126784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_473
timestamp 1698431365
transform 1 0 134624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_474
timestamp 1698431365
transform 1 0 142464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_475
timestamp 1698431365
transform 1 0 150304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_476
timestamp 1698431365
transform 1 0 158144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_477
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_478
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_479
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_480
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_481
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_482
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_483
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_484
timestamp 1698431365
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_485
timestamp 1698431365
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_486
timestamp 1698431365
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_487
timestamp 1698431365
transform 1 0 83664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_488
timestamp 1698431365
transform 1 0 91504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_489
timestamp 1698431365
transform 1 0 99344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_490
timestamp 1698431365
transform 1 0 107184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_491
timestamp 1698431365
transform 1 0 115024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_492
timestamp 1698431365
transform 1 0 122864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_493
timestamp 1698431365
transform 1 0 130704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_494
timestamp 1698431365
transform 1 0 138544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_495
timestamp 1698431365
transform 1 0 146384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_496
timestamp 1698431365
transform 1 0 154224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_497
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_498
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_499
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_500
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_501
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_502
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_503
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_504
timestamp 1698431365
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_505
timestamp 1698431365
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_506
timestamp 1698431365
transform 1 0 79744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_507
timestamp 1698431365
transform 1 0 87584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_508
timestamp 1698431365
transform 1 0 95424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_509
timestamp 1698431365
transform 1 0 103264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_510
timestamp 1698431365
transform 1 0 111104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_511
timestamp 1698431365
transform 1 0 118944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_512
timestamp 1698431365
transform 1 0 126784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_513
timestamp 1698431365
transform 1 0 134624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_514
timestamp 1698431365
transform 1 0 142464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_515
timestamp 1698431365
transform 1 0 150304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_516
timestamp 1698431365
transform 1 0 158144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_517
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_518
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_519
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_520
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_521
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_522
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_523
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_524
timestamp 1698431365
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_525
timestamp 1698431365
transform 1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_526
timestamp 1698431365
transform 1 0 75824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_527
timestamp 1698431365
transform 1 0 83664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_528
timestamp 1698431365
transform 1 0 91504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_529
timestamp 1698431365
transform 1 0 99344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_530
timestamp 1698431365
transform 1 0 107184 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_531
timestamp 1698431365
transform 1 0 115024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_532
timestamp 1698431365
transform 1 0 122864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_533
timestamp 1698431365
transform 1 0 130704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_534
timestamp 1698431365
transform 1 0 138544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_535
timestamp 1698431365
transform 1 0 146384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_536
timestamp 1698431365
transform 1 0 154224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_537
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_538
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_539
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_540
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_541
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_542
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_543
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_544
timestamp 1698431365
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_545
timestamp 1698431365
transform 1 0 71904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_546
timestamp 1698431365
transform 1 0 79744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_547
timestamp 1698431365
transform 1 0 87584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_548
timestamp 1698431365
transform 1 0 95424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_549
timestamp 1698431365
transform 1 0 103264 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_550
timestamp 1698431365
transform 1 0 111104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_551
timestamp 1698431365
transform 1 0 118944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_552
timestamp 1698431365
transform 1 0 126784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_553
timestamp 1698431365
transform 1 0 134624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_554
timestamp 1698431365
transform 1 0 142464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_555
timestamp 1698431365
transform 1 0 150304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_556
timestamp 1698431365
transform 1 0 158144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_557
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_558
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_559
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_560
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_561
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_562
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_563
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_564
timestamp 1698431365
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_565
timestamp 1698431365
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_566
timestamp 1698431365
transform 1 0 75824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_567
timestamp 1698431365
transform 1 0 83664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_568
timestamp 1698431365
transform 1 0 91504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_569
timestamp 1698431365
transform 1 0 99344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_570
timestamp 1698431365
transform 1 0 107184 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_571
timestamp 1698431365
transform 1 0 115024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_572
timestamp 1698431365
transform 1 0 122864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_573
timestamp 1698431365
transform 1 0 130704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_574
timestamp 1698431365
transform 1 0 138544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_575
timestamp 1698431365
transform 1 0 146384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_576
timestamp 1698431365
transform 1 0 154224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_577
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_578
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_579
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_580
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_581
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_582
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_583
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_584
timestamp 1698431365
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_585
timestamp 1698431365
transform 1 0 71904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_586
timestamp 1698431365
transform 1 0 79744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_587
timestamp 1698431365
transform 1 0 87584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_588
timestamp 1698431365
transform 1 0 95424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_589
timestamp 1698431365
transform 1 0 103264 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_590
timestamp 1698431365
transform 1 0 111104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_591
timestamp 1698431365
transform 1 0 118944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_592
timestamp 1698431365
transform 1 0 126784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_593
timestamp 1698431365
transform 1 0 134624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_594
timestamp 1698431365
transform 1 0 142464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_595
timestamp 1698431365
transform 1 0 150304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_596
timestamp 1698431365
transform 1 0 158144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_597
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_598
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_599
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_600
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_601
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_602
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_603
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_604
timestamp 1698431365
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_605
timestamp 1698431365
transform 1 0 67984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_606
timestamp 1698431365
transform 1 0 75824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_607
timestamp 1698431365
transform 1 0 83664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_608
timestamp 1698431365
transform 1 0 91504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_609
timestamp 1698431365
transform 1 0 99344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_610
timestamp 1698431365
transform 1 0 107184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_611
timestamp 1698431365
transform 1 0 115024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_612
timestamp 1698431365
transform 1 0 122864 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_613
timestamp 1698431365
transform 1 0 130704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_614
timestamp 1698431365
transform 1 0 138544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_615
timestamp 1698431365
transform 1 0 146384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_616
timestamp 1698431365
transform 1 0 154224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_617
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_618
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_619
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_620
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_621
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_622
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_623
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_624
timestamp 1698431365
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_625
timestamp 1698431365
transform 1 0 71904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_626
timestamp 1698431365
transform 1 0 79744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_627
timestamp 1698431365
transform 1 0 87584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_628
timestamp 1698431365
transform 1 0 95424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_629
timestamp 1698431365
transform 1 0 103264 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_630
timestamp 1698431365
transform 1 0 111104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_631
timestamp 1698431365
transform 1 0 118944 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_632
timestamp 1698431365
transform 1 0 126784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_633
timestamp 1698431365
transform 1 0 134624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_634
timestamp 1698431365
transform 1 0 142464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_635
timestamp 1698431365
transform 1 0 150304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_636
timestamp 1698431365
transform 1 0 158144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_637
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_638
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_639
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_640
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_641
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_642
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_643
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_644
timestamp 1698431365
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_645
timestamp 1698431365
transform 1 0 67984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_646
timestamp 1698431365
transform 1 0 75824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_647
timestamp 1698431365
transform 1 0 83664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_648
timestamp 1698431365
transform 1 0 91504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_649
timestamp 1698431365
transform 1 0 99344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_650
timestamp 1698431365
transform 1 0 107184 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_651
timestamp 1698431365
transform 1 0 115024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_652
timestamp 1698431365
transform 1 0 122864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_653
timestamp 1698431365
transform 1 0 130704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_654
timestamp 1698431365
transform 1 0 138544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_655
timestamp 1698431365
transform 1 0 146384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_656
timestamp 1698431365
transform 1 0 154224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_657
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_658
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_659
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_660
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_661
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_662
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_663
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_664
timestamp 1698431365
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_665
timestamp 1698431365
transform 1 0 71904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_666
timestamp 1698431365
transform 1 0 79744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_667
timestamp 1698431365
transform 1 0 87584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_668
timestamp 1698431365
transform 1 0 95424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_669
timestamp 1698431365
transform 1 0 103264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_670
timestamp 1698431365
transform 1 0 111104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_671
timestamp 1698431365
transform 1 0 118944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_672
timestamp 1698431365
transform 1 0 126784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_673
timestamp 1698431365
transform 1 0 134624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_674
timestamp 1698431365
transform 1 0 142464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_675
timestamp 1698431365
transform 1 0 150304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_676
timestamp 1698431365
transform 1 0 158144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_677
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_678
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_679
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_680
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_681
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_682
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_683
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_684
timestamp 1698431365
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_685
timestamp 1698431365
transform 1 0 67984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_686
timestamp 1698431365
transform 1 0 75824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_687
timestamp 1698431365
transform 1 0 83664 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_688
timestamp 1698431365
transform 1 0 91504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_689
timestamp 1698431365
transform 1 0 99344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_690
timestamp 1698431365
transform 1 0 107184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_691
timestamp 1698431365
transform 1 0 115024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_692
timestamp 1698431365
transform 1 0 122864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_693
timestamp 1698431365
transform 1 0 130704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_694
timestamp 1698431365
transform 1 0 138544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_695
timestamp 1698431365
transform 1 0 146384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_696
timestamp 1698431365
transform 1 0 154224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_697
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_698
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_699
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_700
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_701
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_702
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_703
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_704
timestamp 1698431365
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_705
timestamp 1698431365
transform 1 0 71904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_706
timestamp 1698431365
transform 1 0 79744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_707
timestamp 1698431365
transform 1 0 87584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_708
timestamp 1698431365
transform 1 0 95424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_709
timestamp 1698431365
transform 1 0 103264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_710
timestamp 1698431365
transform 1 0 111104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_711
timestamp 1698431365
transform 1 0 118944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_712
timestamp 1698431365
transform 1 0 126784 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_713
timestamp 1698431365
transform 1 0 134624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_714
timestamp 1698431365
transform 1 0 142464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_715
timestamp 1698431365
transform 1 0 150304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_716
timestamp 1698431365
transform 1 0 158144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_717
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_718
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_719
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_720
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_721
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_722
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_723
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_724
timestamp 1698431365
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_725
timestamp 1698431365
transform 1 0 67984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_726
timestamp 1698431365
transform 1 0 75824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_727
timestamp 1698431365
transform 1 0 83664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_728
timestamp 1698431365
transform 1 0 91504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_729
timestamp 1698431365
transform 1 0 99344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_730
timestamp 1698431365
transform 1 0 107184 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_731
timestamp 1698431365
transform 1 0 115024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_732
timestamp 1698431365
transform 1 0 122864 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_733
timestamp 1698431365
transform 1 0 130704 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_734
timestamp 1698431365
transform 1 0 138544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_735
timestamp 1698431365
transform 1 0 146384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_736
timestamp 1698431365
transform 1 0 154224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_737
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_738
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_739
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_740
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_741
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_742
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_743
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_744
timestamp 1698431365
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_745
timestamp 1698431365
transform 1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_746
timestamp 1698431365
transform 1 0 79744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_747
timestamp 1698431365
transform 1 0 87584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_748
timestamp 1698431365
transform 1 0 95424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_749
timestamp 1698431365
transform 1 0 103264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_750
timestamp 1698431365
transform 1 0 111104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_751
timestamp 1698431365
transform 1 0 118944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_752
timestamp 1698431365
transform 1 0 126784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_753
timestamp 1698431365
transform 1 0 134624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_754
timestamp 1698431365
transform 1 0 142464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_755
timestamp 1698431365
transform 1 0 150304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_756
timestamp 1698431365
transform 1 0 158144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_757
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_758
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_759
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_760
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_761
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_762
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_763
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_764
timestamp 1698431365
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_765
timestamp 1698431365
transform 1 0 67984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_766
timestamp 1698431365
transform 1 0 75824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_767
timestamp 1698431365
transform 1 0 83664 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_768
timestamp 1698431365
transform 1 0 91504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_769
timestamp 1698431365
transform 1 0 99344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_770
timestamp 1698431365
transform 1 0 107184 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_771
timestamp 1698431365
transform 1 0 115024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_772
timestamp 1698431365
transform 1 0 122864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_773
timestamp 1698431365
transform 1 0 130704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_774
timestamp 1698431365
transform 1 0 138544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_775
timestamp 1698431365
transform 1 0 146384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_776
timestamp 1698431365
transform 1 0 154224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_777
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_778
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_779
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_780
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_781
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_782
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_783
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_784
timestamp 1698431365
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_785
timestamp 1698431365
transform 1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_786
timestamp 1698431365
transform 1 0 79744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_787
timestamp 1698431365
transform 1 0 87584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_788
timestamp 1698431365
transform 1 0 95424 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_789
timestamp 1698431365
transform 1 0 103264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_790
timestamp 1698431365
transform 1 0 111104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_791
timestamp 1698431365
transform 1 0 118944 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_792
timestamp 1698431365
transform 1 0 126784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_793
timestamp 1698431365
transform 1 0 134624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_794
timestamp 1698431365
transform 1 0 142464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_795
timestamp 1698431365
transform 1 0 150304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_796
timestamp 1698431365
transform 1 0 158144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_797
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_798
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_799
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_800
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_801
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_802
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_803
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_804
timestamp 1698431365
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_805
timestamp 1698431365
transform 1 0 67984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_806
timestamp 1698431365
transform 1 0 75824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_807
timestamp 1698431365
transform 1 0 83664 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_808
timestamp 1698431365
transform 1 0 91504 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_809
timestamp 1698431365
transform 1 0 99344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_810
timestamp 1698431365
transform 1 0 107184 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_811
timestamp 1698431365
transform 1 0 115024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_812
timestamp 1698431365
transform 1 0 122864 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_813
timestamp 1698431365
transform 1 0 130704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_814
timestamp 1698431365
transform 1 0 138544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_815
timestamp 1698431365
transform 1 0 146384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_816
timestamp 1698431365
transform 1 0 154224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_817
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_818
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_819
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_820
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_821
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_822
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_823
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_824
timestamp 1698431365
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_825
timestamp 1698431365
transform 1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_826
timestamp 1698431365
transform 1 0 79744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_827
timestamp 1698431365
transform 1 0 87584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_828
timestamp 1698431365
transform 1 0 95424 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_829
timestamp 1698431365
transform 1 0 103264 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_830
timestamp 1698431365
transform 1 0 111104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_831
timestamp 1698431365
transform 1 0 118944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_832
timestamp 1698431365
transform 1 0 126784 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_833
timestamp 1698431365
transform 1 0 134624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_834
timestamp 1698431365
transform 1 0 142464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_835
timestamp 1698431365
transform 1 0 150304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_836
timestamp 1698431365
transform 1 0 158144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_837
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_838
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_839
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_840
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_841
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_842
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_843
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_844
timestamp 1698431365
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_845
timestamp 1698431365
transform 1 0 67984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_846
timestamp 1698431365
transform 1 0 75824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_847
timestamp 1698431365
transform 1 0 83664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_848
timestamp 1698431365
transform 1 0 91504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_849
timestamp 1698431365
transform 1 0 99344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_850
timestamp 1698431365
transform 1 0 107184 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_851
timestamp 1698431365
transform 1 0 115024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_852
timestamp 1698431365
transform 1 0 122864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_853
timestamp 1698431365
transform 1 0 130704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_854
timestamp 1698431365
transform 1 0 138544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_855
timestamp 1698431365
transform 1 0 146384 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_856
timestamp 1698431365
transform 1 0 154224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_857
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_858
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_859
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_860
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_861
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_862
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_863
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_864
timestamp 1698431365
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_865
timestamp 1698431365
transform 1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_866
timestamp 1698431365
transform 1 0 79744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_867
timestamp 1698431365
transform 1 0 87584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_868
timestamp 1698431365
transform 1 0 95424 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_869
timestamp 1698431365
transform 1 0 103264 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_870
timestamp 1698431365
transform 1 0 111104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_871
timestamp 1698431365
transform 1 0 118944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_872
timestamp 1698431365
transform 1 0 126784 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_873
timestamp 1698431365
transform 1 0 134624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_874
timestamp 1698431365
transform 1 0 142464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_875
timestamp 1698431365
transform 1 0 150304 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_876
timestamp 1698431365
transform 1 0 158144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_877
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_878
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_879
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_880
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_881
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_882
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_883
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_884
timestamp 1698431365
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_885
timestamp 1698431365
transform 1 0 67984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_886
timestamp 1698431365
transform 1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_887
timestamp 1698431365
transform 1 0 83664 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_888
timestamp 1698431365
transform 1 0 91504 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_889
timestamp 1698431365
transform 1 0 99344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_890
timestamp 1698431365
transform 1 0 107184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_891
timestamp 1698431365
transform 1 0 115024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_892
timestamp 1698431365
transform 1 0 122864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_893
timestamp 1698431365
transform 1 0 130704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_894
timestamp 1698431365
transform 1 0 138544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_895
timestamp 1698431365
transform 1 0 146384 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_896
timestamp 1698431365
transform 1 0 154224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_897
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_898
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_899
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_900
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_901
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_902
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_903
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_904
timestamp 1698431365
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_905
timestamp 1698431365
transform 1 0 71904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_906
timestamp 1698431365
transform 1 0 79744 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_907
timestamp 1698431365
transform 1 0 87584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_908
timestamp 1698431365
transform 1 0 95424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_909
timestamp 1698431365
transform 1 0 103264 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_910
timestamp 1698431365
transform 1 0 111104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_911
timestamp 1698431365
transform 1 0 118944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_912
timestamp 1698431365
transform 1 0 126784 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_913
timestamp 1698431365
transform 1 0 134624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_914
timestamp 1698431365
transform 1 0 142464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_915
timestamp 1698431365
transform 1 0 150304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_916
timestamp 1698431365
transform 1 0 158144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_917
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_918
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_919
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_920
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_921
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_922
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_923
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_924
timestamp 1698431365
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_925
timestamp 1698431365
transform 1 0 67984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_926
timestamp 1698431365
transform 1 0 75824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_927
timestamp 1698431365
transform 1 0 83664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_928
timestamp 1698431365
transform 1 0 91504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_929
timestamp 1698431365
transform 1 0 99344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_930
timestamp 1698431365
transform 1 0 107184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_931
timestamp 1698431365
transform 1 0 115024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_932
timestamp 1698431365
transform 1 0 122864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_933
timestamp 1698431365
transform 1 0 130704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_934
timestamp 1698431365
transform 1 0 138544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_935
timestamp 1698431365
transform 1 0 146384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_936
timestamp 1698431365
transform 1 0 154224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_937
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_938
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_939
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_940
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_941
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_942
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_943
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_944
timestamp 1698431365
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_945
timestamp 1698431365
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_946
timestamp 1698431365
transform 1 0 79744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_947
timestamp 1698431365
transform 1 0 87584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_948
timestamp 1698431365
transform 1 0 95424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_949
timestamp 1698431365
transform 1 0 103264 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_950
timestamp 1698431365
transform 1 0 111104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_951
timestamp 1698431365
transform 1 0 118944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_952
timestamp 1698431365
transform 1 0 126784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_953
timestamp 1698431365
transform 1 0 134624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_954
timestamp 1698431365
transform 1 0 142464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_955
timestamp 1698431365
transform 1 0 150304 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_956
timestamp 1698431365
transform 1 0 158144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_957
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_958
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_959
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_960
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_961
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_962
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_963
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_964
timestamp 1698431365
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_965
timestamp 1698431365
transform 1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_966
timestamp 1698431365
transform 1 0 75824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_967
timestamp 1698431365
transform 1 0 83664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_968
timestamp 1698431365
transform 1 0 91504 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_969
timestamp 1698431365
transform 1 0 99344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_970
timestamp 1698431365
transform 1 0 107184 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_971
timestamp 1698431365
transform 1 0 115024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_972
timestamp 1698431365
transform 1 0 122864 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_973
timestamp 1698431365
transform 1 0 130704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_974
timestamp 1698431365
transform 1 0 138544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_975
timestamp 1698431365
transform 1 0 146384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_976
timestamp 1698431365
transform 1 0 154224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_977
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_978
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_979
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_980
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_981
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_982
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_983
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_984
timestamp 1698431365
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_985
timestamp 1698431365
transform 1 0 71904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_986
timestamp 1698431365
transform 1 0 79744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_987
timestamp 1698431365
transform 1 0 87584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_988
timestamp 1698431365
transform 1 0 95424 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_989
timestamp 1698431365
transform 1 0 103264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_990
timestamp 1698431365
transform 1 0 111104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_991
timestamp 1698431365
transform 1 0 118944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_992
timestamp 1698431365
transform 1 0 126784 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_993
timestamp 1698431365
transform 1 0 134624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_994
timestamp 1698431365
transform 1 0 142464 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_995
timestamp 1698431365
transform 1 0 150304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_996
timestamp 1698431365
transform 1 0 158144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_997
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_998
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_999
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1000
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1001
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1002
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1003
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1004
timestamp 1698431365
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1005
timestamp 1698431365
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1006
timestamp 1698431365
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1007
timestamp 1698431365
transform 1 0 83664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1008
timestamp 1698431365
transform 1 0 91504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1009
timestamp 1698431365
transform 1 0 99344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1010
timestamp 1698431365
transform 1 0 107184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1011
timestamp 1698431365
transform 1 0 115024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1012
timestamp 1698431365
transform 1 0 122864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1013
timestamp 1698431365
transform 1 0 130704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1014
timestamp 1698431365
transform 1 0 138544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1015
timestamp 1698431365
transform 1 0 146384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1016
timestamp 1698431365
transform 1 0 154224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1017
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1018
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1019
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1020
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1021
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1022
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1023
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1024
timestamp 1698431365
transform 1 0 64064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1025
timestamp 1698431365
transform 1 0 71904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1026
timestamp 1698431365
transform 1 0 79744 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1027
timestamp 1698431365
transform 1 0 87584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1028
timestamp 1698431365
transform 1 0 95424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1029
timestamp 1698431365
transform 1 0 103264 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1030
timestamp 1698431365
transform 1 0 111104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1031
timestamp 1698431365
transform 1 0 118944 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1032
timestamp 1698431365
transform 1 0 126784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1033
timestamp 1698431365
transform 1 0 134624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1034
timestamp 1698431365
transform 1 0 142464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1035
timestamp 1698431365
transform 1 0 150304 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1036
timestamp 1698431365
transform 1 0 158144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1037
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1038
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1039
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1040
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1041
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1042
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1043
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1044
timestamp 1698431365
transform 1 0 60144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1045
timestamp 1698431365
transform 1 0 67984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1046
timestamp 1698431365
transform 1 0 75824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1047
timestamp 1698431365
transform 1 0 83664 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1048
timestamp 1698431365
transform 1 0 91504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1049
timestamp 1698431365
transform 1 0 99344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1050
timestamp 1698431365
transform 1 0 107184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1051
timestamp 1698431365
transform 1 0 115024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1052
timestamp 1698431365
transform 1 0 122864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1053
timestamp 1698431365
transform 1 0 130704 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1054
timestamp 1698431365
transform 1 0 138544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1055
timestamp 1698431365
transform 1 0 146384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1056
timestamp 1698431365
transform 1 0 154224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1057
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1058
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1059
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1060
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1061
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1062
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1063
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1064
timestamp 1698431365
transform 1 0 64064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1065
timestamp 1698431365
transform 1 0 71904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1066
timestamp 1698431365
transform 1 0 79744 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1067
timestamp 1698431365
transform 1 0 87584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1068
timestamp 1698431365
transform 1 0 95424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1069
timestamp 1698431365
transform 1 0 103264 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1070
timestamp 1698431365
transform 1 0 111104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1071
timestamp 1698431365
transform 1 0 118944 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1072
timestamp 1698431365
transform 1 0 126784 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1073
timestamp 1698431365
transform 1 0 134624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1074
timestamp 1698431365
transform 1 0 142464 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1075
timestamp 1698431365
transform 1 0 150304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1076
timestamp 1698431365
transform 1 0 158144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1077
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1078
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1079
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1080
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1081
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1082
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1083
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1084
timestamp 1698431365
transform 1 0 60144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1085
timestamp 1698431365
transform 1 0 67984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1086
timestamp 1698431365
transform 1 0 75824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1087
timestamp 1698431365
transform 1 0 83664 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1088
timestamp 1698431365
transform 1 0 91504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1089
timestamp 1698431365
transform 1 0 99344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1090
timestamp 1698431365
transform 1 0 107184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1091
timestamp 1698431365
transform 1 0 115024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1092
timestamp 1698431365
transform 1 0 122864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1093
timestamp 1698431365
transform 1 0 130704 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1094
timestamp 1698431365
transform 1 0 138544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1095
timestamp 1698431365
transform 1 0 146384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1096
timestamp 1698431365
transform 1 0 154224 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1097
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1098
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1099
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1100
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1101
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1102
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1103
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1104
timestamp 1698431365
transform 1 0 64064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1105
timestamp 1698431365
transform 1 0 71904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1106
timestamp 1698431365
transform 1 0 79744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1107
timestamp 1698431365
transform 1 0 87584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1108
timestamp 1698431365
transform 1 0 95424 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1109
timestamp 1698431365
transform 1 0 103264 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1110
timestamp 1698431365
transform 1 0 111104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1111
timestamp 1698431365
transform 1 0 118944 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1112
timestamp 1698431365
transform 1 0 126784 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1113
timestamp 1698431365
transform 1 0 134624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1114
timestamp 1698431365
transform 1 0 142464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1115
timestamp 1698431365
transform 1 0 150304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1116
timestamp 1698431365
transform 1 0 158144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1117
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1118
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1119
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1120
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1121
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1122
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1123
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1124
timestamp 1698431365
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1125
timestamp 1698431365
transform 1 0 67984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1126
timestamp 1698431365
transform 1 0 75824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1127
timestamp 1698431365
transform 1 0 83664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1128
timestamp 1698431365
transform 1 0 91504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1129
timestamp 1698431365
transform 1 0 99344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1130
timestamp 1698431365
transform 1 0 107184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1131
timestamp 1698431365
transform 1 0 115024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1132
timestamp 1698431365
transform 1 0 122864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1133
timestamp 1698431365
transform 1 0 130704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1134
timestamp 1698431365
transform 1 0 138544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1135
timestamp 1698431365
transform 1 0 146384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1136
timestamp 1698431365
transform 1 0 154224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1137
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1138
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1139
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1140
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1141
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1142
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1143
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1144
timestamp 1698431365
transform 1 0 64064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1145
timestamp 1698431365
transform 1 0 71904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1146
timestamp 1698431365
transform 1 0 79744 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1147
timestamp 1698431365
transform 1 0 87584 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1148
timestamp 1698431365
transform 1 0 95424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1149
timestamp 1698431365
transform 1 0 103264 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1150
timestamp 1698431365
transform 1 0 111104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1151
timestamp 1698431365
transform 1 0 118944 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1152
timestamp 1698431365
transform 1 0 126784 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1153
timestamp 1698431365
transform 1 0 134624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1154
timestamp 1698431365
transform 1 0 142464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1155
timestamp 1698431365
transform 1 0 150304 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1156
timestamp 1698431365
transform 1 0 158144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1157
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1158
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1159
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1160
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1161
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1162
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1163
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1164
timestamp 1698431365
transform 1 0 60144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1165
timestamp 1698431365
transform 1 0 67984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1166
timestamp 1698431365
transform 1 0 75824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1167
timestamp 1698431365
transform 1 0 83664 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1168
timestamp 1698431365
transform 1 0 91504 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1169
timestamp 1698431365
transform 1 0 99344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1170
timestamp 1698431365
transform 1 0 107184 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1171
timestamp 1698431365
transform 1 0 115024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1172
timestamp 1698431365
transform 1 0 122864 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1173
timestamp 1698431365
transform 1 0 130704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1174
timestamp 1698431365
transform 1 0 138544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1175
timestamp 1698431365
transform 1 0 146384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1176
timestamp 1698431365
transform 1 0 154224 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1177
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1178
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1179
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1180
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1181
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1182
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1183
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1184
timestamp 1698431365
transform 1 0 64064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1185
timestamp 1698431365
transform 1 0 71904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1186
timestamp 1698431365
transform 1 0 79744 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1187
timestamp 1698431365
transform 1 0 87584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1188
timestamp 1698431365
transform 1 0 95424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1189
timestamp 1698431365
transform 1 0 103264 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1190
timestamp 1698431365
transform 1 0 111104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1191
timestamp 1698431365
transform 1 0 118944 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1192
timestamp 1698431365
transform 1 0 126784 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1193
timestamp 1698431365
transform 1 0 134624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1194
timestamp 1698431365
transform 1 0 142464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1195
timestamp 1698431365
transform 1 0 150304 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1196
timestamp 1698431365
transform 1 0 158144 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1197
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1198
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1199
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1200
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1201
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1202
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1203
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1204
timestamp 1698431365
transform 1 0 60144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1205
timestamp 1698431365
transform 1 0 67984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1206
timestamp 1698431365
transform 1 0 75824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1207
timestamp 1698431365
transform 1 0 83664 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1208
timestamp 1698431365
transform 1 0 91504 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1209
timestamp 1698431365
transform 1 0 99344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1210
timestamp 1698431365
transform 1 0 107184 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1211
timestamp 1698431365
transform 1 0 115024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1212
timestamp 1698431365
transform 1 0 122864 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1213
timestamp 1698431365
transform 1 0 130704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1214
timestamp 1698431365
transform 1 0 138544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1215
timestamp 1698431365
transform 1 0 146384 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1216
timestamp 1698431365
transform 1 0 154224 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1217
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1218
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1219
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1220
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1221
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1222
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1223
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1224
timestamp 1698431365
transform 1 0 64064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1225
timestamp 1698431365
transform 1 0 71904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1226
timestamp 1698431365
transform 1 0 79744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1227
timestamp 1698431365
transform 1 0 87584 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1228
timestamp 1698431365
transform 1 0 95424 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1229
timestamp 1698431365
transform 1 0 103264 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1230
timestamp 1698431365
transform 1 0 111104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1231
timestamp 1698431365
transform 1 0 118944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1232
timestamp 1698431365
transform 1 0 126784 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1233
timestamp 1698431365
transform 1 0 134624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1234
timestamp 1698431365
transform 1 0 142464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1235
timestamp 1698431365
transform 1 0 150304 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1236
timestamp 1698431365
transform 1 0 158144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1237
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1238
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1239
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1240
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1241
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1242
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1243
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1244
timestamp 1698431365
transform 1 0 60144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1245
timestamp 1698431365
transform 1 0 67984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1246
timestamp 1698431365
transform 1 0 75824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1247
timestamp 1698431365
transform 1 0 83664 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1248
timestamp 1698431365
transform 1 0 91504 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1249
timestamp 1698431365
transform 1 0 99344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1250
timestamp 1698431365
transform 1 0 107184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1251
timestamp 1698431365
transform 1 0 115024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1252
timestamp 1698431365
transform 1 0 122864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1253
timestamp 1698431365
transform 1 0 130704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1254
timestamp 1698431365
transform 1 0 138544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1255
timestamp 1698431365
transform 1 0 146384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1256
timestamp 1698431365
transform 1 0 154224 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1257
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1258
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1259
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1260
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1261
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1262
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1263
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1264
timestamp 1698431365
transform 1 0 64064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1265
timestamp 1698431365
transform 1 0 71904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1266
timestamp 1698431365
transform 1 0 79744 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1267
timestamp 1698431365
transform 1 0 87584 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1268
timestamp 1698431365
transform 1 0 95424 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1269
timestamp 1698431365
transform 1 0 103264 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1270
timestamp 1698431365
transform 1 0 111104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1271
timestamp 1698431365
transform 1 0 118944 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1272
timestamp 1698431365
transform 1 0 126784 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1273
timestamp 1698431365
transform 1 0 134624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1274
timestamp 1698431365
transform 1 0 142464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1275
timestamp 1698431365
transform 1 0 150304 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1276
timestamp 1698431365
transform 1 0 158144 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1277
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1278
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1279
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1280
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1281
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1282
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1283
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1284
timestamp 1698431365
transform 1 0 60144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1285
timestamp 1698431365
transform 1 0 67984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1286
timestamp 1698431365
transform 1 0 75824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1287
timestamp 1698431365
transform 1 0 83664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1288
timestamp 1698431365
transform 1 0 91504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1289
timestamp 1698431365
transform 1 0 99344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1290
timestamp 1698431365
transform 1 0 107184 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1291
timestamp 1698431365
transform 1 0 115024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1292
timestamp 1698431365
transform 1 0 122864 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1293
timestamp 1698431365
transform 1 0 130704 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1294
timestamp 1698431365
transform 1 0 138544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1295
timestamp 1698431365
transform 1 0 146384 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1296
timestamp 1698431365
transform 1 0 154224 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1297
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1298
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1299
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1300
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1301
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1302
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1303
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1304
timestamp 1698431365
transform 1 0 64064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1305
timestamp 1698431365
transform 1 0 71904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1306
timestamp 1698431365
transform 1 0 79744 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1307
timestamp 1698431365
transform 1 0 87584 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1308
timestamp 1698431365
transform 1 0 95424 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1309
timestamp 1698431365
transform 1 0 103264 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1310
timestamp 1698431365
transform 1 0 111104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1311
timestamp 1698431365
transform 1 0 118944 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1312
timestamp 1698431365
transform 1 0 126784 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1313
timestamp 1698431365
transform 1 0 134624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1314
timestamp 1698431365
transform 1 0 142464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1315
timestamp 1698431365
transform 1 0 150304 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1316
timestamp 1698431365
transform 1 0 158144 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1317
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1318
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1319
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1320
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1321
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1322
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1323
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1324
timestamp 1698431365
transform 1 0 60144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1325
timestamp 1698431365
transform 1 0 67984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1326
timestamp 1698431365
transform 1 0 75824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1327
timestamp 1698431365
transform 1 0 83664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1328
timestamp 1698431365
transform 1 0 91504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1329
timestamp 1698431365
transform 1 0 99344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1330
timestamp 1698431365
transform 1 0 107184 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1331
timestamp 1698431365
transform 1 0 115024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1332
timestamp 1698431365
transform 1 0 122864 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1333
timestamp 1698431365
transform 1 0 130704 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1334
timestamp 1698431365
transform 1 0 138544 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1335
timestamp 1698431365
transform 1 0 146384 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1336
timestamp 1698431365
transform 1 0 154224 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1337
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1338
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1339
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1340
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1341
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1342
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1343
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1344
timestamp 1698431365
transform 1 0 64064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1345
timestamp 1698431365
transform 1 0 71904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1346
timestamp 1698431365
transform 1 0 79744 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1347
timestamp 1698431365
transform 1 0 87584 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1348
timestamp 1698431365
transform 1 0 95424 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1349
timestamp 1698431365
transform 1 0 103264 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1350
timestamp 1698431365
transform 1 0 111104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1351
timestamp 1698431365
transform 1 0 118944 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1352
timestamp 1698431365
transform 1 0 126784 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1353
timestamp 1698431365
transform 1 0 134624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1354
timestamp 1698431365
transform 1 0 142464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1355
timestamp 1698431365
transform 1 0 150304 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1356
timestamp 1698431365
transform 1 0 158144 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1357
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1358
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1359
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1360
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1361
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1362
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1363
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1364
timestamp 1698431365
transform 1 0 60144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1365
timestamp 1698431365
transform 1 0 67984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1366
timestamp 1698431365
transform 1 0 75824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1367
timestamp 1698431365
transform 1 0 83664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1368
timestamp 1698431365
transform 1 0 91504 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1369
timestamp 1698431365
transform 1 0 99344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1370
timestamp 1698431365
transform 1 0 107184 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1371
timestamp 1698431365
transform 1 0 115024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1372
timestamp 1698431365
transform 1 0 122864 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1373
timestamp 1698431365
transform 1 0 130704 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1374
timestamp 1698431365
transform 1 0 138544 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1375
timestamp 1698431365
transform 1 0 146384 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1376
timestamp 1698431365
transform 1 0 154224 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1377
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1378
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1379
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1380
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1381
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1382
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1383
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1384
timestamp 1698431365
transform 1 0 64064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1385
timestamp 1698431365
transform 1 0 71904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1386
timestamp 1698431365
transform 1 0 79744 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1387
timestamp 1698431365
transform 1 0 87584 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1388
timestamp 1698431365
transform 1 0 95424 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1389
timestamp 1698431365
transform 1 0 103264 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1390
timestamp 1698431365
transform 1 0 111104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1391
timestamp 1698431365
transform 1 0 118944 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1392
timestamp 1698431365
transform 1 0 126784 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1393
timestamp 1698431365
transform 1 0 134624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1394
timestamp 1698431365
transform 1 0 142464 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1395
timestamp 1698431365
transform 1 0 150304 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1396
timestamp 1698431365
transform 1 0 158144 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1397
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1398
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1399
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1400
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1401
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1402
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1403
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1404
timestamp 1698431365
transform 1 0 60144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1405
timestamp 1698431365
transform 1 0 67984 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1406
timestamp 1698431365
transform 1 0 75824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1407
timestamp 1698431365
transform 1 0 83664 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1408
timestamp 1698431365
transform 1 0 91504 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1409
timestamp 1698431365
transform 1 0 99344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1410
timestamp 1698431365
transform 1 0 107184 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1411
timestamp 1698431365
transform 1 0 115024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1412
timestamp 1698431365
transform 1 0 122864 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1413
timestamp 1698431365
transform 1 0 130704 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1414
timestamp 1698431365
transform 1 0 138544 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1415
timestamp 1698431365
transform 1 0 146384 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1416
timestamp 1698431365
transform 1 0 154224 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1417
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1418
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1419
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1420
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1421
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1422
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1423
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1424
timestamp 1698431365
transform 1 0 64064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1425
timestamp 1698431365
transform 1 0 71904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1426
timestamp 1698431365
transform 1 0 79744 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1427
timestamp 1698431365
transform 1 0 87584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1428
timestamp 1698431365
transform 1 0 95424 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1429
timestamp 1698431365
transform 1 0 103264 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1430
timestamp 1698431365
transform 1 0 111104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1431
timestamp 1698431365
transform 1 0 118944 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1432
timestamp 1698431365
transform 1 0 126784 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1433
timestamp 1698431365
transform 1 0 134624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1434
timestamp 1698431365
transform 1 0 142464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1435
timestamp 1698431365
transform 1 0 150304 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1436
timestamp 1698431365
transform 1 0 158144 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1437
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1438
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1439
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1440
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1441
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1442
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1443
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1444
timestamp 1698431365
transform 1 0 60144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1445
timestamp 1698431365
transform 1 0 67984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1446
timestamp 1698431365
transform 1 0 75824 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1447
timestamp 1698431365
transform 1 0 83664 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1448
timestamp 1698431365
transform 1 0 91504 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1449
timestamp 1698431365
transform 1 0 99344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1450
timestamp 1698431365
transform 1 0 107184 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1451
timestamp 1698431365
transform 1 0 115024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1452
timestamp 1698431365
transform 1 0 122864 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1453
timestamp 1698431365
transform 1 0 130704 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1454
timestamp 1698431365
transform 1 0 138544 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1455
timestamp 1698431365
transform 1 0 146384 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1456
timestamp 1698431365
transform 1 0 154224 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1457
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1458
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1459
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1460
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1461
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1462
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1463
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1464
timestamp 1698431365
transform 1 0 64064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1465
timestamp 1698431365
transform 1 0 71904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1466
timestamp 1698431365
transform 1 0 79744 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1467
timestamp 1698431365
transform 1 0 87584 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1468
timestamp 1698431365
transform 1 0 95424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1469
timestamp 1698431365
transform 1 0 103264 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1470
timestamp 1698431365
transform 1 0 111104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1471
timestamp 1698431365
transform 1 0 118944 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1472
timestamp 1698431365
transform 1 0 126784 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1473
timestamp 1698431365
transform 1 0 134624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1474
timestamp 1698431365
transform 1 0 142464 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1475
timestamp 1698431365
transform 1 0 150304 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1476
timestamp 1698431365
transform 1 0 158144 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1477
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1478
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1479
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1480
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1481
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1482
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1483
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1484
timestamp 1698431365
transform 1 0 60144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1485
timestamp 1698431365
transform 1 0 67984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1486
timestamp 1698431365
transform 1 0 75824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1487
timestamp 1698431365
transform 1 0 83664 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1488
timestamp 1698431365
transform 1 0 91504 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1489
timestamp 1698431365
transform 1 0 99344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1490
timestamp 1698431365
transform 1 0 107184 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1491
timestamp 1698431365
transform 1 0 115024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1492
timestamp 1698431365
transform 1 0 122864 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1493
timestamp 1698431365
transform 1 0 130704 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1494
timestamp 1698431365
transform 1 0 138544 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1495
timestamp 1698431365
transform 1 0 146384 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1496
timestamp 1698431365
transform 1 0 154224 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1497
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1498
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1499
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1500
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1501
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1502
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1503
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1504
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1505
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1506
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1507
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1508
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1509
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1510
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1511
timestamp 1698431365
transform 1 0 58464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1512
timestamp 1698431365
transform 1 0 62272 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1513
timestamp 1698431365
transform 1 0 66080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1514
timestamp 1698431365
transform 1 0 69888 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1515
timestamp 1698431365
transform 1 0 73696 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1516
timestamp 1698431365
transform 1 0 77504 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1517
timestamp 1698431365
transform 1 0 81312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1518
timestamp 1698431365
transform 1 0 85120 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1519
timestamp 1698431365
transform 1 0 88928 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1520
timestamp 1698431365
transform 1 0 92736 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1521
timestamp 1698431365
transform 1 0 96544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1522
timestamp 1698431365
transform 1 0 100352 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1523
timestamp 1698431365
transform 1 0 104160 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1524
timestamp 1698431365
transform 1 0 107968 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1525
timestamp 1698431365
transform 1 0 111776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1526
timestamp 1698431365
transform 1 0 115584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1527
timestamp 1698431365
transform 1 0 119392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1528
timestamp 1698431365
transform 1 0 123200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1529
timestamp 1698431365
transform 1 0 127008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1530
timestamp 1698431365
transform 1 0 130816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1531
timestamp 1698431365
transform 1 0 134624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1532
timestamp 1698431365
transform 1 0 138432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1533
timestamp 1698431365
transform 1 0 142240 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1534
timestamp 1698431365
transform 1 0 146048 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1535
timestamp 1698431365
transform 1 0 149856 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1536
timestamp 1698431365
transform 1 0 153664 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1537
timestamp 1698431365
transform 1 0 157472 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  wire140
timestamp 1698431365
transform -1 0 137536 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_wb_hyperram_141 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_wb_hyperram_142
timestamp 1698431365
transform -1 0 25200 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_wb_hyperram_143
timestamp 1698431365
transform -1 0 36624 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_wb_hyperram_144
timestamp 1698431365
transform -1 0 48048 0 -1 56448
box -86 -86 534 870
<< labels >>
flabel metal2 s 9408 59200 9520 60000 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 123648 59200 123760 60000 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 135072 59200 135184 60000 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 146496 59200 146608 60000 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 20832 59200 20944 60000 0 FreeSans 448 90 0 0 io_in[1]
port 4 nsew signal input
flabel metal2 s 32256 59200 32368 60000 0 FreeSans 448 90 0 0 io_in[2]
port 5 nsew signal input
flabel metal2 s 43680 59200 43792 60000 0 FreeSans 448 90 0 0 io_in[3]
port 6 nsew signal input
flabel metal2 s 55104 59200 55216 60000 0 FreeSans 448 90 0 0 io_in[4]
port 7 nsew signal input
flabel metal2 s 66528 59200 66640 60000 0 FreeSans 448 90 0 0 io_in[5]
port 8 nsew signal input
flabel metal2 s 77952 59200 78064 60000 0 FreeSans 448 90 0 0 io_in[6]
port 9 nsew signal input
flabel metal2 s 89376 59200 89488 60000 0 FreeSans 448 90 0 0 io_in[7]
port 10 nsew signal input
flabel metal2 s 100800 59200 100912 60000 0 FreeSans 448 90 0 0 io_in[8]
port 11 nsew signal input
flabel metal2 s 112224 59200 112336 60000 0 FreeSans 448 90 0 0 io_in[9]
port 12 nsew signal input
flabel metal2 s 13216 59200 13328 60000 0 FreeSans 448 90 0 0 io_oeb[0]
port 13 nsew signal tristate
flabel metal2 s 127456 59200 127568 60000 0 FreeSans 448 90 0 0 io_oeb[10]
port 14 nsew signal tristate
flabel metal2 s 138880 59200 138992 60000 0 FreeSans 448 90 0 0 io_oeb[11]
port 15 nsew signal tristate
flabel metal2 s 150304 59200 150416 60000 0 FreeSans 448 90 0 0 io_oeb[12]
port 16 nsew signal tristate
flabel metal2 s 24640 59200 24752 60000 0 FreeSans 448 90 0 0 io_oeb[1]
port 17 nsew signal tristate
flabel metal2 s 36064 59200 36176 60000 0 FreeSans 448 90 0 0 io_oeb[2]
port 18 nsew signal tristate
flabel metal2 s 47488 59200 47600 60000 0 FreeSans 448 90 0 0 io_oeb[3]
port 19 nsew signal tristate
flabel metal2 s 58912 59200 59024 60000 0 FreeSans 448 90 0 0 io_oeb[4]
port 20 nsew signal tristate
flabel metal2 s 70336 59200 70448 60000 0 FreeSans 448 90 0 0 io_oeb[5]
port 21 nsew signal tristate
flabel metal2 s 81760 59200 81872 60000 0 FreeSans 448 90 0 0 io_oeb[6]
port 22 nsew signal tristate
flabel metal2 s 93184 59200 93296 60000 0 FreeSans 448 90 0 0 io_oeb[7]
port 23 nsew signal tristate
flabel metal2 s 104608 59200 104720 60000 0 FreeSans 448 90 0 0 io_oeb[8]
port 24 nsew signal tristate
flabel metal2 s 116032 59200 116144 60000 0 FreeSans 448 90 0 0 io_oeb[9]
port 25 nsew signal tristate
flabel metal2 s 17024 59200 17136 60000 0 FreeSans 448 90 0 0 io_out[0]
port 26 nsew signal tristate
flabel metal2 s 131264 59200 131376 60000 0 FreeSans 448 90 0 0 io_out[10]
port 27 nsew signal tristate
flabel metal2 s 142688 59200 142800 60000 0 FreeSans 448 90 0 0 io_out[11]
port 28 nsew signal tristate
flabel metal2 s 154112 59200 154224 60000 0 FreeSans 448 90 0 0 io_out[12]
port 29 nsew signal tristate
flabel metal2 s 28448 59200 28560 60000 0 FreeSans 448 90 0 0 io_out[1]
port 30 nsew signal tristate
flabel metal2 s 39872 59200 39984 60000 0 FreeSans 448 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 51296 59200 51408 60000 0 FreeSans 448 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 62720 59200 62832 60000 0 FreeSans 448 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 74144 59200 74256 60000 0 FreeSans 448 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 85568 59200 85680 60000 0 FreeSans 448 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 96992 59200 97104 60000 0 FreeSans 448 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 108416 59200 108528 60000 0 FreeSans 448 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 119840 59200 119952 60000 0 FreeSans 448 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal2 s 5600 59200 5712 60000 0 FreeSans 448 90 0 0 rst_i
port 39 nsew signal input
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 65888 3076 66208 56508 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 96608 3076 96928 56508 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 127328 3076 127648 56508 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 158048 3076 158368 56508 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 81248 3076 81568 56508 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 111968 3076 112288 56508 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 142688 3076 143008 56508 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal2 s 9184 0 9296 800 0 FreeSans 448 90 0 0 wb_clk_i
port 42 nsew signal input
flabel metal2 s 10528 0 10640 800 0 FreeSans 448 90 0 0 wb_rst_i
port 43 nsew signal input
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 wbs_ack_o
port 44 nsew signal tristate
flabel metal2 s 17248 0 17360 800 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 45 nsew signal input
flabel metal2 s 62944 0 63056 800 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 46 nsew signal input
flabel metal2 s 66976 0 67088 800 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 47 nsew signal input
flabel metal2 s 71008 0 71120 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 48 nsew signal input
flabel metal2 s 75040 0 75152 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 49 nsew signal input
flabel metal2 s 79072 0 79184 800 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 50 nsew signal input
flabel metal2 s 83104 0 83216 800 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 51 nsew signal input
flabel metal2 s 87136 0 87248 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 52 nsew signal input
flabel metal2 s 91168 0 91280 800 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 53 nsew signal input
flabel metal2 s 95200 0 95312 800 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 54 nsew signal input
flabel metal2 s 99232 0 99344 800 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 55 nsew signal input
flabel metal2 s 22624 0 22736 800 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 56 nsew signal input
flabel metal2 s 103264 0 103376 800 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 57 nsew signal input
flabel metal2 s 107296 0 107408 800 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 58 nsew signal input
flabel metal2 s 111328 0 111440 800 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 59 nsew signal input
flabel metal2 s 115360 0 115472 800 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 60 nsew signal input
flabel metal2 s 119392 0 119504 800 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 61 nsew signal input
flabel metal2 s 123424 0 123536 800 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 62 nsew signal input
flabel metal2 s 127456 0 127568 800 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 63 nsew signal input
flabel metal2 s 131488 0 131600 800 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 64 nsew signal input
flabel metal2 s 135520 0 135632 800 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 65 nsew signal input
flabel metal2 s 139552 0 139664 800 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 66 nsew signal input
flabel metal2 s 28000 0 28112 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 67 nsew signal input
flabel metal2 s 143584 0 143696 800 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 68 nsew signal input
flabel metal2 s 147616 0 147728 800 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 69 nsew signal input
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 70 nsew signal input
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 71 nsew signal input
flabel metal2 s 42784 0 42896 800 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 72 nsew signal input
flabel metal2 s 46816 0 46928 800 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 73 nsew signal input
flabel metal2 s 50848 0 50960 800 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 74 nsew signal input
flabel metal2 s 54880 0 54992 800 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 75 nsew signal input
flabel metal2 s 58912 0 59024 800 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 76 nsew signal input
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 77 nsew signal input
flabel metal2 s 18592 0 18704 800 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 78 nsew signal input
flabel metal2 s 64288 0 64400 800 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 79 nsew signal input
flabel metal2 s 68320 0 68432 800 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 80 nsew signal input
flabel metal2 s 72352 0 72464 800 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 81 nsew signal input
flabel metal2 s 76384 0 76496 800 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 82 nsew signal input
flabel metal2 s 80416 0 80528 800 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 83 nsew signal input
flabel metal2 s 84448 0 84560 800 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 84 nsew signal input
flabel metal2 s 88480 0 88592 800 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 85 nsew signal input
flabel metal2 s 92512 0 92624 800 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 86 nsew signal input
flabel metal2 s 96544 0 96656 800 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 87 nsew signal input
flabel metal2 s 100576 0 100688 800 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 88 nsew signal input
flabel metal2 s 23968 0 24080 800 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 89 nsew signal input
flabel metal2 s 104608 0 104720 800 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 90 nsew signal input
flabel metal2 s 108640 0 108752 800 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 91 nsew signal input
flabel metal2 s 112672 0 112784 800 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 92 nsew signal input
flabel metal2 s 116704 0 116816 800 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 93 nsew signal input
flabel metal2 s 120736 0 120848 800 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 94 nsew signal input
flabel metal2 s 124768 0 124880 800 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 95 nsew signal input
flabel metal2 s 128800 0 128912 800 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 96 nsew signal input
flabel metal2 s 132832 0 132944 800 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 97 nsew signal input
flabel metal2 s 136864 0 136976 800 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 98 nsew signal input
flabel metal2 s 140896 0 141008 800 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 99 nsew signal input
flabel metal2 s 29344 0 29456 800 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 100 nsew signal input
flabel metal2 s 144928 0 145040 800 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 101 nsew signal input
flabel metal2 s 148960 0 149072 800 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 102 nsew signal input
flabel metal2 s 34720 0 34832 800 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 103 nsew signal input
flabel metal2 s 40096 0 40208 800 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 104 nsew signal input
flabel metal2 s 44128 0 44240 800 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 105 nsew signal input
flabel metal2 s 48160 0 48272 800 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 106 nsew signal input
flabel metal2 s 52192 0 52304 800 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 107 nsew signal input
flabel metal2 s 56224 0 56336 800 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 108 nsew signal input
flabel metal2 s 60256 0 60368 800 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 109 nsew signal input
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 110 nsew signal tristate
flabel metal2 s 65632 0 65744 800 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 111 nsew signal tristate
flabel metal2 s 69664 0 69776 800 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 112 nsew signal tristate
flabel metal2 s 73696 0 73808 800 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 113 nsew signal tristate
flabel metal2 s 77728 0 77840 800 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 114 nsew signal tristate
flabel metal2 s 81760 0 81872 800 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 115 nsew signal tristate
flabel metal2 s 85792 0 85904 800 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 116 nsew signal tristate
flabel metal2 s 89824 0 89936 800 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 117 nsew signal tristate
flabel metal2 s 93856 0 93968 800 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 118 nsew signal tristate
flabel metal2 s 97888 0 98000 800 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 119 nsew signal tristate
flabel metal2 s 101920 0 102032 800 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 120 nsew signal tristate
flabel metal2 s 25312 0 25424 800 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 121 nsew signal tristate
flabel metal2 s 105952 0 106064 800 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 122 nsew signal tristate
flabel metal2 s 109984 0 110096 800 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 123 nsew signal tristate
flabel metal2 s 114016 0 114128 800 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 124 nsew signal tristate
flabel metal2 s 118048 0 118160 800 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 125 nsew signal tristate
flabel metal2 s 122080 0 122192 800 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 126 nsew signal tristate
flabel metal2 s 126112 0 126224 800 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 127 nsew signal tristate
flabel metal2 s 130144 0 130256 800 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 128 nsew signal tristate
flabel metal2 s 134176 0 134288 800 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 129 nsew signal tristate
flabel metal2 s 138208 0 138320 800 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 130 nsew signal tristate
flabel metal2 s 142240 0 142352 800 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 131 nsew signal tristate
flabel metal2 s 30688 0 30800 800 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 132 nsew signal tristate
flabel metal2 s 146272 0 146384 800 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 133 nsew signal tristate
flabel metal2 s 150304 0 150416 800 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 134 nsew signal tristate
flabel metal2 s 36064 0 36176 800 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 135 nsew signal tristate
flabel metal2 s 41440 0 41552 800 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 136 nsew signal tristate
flabel metal2 s 45472 0 45584 800 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 137 nsew signal tristate
flabel metal2 s 49504 0 49616 800 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 138 nsew signal tristate
flabel metal2 s 53536 0 53648 800 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 139 nsew signal tristate
flabel metal2 s 57568 0 57680 800 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 140 nsew signal tristate
flabel metal2 s 61600 0 61712 800 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 141 nsew signal tristate
flabel metal2 s 21280 0 21392 800 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 142 nsew signal input
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 143 nsew signal input
flabel metal2 s 32032 0 32144 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 144 nsew signal input
flabel metal2 s 37408 0 37520 800 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 145 nsew signal input
flabel metal2 s 14560 0 14672 800 0 FreeSans 448 90 0 0 wbs_stb_i
port 146 nsew signal input
flabel metal2 s 15904 0 16016 800 0 FreeSans 448 90 0 0 wbs_we_i
port 147 nsew signal input
rlabel metal1 79968 55664 79968 55664 0 vdd
rlabel metal1 79968 56448 79968 56448 0 vss
rlabel metal2 112392 20468 112392 20468 0 _0000_
rlabel metal2 109032 20496 109032 20496 0 _0001_
rlabel metal2 112840 17584 112840 17584 0 _0002_
rlabel metal2 109816 17976 109816 17976 0 _0003_
rlabel metal3 107408 14280 107408 14280 0 _0004_
rlabel metal2 108248 14616 108248 14616 0 _0005_
rlabel metal2 106344 17136 106344 17136 0 _0006_
rlabel metal2 104776 20496 104776 20496 0 _0007_
rlabel metal2 95368 22680 95368 22680 0 _0008_
rlabel metal2 91112 21504 91112 21504 0 _0009_
rlabel metal2 90496 23128 90496 23128 0 _0010_
rlabel metal2 86408 22344 86408 22344 0 _0011_
rlabel metal2 86072 16856 86072 16856 0 _0012_
rlabel metal2 88200 18088 88200 18088 0 _0013_
rlabel metal2 86296 20496 86296 20496 0 _0014_
rlabel metal2 90888 19656 90888 19656 0 _0015_
rlabel metal2 100856 20048 100856 20048 0 _0016_
rlabel metal2 96600 20272 96600 20272 0 _0017_
rlabel metal2 94920 17976 94920 17976 0 _0018_
rlabel metal2 96488 16352 96488 16352 0 _0019_
rlabel metal2 100296 15008 100296 15008 0 _0020_
rlabel metal2 103768 14224 103768 14224 0 _0021_
rlabel metal2 104216 15792 104216 15792 0 _0022_
rlabel metal2 101920 16072 101920 16072 0 _0023_
rlabel metal3 42728 4200 42728 4200 0 _0024_
rlabel metal2 69496 14168 69496 14168 0 _0025_
rlabel metal2 73192 16464 73192 16464 0 _0026_
rlabel metal2 75880 15624 75880 15624 0 _0027_
rlabel metal2 70392 12600 70392 12600 0 _0028_
rlabel metal2 68376 15736 68376 15736 0 _0029_
rlabel metal2 65240 14728 65240 14728 0 _0030_
rlabel metal2 64008 8400 64008 8400 0 _0031_
rlabel metal2 66248 11312 66248 11312 0 _0032_
rlabel metal2 64736 12376 64736 12376 0 _0033_
rlabel metal2 67816 7616 67816 7616 0 _0034_
rlabel metal2 70280 10192 70280 10192 0 _0035_
rlabel metal2 74648 8288 74648 8288 0 _0036_
rlabel metal2 72968 8680 72968 8680 0 _0037_
rlabel metal2 74536 10696 74536 10696 0 _0038_
rlabel metal2 88760 9352 88760 9352 0 _0039_
rlabel metal2 89432 16240 89432 16240 0 _0040_
rlabel metal2 92456 11200 92456 11200 0 _0041_
rlabel metal3 92848 9128 92848 9128 0 _0042_
rlabel metal2 85904 10808 85904 10808 0 _0043_
rlabel metal2 83384 9352 83384 9352 0 _0044_
rlabel metal2 80360 8344 80360 8344 0 _0045_
rlabel metal3 80080 9912 80080 9912 0 _0046_
rlabel metal2 80920 15456 80920 15456 0 _0047_
rlabel metal2 64848 23016 64848 23016 0 _0048_
rlabel metal2 70504 21728 70504 21728 0 _0049_
rlabel metal3 64232 28056 64232 28056 0 _0050_
rlabel metal2 25816 25816 25816 25816 0 _0051_
rlabel metal3 76888 27160 76888 27160 0 _0052_
rlabel metal2 69720 27608 69720 27608 0 _0053_
rlabel metal2 65464 23464 65464 23464 0 _0054_
rlabel metal2 40824 6272 40824 6272 0 _0055_
rlabel metal2 73080 23072 73080 23072 0 _0056_
rlabel metal2 72856 21112 72856 21112 0 _0057_
rlabel metal2 77224 21224 77224 21224 0 _0058_
rlabel metal2 78680 24416 78680 24416 0 _0059_
rlabel metal2 82936 22512 82936 22512 0 _0060_
rlabel metal2 82600 24024 82600 24024 0 _0061_
rlabel metal2 82152 17360 82152 17360 0 _0062_
rlabel metal2 81144 18816 81144 18816 0 _0063_
rlabel metal2 33992 21392 33992 21392 0 _0064_
rlabel metal3 32312 22456 32312 22456 0 _0065_
rlabel metal2 23352 21168 23352 21168 0 _0066_
rlabel metal2 32088 18200 32088 18200 0 _0067_
rlabel metal2 30240 28504 30240 28504 0 _0068_
rlabel metal2 27608 27300 27608 27300 0 _0069_
rlabel metal2 27832 24304 27832 24304 0 _0070_
rlabel metal3 29904 19880 29904 19880 0 _0071_
rlabel metal2 37128 19600 37128 19600 0 _0072_
rlabel metal2 37240 21392 37240 21392 0 _0073_
rlabel metal2 27496 21728 27496 21728 0 _0074_
rlabel metal2 41776 15400 41776 15400 0 _0075_
rlabel metal2 38136 17696 38136 17696 0 _0076_
rlabel metal3 41328 16184 41328 16184 0 _0077_
rlabel metal2 26264 18872 26264 18872 0 _0078_
rlabel metal2 37352 15736 37352 15736 0 _0079_
rlabel metal2 23352 22736 23352 22736 0 _0080_
rlabel metal2 23240 18088 23240 18088 0 _0081_
rlabel metal2 22792 19656 22792 19656 0 _0082_
rlabel metal3 52304 11480 52304 11480 0 _0083_
rlabel metal2 53592 10360 53592 10360 0 _0084_
rlabel metal2 55048 9184 55048 9184 0 _0085_
rlabel metal2 57624 12320 57624 12320 0 _0086_
rlabel metal2 54936 12600 54936 12600 0 _0087_
rlabel metal2 60872 10192 60872 10192 0 _0088_
rlabel metal2 58744 7616 58744 7616 0 _0089_
rlabel metal2 60648 13104 60648 13104 0 _0090_
rlabel metal3 54320 5096 54320 5096 0 _0091_
rlabel metal2 57176 4144 57176 4144 0 _0092_
rlabel metal2 61096 5544 61096 5544 0 _0093_
rlabel metal3 68376 5880 68376 5880 0 _0094_
rlabel metal2 73752 5208 73752 5208 0 _0095_
rlabel metal3 67760 3640 67760 3640 0 _0096_
rlabel metal3 84560 5768 84560 5768 0 _0097_
rlabel metal2 83720 4480 83720 4480 0 _0098_
rlabel metal2 87304 4760 87304 4760 0 _0099_
rlabel metal2 88704 7560 88704 7560 0 _0100_
rlabel metal3 101304 9912 101304 9912 0 _0101_
rlabel metal3 101248 11480 101248 11480 0 _0102_
rlabel metal2 104888 10584 104888 10584 0 _0103_
rlabel metal2 108360 9632 108360 9632 0 _0104_
rlabel metal2 113120 9128 113120 9128 0 _0105_
rlabel metal3 113232 8344 113232 8344 0 _0106_
rlabel metal2 114520 7560 114520 7560 0 _0107_
rlabel metal2 113680 9576 113680 9576 0 _0108_
rlabel metal2 106344 8008 106344 8008 0 _0109_
rlabel metal2 109760 6664 109760 6664 0 _0110_
rlabel metal3 103936 6664 103936 6664 0 _0111_
rlabel metal2 102648 6664 102648 6664 0 _0112_
rlabel metal3 96600 8176 96600 8176 0 _0113_
rlabel metal2 98168 7784 98168 7784 0 _0114_
rlabel metal2 54152 6944 54152 6944 0 _0115_
rlabel metal3 52360 5992 52360 5992 0 _0116_
rlabel metal2 45640 7056 45640 7056 0 _0117_
rlabel metal2 42840 7784 42840 7784 0 _0118_
rlabel metal2 46088 16128 46088 16128 0 _0119_
rlabel metal2 53032 14728 53032 14728 0 _0120_
rlabel metal2 46760 29232 46760 29232 0 _0121_
rlabel metal2 50904 28672 50904 28672 0 _0122_
rlabel metal2 50008 29456 50008 29456 0 _0123_
rlabel metal2 45192 28952 45192 28952 0 _0124_
rlabel metal2 53536 16968 53536 16968 0 _0125_
rlabel metal2 70616 19712 70616 19712 0 _0126_
rlabel metal3 55720 17752 55720 17752 0 _0127_
rlabel metal2 67144 19432 67144 19432 0 _0128_
rlabel metal2 64456 20720 64456 20720 0 _0129_
rlabel metal2 60648 22736 60648 22736 0 _0130_
rlabel metal2 17752 11816 17752 11816 0 _0131_
rlabel metal2 17864 13720 17864 13720 0 _0132_
rlabel metal2 22400 15512 22400 15512 0 _0133_
rlabel metal2 18200 10920 18200 10920 0 _0134_
rlabel metal3 19712 15512 19712 15512 0 _0135_
rlabel metal2 23016 10360 23016 10360 0 _0136_
rlabel metal2 26376 15540 26376 15540 0 _0137_
rlabel metal3 23688 12376 23688 12376 0 _0138_
rlabel metal2 26264 10192 26264 10192 0 _0139_
rlabel metal2 34328 13104 34328 13104 0 _0140_
rlabel metal2 31864 13552 31864 13552 0 _0141_
rlabel metal3 28840 13608 28840 13608 0 _0142_
rlabel metal2 40712 8624 40712 8624 0 _0143_
rlabel metal2 41832 12600 41832 12600 0 _0144_
rlabel metal2 44520 9464 44520 9464 0 _0145_
rlabel metal2 38248 13328 38248 13328 0 _0146_
rlabel metal2 46984 12600 46984 12600 0 _0147_
rlabel metal2 21784 5040 21784 5040 0 _0148_
rlabel metal2 23688 5880 23688 5880 0 _0149_
rlabel metal2 25088 6776 25088 6776 0 _0150_
rlabel metal2 29456 7672 29456 7672 0 _0151_
rlabel metal3 19264 8120 19264 8120 0 _0152_
rlabel metal2 22904 7392 22904 7392 0 _0153_
rlabel metal2 34328 4984 34328 4984 0 _0154_
rlabel metal2 31976 17696 31976 17696 0 _0155_
rlabel metal2 24080 20552 24080 20552 0 _0156_
rlabel metal2 26096 21784 26096 21784 0 _0157_
rlabel metal2 23464 19600 23464 19600 0 _0158_
rlabel metal2 23800 20832 23800 20832 0 _0159_
rlabel metal3 32032 20104 32032 20104 0 _0160_
rlabel metal3 33656 19992 33656 19992 0 _0161_
rlabel metal2 31080 18312 31080 18312 0 _0162_
rlabel metal2 69160 20832 69160 20832 0 _0163_
rlabel metal3 23464 17640 23464 17640 0 _0164_
rlabel metal2 29792 18424 29792 18424 0 _0165_
rlabel metal2 31752 27440 31752 27440 0 _0166_
rlabel metal2 35728 21560 35728 21560 0 _0167_
rlabel metal2 32200 16856 32200 16856 0 _0168_
rlabel metal3 32648 18424 32648 18424 0 _0169_
rlabel metal3 23688 22344 23688 22344 0 _0170_
rlabel metal2 34216 27888 34216 27888 0 _0171_
rlabel metal2 39480 25312 39480 25312 0 _0172_
rlabel metal2 27832 23016 27832 23016 0 _0173_
rlabel metal2 27160 8512 27160 8512 0 _0174_
rlabel metal2 27608 17472 27608 17472 0 _0175_
rlabel metal2 35784 25648 35784 25648 0 _0176_
rlabel metal3 34944 24920 34944 24920 0 _0177_
rlabel metal2 28280 20440 28280 20440 0 _0178_
rlabel metal2 31416 20832 31416 20832 0 _0179_
rlabel metal2 30128 17080 30128 17080 0 _0180_
rlabel metal2 38472 19544 38472 19544 0 _0181_
rlabel metal3 37128 15288 37128 15288 0 _0182_
rlabel metal2 36008 16184 36008 16184 0 _0183_
rlabel metal2 37352 20832 37352 20832 0 _0184_
rlabel metal2 36680 15512 36680 15512 0 _0185_
rlabel metal3 28560 20328 28560 20328 0 _0186_
rlabel metal3 28560 22232 28560 22232 0 _0187_
rlabel metal3 40320 17528 40320 17528 0 _0188_
rlabel metal2 41944 16072 41944 16072 0 _0189_
rlabel metal3 41720 15624 41720 15624 0 _0190_
rlabel metal2 43400 15960 43400 15960 0 _0191_
rlabel metal2 41384 16184 41384 16184 0 _0192_
rlabel metal3 43008 19096 43008 19096 0 _0193_
rlabel metal2 38248 17192 38248 17192 0 _0194_
rlabel metal3 23744 15400 23744 15400 0 _0195_
rlabel metal2 26040 16184 26040 16184 0 _0196_
rlabel metal3 30184 16072 30184 16072 0 _0197_
rlabel metal2 31192 16688 31192 16688 0 _0198_
rlabel metal2 41384 19656 41384 19656 0 _0199_
rlabel metal2 41216 16072 41216 16072 0 _0200_
rlabel metal2 40824 15848 40824 15848 0 _0201_
rlabel metal3 26488 18480 26488 18480 0 _0202_
rlabel metal2 26712 19208 26712 19208 0 _0203_
rlabel metal2 26600 17584 26600 17584 0 _0204_
rlabel metal2 37240 16072 37240 16072 0 _0205_
rlabel metal2 37016 15568 37016 15568 0 _0206_
rlabel metal2 22792 16128 22792 16128 0 _0207_
rlabel metal2 23800 22568 23800 22568 0 _0208_
rlabel metal2 23408 17640 23408 17640 0 _0209_
rlabel metal2 22792 17864 22792 17864 0 _0210_
rlabel metal2 23128 19600 23128 19600 0 _0211_
rlabel metal2 23800 17752 23800 17752 0 _0212_
rlabel metal2 20328 5992 20328 5992 0 _0213_
rlabel metal2 24472 10528 24472 10528 0 _0214_
rlabel metal2 58408 12712 58408 12712 0 _0215_
rlabel metal2 56672 10808 56672 10808 0 _0216_
rlabel metal2 53256 12152 53256 12152 0 _0217_
rlabel metal2 21448 13440 21448 13440 0 _0218_
rlabel metal2 62440 10976 62440 10976 0 _0219_
rlabel metal2 55608 11032 55608 11032 0 _0220_
rlabel metal2 51912 7728 51912 7728 0 _0221_
rlabel metal3 56280 9016 56280 9016 0 _0222_
rlabel metal2 25592 4200 25592 4200 0 _0223_
rlabel metal2 56504 9688 56504 9688 0 _0224_
rlabel metal2 57288 5600 57288 5600 0 _0225_
rlabel metal2 26712 4592 26712 4592 0 _0226_
rlabel metal2 26152 9856 26152 9856 0 _0227_
rlabel metal2 56840 11816 56840 11816 0 _0228_
rlabel metal2 44072 12096 44072 12096 0 _0229_
rlabel metal2 55272 12936 55272 12936 0 _0230_
rlabel metal4 44632 6944 44632 6944 0 _0231_
rlabel metal2 61320 10080 61320 10080 0 _0232_
rlabel metal2 57400 8400 57400 8400 0 _0233_
rlabel metal2 56952 7840 56952 7840 0 _0234_
rlabel metal2 45192 11648 45192 11648 0 _0235_
rlabel metal2 61096 13160 61096 13160 0 _0236_
rlabel metal2 53480 5768 53480 5768 0 _0237_
rlabel metal3 67536 9016 67536 9016 0 _0238_
rlabel metal2 53816 7616 53816 7616 0 _0239_
rlabel metal2 52808 5376 52808 5376 0 _0240_
rlabel metal3 55104 5992 55104 5992 0 _0241_
rlabel metal2 73248 11928 73248 11928 0 _0242_
rlabel metal2 66584 7448 66584 7448 0 _0243_
rlabel metal2 60592 5320 60592 5320 0 _0244_
rlabel metal2 56896 4424 56896 4424 0 _0245_
rlabel metal2 72968 6720 72968 6720 0 _0246_
rlabel metal2 67704 6104 67704 6104 0 _0247_
rlabel metal2 67368 7336 67368 7336 0 _0248_
rlabel metal2 73192 7840 73192 7840 0 _0249_
rlabel metal2 121912 3976 121912 3976 0 _0250_
rlabel metal3 85848 15288 85848 15288 0 _0251_
rlabel metal2 73640 7336 73640 7336 0 _0252_
rlabel metal2 66584 6944 66584 6944 0 _0253_
rlabel metal2 72520 5320 72520 5320 0 _0254_
rlabel metal2 92176 4984 92176 4984 0 _0255_
rlabel metal3 87192 5880 87192 5880 0 _0256_
rlabel metal2 85848 3752 85848 3752 0 _0257_
rlabel metal2 86744 5824 86744 5824 0 _0258_
rlabel metal2 86408 5936 86408 5936 0 _0259_
rlabel metal2 83608 7056 83608 7056 0 _0260_
rlabel metal2 87192 4592 87192 4592 0 _0261_
rlabel metal2 91000 11088 91000 11088 0 _0262_
rlabel metal2 87528 5880 87528 5880 0 _0263_
rlabel metal2 94696 7896 94696 7896 0 _0264_
rlabel metal2 88872 9688 88872 9688 0 _0265_
rlabel metal2 101304 12096 101304 12096 0 _0266_
rlabel metal2 100632 10696 100632 10696 0 _0267_
rlabel metal3 102200 6552 102200 6552 0 _0268_
rlabel metal2 71344 17752 71344 17752 0 _0269_
rlabel metal3 106904 11256 106904 11256 0 _0270_
rlabel metal2 100408 12264 100408 12264 0 _0271_
rlabel metal2 103544 5768 103544 5768 0 _0272_
rlabel metal2 104664 10304 104664 10304 0 _0273_
rlabel metal2 110936 4480 110936 4480 0 _0274_
rlabel metal2 104888 8960 104888 8960 0 _0275_
rlabel metal2 107800 11760 107800 11760 0 _0276_
rlabel metal2 108136 7784 108136 7784 0 _0277_
rlabel metal2 111496 11144 111496 11144 0 _0278_
rlabel metal2 113288 9576 113288 9576 0 _0279_
rlabel metal2 112896 9016 112896 9016 0 _0280_
rlabel metal2 112504 9632 112504 9632 0 _0281_
rlabel metal3 114072 9240 114072 9240 0 _0282_
rlabel metal2 114912 8120 114912 8120 0 _0283_
rlabel metal3 114744 9128 114744 9128 0 _0284_
rlabel metal2 109480 11816 109480 11816 0 _0285_
rlabel metal2 117544 8288 117544 8288 0 _0286_
rlabel metal2 113736 9856 113736 9856 0 _0287_
rlabel metal2 115976 9464 115976 9464 0 _0288_
rlabel metal2 107576 13272 107576 13272 0 _0289_
rlabel metal3 107856 6104 107856 6104 0 _0290_
rlabel metal2 109368 11760 109368 11760 0 _0291_
rlabel metal2 105224 8904 105224 8904 0 _0292_
rlabel metal2 109704 11704 109704 11704 0 _0293_
rlabel metal2 117320 7336 117320 7336 0 _0294_
rlabel metal2 105000 12824 105000 12824 0 _0295_
rlabel metal2 108136 12040 108136 12040 0 _0296_
rlabel metal3 106848 9128 106848 9128 0 _0297_
rlabel metal2 102872 6104 102872 6104 0 _0298_
rlabel metal2 102536 6496 102536 6496 0 _0299_
rlabel metal2 49392 9240 49392 9240 0 _0300_
rlabel metal2 95592 9128 95592 9128 0 _0301_
rlabel metal3 104384 12040 104384 12040 0 _0302_
rlabel metal3 93576 10472 93576 10472 0 _0303_
rlabel metal2 99064 5544 99064 5544 0 _0304_
rlabel metal2 102312 10136 102312 10136 0 _0305_
rlabel metal2 54488 7784 54488 7784 0 _0306_
rlabel metal2 44016 6552 44016 6552 0 _0307_
rlabel metal2 47208 6776 47208 6776 0 _0308_
rlabel metal2 49560 7896 49560 7896 0 _0309_
rlabel metal2 48328 5320 48328 5320 0 _0310_
rlabel metal2 45864 6888 45864 6888 0 _0311_
rlabel metal2 45416 6608 45416 6608 0 _0312_
rlabel metal2 47432 17080 47432 17080 0 _0313_
rlabel metal2 45528 8792 45528 8792 0 _0314_
rlabel metal3 44744 8232 44744 8232 0 _0315_
rlabel metal2 48720 16744 48720 16744 0 _0316_
rlabel metal3 50008 27832 50008 27832 0 _0317_
rlabel metal2 45976 27328 45976 27328 0 _0318_
rlabel metal2 46200 27328 46200 27328 0 _0319_
rlabel metal2 49896 16296 49896 16296 0 _0320_
rlabel metal2 49560 16464 49560 16464 0 _0321_
rlabel metal2 55440 21560 55440 21560 0 _0322_
rlabel metal3 53592 15176 53592 15176 0 _0323_
rlabel metal2 53144 16184 53144 16184 0 _0324_
rlabel metal3 52360 23576 52360 23576 0 _0325_
rlabel metal2 62440 19096 62440 19096 0 _0326_
rlabel metal2 56840 19768 56840 19768 0 _0327_
rlabel metal2 57176 21952 57176 21952 0 _0328_
rlabel metal2 47208 24024 47208 24024 0 _0329_
rlabel metal2 47768 22344 47768 22344 0 _0330_
rlabel metal2 43736 22512 43736 22512 0 _0331_
rlabel metal3 56448 26264 56448 26264 0 _0332_
rlabel metal3 58296 24696 58296 24696 0 _0333_
rlabel metal2 54264 24304 54264 24304 0 _0334_
rlabel metal2 53592 24304 53592 24304 0 _0335_
rlabel metal2 51912 26096 51912 26096 0 _0336_
rlabel metal2 56840 25648 56840 25648 0 _0337_
rlabel metal2 53144 25816 53144 25816 0 _0338_
rlabel metal2 49896 28560 49896 28560 0 _0339_
rlabel metal2 46480 25256 46480 25256 0 _0340_
rlabel metal3 47320 26936 47320 26936 0 _0341_
rlabel metal2 49336 18256 49336 18256 0 _0342_
rlabel metal2 49504 18648 49504 18648 0 _0343_
rlabel metal2 43232 24920 43232 24920 0 _0344_
rlabel metal3 39872 26376 39872 26376 0 _0345_
rlabel metal3 44464 26264 44464 26264 0 _0346_
rlabel metal2 44856 25872 44856 25872 0 _0347_
rlabel metal2 48104 25648 48104 25648 0 _0348_
rlabel metal3 49112 28504 49112 28504 0 _0349_
rlabel metal3 50148 17528 50148 17528 0 _0350_
rlabel metal2 49448 25928 49448 25928 0 _0351_
rlabel metal2 49224 25984 49224 25984 0 _0352_
rlabel metal3 51520 27272 51520 27272 0 _0353_
rlabel metal2 50120 27104 50120 27104 0 _0354_
rlabel metal2 48888 25760 48888 25760 0 _0355_
rlabel metal3 47152 25592 47152 25592 0 _0356_
rlabel metal2 44744 28280 44744 28280 0 _0357_
rlabel metal2 64120 20608 64120 20608 0 _0358_
rlabel metal2 45192 14056 45192 14056 0 _0359_
rlabel metal2 51240 17304 51240 17304 0 _0360_
rlabel metal2 51016 18144 51016 18144 0 _0361_
rlabel metal2 43960 22176 43960 22176 0 _0362_
rlabel metal2 44688 23352 44688 23352 0 _0363_
rlabel metal2 46872 21504 46872 21504 0 _0364_
rlabel metal2 55160 22680 55160 22680 0 _0365_
rlabel metal4 50120 24024 50120 24024 0 _0366_
rlabel metal2 50904 25816 50904 25816 0 _0367_
rlabel metal2 51016 23240 51016 23240 0 _0368_
rlabel metal2 52640 19320 52640 19320 0 _0369_
rlabel metal2 68600 23576 68600 23576 0 _0370_
rlabel metal2 54040 22344 54040 22344 0 _0371_
rlabel metal2 47432 20944 47432 20944 0 _0372_
rlabel metal2 62552 19376 62552 19376 0 _0373_
rlabel metal2 52472 18760 52472 18760 0 _0374_
rlabel metal2 48440 18984 48440 18984 0 _0375_
rlabel metal3 39704 25368 39704 25368 0 _0376_
rlabel metal2 41496 26488 41496 26488 0 _0377_
rlabel metal2 40376 27328 40376 27328 0 _0378_
rlabel metal2 39032 26208 39032 26208 0 _0379_
rlabel metal3 40488 26936 40488 26936 0 _0380_
rlabel metal2 40712 26544 40712 26544 0 _0381_
rlabel metal2 44744 25816 44744 25816 0 _0382_
rlabel metal3 45752 24920 45752 24920 0 _0383_
rlabel metal2 43400 23464 43400 23464 0 _0384_
rlabel metal2 46088 23744 46088 23744 0 _0385_
rlabel metal2 45192 23576 45192 23576 0 _0386_
rlabel metal3 47040 23912 47040 23912 0 _0387_
rlabel metal2 46984 24416 46984 24416 0 _0388_
rlabel metal2 46536 24304 46536 24304 0 _0389_
rlabel metal3 49784 18984 49784 18984 0 _0390_
rlabel metal2 41720 23520 41720 23520 0 _0391_
rlabel metal2 47656 17808 47656 17808 0 _0392_
rlabel metal3 47152 18424 47152 18424 0 _0393_
rlabel metal2 48216 18536 48216 18536 0 _0394_
rlabel metal2 49224 21896 49224 21896 0 _0395_
rlabel metal2 49784 29008 49784 29008 0 _0396_
rlabel metal2 62888 18088 62888 18088 0 _0397_
rlabel metal2 70168 19320 70168 19320 0 _0398_
rlabel metal3 53984 19208 53984 19208 0 _0399_
rlabel metal3 39228 26264 39228 26264 0 _0400_
rlabel metal2 40040 26544 40040 26544 0 _0401_
rlabel metal3 40824 25480 40824 25480 0 _0402_
rlabel metal2 40040 25592 40040 25592 0 _0403_
rlabel metal3 40600 25256 40600 25256 0 _0404_
rlabel metal2 41160 24976 41160 24976 0 _0405_
rlabel metal2 43176 21784 43176 21784 0 _0406_
rlabel metal2 43400 22176 43400 22176 0 _0407_
rlabel metal2 51464 22624 51464 22624 0 _0408_
rlabel metal2 50904 24248 50904 24248 0 _0409_
rlabel metal2 50680 21392 50680 21392 0 _0410_
rlabel metal2 52808 20328 52808 20328 0 _0411_
rlabel metal2 51800 21504 51800 21504 0 _0412_
rlabel metal2 53088 21784 53088 21784 0 _0413_
rlabel metal3 46648 21560 46648 21560 0 _0414_
rlabel metal2 52808 21644 52808 21644 0 _0415_
rlabel metal2 52360 21392 52360 21392 0 _0416_
rlabel metal2 52640 20216 52640 20216 0 _0417_
rlabel metal2 38808 13104 38808 13104 0 _0418_
rlabel metal2 51352 19264 51352 19264 0 _0419_
rlabel metal2 55160 19320 55160 19320 0 _0420_
rlabel metal3 55552 19096 55552 19096 0 _0421_
rlabel metal2 50008 16968 50008 16968 0 _0422_
rlabel metal2 60088 19376 60088 19376 0 _0423_
rlabel metal2 51576 20496 51576 20496 0 _0424_
rlabel metal3 52416 18312 52416 18312 0 _0425_
rlabel metal2 37576 25872 37576 25872 0 _0426_
rlabel metal2 34440 27384 34440 27384 0 _0427_
rlabel metal3 36512 26264 36512 26264 0 _0428_
rlabel metal2 37408 25256 37408 25256 0 _0429_
rlabel metal2 36792 25032 36792 25032 0 _0430_
rlabel metal2 38528 26040 38528 26040 0 _0431_
rlabel metal2 39032 25368 39032 25368 0 _0432_
rlabel metal3 42952 23688 42952 23688 0 _0433_
rlabel metal2 43400 18816 43400 18816 0 _0434_
rlabel metal2 42840 21168 42840 21168 0 _0435_
rlabel metal2 42728 22512 42728 22512 0 _0436_
rlabel metal2 47656 21728 47656 21728 0 _0437_
rlabel metal2 47992 22512 47992 22512 0 _0438_
rlabel metal2 46760 21952 46760 21952 0 _0439_
rlabel metal3 48748 20552 48748 20552 0 _0440_
rlabel metal2 52584 20832 52584 20832 0 _0441_
rlabel metal2 57512 19936 57512 19936 0 _0442_
rlabel metal2 64400 20216 64400 20216 0 _0443_
rlabel metal3 60032 20776 60032 20776 0 _0444_
rlabel metal3 60256 20888 60256 20888 0 _0445_
rlabel metal2 59864 21000 59864 21000 0 _0446_
rlabel metal2 59080 22120 59080 22120 0 _0447_
rlabel metal2 42280 18256 42280 18256 0 _0448_
rlabel metal2 44296 20440 44296 20440 0 _0449_
rlabel metal2 46480 21000 46480 21000 0 _0450_
rlabel metal2 63672 21280 63672 21280 0 _0451_
rlabel metal2 34664 25984 34664 25984 0 _0452_
rlabel metal2 31080 25816 31080 25816 0 _0453_
rlabel metal3 33432 25480 33432 25480 0 _0454_
rlabel metal3 35784 25704 35784 25704 0 _0455_
rlabel metal2 35784 26208 35784 26208 0 _0456_
rlabel metal2 35616 25704 35616 25704 0 _0457_
rlabel metal2 49504 29064 49504 29064 0 _0458_
rlabel metal2 63336 20888 63336 20888 0 _0459_
rlabel metal2 59640 22008 59640 22008 0 _0460_
rlabel metal2 60088 23072 60088 23072 0 _0461_
rlabel metal2 60872 22568 60872 22568 0 _0462_
rlabel metal3 33712 24696 33712 24696 0 _0463_
rlabel metal2 35448 24528 35448 24528 0 _0464_
rlabel metal2 43848 24248 43848 24248 0 _0465_
rlabel metal2 40824 21224 40824 21224 0 _0466_
rlabel metal3 41608 23240 41608 23240 0 _0467_
rlabel metal3 42392 23296 42392 23296 0 _0468_
rlabel metal2 42616 23408 42616 23408 0 _0469_
rlabel metal3 46536 23856 46536 23856 0 _0470_
rlabel metal2 60424 22680 60424 22680 0 _0471_
rlabel metal2 30744 4760 30744 4760 0 _0472_
rlabel metal2 34776 6384 34776 6384 0 _0473_
rlabel metal2 22120 11088 22120 11088 0 _0474_
rlabel metal3 21560 15288 21560 15288 0 _0475_
rlabel metal3 21392 12152 21392 12152 0 _0476_
rlabel metal3 19488 12040 19488 12040 0 _0477_
rlabel metal3 24360 10584 24360 10584 0 _0478_
rlabel metal2 25816 12320 25816 12320 0 _0479_
rlabel metal2 24416 11144 24416 11144 0 _0480_
rlabel metal2 20216 13384 20216 13384 0 _0481_
rlabel metal3 22008 12264 22008 12264 0 _0482_
rlabel metal2 22008 13888 22008 13888 0 _0483_
rlabel metal2 21336 11536 21336 11536 0 _0484_
rlabel metal2 21224 13832 21224 13832 0 _0485_
rlabel metal2 32200 8736 32200 8736 0 _0486_
rlabel metal2 27832 8736 27832 8736 0 _0487_
rlabel metal2 24696 11256 24696 11256 0 _0488_
rlabel metal3 26208 10360 26208 10360 0 _0489_
rlabel metal3 24752 10360 24752 10360 0 _0490_
rlabel metal2 27272 12768 27272 12768 0 _0491_
rlabel metal2 32032 12936 32032 12936 0 _0492_
rlabel metal3 24976 12152 24976 12152 0 _0493_
rlabel metal2 27608 10360 27608 10360 0 _0494_
rlabel metal2 37800 9016 37800 9016 0 _0495_
rlabel metal2 31416 13328 31416 13328 0 _0496_
rlabel metal2 32872 12544 32872 12544 0 _0497_
rlabel metal2 35112 13552 35112 13552 0 _0498_
rlabel metal2 32424 13160 32424 13160 0 _0499_
rlabel metal2 29512 12656 29512 12656 0 _0500_
rlabel metal3 40936 10696 40936 10696 0 _0501_
rlabel metal2 45024 10024 45024 10024 0 _0502_
rlabel metal2 40264 10416 40264 10416 0 _0503_
rlabel metal3 40040 10584 40040 10584 0 _0504_
rlabel metal2 42952 11760 42952 11760 0 _0505_
rlabel metal3 45024 9912 45024 9912 0 _0506_
rlabel metal2 37800 12656 37800 12656 0 _0507_
rlabel metal2 45472 11928 45472 11928 0 _0508_
rlabel metal2 28392 6944 28392 6944 0 _0509_
rlabel metal2 26264 7896 26264 7896 0 _0510_
rlabel metal2 22568 8288 22568 8288 0 _0511_
rlabel metal2 21672 6048 21672 6048 0 _0512_
rlabel metal3 19208 5096 19208 5096 0 _0513_
rlabel metal2 25928 7336 25928 7336 0 _0514_
rlabel metal2 24192 7560 24192 7560 0 _0515_
rlabel metal2 23912 5992 23912 5992 0 _0516_
rlabel metal2 25256 8232 25256 8232 0 _0517_
rlabel metal2 25368 6328 25368 6328 0 _0518_
rlabel metal3 28840 7448 28840 7448 0 _0519_
rlabel metal2 20664 7952 20664 7952 0 _0520_
rlabel metal2 20776 8344 20776 8344 0 _0521_
rlabel metal2 23128 7840 23128 7840 0 _0522_
rlabel metal3 22792 7448 22792 7448 0 _0523_
rlabel metal2 46536 17304 46536 17304 0 _0524_
rlabel metal2 73304 18088 73304 18088 0 _0525_
rlabel metal2 72968 18144 72968 18144 0 _0526_
rlabel metal2 45416 18704 45416 18704 0 _0527_
rlabel metal3 54768 27832 54768 27832 0 _0528_
rlabel metal2 49448 28224 49448 28224 0 _0529_
rlabel metal2 57176 25592 57176 25592 0 _0530_
rlabel metal2 57176 25200 57176 25200 0 _0531_
rlabel metal2 59528 28392 59528 28392 0 _0532_
rlabel metal2 28504 55104 28504 55104 0 _0533_
rlabel metal2 55888 25592 55888 25592 0 _0534_
rlabel metal2 59416 26572 59416 26572 0 _0535_
rlabel metal2 60536 25872 60536 25872 0 _0536_
rlabel metal2 68040 22400 68040 22400 0 _0537_
rlabel metal2 59976 28616 59976 28616 0 _0538_
rlabel metal3 47992 21448 47992 21448 0 _0539_
rlabel metal3 54208 27048 54208 27048 0 _0540_
rlabel metal2 57176 27384 57176 27384 0 _0541_
rlabel metal3 58576 28392 58576 28392 0 _0542_
rlabel metal3 61656 26824 61656 26824 0 _0543_
rlabel metal2 48664 27272 48664 27272 0 _0544_
rlabel metal3 28168 2520 28168 2520 0 _0545_
rlabel metal2 41160 6944 41160 6944 0 _0546_
rlabel metal2 141512 4592 141512 4592 0 _0547_
rlabel metal3 140504 4312 140504 4312 0 _0548_
rlabel metal2 141400 4704 141400 4704 0 _0549_
rlabel metal2 122920 4984 122920 4984 0 _0550_
rlabel metal2 94192 8456 94192 8456 0 _0551_
rlabel via2 94024 7560 94024 7560 0 _0552_
rlabel metal2 94360 5320 94360 5320 0 _0553_
rlabel metal3 48328 13944 48328 13944 0 _0554_
rlabel metal3 43120 5208 43120 5208 0 _0555_
rlabel metal2 48720 11256 48720 11256 0 _0556_
rlabel metal2 48216 7784 48216 7784 0 _0557_
rlabel metal2 15960 6552 15960 6552 0 _0558_
rlabel metal2 39144 9520 39144 9520 0 _0559_
rlabel metal2 93688 5936 93688 5936 0 _0560_
rlabel metal2 94024 5656 94024 5656 0 _0561_
rlabel metal2 91168 16856 91168 16856 0 _0562_
rlabel metal2 95312 4984 95312 4984 0 _0563_
rlabel metal2 69496 3276 69496 3276 0 _0564_
rlabel metal2 38920 6832 38920 6832 0 _0565_
rlabel metal2 26040 8176 26040 8176 0 _0566_
rlabel metal2 43176 13048 43176 13048 0 _0567_
rlabel metal3 37912 5992 37912 5992 0 _0568_
rlabel metal2 38696 5600 38696 5600 0 _0569_
rlabel metal2 66808 5600 66808 5600 0 _0570_
rlabel metal2 64456 5544 64456 5544 0 _0571_
rlabel metal2 65016 6216 65016 6216 0 _0572_
rlabel metal2 41496 5376 41496 5376 0 _0573_
rlabel metal2 39816 6160 39816 6160 0 _0574_
rlabel metal2 38136 10080 38136 10080 0 _0575_
rlabel metal2 45864 9576 45864 9576 0 _0576_
rlabel metal2 34328 9352 34328 9352 0 _0577_
rlabel metal2 39256 8624 39256 8624 0 _0578_
rlabel metal2 72072 16408 72072 16408 0 _0579_
rlabel metal2 38080 5768 38080 5768 0 _0580_
rlabel metal2 50344 5936 50344 5936 0 _0581_
rlabel metal2 50456 4816 50456 4816 0 _0582_
rlabel metal2 70728 3864 70728 3864 0 _0583_
rlabel metal3 64568 4704 64568 4704 0 _0584_
rlabel metal2 24808 8904 24808 8904 0 _0585_
rlabel metal3 29848 6888 29848 6888 0 _0586_
rlabel metal2 33880 8176 33880 8176 0 _0587_
rlabel metal2 38024 10864 38024 10864 0 _0588_
rlabel metal2 65296 18872 65296 18872 0 _0589_
rlabel metal3 76104 2968 76104 2968 0 _0590_
rlabel metal2 89768 21000 89768 21000 0 _0591_
rlabel metal2 90104 12880 90104 12880 0 _0592_
rlabel metal3 41832 10472 41832 10472 0 _0593_
rlabel metal2 39032 6832 39032 6832 0 _0594_
rlabel metal3 40712 7672 40712 7672 0 _0595_
rlabel metal2 39536 5880 39536 5880 0 _0596_
rlabel metal2 40712 10248 40712 10248 0 _0597_
rlabel metal2 40488 10528 40488 10528 0 _0598_
rlabel metal2 33768 7896 33768 7896 0 _0599_
rlabel metal2 80584 1904 80584 1904 0 _0600_
rlabel metal2 36344 10136 36344 10136 0 _0601_
rlabel metal3 30072 6776 30072 6776 0 _0602_
rlabel metal2 30520 9968 30520 9968 0 _0603_
rlabel metal3 44072 12152 44072 12152 0 _0604_
rlabel metal2 91056 21784 91056 21784 0 _0605_
rlabel metal3 32984 10696 32984 10696 0 _0606_
rlabel metal3 30464 12824 30464 12824 0 _0607_
rlabel metal2 30632 12656 30632 12656 0 _0608_
rlabel metal2 30744 12544 30744 12544 0 _0609_
rlabel metal2 25816 8176 25816 8176 0 _0610_
rlabel metal2 91728 7224 91728 7224 0 _0611_
rlabel metal2 31416 9688 31416 9688 0 _0612_
rlabel metal2 29792 12712 29792 12712 0 _0613_
rlabel metal2 30464 17080 30464 17080 0 _0614_
rlabel metal2 88032 7112 88032 7112 0 _0615_
rlabel metal3 34160 9688 34160 9688 0 _0616_
rlabel metal2 35336 10416 35336 10416 0 _0617_
rlabel metal3 40320 11256 40320 11256 0 _0618_
rlabel metal3 47880 12152 47880 12152 0 _0619_
rlabel metal3 45584 12264 45584 12264 0 _0620_
rlabel metal2 41160 11872 41160 11872 0 _0621_
rlabel metal2 43176 10136 43176 10136 0 _0622_
rlabel metal2 46200 11032 46200 11032 0 _0623_
rlabel metal2 46032 10024 46032 10024 0 _0624_
rlabel metal2 48944 13048 48944 13048 0 _0625_
rlabel metal2 49672 12544 49672 12544 0 _0626_
rlabel metal2 74816 3640 74816 3640 0 _0627_
rlabel metal3 71792 15736 71792 15736 0 _0628_
rlabel metal2 77728 4984 77728 4984 0 _0629_
rlabel metal2 75992 16184 75992 16184 0 _0630_
rlabel metal2 77840 17416 77840 17416 0 _0631_
rlabel metal2 78960 22120 78960 22120 0 _0632_
rlabel metal2 82264 7448 82264 7448 0 _0633_
rlabel metal2 80416 16744 80416 16744 0 _0634_
rlabel metal2 81480 8176 81480 8176 0 _0635_
rlabel metal3 78232 15736 78232 15736 0 _0636_
rlabel metal3 82152 15624 82152 15624 0 _0637_
rlabel metal3 84784 8008 84784 8008 0 _0638_
rlabel metal2 109704 8736 109704 8736 0 _0639_
rlabel metal4 85456 17010 85456 17010 0 _0640_
rlabel metal3 102592 17304 102592 17304 0 _0641_
rlabel metal3 111104 10584 111104 10584 0 _0642_
rlabel metal2 109592 4872 109592 4872 0 _0643_
rlabel metal3 98392 14504 98392 14504 0 _0644_
rlabel metal2 98336 12936 98336 12936 0 _0645_
rlabel metal2 122360 4032 122360 4032 0 _0646_
rlabel metal2 109256 5376 109256 5376 0 _0647_
rlabel metal2 103096 10948 103096 10948 0 _0648_
rlabel metal2 112056 7168 112056 7168 0 _0649_
rlabel metal2 108248 11088 108248 11088 0 _0650_
rlabel metal2 105168 13496 105168 13496 0 _0651_
rlabel metal2 121688 5656 121688 5656 0 _0652_
rlabel metal2 117880 5712 117880 5712 0 _0653_
rlabel metal3 117600 18200 117600 18200 0 _0654_
rlabel metal2 117656 5712 117656 5712 0 _0655_
rlabel metal3 115976 18648 115976 18648 0 _0656_
rlabel metal2 115752 15876 115752 15876 0 _0657_
rlabel metal3 113736 15848 113736 15848 0 _0658_
rlabel metal2 112616 6384 112616 6384 0 _0659_
rlabel metal3 111720 3640 111720 3640 0 _0660_
rlabel metal2 111384 5096 111384 5096 0 _0661_
rlabel metal2 113064 6888 113064 6888 0 _0662_
rlabel metal3 110768 13496 110768 13496 0 _0663_
rlabel metal4 110152 12488 110152 12488 0 _0664_
rlabel metal3 94472 15176 94472 15176 0 _0665_
rlabel metal2 62384 16856 62384 16856 0 _0666_
rlabel metal2 62216 17248 62216 17248 0 _0667_
rlabel metal2 61992 18032 61992 18032 0 _0668_
rlabel metal2 64288 17752 64288 17752 0 _0669_
rlabel metal2 61320 18704 61320 18704 0 _0670_
rlabel metal2 62104 17472 62104 17472 0 _0671_
rlabel metal2 63112 16688 63112 16688 0 _0672_
rlabel metal2 86184 13216 86184 13216 0 _0673_
rlabel metal2 89208 11760 89208 11760 0 _0674_
rlabel metal2 59192 17136 59192 17136 0 _0675_
rlabel metal2 73752 12432 73752 12432 0 _0676_
rlabel metal2 94584 11480 94584 11480 0 _0677_
rlabel metal2 90216 10808 90216 10808 0 _0678_
rlabel metal2 57288 17696 57288 17696 0 _0679_
rlabel metal2 61096 16800 61096 16800 0 _0680_
rlabel metal2 49224 15960 49224 15960 0 _0681_
rlabel metal2 43064 20160 43064 20160 0 _0682_
rlabel metal2 58408 14560 58408 14560 0 _0683_
rlabel metal2 64568 16464 64568 16464 0 _0684_
rlabel metal3 64792 17640 64792 17640 0 _0685_
rlabel metal2 64008 15848 64008 15848 0 _0686_
rlabel metal2 65912 10416 65912 10416 0 _0687_
rlabel metal2 59080 10192 59080 10192 0 _0688_
rlabel metal2 89656 9912 89656 9912 0 _0689_
rlabel metal2 88928 13160 88928 13160 0 _0690_
rlabel metal2 67592 11144 67592 11144 0 _0691_
rlabel metal2 50064 20664 50064 20664 0 _0692_
rlabel metal2 87752 12040 87752 12040 0 _0693_
rlabel metal2 64512 19880 64512 19880 0 _0694_
rlabel metal3 66584 18312 66584 18312 0 _0695_
rlabel metal3 65576 19096 65576 19096 0 _0696_
rlabel metal2 67704 19152 67704 19152 0 _0697_
rlabel metal2 66808 16884 66808 16884 0 _0698_
rlabel metal2 77168 10808 77168 10808 0 _0699_
rlabel metal2 76328 12432 76328 12432 0 _0700_
rlabel metal2 86688 16072 86688 16072 0 _0701_
rlabel metal2 54488 26320 54488 26320 0 _0702_
rlabel metal3 57568 26600 57568 26600 0 _0703_
rlabel metal2 47768 25368 47768 25368 0 _0704_
rlabel metal2 46536 26040 46536 26040 0 _0705_
rlabel metal2 92904 14784 92904 14784 0 _0706_
rlabel metal2 58296 10584 58296 10584 0 _0707_
rlabel metal2 90104 11144 90104 11144 0 _0708_
rlabel metal2 88368 10808 88368 10808 0 _0709_
rlabel metal2 75208 12152 75208 12152 0 _0710_
rlabel metal2 75376 14280 75376 14280 0 _0711_
rlabel metal2 86856 14672 86856 14672 0 _0712_
rlabel metal2 97048 10584 97048 10584 0 _0713_
rlabel metal2 96376 8344 96376 8344 0 _0714_
rlabel metal2 59304 5040 59304 5040 0 _0715_
rlabel metal3 95928 8624 95928 8624 0 _0716_
rlabel metal2 95704 12712 95704 12712 0 _0717_
rlabel metal3 59836 16072 59836 16072 0 _0718_
rlabel metal2 84448 12264 84448 12264 0 _0719_
rlabel metal2 77112 11648 77112 11648 0 _0720_
rlabel metal2 79240 14224 79240 14224 0 _0721_
rlabel metal2 81256 14392 81256 14392 0 _0722_
rlabel metal3 67816 19320 67816 19320 0 _0723_
rlabel metal3 83720 9576 83720 9576 0 _0724_
rlabel metal2 83272 12208 83272 12208 0 _0725_
rlabel metal2 84280 8008 84280 8008 0 _0726_
rlabel metal2 86072 12264 86072 12264 0 _0727_
rlabel metal2 87976 13160 87976 13160 0 _0728_
rlabel metal2 89096 12600 89096 12600 0 _0729_
rlabel metal2 96376 13160 96376 13160 0 _0730_
rlabel metal2 85176 9408 85176 9408 0 _0731_
rlabel metal2 85064 11088 85064 11088 0 _0732_
rlabel metal2 96264 12432 96264 12432 0 _0733_
rlabel metal3 92456 12376 92456 12376 0 _0734_
rlabel metal3 95536 15176 95536 15176 0 _0735_
rlabel metal3 74536 2464 74536 2464 0 _0736_
rlabel metal2 97384 10360 97384 10360 0 _0737_
rlabel metal2 98168 10584 98168 10584 0 _0738_
rlabel metal2 67032 15176 67032 15176 0 _0739_
rlabel metal3 91056 13944 91056 13944 0 _0740_
rlabel metal2 95816 7616 95816 7616 0 _0741_
rlabel metal2 95984 7672 95984 7672 0 _0742_
rlabel metal2 97608 15204 97608 15204 0 _0743_
rlabel metal2 71008 28392 71008 28392 0 _0744_
rlabel metal2 96040 15456 96040 15456 0 _0745_
rlabel metal2 84728 9072 84728 9072 0 _0746_
rlabel metal2 97944 6776 97944 6776 0 _0747_
rlabel metal2 98056 10584 98056 10584 0 _0748_
rlabel metal2 42840 23632 42840 23632 0 _0749_
rlabel metal2 43512 22008 43512 22008 0 _0750_
rlabel metal2 48272 20664 48272 20664 0 _0751_
rlabel metal3 87752 13552 87752 13552 0 _0752_
rlabel metal2 51016 49364 51016 49364 0 _0753_
rlabel metal3 57456 23128 57456 23128 0 _0754_
rlabel metal2 63336 27664 63336 27664 0 _0755_
rlabel metal2 72856 27888 72856 27888 0 _0756_
rlabel metal2 64344 27104 64344 27104 0 _0757_
rlabel metal2 71512 27272 71512 27272 0 _0758_
rlabel metal2 65688 27272 65688 27272 0 _0759_
rlabel metal2 73864 25032 73864 25032 0 _0760_
rlabel metal2 72744 25424 72744 25424 0 _0761_
rlabel metal2 69608 25032 69608 25032 0 _0762_
rlabel metal3 68096 24696 68096 24696 0 _0763_
rlabel metal2 71288 24864 71288 24864 0 _0764_
rlabel metal2 50344 23184 50344 23184 0 _0765_
rlabel metal2 74760 25872 74760 25872 0 _0766_
rlabel metal2 74872 25536 74872 25536 0 _0767_
rlabel metal3 112728 18424 112728 18424 0 _0768_
rlabel metal3 50848 25480 50848 25480 0 _0769_
rlabel metal2 64456 24472 64456 24472 0 _0770_
rlabel metal3 67984 24808 67984 24808 0 _0771_
rlabel metal2 70728 27720 70728 27720 0 _0772_
rlabel metal3 75096 27720 75096 27720 0 _0773_
rlabel metal2 109816 19600 109816 19600 0 _0774_
rlabel metal2 110264 19656 110264 19656 0 _0775_
rlabel metal3 112728 19880 112728 19880 0 _0776_
rlabel metal3 92120 20832 92120 20832 0 _0777_
rlabel metal2 109928 20132 109928 20132 0 _0778_
rlabel metal3 89376 25480 89376 25480 0 _0779_
rlabel metal2 111048 18088 111048 18088 0 _0780_
rlabel metal2 112392 18536 112392 18536 0 _0781_
rlabel metal2 96432 17080 96432 17080 0 _0782_
rlabel metal2 109256 17248 109256 17248 0 _0783_
rlabel metal2 109760 17080 109760 17080 0 _0784_
rlabel metal2 105896 19208 105896 19208 0 _0785_
rlabel metal2 86408 17024 86408 17024 0 _0786_
rlabel metal2 106792 19992 106792 19992 0 _0787_
rlabel metal3 107968 15400 107968 15400 0 _0788_
rlabel metal2 108696 15848 108696 15848 0 _0789_
rlabel metal2 108024 15568 108024 15568 0 _0790_
rlabel metal2 72184 26656 72184 26656 0 _0791_
rlabel metal3 91112 17136 91112 17136 0 _0792_
rlabel metal3 107240 17528 107240 17528 0 _0793_
rlabel metal2 92008 18424 92008 18424 0 _0794_
rlabel metal2 94472 21504 94472 21504 0 _0795_
rlabel metal3 105616 19992 105616 19992 0 _0796_
rlabel metal2 73304 27720 73304 27720 0 _0797_
rlabel metal2 74200 27104 74200 27104 0 _0798_
rlabel metal2 74536 25368 74536 25368 0 _0799_
rlabel metal2 86856 23856 86856 23856 0 _0800_
rlabel metal2 86408 23464 86408 23464 0 _0801_
rlabel metal3 87864 21672 87864 21672 0 _0802_
rlabel metal2 93912 22456 93912 22456 0 _0803_
rlabel metal3 92680 20776 92680 20776 0 _0804_
rlabel metal3 91616 22456 91616 22456 0 _0805_
rlabel metal2 87304 17584 87304 17584 0 _0806_
rlabel metal2 87696 19096 87696 19096 0 _0807_
rlabel metal3 87696 21784 87696 21784 0 _0808_
rlabel metal2 86128 20104 86128 20104 0 _0809_
rlabel metal3 88088 18928 88088 18928 0 _0810_
rlabel metal2 86296 17976 86296 17976 0 _0811_
rlabel metal2 87864 18088 87864 18088 0 _0812_
rlabel metal2 86744 19656 86744 19656 0 _0813_
rlabel metal2 97272 19040 97272 19040 0 _0814_
rlabel metal2 91672 18872 91672 18872 0 _0815_
rlabel metal3 69104 23800 69104 23800 0 _0816_
rlabel metal3 68544 28392 68544 28392 0 _0817_
rlabel metal2 73416 25368 73416 25368 0 _0818_
rlabel metal2 95256 21000 95256 21000 0 _0819_
rlabel metal2 96600 19992 96600 19992 0 _0820_
rlabel metal2 97384 18032 97384 18032 0 _0821_
rlabel metal2 98224 19320 98224 19320 0 _0822_
rlabel metal3 97272 19992 97272 19992 0 _0823_
rlabel metal2 96376 18592 96376 18592 0 _0824_
rlabel metal2 94472 17080 94472 17080 0 _0825_
rlabel metal2 97048 16800 97048 16800 0 _0826_
rlabel metal2 101976 17808 101976 17808 0 _0827_
rlabel metal2 101080 16800 101080 16800 0 _0828_
rlabel metal2 100632 15204 100632 15204 0 _0829_
rlabel metal3 102984 15400 102984 15400 0 _0830_
rlabel metal2 102200 16184 102200 16184 0 _0831_
rlabel metal2 91112 16184 91112 16184 0 _0832_
rlabel metal2 100968 17752 100968 17752 0 _0833_
rlabel metal3 49224 17640 49224 17640 0 _0834_
rlabel metal2 45752 27440 45752 27440 0 _0835_
rlabel metal2 49448 15568 49448 15568 0 _0836_
rlabel metal2 48776 9184 48776 9184 0 _0837_
rlabel metal2 48104 15904 48104 15904 0 _0838_
rlabel metal2 50120 11536 50120 11536 0 _0839_
rlabel metal2 72744 9184 72744 9184 0 _0840_
rlabel metal2 71064 15204 71064 15204 0 _0841_
rlabel metal3 70336 13720 70336 13720 0 _0842_
rlabel metal3 49504 9800 49504 9800 0 _0843_
rlabel metal2 68488 6272 68488 6272 0 _0844_
rlabel metal2 63448 8680 63448 8680 0 _0845_
rlabel metal3 62300 9240 62300 9240 0 _0846_
rlabel metal2 69160 13440 69160 13440 0 _0847_
rlabel metal3 71400 17640 71400 17640 0 _0848_
rlabel metal3 65072 17976 65072 17976 0 _0849_
rlabel metal2 69832 13216 69832 13216 0 _0850_
rlabel metal2 61600 11256 61600 11256 0 _0851_
rlabel metal3 70392 15400 70392 15400 0 _0852_
rlabel metal2 88144 18760 88144 18760 0 _0853_
rlabel metal2 87976 15792 87976 15792 0 _0854_
rlabel metal2 73640 16408 73640 16408 0 _0855_
rlabel metal2 76888 16072 76888 16072 0 _0856_
rlabel metal2 70280 12824 70280 12824 0 _0857_
rlabel metal3 61264 9800 61264 9800 0 _0858_
rlabel metal3 66808 12152 66808 12152 0 _0859_
rlabel metal3 69608 15288 69608 15288 0 _0860_
rlabel metal3 65576 15176 65576 15176 0 _0861_
rlabel metal2 50344 11088 50344 11088 0 _0862_
rlabel metal2 65800 13944 65800 13944 0 _0863_
rlabel metal3 65912 14392 65912 14392 0 _0864_
rlabel metal2 65016 12264 65016 12264 0 _0865_
rlabel metal2 64680 9800 64680 9800 0 _0866_
rlabel metal2 64344 9296 64344 9296 0 _0867_
rlabel metal2 65016 8624 65016 8624 0 _0868_
rlabel metal2 67032 11648 67032 11648 0 _0869_
rlabel metal3 64736 9688 64736 9688 0 _0870_
rlabel metal2 66080 9240 66080 9240 0 _0871_
rlabel metal2 65128 12992 65128 12992 0 _0872_
rlabel metal2 64120 10976 64120 10976 0 _0873_
rlabel metal2 66472 9520 66472 9520 0 _0874_
rlabel metal2 69496 9632 69496 9632 0 _0875_
rlabel metal2 67088 8232 67088 8232 0 _0876_
rlabel metal2 67256 8512 67256 8512 0 _0877_
rlabel metal3 70728 9688 70728 9688 0 _0878_
rlabel metal2 66696 9464 66696 9464 0 _0879_
rlabel metal3 74368 9800 74368 9800 0 _0880_
rlabel metal2 75768 8288 75768 8288 0 _0881_
rlabel metal2 71904 6104 71904 6104 0 _0882_
rlabel metal2 69384 11032 69384 11032 0 _0883_
rlabel metal2 73080 8792 73080 8792 0 _0884_
rlabel metal2 73416 9856 73416 9856 0 _0885_
rlabel metal2 67480 8288 67480 8288 0 _0886_
rlabel metal2 73416 11928 73416 11928 0 _0887_
rlabel metal3 75488 11368 75488 11368 0 _0888_
rlabel metal3 73752 11368 73752 11368 0 _0889_
rlabel metal2 89040 8232 89040 8232 0 _0890_
rlabel metal2 86184 9520 86184 9520 0 _0891_
rlabel metal2 69720 20272 69720 20272 0 _0892_
rlabel metal2 85960 15736 85960 15736 0 _0893_
rlabel metal3 90384 16184 90384 16184 0 _0894_
rlabel metal2 92400 11368 92400 11368 0 _0895_
rlabel metal2 93072 9688 93072 9688 0 _0896_
rlabel metal2 92680 11480 92680 11480 0 _0897_
rlabel metal2 92232 9912 92232 9912 0 _0898_
rlabel metal2 92568 10472 92568 10472 0 _0899_
rlabel metal2 87304 6328 87304 6328 0 _0900_
rlabel metal2 85736 11256 85736 11256 0 _0901_
rlabel metal3 94808 5152 94808 5152 0 _0902_
rlabel metal2 83272 10080 83272 10080 0 _0903_
rlabel metal3 88144 9800 88144 9800 0 _0904_
rlabel metal3 80192 16072 80192 16072 0 _0905_
rlabel metal2 86968 5432 86968 5432 0 _0906_
rlabel metal2 50344 9408 50344 9408 0 _0907_
rlabel metal2 80808 6272 80808 6272 0 _0908_
rlabel metal2 79240 11424 79240 11424 0 _0909_
rlabel metal2 79688 10640 79688 10640 0 _0910_
rlabel metal2 80528 16072 80528 16072 0 _0911_
rlabel metal2 49224 18368 49224 18368 0 _0912_
rlabel metal3 63224 8288 63224 8288 0 _0913_
rlabel metal2 64960 20104 64960 20104 0 _0914_
rlabel metal2 75992 19208 75992 19208 0 _0915_
rlabel metal2 75208 22400 75208 22400 0 _0916_
rlabel metal2 74648 18648 74648 18648 0 _0917_
rlabel metal2 64344 28056 64344 28056 0 _0918_
rlabel metal3 65520 27832 65520 27832 0 _0919_
rlabel metal2 68768 26936 68768 26936 0 _0920_
rlabel metal2 58520 24808 58520 24808 0 _0921_
rlabel metal3 57680 24808 57680 24808 0 _0922_
rlabel metal2 49000 28224 49000 28224 0 _0923_
rlabel metal2 48104 26320 48104 26320 0 _0924_
rlabel metal2 48216 26040 48216 26040 0 _0925_
rlabel metal2 25816 26656 25816 26656 0 _0926_
rlabel metal2 45416 26376 45416 26376 0 _0927_
rlabel metal3 25200 26264 25200 26264 0 _0928_
rlabel metal2 69496 25928 69496 25928 0 _0929_
rlabel metal3 65632 26600 65632 26600 0 _0930_
rlabel metal2 71176 27608 71176 27608 0 _0931_
rlabel metal3 72520 26936 72520 26936 0 _0932_
rlabel metal2 74984 26992 74984 26992 0 _0933_
rlabel metal2 75488 26488 75488 26488 0 _0934_
rlabel metal2 72296 27384 72296 27384 0 _0935_
rlabel metal2 71960 27440 71960 27440 0 _0936_
rlabel metal2 70280 27216 70280 27216 0 _0937_
rlabel metal2 69832 26992 69832 26992 0 _0938_
rlabel metal2 70784 24584 70784 24584 0 _0939_
rlabel metal2 71008 24920 71008 24920 0 _0940_
rlabel metal2 70056 25032 70056 25032 0 _0941_
rlabel metal2 65800 23912 65800 23912 0 _0942_
rlabel metal2 38360 6944 38360 6944 0 _0943_
rlabel metal3 40600 5880 40600 5880 0 _0944_
rlabel metal2 39984 6104 39984 6104 0 _0945_
rlabel metal3 73360 26264 73360 26264 0 _0946_
rlabel metal2 76552 24976 76552 24976 0 _0947_
rlabel metal2 73864 21952 73864 21952 0 _0948_
rlabel metal2 78232 24136 78232 24136 0 _0949_
rlabel metal2 74648 22568 74648 22568 0 _0950_
rlabel metal4 74648 20216 74648 20216 0 _0951_
rlabel metal2 78792 20720 78792 20720 0 _0952_
rlabel metal2 78456 20944 78456 20944 0 _0953_
rlabel metal2 79016 23184 79016 23184 0 _0954_
rlabel metal2 81256 19824 81256 19824 0 _0955_
rlabel metal2 82152 19544 82152 19544 0 _0956_
rlabel metal2 82208 21784 82208 21784 0 _0957_
rlabel metal2 82152 23016 82152 23016 0 _0958_
rlabel metal2 42392 16184 42392 16184 0 _0959_
rlabel metal2 81704 17024 81704 17024 0 _0960_
rlabel metal3 82040 20104 82040 20104 0 _0961_
rlabel metal2 48440 17136 48440 17136 0 _0962_
rlabel metal2 33208 17920 33208 17920 0 _0963_
rlabel metal2 26656 20776 26656 20776 0 _0964_
rlabel metal2 25480 22736 25480 22736 0 _0965_
rlabel metal2 34104 22232 34104 22232 0 _0966_
rlabel metal3 32144 16856 32144 16856 0 _0967_
rlabel metal3 30352 16856 30352 16856 0 _0968_
rlabel metal3 32200 16072 32200 16072 0 _0969_
rlabel metal2 32648 17136 32648 17136 0 _0970_
rlabel metal2 32984 22736 32984 22736 0 _0971_
rlabel metal3 68936 16912 68936 16912 0 clknet_0_wb_clk_i
rlabel metal2 34440 10192 34440 10192 0 clknet_3_0_0_wb_clk_i
rlabel metal2 54600 10976 54600 10976 0 clknet_3_1_0_wb_clk_i
rlabel metal2 33880 18088 33880 18088 0 clknet_3_2_0_wb_clk_i
rlabel metal3 51856 22344 51856 22344 0 clknet_3_3_0_wb_clk_i
rlabel metal2 81928 10920 81928 10920 0 clknet_3_4_0_wb_clk_i
rlabel metal2 102424 11760 102424 11760 0 clknet_3_5_0_wb_clk_i
rlabel metal2 77224 19656 77224 19656 0 clknet_3_6_0_wb_clk_i
rlabel metal2 98952 18368 98952 18368 0 clknet_3_7_0_wb_clk_i
rlabel metal2 25480 10472 25480 10472 0 clknet_4_0__leaf_wb_clk_i
rlabel metal2 113848 12544 113848 12544 0 clknet_4_10__leaf_wb_clk_i
rlabel metal2 110376 12712 110376 12712 0 clknet_4_11__leaf_wb_clk_i
rlabel metal2 72520 16912 72520 16912 0 clknet_4_12__leaf_wb_clk_i
rlabel metal2 70392 28112 70392 28112 0 clknet_4_13__leaf_wb_clk_i
rlabel metal2 112056 16856 112056 16856 0 clknet_4_14__leaf_wb_clk_i
rlabel metal2 111720 20664 111720 20664 0 clknet_4_15__leaf_wb_clk_i
rlabel metal2 26712 14000 26712 14000 0 clknet_4_1__leaf_wb_clk_i
rlabel metal2 43848 8680 43848 8680 0 clknet_4_2__leaf_wb_clk_i
rlabel metal2 47768 12656 47768 12656 0 clknet_4_3__leaf_wb_clk_i
rlabel metal2 20440 15792 20440 15792 0 clknet_4_4__leaf_wb_clk_i
rlabel metal3 28560 27720 28560 27720 0 clknet_4_5__leaf_wb_clk_i
rlabel metal2 47208 29288 47208 29288 0 clknet_4_6__leaf_wb_clk_i
rlabel metal2 49336 30072 49336 30072 0 clknet_4_7__leaf_wb_clk_i
rlabel metal2 89656 18032 89656 18032 0 clknet_4_8__leaf_wb_clk_i
rlabel metal2 88648 15848 88648 15848 0 clknet_4_9__leaf_wb_clk_i
rlabel metal2 124152 56000 124152 56000 0 io_in[10]
rlabel metal2 135240 56280 135240 56280 0 io_in[11]
rlabel metal2 146888 55412 146888 55412 0 io_in[12]
rlabel metal2 55272 56280 55272 56280 0 io_in[4]
rlabel metal2 66696 56280 66696 56280 0 io_in[5]
rlabel metal2 78120 56168 78120 56168 0 io_in[6]
rlabel metal2 89544 56280 89544 56280 0 io_in[7]
rlabel metal2 100968 56280 100968 56280 0 io_in[8]
rlabel metal2 112280 55412 112280 55412 0 io_in[9]
rlabel metal2 127512 57778 127512 57778 0 io_oeb[10]
rlabel metal2 138936 57778 138936 57778 0 io_oeb[11]
rlabel metal2 150360 57778 150360 57778 0 io_oeb[12]
rlabel metal2 58968 57610 58968 57610 0 io_oeb[4]
rlabel metal2 70392 57778 70392 57778 0 io_oeb[5]
rlabel metal2 81816 57778 81816 57778 0 io_oeb[6]
rlabel metal2 93240 57778 93240 57778 0 io_oeb[7]
rlabel metal2 104664 57778 104664 57778 0 io_oeb[8]
rlabel metal2 116088 57778 116088 57778 0 io_oeb[9]
rlabel metal2 17080 57610 17080 57610 0 io_out[0]
rlabel metal2 131320 57778 131320 57778 0 io_out[10]
rlabel metal2 142744 58170 142744 58170 0 io_out[11]
rlabel metal2 154168 57778 154168 57778 0 io_out[12]
rlabel metal2 28504 57778 28504 57778 0 io_out[1]
rlabel metal2 39928 57610 39928 57610 0 io_out[2]
rlabel metal2 51352 57778 51352 57778 0 io_out[3]
rlabel metal2 62776 57778 62776 57778 0 io_out[4]
rlabel metal2 74200 57610 74200 57610 0 io_out[5]
rlabel metal2 85624 57610 85624 57610 0 io_out[6]
rlabel metal2 97048 57778 97048 57778 0 io_out[7]
rlabel metal2 108472 57778 108472 57778 0 io_out[8]
rlabel metal2 119896 57778 119896 57778 0 io_out[9]
rlabel metal3 119504 56168 119504 56168 0 net1
rlabel metal3 7728 56168 7728 56168 0 net10
rlabel metal2 77224 42224 77224 42224 0 net100
rlabel metal2 88648 49364 88648 49364 0 net101
rlabel metal3 95760 55048 95760 55048 0 net102
rlabel metal3 98784 29400 98784 29400 0 net103
rlabel metal2 119784 55244 119784 55244 0 net104
rlabel metal2 15064 3864 15064 3864 0 net105
rlabel metal3 28616 3080 28616 3080 0 net106
rlabel metal2 65912 3640 65912 3640 0 net107
rlabel metal2 72408 4704 72408 4704 0 net108
rlabel metal2 76440 6160 76440 6160 0 net109
rlabel metal2 11368 4368 11368 4368 0 net11
rlabel metal2 77448 6888 77448 6888 0 net110
rlabel metal2 82040 5768 82040 5768 0 net111
rlabel metal2 86072 4032 86072 4032 0 net112
rlabel metal2 92344 3640 92344 3640 0 net113
rlabel metal2 98448 4312 98448 4312 0 net114
rlabel metal2 99680 3528 99680 3528 0 net115
rlabel metal2 109256 3808 109256 3808 0 net116
rlabel metal2 27832 3864 27832 3864 0 net117
rlabel metal2 106456 6160 106456 6160 0 net118
rlabel metal2 108920 9016 108920 9016 0 net119
rlabel metal2 22568 5992 22568 5992 0 net12
rlabel metal2 116312 5208 116312 5208 0 net120
rlabel metal2 119784 3808 119784 3808 0 net121
rlabel metal2 120680 4704 120680 4704 0 net122
rlabel metal2 127176 4592 127176 4592 0 net123
rlabel metal2 131208 4144 131208 4144 0 net124
rlabel metal2 135016 3248 135016 3248 0 net125
rlabel metal2 139272 3864 139272 3864 0 net126
rlabel metal2 142520 3528 142520 3528 0 net127
rlabel metal2 31192 6720 31192 6720 0 net128
rlabel metal2 146552 3584 146552 3584 0 net129
rlabel metal2 67816 4760 67816 4760 0 net13
rlabel metal3 137760 4928 137760 4928 0 net130
rlabel metal2 40040 4592 40040 4592 0 net131
rlabel metal2 43736 6272 43736 6272 0 net132
rlabel metal2 46872 7168 46872 7168 0 net133
rlabel metal2 48552 6048 48552 6048 0 net134
rlabel metal2 50568 10360 50568 10360 0 net135
rlabel metal2 74312 2912 74312 2912 0 net136
rlabel metal2 63672 4984 63672 4984 0 net137
rlabel metal3 71120 55160 71120 55160 0 net138
rlabel metal2 115864 54432 115864 54432 0 net139
rlabel metal2 65800 5040 65800 5040 0 net14
rlabel metal2 136248 4872 136248 4872 0 net140
rlabel metal2 13384 56280 13384 56280 0 net141
rlabel metal2 24808 56280 24808 56280 0 net142
rlabel metal2 36232 56280 36232 56280 0 net143
rlabel metal2 47656 56280 47656 56280 0 net144
rlabel metal2 89656 3864 89656 3864 0 net145
rlabel metal2 47656 4256 47656 4256 0 net146
rlabel metal2 68824 5376 68824 5376 0 net147
rlabel metal2 55832 5432 55832 5432 0 net148
rlabel metal2 79800 6664 79800 6664 0 net149
rlabel metal2 71792 8344 71792 8344 0 net15
rlabel metal2 115192 8848 115192 8848 0 net150
rlabel metal2 104384 5768 104384 5768 0 net151
rlabel metal2 74088 8232 74088 8232 0 net152
rlabel metal2 62888 3864 62888 3864 0 net153
rlabel metal2 109312 11368 109312 11368 0 net154
rlabel metal2 108696 4368 108696 4368 0 net155
rlabel metal2 84168 5712 84168 5712 0 net156
rlabel metal2 97272 4144 97272 4144 0 net157
rlabel metal2 101808 10584 101808 10584 0 net158
rlabel metal2 121464 4704 121464 4704 0 net159
rlabel metal2 71176 5936 71176 5936 0 net16
rlabel metal2 107576 3864 107576 3864 0 net160
rlabel metal2 61992 4312 61992 4312 0 net161
rlabel metal2 86296 4928 86296 4928 0 net162
rlabel metal3 22568 5880 22568 5880 0 net163
rlabel metal2 122920 3864 122920 3864 0 net164
rlabel metal3 44576 4536 44576 4536 0 net165
rlabel metal2 16632 4760 16632 4760 0 net166
rlabel metal2 21560 4928 21560 4928 0 net167
rlabel metal3 70840 7336 70840 7336 0 net168
rlabel metal2 43288 7336 43288 7336 0 net169
rlabel metal3 70504 15512 70504 15512 0 net17
rlabel metal2 73528 4368 73528 4368 0 net170
rlabel metal3 29904 3528 29904 3528 0 net171
rlabel metal3 28840 4424 28840 4424 0 net172
rlabel metal2 100968 4032 100968 4032 0 net173
rlabel metal2 119112 4760 119112 4760 0 net174
rlabel metal2 115304 4424 115304 4424 0 net175
rlabel metal2 126672 3528 126672 3528 0 net176
rlabel metal2 81704 6552 81704 6552 0 net177
rlabel metal2 62888 8008 62888 8008 0 net178
rlabel metal2 26824 5600 26824 5600 0 net179
rlabel metal3 70504 15624 70504 15624 0 net18
rlabel metal2 77112 7448 77112 7448 0 net180
rlabel metal3 88368 7448 88368 7448 0 net181
rlabel metal2 129192 4648 129192 4648 0 net182
rlabel metal2 100744 7840 100744 7840 0 net183
rlabel metal2 93352 7224 93352 7224 0 net184
rlabel metal2 53592 8568 53592 8568 0 net185
rlabel metal2 69272 8512 69272 8512 0 net186
rlabel metal2 58296 5040 58296 5040 0 net187
rlabel metal2 134344 4368 134344 4368 0 net188
rlabel metal2 35000 6328 35000 6328 0 net189
rlabel metal2 91224 5544 91224 5544 0 net19
rlabel metal2 55160 5824 55160 5824 0 net190
rlabel metal3 28280 4424 28280 4424 0 net191
rlabel metal3 28952 3192 28952 3192 0 net192
rlabel metal2 19320 6104 19320 6104 0 net193
rlabel metal2 39480 10304 39480 10304 0 net194
rlabel metal2 22680 6328 22680 6328 0 net195
rlabel metal2 138264 3864 138264 3864 0 net196
rlabel metal2 51184 3528 51184 3528 0 net197
rlabel metal2 23800 3696 23800 3696 0 net198
rlabel metal2 142128 3528 142128 3528 0 net199
rlabel metal2 125160 44352 125160 44352 0 net2
rlabel metal2 93912 7448 93912 7448 0 net20
rlabel metal2 150024 4872 150024 4872 0 net200
rlabel metal2 22904 4368 22904 4368 0 net201
rlabel metal3 146832 3528 146832 3528 0 net202
rlabel metal2 47600 3528 47600 3528 0 net203
rlabel metal2 38472 6440 38472 6440 0 net204
rlabel metal2 43680 3528 43680 3528 0 net205
rlabel metal3 18368 3640 18368 3640 0 net206
rlabel metal2 121016 5544 121016 5544 0 net207
rlabel metal2 95592 5488 95592 5488 0 net208
rlabel metal2 41608 7056 41608 7056 0 net209
rlabel metal3 92344 11144 92344 11144 0 net21
rlabel metal3 117600 7336 117600 7336 0 net210
rlabel metal2 145096 4592 145096 4592 0 net211
rlabel metal2 137368 4760 137368 4760 0 net212
rlabel metal3 107240 4984 107240 4984 0 net213
rlabel metal2 53928 4480 53928 4480 0 net214
rlabel metal2 98896 5992 98896 5992 0 net215
rlabel metal2 92008 7448 92008 7448 0 net216
rlabel metal2 46312 4816 46312 4816 0 net217
rlabel metal2 71512 5880 71512 5880 0 net218
rlabel metal2 24864 5992 24864 5992 0 net219
rlabel metal2 94360 10024 94360 10024 0 net22
rlabel metal2 80360 5600 80360 5600 0 net220
rlabel metal2 90664 5544 90664 5544 0 net221
rlabel metal2 90888 5712 90888 5712 0 net222
rlabel metal2 41944 8736 41944 8736 0 net223
rlabel metal2 47880 6384 47880 6384 0 net224
rlabel metal2 61544 7728 61544 7728 0 net225
rlabel metal2 57400 4648 57400 4648 0 net226
rlabel metal2 102088 7168 102088 7168 0 net227
rlabel metal2 108920 7784 108920 7784 0 net228
rlabel metal2 24808 7616 24808 7616 0 net23
rlabel metal2 67816 6944 67816 6944 0 net230
rlabel metal2 78456 6832 78456 6832 0 net231
rlabel metal3 31696 7560 31696 7560 0 net232
rlabel metal3 115136 6552 115136 6552 0 net233
rlabel metal2 36232 7560 36232 7560 0 net234
rlabel metal2 63784 5096 63784 5096 0 net235
rlabel metal2 116648 7560 116648 7560 0 net236
rlabel metal2 69944 6832 69944 6832 0 net237
rlabel metal2 80136 5376 80136 5376 0 net238
rlabel metal2 123256 5600 123256 5600 0 net239
rlabel metal2 95368 16744 95368 16744 0 net24
rlabel metal2 57736 8736 57736 8736 0 net240
rlabel metal2 105616 5992 105616 5992 0 net241
rlabel metal2 58632 6160 58632 6160 0 net242
rlabel metal3 86856 6552 86856 6552 0 net243
rlabel metal3 94248 4424 94248 4424 0 net244
rlabel metal2 75544 4760 75544 4760 0 net245
rlabel metal2 127736 4312 127736 4312 0 net246
rlabel metal2 118216 6944 118216 6944 0 net247
rlabel metal3 100240 5320 100240 5320 0 net248
rlabel metal3 111048 5992 111048 5992 0 net249
rlabel metal2 115080 2968 115080 2968 0 net25
rlabel metal2 125608 5712 125608 5712 0 net250
rlabel metal2 75432 8848 75432 8848 0 net251
rlabel metal2 119784 4816 119784 4816 0 net252
rlabel metal2 101472 4424 101472 4424 0 net253
rlabel metal2 104776 4032 104776 4032 0 net254
rlabel metal3 86968 14280 86968 14280 0 net26
rlabel metal2 93576 18760 93576 18760 0 net27
rlabel metal2 121240 5208 121240 5208 0 net28
rlabel metal2 124936 5152 124936 5152 0 net29
rlabel metal2 105784 27440 105784 27440 0 net3
rlabel metal2 124600 4368 124600 4368 0 net30
rlabel metal2 126112 4424 126112 4424 0 net31
rlabel metal2 135800 4760 135800 4760 0 net32
rlabel metal2 142968 4536 142968 4536 0 net33
rlabel metal2 26376 5544 26376 5544 0 net34
rlabel metal2 141736 4704 141736 4704 0 net35
rlabel metal2 142072 4816 142072 4816 0 net36
rlabel metal2 24696 4200 24696 4200 0 net37
rlabel metal2 42392 6216 42392 6216 0 net38
rlabel metal2 49672 5096 49672 5096 0 net39
rlabel metal2 63224 27608 63224 27608 0 net4
rlabel metal2 42168 4088 42168 4088 0 net40
rlabel metal2 47544 10528 47544 10528 0 net41
rlabel metal2 64680 6440 64680 6440 0 net42
rlabel metal2 64904 5488 64904 5488 0 net43
rlabel metal2 15456 5096 15456 5096 0 net44
rlabel metal3 17920 4424 17920 4424 0 net45
rlabel metal2 62552 3920 62552 3920 0 net46
rlabel metal2 68600 6552 68600 6552 0 net47
rlabel metal2 72744 6272 72744 6272 0 net48
rlabel metal2 73136 3416 73136 3416 0 net49
rlabel metal2 73416 29624 73416 29624 0 net5
rlabel metal2 85624 3808 85624 3808 0 net50
rlabel metal2 84392 5600 84392 5600 0 net51
rlabel metal2 89320 4816 89320 4816 0 net52
rlabel metal2 96936 3528 96936 3528 0 net53
rlabel metal2 107352 4144 107352 4144 0 net54
rlabel metal3 102984 4984 102984 4984 0 net55
rlabel metal2 22904 6328 22904 6328 0 net56
rlabel metal2 110936 9240 110936 9240 0 net57
rlabel metal2 110824 5152 110824 5152 0 net58
rlabel metal2 114856 9800 114856 9800 0 net59
rlabel metal2 78232 28000 78232 28000 0 net6
rlabel metal2 122696 5432 122696 5432 0 net60
rlabel metal2 121128 4312 121128 4312 0 net61
rlabel metal2 126504 6272 126504 6272 0 net62
rlabel metal2 121800 10584 121800 10584 0 net63
rlabel metal2 134120 4928 134120 4928 0 net64
rlabel metal2 122696 10584 122696 10584 0 net65
rlabel metal3 141400 3416 141400 3416 0 net66
rlabel metal2 24472 8120 24472 8120 0 net67
rlabel metal2 145544 7728 145544 7728 0 net68
rlabel metal2 149688 3024 149688 3024 0 net69
rlabel metal2 90160 55440 90160 55440 0 net7
rlabel metal2 28392 4312 28392 4312 0 net70
rlabel metal2 21896 13272 21896 13272 0 net71
rlabel metal2 22008 9464 22008 9464 0 net72
rlabel metal2 39312 12712 39312 12712 0 net73
rlabel metal3 55272 7560 55272 7560 0 net74
rlabel metal2 56056 5488 56056 5488 0 net75
rlabel metal3 57456 3416 57456 3416 0 net76
rlabel metal3 39200 15176 39200 15176 0 net77
rlabel metal3 35616 2968 35616 2968 0 net78
rlabel metal3 34048 3304 34048 3304 0 net79
rlabel metal2 101640 55440 101640 55440 0 net8
rlabel metal2 44184 9744 44184 9744 0 net80
rlabel metal2 16016 4312 16016 4312 0 net81
rlabel metal3 88424 2408 88424 2408 0 net82
rlabel metal2 127512 55300 127512 55300 0 net83
rlabel metal2 139272 55608 139272 55608 0 net84
rlabel metal3 70448 55272 70448 55272 0 net85
rlabel metal3 61376 55272 61376 55272 0 net86
rlabel metal2 70448 55160 70448 55160 0 net87
rlabel metal2 81816 55300 81816 55300 0 net88
rlabel metal2 93240 55300 93240 55300 0 net89
rlabel metal3 111272 56168 111272 56168 0 net9
rlabel metal2 104664 55300 104664 55300 0 net90
rlabel metal2 116088 55076 116088 55076 0 net91
rlabel metal2 28168 55048 28168 55048 0 net92
rlabel metal2 131208 34720 131208 34720 0 net93
rlabel metal2 142632 35616 142632 35616 0 net94
rlabel metal2 154056 35560 154056 35560 0 net95
rlabel metal2 28392 55776 28392 55776 0 net96
rlabel metal2 44184 28784 44184 28784 0 net97
rlabel metal3 50848 56056 50848 56056 0 net98
rlabel metal3 62160 56056 62160 56056 0 net99
rlabel metal2 5768 56280 5768 56280 0 rst_i
rlabel metal2 9240 8358 9240 8358 0 wb_clk_i
rlabel metal2 38864 3640 38864 3640 0 wb_hyperram.csr_ack_r
rlabel metal2 32200 3920 32200 3920 0 wb_hyperram.csr_valid_prev_r
rlabel metal2 23968 17528 23968 17528 0 wb_hyperram.double_latency
rlabel metal2 22680 17304 22680 17304 0 wb_hyperram.fixed_latency
rlabel metal2 92960 22120 92960 22120 0 wb_hyperram.hb_data_out\[0\]
rlabel metal2 78568 21112 78568 21112 0 wb_hyperram.hb_data_out\[10\]
rlabel metal3 79464 24920 79464 24920 0 wb_hyperram.hb_data_out\[11\]
rlabel metal3 81256 21784 81256 21784 0 wb_hyperram.hb_data_out\[12\]
rlabel metal2 81648 23352 81648 23352 0 wb_hyperram.hb_data_out\[13\]
rlabel metal2 82712 17192 82712 17192 0 wb_hyperram.hb_data_out\[14\]
rlabel metal3 82936 18424 82936 18424 0 wb_hyperram.hb_data_out\[15\]
rlabel metal2 98056 18872 98056 18872 0 wb_hyperram.hb_data_out\[16\]
rlabel metal2 97608 20328 97608 20328 0 wb_hyperram.hb_data_out\[17\]
rlabel metal2 97272 18088 97272 18088 0 wb_hyperram.hb_data_out\[18\]
rlabel metal3 98224 16184 98224 16184 0 wb_hyperram.hb_data_out\[19\]
rlabel metal2 93016 20384 93016 20384 0 wb_hyperram.hb_data_out\[1\]
rlabel metal2 102984 12264 102984 12264 0 wb_hyperram.hb_data_out\[20\]
rlabel metal2 106120 14672 106120 14672 0 wb_hyperram.hb_data_out\[21\]
rlabel metal3 103544 15288 103544 15288 0 wb_hyperram.hb_data_out\[22\]
rlabel metal2 104440 16352 104440 16352 0 wb_hyperram.hb_data_out\[23\]
rlabel metal2 114856 20356 114856 20356 0 wb_hyperram.hb_data_out\[24\]
rlabel metal3 112728 19320 112728 19320 0 wb_hyperram.hb_data_out\[25\]
rlabel metal2 115640 17024 115640 17024 0 wb_hyperram.hb_data_out\[26\]
rlabel metal3 110936 17416 110936 17416 0 wb_hyperram.hb_data_out\[27\]
rlabel metal2 110712 13776 110712 13776 0 wb_hyperram.hb_data_out\[28\]
rlabel metal2 110544 13944 110544 13944 0 wb_hyperram.hb_data_out\[29\]
rlabel metal2 92120 22064 92120 22064 0 wb_hyperram.hb_data_out\[2\]
rlabel metal2 110264 16408 110264 16408 0 wb_hyperram.hb_data_out\[30\]
rlabel metal2 106680 20328 106680 20328 0 wb_hyperram.hb_data_out\[31\]
rlabel metal2 88312 20160 88312 20160 0 wb_hyperram.hb_data_out\[3\]
rlabel metal2 62776 16016 62776 16016 0 wb_hyperram.hb_data_out\[4\]
rlabel metal2 87976 18144 87976 18144 0 wb_hyperram.hb_data_out\[5\]
rlabel metal3 68040 18928 68040 18928 0 wb_hyperram.hb_data_out\[6\]
rlabel metal3 68264 18816 68264 18816 0 wb_hyperram.hb_data_out\[7\]
rlabel metal2 74872 22344 74872 22344 0 wb_hyperram.hb_data_out\[8\]
rlabel metal2 74760 20384 74760 20384 0 wb_hyperram.hb_data_out\[9\]
rlabel metal3 40656 7448 40656 7448 0 wb_hyperram.hb_read_timeout
rlabel metal3 46704 5320 46704 5320 0 wb_hyperram.hb_valid_prev_r
rlabel metal2 71848 14280 71848 14280 0 wb_hyperram.hram.CA_r\[0\]
rlabel metal2 72744 12600 72744 12600 0 wb_hyperram.hram.CA_r\[16\]
rlabel metal2 70952 15344 70952 15344 0 wb_hyperram.hram.CA_r\[17\]
rlabel metal2 66696 14728 66696 14728 0 wb_hyperram.hram.CA_r\[18\]
rlabel metal2 64904 10640 64904 10640 0 wb_hyperram.hram.CA_r\[19\]
rlabel metal2 76440 16576 76440 16576 0 wb_hyperram.hram.CA_r\[1\]
rlabel metal2 67088 11256 67088 11256 0 wb_hyperram.hram.CA_r\[20\]
rlabel metal2 66304 13720 66304 13720 0 wb_hyperram.hram.CA_r\[21\]
rlabel metal2 67928 11088 67928 11088 0 wb_hyperram.hram.CA_r\[22\]
rlabel metal2 71904 11928 71904 11928 0 wb_hyperram.hram.CA_r\[23\]
rlabel metal3 77000 7336 77000 7336 0 wb_hyperram.hram.CA_r\[24\]
rlabel metal2 75096 8960 75096 8960 0 wb_hyperram.hram.CA_r\[25\]
rlabel metal2 76328 11312 76328 11312 0 wb_hyperram.hram.CA_r\[26\]
rlabel metal2 90888 9184 90888 9184 0 wb_hyperram.hram.CA_r\[27\]
rlabel via2 90888 15176 90888 15176 0 wb_hyperram.hram.CA_r\[28\]
rlabel metal2 91896 12264 91896 12264 0 wb_hyperram.hram.CA_r\[29\]
rlabel metal3 77616 15176 77616 15176 0 wb_hyperram.hram.CA_r\[2\]
rlabel metal2 91224 8848 91224 8848 0 wb_hyperram.hram.CA_r\[30\]
rlabel metal2 83944 15148 83944 15148 0 wb_hyperram.hram.CA_r\[31\]
rlabel metal2 84448 10696 84448 10696 0 wb_hyperram.hram.CA_r\[32\]
rlabel metal2 78120 8176 78120 8176 0 wb_hyperram.hram.CA_r\[33\]
rlabel metal2 77448 11816 77448 11816 0 wb_hyperram.hram.CA_r\[34\]
rlabel metal2 82600 14056 82600 14056 0 wb_hyperram.hram.CA_r\[45\]
rlabel metal2 45080 27272 45080 27272 0 wb_hyperram.hram.CA_r\[46\]
rlabel metal2 43232 24696 43232 24696 0 wb_hyperram.hram.CA_r\[47\]
rlabel metal2 49336 28784 49336 28784 0 wb_hyperram.hram.bus_state_r\[0\]
rlabel metal2 55272 29736 55272 29736 0 wb_hyperram.hram.bus_state_r\[1\]
rlabel metal3 53368 29512 53368 29512 0 wb_hyperram.hram.bus_state_r\[2\]
rlabel metal3 49224 16072 49224 16072 0 wb_hyperram.hram.busy_r
rlabel metal3 56392 16856 56392 16856 0 wb_hyperram.hram.cycle_cnt_r\[0\]
rlabel metal3 66528 17080 66528 17080 0 wb_hyperram.hram.cycle_cnt_r\[1\]
rlabel metal2 58744 19376 58744 19376 0 wb_hyperram.hram.cycle_cnt_r\[2\]
rlabel metal2 65016 19824 65016 19824 0 wb_hyperram.hram.cycle_cnt_r\[3\]
rlabel metal2 63784 18648 63784 18648 0 wb_hyperram.hram.cycle_cnt_r\[4\]
rlabel metal2 63448 20720 63448 20720 0 wb_hyperram.hram.cycle_cnt_r\[5\]
rlabel metal2 53928 11984 53928 11984 0 wb_hyperram.hram.dataw_r\[0\]
rlabel metal2 60536 4984 60536 4984 0 wb_hyperram.hram.dataw_r\[10\]
rlabel metal3 70280 11144 70280 11144 0 wb_hyperram.hram.dataw_r\[11\]
rlabel metal3 72184 9688 72184 9688 0 wb_hyperram.hram.dataw_r\[12\]
rlabel metal2 66472 7672 66472 7672 0 wb_hyperram.hram.dataw_r\[13\]
rlabel metal2 86856 8120 86856 8120 0 wb_hyperram.hram.dataw_r\[14\]
rlabel metal2 87416 7952 87416 7952 0 wb_hyperram.hram.dataw_r\[15\]
rlabel metal2 89600 5208 89600 5208 0 wb_hyperram.hram.dataw_r\[16\]
rlabel metal3 90216 7336 90216 7336 0 wb_hyperram.hram.dataw_r\[17\]
rlabel metal2 99848 10752 99848 10752 0 wb_hyperram.hram.dataw_r\[18\]
rlabel metal2 88312 12992 88312 12992 0 wb_hyperram.hram.dataw_r\[19\]
rlabel metal2 55720 9856 55720 9856 0 wb_hyperram.hram.dataw_r\[1\]
rlabel metal2 102984 11424 102984 11424 0 wb_hyperram.hram.dataw_r\[20\]
rlabel metal2 106232 9072 106232 9072 0 wb_hyperram.hram.dataw_r\[21\]
rlabel metal2 111496 10360 111496 10360 0 wb_hyperram.hram.dataw_r\[22\]
rlabel metal2 111384 8232 111384 8232 0 wb_hyperram.hram.dataw_r\[23\]
rlabel metal2 90832 2968 90832 2968 0 wb_hyperram.hram.dataw_r\[24\]
rlabel metal3 94136 10640 94136 10640 0 wb_hyperram.hram.dataw_r\[25\]
rlabel metal2 96152 9464 96152 9464 0 wb_hyperram.hram.dataw_r\[26\]
rlabel metal2 107632 3304 107632 3304 0 wb_hyperram.hram.dataw_r\[27\]
rlabel metal3 92456 6720 92456 6720 0 wb_hyperram.hram.dataw_r\[28\]
rlabel metal2 96600 8904 96600 8904 0 wb_hyperram.hram.dataw_r\[29\]
rlabel metal2 57176 8736 57176 8736 0 wb_hyperram.hram.dataw_r\[2\]
rlabel metal2 95256 10304 95256 10304 0 wb_hyperram.hram.dataw_r\[30\]
rlabel metal2 96040 5880 96040 5880 0 wb_hyperram.hram.dataw_r\[31\]
rlabel metal2 85848 13720 85848 13720 0 wb_hyperram.hram.dataw_r\[3\]
rlabel metal3 70728 12208 70728 12208 0 wb_hyperram.hram.dataw_r\[4\]
rlabel metal2 63000 10584 63000 10584 0 wb_hyperram.hram.dataw_r\[5\]
rlabel metal2 63336 5712 63336 5712 0 wb_hyperram.hram.dataw_r\[6\]
rlabel metal2 63560 18732 63560 18732 0 wb_hyperram.hram.dataw_r\[7\]
rlabel metal3 56840 5208 56840 5208 0 wb_hyperram.hram.dataw_r\[8\]
rlabel metal2 55048 4312 55048 4312 0 wb_hyperram.hram.dataw_r\[9\]
rlabel metal2 23352 20384 23352 20384 0 wb_hyperram.hram.double_latency_r
rlabel metal2 23800 19712 23800 19712 0 wb_hyperram.hram.fixed_latency_r
rlabel metal3 74760 27048 74760 27048 0 wb_hyperram.hram.read_cnt_r\[0\]
rlabel metal2 69160 27888 69160 27888 0 wb_hyperram.hram.read_cnt_r\[1\]
rlabel metal3 69160 24024 69160 24024 0 wb_hyperram.hram.read_cnt_r\[2\]
rlabel metal2 24584 25592 24584 25592 0 wb_hyperram.hram.rwds_2x_latency_r
rlabel metal3 65688 27944 65688 27944 0 wb_hyperram.hram.rwds_r
rlabel metal2 53592 7112 53592 7112 0 wb_hyperram.hram.sel_r\[0\]
rlabel metal2 49336 7504 49336 7504 0 wb_hyperram.hram.sel_r\[1\]
rlabel metal3 47936 7336 47936 7336 0 wb_hyperram.hram.sel_r\[2\]
rlabel metal2 46648 9576 46648 9576 0 wb_hyperram.hram.sel_r\[3\]
rlabel metal2 24360 7952 24360 7952 0 wb_hyperram.hram.tacc_i\[0\]
rlabel metal2 25816 6440 25816 6440 0 wb_hyperram.hram.tacc_i\[1\]
rlabel metal2 27328 8120 27328 8120 0 wb_hyperram.hram.tacc_i\[2\]
rlabel metal2 27048 8568 27048 8568 0 wb_hyperram.hram.tacc_i\[3\]
rlabel metal2 33432 27944 33432 27944 0 wb_hyperram.hram.tacc_r\[0\]
rlabel metal2 30744 27440 30744 27440 0 wb_hyperram.hram.tacc_r\[1\]
rlabel metal2 30240 26264 30240 26264 0 wb_hyperram.hram.tacc_r\[2\]
rlabel metal3 31192 21672 31192 21672 0 wb_hyperram.hram.tacc_r\[3\]
rlabel metal2 25368 10304 25368 10304 0 wb_hyperram.hram.tcsh_i\[0\]
rlabel metal2 28504 15652 28504 15652 0 wb_hyperram.hram.tcsh_i\[1\]
rlabel metal2 25480 12544 25480 12544 0 wb_hyperram.hram.tcsh_i\[2\]
rlabel metal3 29344 17416 29344 17416 0 wb_hyperram.hram.tcsh_i\[3\]
rlabel metal3 49896 22400 49896 22400 0 wb_hyperram.hram.tcsh_r\[0\]
rlabel metal2 33544 23184 33544 23184 0 wb_hyperram.hram.tcsh_r\[1\]
rlabel metal2 24472 21504 24472 21504 0 wb_hyperram.hram.tcsh_r\[2\]
rlabel metal2 46312 20608 46312 20608 0 wb_hyperram.hram.tcsh_r\[3\]
rlabel metal2 35784 15260 35784 15260 0 wb_hyperram.hram.tpost_i\[0\]
rlabel metal3 35168 15400 35168 15400 0 wb_hyperram.hram.tpost_i\[1\]
rlabel metal2 29512 14000 29512 14000 0 wb_hyperram.hram.tpost_i\[2\]
rlabel metal2 40040 10976 40040 10976 0 wb_hyperram.hram.tpost_i\[3\]
rlabel metal2 49112 22960 49112 22960 0 wb_hyperram.hram.tpost_r\[0\]
rlabel metal2 47432 23240 47432 23240 0 wb_hyperram.hram.tpost_r\[1\]
rlabel metal2 50344 21840 50344 21840 0 wb_hyperram.hram.tpost_r\[2\]
rlabel metal2 43848 15512 43848 15512 0 wb_hyperram.hram.tpost_r\[3\]
rlabel metal2 43960 13272 43960 13272 0 wb_hyperram.hram.tpre_i\[0\]
rlabel metal2 46872 15596 46872 15596 0 wb_hyperram.hram.tpre_i\[1\]
rlabel metal3 44296 13608 44296 13608 0 wb_hyperram.hram.tpre_i\[2\]
rlabel metal2 45864 13272 45864 13272 0 wb_hyperram.hram.tpre_i\[3\]
rlabel metal3 19600 12376 19600 12376 0 wb_hyperram.hram.trmax_i\[0\]
rlabel metal2 20104 13832 20104 13832 0 wb_hyperram.hram.trmax_i\[1\]
rlabel metal2 26712 16072 26712 16072 0 wb_hyperram.hram.trmax_i\[2\]
rlabel metal2 26152 15456 26152 15456 0 wb_hyperram.hram.trmax_i\[3\]
rlabel metal2 22904 15792 22904 15792 0 wb_hyperram.hram.trmax_i\[4\]
rlabel metal2 41048 19768 41048 19768 0 wb_hyperram.hram.trmax_r\[0\]
rlabel metal2 43624 17584 43624 17584 0 wb_hyperram.hram.trmax_r\[1\]
rlabel metal2 39144 19320 39144 19320 0 wb_hyperram.hram.trmax_r\[2\]
rlabel metal2 39816 19152 39816 19152 0 wb_hyperram.hram.trmax_r\[3\]
rlabel metal2 24696 23184 24696 23184 0 wb_hyperram.hram.trmax_r\[4\]
rlabel metal2 10584 2086 10584 2086 0 wb_rst_i
rlabel metal2 11928 2198 11928 2198 0 wbs_ack_o
rlabel metal2 17920 728 17920 728 0 wbs_adr_i[0]
rlabel metal2 63000 854 63000 854 0 wbs_adr_i[10]
rlabel metal3 67424 9128 67424 9128 0 wbs_adr_i[11]
rlabel metal2 69496 4592 69496 4592 0 wbs_adr_i[12]
rlabel metal2 64792 6496 64792 6496 0 wbs_adr_i[13]
rlabel metal2 79128 2422 79128 2422 0 wbs_adr_i[14]
rlabel metal2 86632 6440 86632 6440 0 wbs_adr_i[15]
rlabel metal2 92792 4704 92792 4704 0 wbs_adr_i[16]
rlabel metal2 94248 6888 94248 6888 0 wbs_adr_i[17]
rlabel metal2 95256 2058 95256 2058 0 wbs_adr_i[18]
rlabel metal2 99848 728 99848 728 0 wbs_adr_i[19]
rlabel metal2 22680 2058 22680 2058 0 wbs_adr_i[1]
rlabel metal2 116648 4928 116648 4928 0 wbs_adr_i[20]
rlabel metal2 107408 3192 107408 3192 0 wbs_adr_i[21]
rlabel metal3 113064 6552 113064 6552 0 wbs_adr_i[22]
rlabel metal2 115584 2744 115584 2744 0 wbs_adr_i[23]
rlabel metal2 122136 4480 122136 4480 0 wbs_adr_i[24]
rlabel metal2 124040 4984 124040 4984 0 wbs_adr_i[25]
rlabel metal2 127736 5152 127736 5152 0 wbs_adr_i[26]
rlabel metal3 132160 4312 132160 4312 0 wbs_adr_i[27]
rlabel metal2 135576 2534 135576 2534 0 wbs_adr_i[28]
rlabel metal2 143080 3920 143080 3920 0 wbs_adr_i[29]
rlabel metal2 29848 4872 29848 4872 0 wbs_adr_i[2]
rlabel metal2 144200 3920 144200 3920 0 wbs_adr_i[30]
rlabel metal2 147672 2926 147672 2926 0 wbs_adr_i[31]
rlabel metal2 26264 4312 26264 4312 0 wbs_adr_i[3]
rlabel metal2 41720 7616 41720 7616 0 wbs_adr_i[4]
rlabel metal2 42840 854 42840 854 0 wbs_adr_i[5]
rlabel metal2 46872 2058 46872 2058 0 wbs_adr_i[6]
rlabel metal3 47768 4984 47768 4984 0 wbs_adr_i[7]
rlabel metal2 54936 2058 54936 2058 0 wbs_adr_i[8]
rlabel metal2 58968 854 58968 854 0 wbs_adr_i[9]
rlabel metal2 13272 2478 13272 2478 0 wbs_cyc_i
rlabel metal2 18648 1750 18648 1750 0 wbs_dat_i[0]
rlabel metal2 64344 2702 64344 2702 0 wbs_dat_i[10]
rlabel metal2 68376 2058 68376 2058 0 wbs_dat_i[11]
rlabel metal2 72408 854 72408 854 0 wbs_dat_i[12]
rlabel metal3 75376 4648 75376 4648 0 wbs_dat_i[13]
rlabel metal2 85848 18816 85848 18816 0 wbs_dat_i[14]
rlabel metal2 86520 15484 86520 15484 0 wbs_dat_i[15]
rlabel metal3 92288 5992 92288 5992 0 wbs_dat_i[16]
rlabel metal2 96264 4648 96264 4648 0 wbs_dat_i[17]
rlabel metal2 96600 2086 96600 2086 0 wbs_dat_i[18]
rlabel metal3 113904 2856 113904 2856 0 wbs_dat_i[19]
rlabel metal2 24080 3192 24080 3192 0 wbs_dat_i[1]
rlabel metal2 117096 7672 117096 7672 0 wbs_dat_i[20]
rlabel metal2 108640 3304 108640 3304 0 wbs_dat_i[21]
rlabel metal2 115192 6048 115192 6048 0 wbs_dat_i[22]
rlabel metal2 118832 4984 118832 4984 0 wbs_dat_i[23]
rlabel metal2 122584 4928 122584 4928 0 wbs_dat_i[24]
rlabel metal2 124824 2870 124824 2870 0 wbs_dat_i[25]
rlabel metal3 129640 3528 129640 3528 0 wbs_dat_i[26]
rlabel metal2 133560 2800 133560 2800 0 wbs_dat_i[27]
rlabel metal3 137312 4424 137312 4424 0 wbs_dat_i[28]
rlabel metal2 142744 4984 142744 4984 0 wbs_dat_i[29]
rlabel metal2 29400 2058 29400 2058 0 wbs_dat_i[2]
rlabel metal3 146272 4200 146272 4200 0 wbs_dat_i[30]
rlabel metal2 149016 2870 149016 2870 0 wbs_dat_i[31]
rlabel metal2 20664 5320 20664 5320 0 wbs_dat_i[3]
rlabel metal2 39256 6608 39256 6608 0 wbs_dat_i[4]
rlabel metal2 44184 854 44184 854 0 wbs_dat_i[5]
rlabel metal2 48216 2058 48216 2058 0 wbs_dat_i[6]
rlabel metal2 48216 9352 48216 9352 0 wbs_dat_i[7]
rlabel metal2 56280 854 56280 854 0 wbs_dat_i[8]
rlabel metal2 63896 8960 63896 8960 0 wbs_dat_i[9]
rlabel metal2 19992 1862 19992 1862 0 wbs_dat_o[0]
rlabel metal3 65296 3640 65296 3640 0 wbs_dat_o[10]
rlabel metal3 70112 3640 70112 3640 0 wbs_dat_o[11]
rlabel metal2 73752 2086 73752 2086 0 wbs_dat_o[12]
rlabel metal3 78400 3640 78400 3640 0 wbs_dat_o[13]
rlabel metal3 82432 3640 82432 3640 0 wbs_dat_o[14]
rlabel metal2 85848 854 85848 854 0 wbs_dat_o[15]
rlabel metal2 89880 2058 89880 2058 0 wbs_dat_o[16]
rlabel metal3 94976 4088 94976 4088 0 wbs_dat_o[17]
rlabel metal2 97944 2198 97944 2198 0 wbs_dat_o[18]
rlabel metal2 101976 2198 101976 2198 0 wbs_dat_o[19]
rlabel metal2 25368 2058 25368 2058 0 wbs_dat_o[1]
rlabel metal3 106624 4088 106624 4088 0 wbs_dat_o[20]
rlabel metal2 110040 2030 110040 2030 0 wbs_dat_o[21]
rlabel metal3 115864 3416 115864 3416 0 wbs_dat_o[22]
rlabel metal2 118104 2198 118104 2198 0 wbs_dat_o[23]
rlabel metal2 122136 2198 122136 2198 0 wbs_dat_o[24]
rlabel metal2 126168 2198 126168 2198 0 wbs_dat_o[25]
rlabel metal2 130200 2086 130200 2086 0 wbs_dat_o[26]
rlabel metal2 134232 2198 134232 2198 0 wbs_dat_o[27]
rlabel metal2 138264 854 138264 854 0 wbs_dat_o[28]
rlabel metal2 142296 2198 142296 2198 0 wbs_dat_o[29]
rlabel metal2 30744 2030 30744 2030 0 wbs_dat_o[2]
rlabel metal2 146328 2086 146328 2086 0 wbs_dat_o[30]
rlabel metal2 150360 2198 150360 2198 0 wbs_dat_o[31]
rlabel metal2 36120 1190 36120 1190 0 wbs_dat_o[3]
rlabel metal3 43064 4424 43064 4424 0 wbs_dat_o[4]
rlabel metal2 45528 2198 45528 2198 0 wbs_dat_o[5]
rlabel metal2 49560 2058 49560 2058 0 wbs_dat_o[6]
rlabel metal2 53592 2086 53592 2086 0 wbs_dat_o[7]
rlabel metal3 58352 3640 58352 3640 0 wbs_dat_o[8]
rlabel metal2 61656 2982 61656 2982 0 wbs_dat_o[9]
rlabel metal3 18928 3416 18928 3416 0 wbs_sel_i[0]
rlabel metal2 26712 854 26712 854 0 wbs_sel_i[1]
rlabel metal2 26712 7560 26712 7560 0 wbs_sel_i[2]
rlabel metal2 36120 8680 36120 8680 0 wbs_sel_i[3]
rlabel metal2 14616 2086 14616 2086 0 wbs_stb_i
rlabel metal2 16072 2632 16072 2632 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 160000 60000
<< end >>
