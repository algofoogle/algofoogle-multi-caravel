magic
tech gf180mcuD
magscale 1 10
timestamp 1702289092
<< metal1 >>
rect 12562 57038 12574 57090
rect 12626 57087 12638 57090
rect 13122 57087 13134 57090
rect 12626 57041 13134 57087
rect 12626 57038 12638 57041
rect 13122 57038 13134 57041
rect 13186 57038 13198 57090
rect 54226 56814 54238 56866
rect 54290 56863 54302 56866
rect 55010 56863 55022 56866
rect 54290 56817 55022 56863
rect 54290 56814 54302 56817
rect 55010 56814 55022 56817
rect 55074 56814 55086 56866
rect 16034 56702 16046 56754
rect 16098 56751 16110 56754
rect 17042 56751 17054 56754
rect 16098 56705 17054 56751
rect 16098 56702 16110 56705
rect 17042 56702 17054 56705
rect 17106 56702 17118 56754
rect 17154 56590 17166 56642
rect 17218 56639 17230 56642
rect 17938 56639 17950 56642
rect 17218 56593 17950 56639
rect 17218 56590 17230 56593
rect 17938 56590 17950 56593
rect 18002 56590 18014 56642
rect 18498 56590 18510 56642
rect 18562 56639 18574 56642
rect 18946 56639 18958 56642
rect 18562 56593 18958 56639
rect 18562 56590 18574 56593
rect 18946 56590 18958 56593
rect 19010 56590 19022 56642
rect 24210 56590 24222 56642
rect 24274 56639 24286 56642
rect 24994 56639 25006 56642
rect 24274 56593 25006 56639
rect 24274 56590 24286 56593
rect 24994 56590 25006 56593
rect 25058 56590 25070 56642
rect 28690 56590 28702 56642
rect 28754 56639 28766 56642
rect 29362 56639 29374 56642
rect 28754 56593 29374 56639
rect 28754 56590 28766 56593
rect 29362 56590 29374 56593
rect 29426 56590 29438 56642
rect 44370 56590 44382 56642
rect 44434 56639 44446 56642
rect 44930 56639 44942 56642
rect 44434 56593 44942 56639
rect 44434 56590 44446 56593
rect 44930 56590 44942 56593
rect 44994 56590 45006 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 4622 56306 4674 56318
rect 4622 56242 4674 56254
rect 6190 56306 6242 56318
rect 6190 56242 6242 56254
rect 7422 56306 7474 56318
rect 7422 56242 7474 56254
rect 8654 56306 8706 56318
rect 8654 56242 8706 56254
rect 10110 56306 10162 56318
rect 10110 56242 10162 56254
rect 11454 56306 11506 56318
rect 11454 56242 11506 56254
rect 13134 56306 13186 56318
rect 13134 56242 13186 56254
rect 14030 56306 14082 56318
rect 14030 56242 14082 56254
rect 15038 56306 15090 56318
rect 15038 56242 15090 56254
rect 17166 56306 17218 56318
rect 17166 56242 17218 56254
rect 19406 56306 19458 56318
rect 19406 56242 19458 56254
rect 20750 56306 20802 56318
rect 20750 56242 20802 56254
rect 23214 56306 23266 56318
rect 23214 56242 23266 56254
rect 30718 56306 30770 56318
rect 30718 56242 30770 56254
rect 35310 56306 35362 56318
rect 35310 56242 35362 56254
rect 39118 56306 39170 56318
rect 39118 56242 39170 56254
rect 44046 56306 44098 56318
rect 44046 56242 44098 56254
rect 45390 56306 45442 56318
rect 45390 56242 45442 56254
rect 46398 56306 46450 56318
rect 46398 56242 46450 56254
rect 47854 56306 47906 56318
rect 47854 56242 47906 56254
rect 49086 56306 49138 56318
rect 49086 56242 49138 56254
rect 50430 56306 50482 56318
rect 50430 56242 50482 56254
rect 51774 56306 51826 56318
rect 51774 56242 51826 56254
rect 53118 56306 53170 56318
rect 53118 56242 53170 56254
rect 55022 56306 55074 56318
rect 55022 56242 55074 56254
rect 55918 56306 55970 56318
rect 55918 56242 55970 56254
rect 5518 56194 5570 56206
rect 5518 56130 5570 56142
rect 5854 56194 5906 56206
rect 16046 56194 16098 56206
rect 15698 56142 15710 56194
rect 15762 56142 15774 56194
rect 5854 56130 5906 56142
rect 16046 56130 16098 56142
rect 16382 56194 16434 56206
rect 16382 56130 16434 56142
rect 17614 56194 17666 56206
rect 17614 56130 17666 56142
rect 18622 56194 18674 56206
rect 18622 56130 18674 56142
rect 18958 56194 19010 56206
rect 18958 56130 19010 56142
rect 19854 56194 19906 56206
rect 19854 56130 19906 56142
rect 20190 56194 20242 56206
rect 20190 56130 20242 56142
rect 21310 56194 21362 56206
rect 21310 56130 21362 56142
rect 22430 56082 22482 56094
rect 15474 56030 15486 56082
rect 15538 56030 15550 56082
rect 22430 56018 22482 56030
rect 23998 56082 24050 56094
rect 32174 56082 32226 56094
rect 27346 56030 27358 56082
rect 27410 56030 27422 56082
rect 28690 56030 28702 56082
rect 28754 56030 28766 56082
rect 31378 56030 31390 56082
rect 31442 56030 31454 56082
rect 23998 56018 24050 56030
rect 32174 56018 32226 56030
rect 33742 56082 33794 56094
rect 33742 56018 33794 56030
rect 35982 56082 36034 56094
rect 35982 56018 36034 56030
rect 37550 56082 37602 56094
rect 37550 56018 37602 56030
rect 39790 56082 39842 56094
rect 42466 56030 42478 56082
rect 42530 56030 42542 56082
rect 39790 56018 39842 56030
rect 4958 55970 5010 55982
rect 4958 55906 5010 55918
rect 6974 55970 7026 55982
rect 6974 55906 7026 55918
rect 8206 55970 8258 55982
rect 8206 55906 8258 55918
rect 9662 55970 9714 55982
rect 9662 55906 9714 55918
rect 11006 55970 11058 55982
rect 11006 55906 11058 55918
rect 12350 55970 12402 55982
rect 12350 55906 12402 55918
rect 13582 55970 13634 55982
rect 13582 55906 13634 55918
rect 14590 55970 14642 55982
rect 14590 55906 14642 55918
rect 17726 55970 17778 55982
rect 30494 55970 30546 55982
rect 42926 55970 42978 55982
rect 21970 55918 21982 55970
rect 22034 55918 22046 55970
rect 24546 55918 24558 55970
rect 24610 55918 24622 55970
rect 26674 55918 26686 55970
rect 26738 55918 26750 55970
rect 29362 55918 29374 55970
rect 29426 55918 29438 55970
rect 32610 55918 32622 55970
rect 32674 55918 32686 55970
rect 34178 55918 34190 55970
rect 34242 55918 34254 55970
rect 36418 55918 36430 55970
rect 36482 55918 36494 55970
rect 37986 55918 37998 55970
rect 38050 55918 38062 55970
rect 40338 55918 40350 55970
rect 40402 55918 40414 55970
rect 42018 55918 42030 55970
rect 42082 55918 42094 55970
rect 17726 55906 17778 55918
rect 30494 55906 30546 55918
rect 42926 55906 42978 55918
rect 43598 55970 43650 55982
rect 43598 55906 43650 55918
rect 44494 55970 44546 55982
rect 44494 55906 44546 55918
rect 44942 55970 44994 55982
rect 44942 55906 44994 55918
rect 45950 55970 46002 55982
rect 45950 55906 46002 55918
rect 47406 55970 47458 55982
rect 47406 55906 47458 55918
rect 48638 55970 48690 55982
rect 48638 55906 48690 55918
rect 49982 55970 50034 55982
rect 49982 55906 50034 55918
rect 51326 55970 51378 55982
rect 51326 55906 51378 55918
rect 52670 55970 52722 55982
rect 52670 55906 52722 55918
rect 54014 55970 54066 55982
rect 54014 55906 54066 55918
rect 55470 55970 55522 55982
rect 55470 55906 55522 55918
rect 17838 55858 17890 55870
rect 17838 55794 17890 55806
rect 18286 55858 18338 55870
rect 18286 55794 18338 55806
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 15934 55522 15986 55534
rect 15934 55458 15986 55470
rect 17838 55522 17890 55534
rect 17838 55458 17890 55470
rect 18510 55522 18562 55534
rect 18510 55458 18562 55470
rect 19406 55522 19458 55534
rect 19406 55458 19458 55470
rect 20414 55522 20466 55534
rect 20414 55458 20466 55470
rect 15598 55410 15650 55422
rect 4610 55358 4622 55410
rect 4674 55358 4686 55410
rect 5954 55358 5966 55410
rect 6018 55358 6030 55410
rect 15598 55346 15650 55358
rect 18846 55410 18898 55422
rect 25218 55358 25230 55410
rect 25282 55358 25294 55410
rect 28578 55358 28590 55410
rect 28642 55358 28654 55410
rect 32050 55358 32062 55410
rect 32114 55358 32126 55410
rect 35746 55358 35758 55410
rect 35810 55358 35822 55410
rect 37426 55358 37438 55410
rect 37490 55358 37502 55410
rect 39330 55358 39342 55410
rect 39394 55358 39406 55410
rect 18846 55346 18898 55358
rect 16942 55298 16994 55310
rect 1810 55246 1822 55298
rect 1874 55246 1886 55298
rect 8866 55246 8878 55298
rect 8930 55246 8942 55298
rect 16942 55234 16994 55246
rect 17502 55298 17554 55310
rect 17502 55234 17554 55246
rect 18062 55298 18114 55310
rect 22306 55246 22318 55298
rect 22370 55246 22382 55298
rect 25778 55246 25790 55298
rect 25842 55246 25854 55298
rect 29138 55246 29150 55298
rect 29202 55246 29214 55298
rect 32946 55246 32958 55298
rect 33010 55246 33022 55298
rect 38098 55246 38110 55298
rect 38162 55246 38174 55298
rect 42130 55246 42142 55298
rect 42194 55246 42206 55298
rect 18062 55234 18114 55246
rect 16382 55186 16434 55198
rect 2482 55134 2494 55186
rect 2546 55134 2558 55186
rect 8082 55134 8094 55186
rect 8146 55134 8158 55186
rect 16382 55122 16434 55134
rect 16830 55186 16882 55198
rect 16830 55122 16882 55134
rect 17278 55186 17330 55198
rect 17278 55122 17330 55134
rect 17614 55186 17666 55198
rect 17614 55122 17666 55134
rect 19070 55186 19122 55198
rect 19070 55122 19122 55134
rect 21758 55186 21810 55198
rect 32398 55186 32450 55198
rect 36094 55186 36146 55198
rect 23090 55134 23102 55186
rect 23154 55134 23166 55186
rect 26450 55134 26462 55186
rect 26514 55134 26526 55186
rect 29922 55134 29934 55186
rect 29986 55134 29998 55186
rect 33618 55134 33630 55186
rect 33682 55134 33694 55186
rect 21758 55122 21810 55134
rect 32398 55122 32450 55134
rect 36094 55122 36146 55134
rect 38558 55186 38610 55198
rect 42590 55186 42642 55198
rect 41458 55134 41470 55186
rect 41522 55134 41534 55186
rect 38558 55122 38610 55134
rect 42590 55122 42642 55134
rect 42702 55186 42754 55198
rect 42702 55122 42754 55134
rect 43262 55186 43314 55198
rect 43262 55122 43314 55134
rect 43934 55186 43986 55198
rect 43934 55122 43986 55134
rect 5070 55074 5122 55086
rect 5070 55010 5122 55022
rect 9326 55074 9378 55086
rect 9326 55010 9378 55022
rect 16606 55074 16658 55086
rect 16606 55010 16658 55022
rect 19966 55074 20018 55086
rect 19966 55010 20018 55022
rect 21422 55074 21474 55086
rect 21422 55010 21474 55022
rect 43598 55074 43650 55086
rect 43598 55010 43650 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 2494 54738 2546 54750
rect 2494 54674 2546 54686
rect 15934 54738 15986 54750
rect 15934 54674 15986 54686
rect 16606 54738 16658 54750
rect 16606 54674 16658 54686
rect 16830 54738 16882 54750
rect 16830 54674 16882 54686
rect 22990 54738 23042 54750
rect 22990 54674 23042 54686
rect 23886 54738 23938 54750
rect 23886 54674 23938 54686
rect 25566 54738 25618 54750
rect 25566 54674 25618 54686
rect 26462 54738 26514 54750
rect 26462 54674 26514 54686
rect 27694 54738 27746 54750
rect 27694 54674 27746 54686
rect 28030 54738 28082 54750
rect 28030 54674 28082 54686
rect 29150 54738 29202 54750
rect 29150 54674 29202 54686
rect 29822 54738 29874 54750
rect 29822 54674 29874 54686
rect 31166 54738 31218 54750
rect 31166 54674 31218 54686
rect 39230 54738 39282 54750
rect 39230 54674 39282 54686
rect 40462 54738 40514 54750
rect 40462 54674 40514 54686
rect 41582 54738 41634 54750
rect 41582 54674 41634 54686
rect 2382 54626 2434 54638
rect 2382 54562 2434 54574
rect 7646 54626 7698 54638
rect 7646 54562 7698 54574
rect 16382 54626 16434 54638
rect 16382 54562 16434 54574
rect 40910 54626 40962 54638
rect 40910 54562 40962 54574
rect 41246 54626 41298 54638
rect 44594 54574 44606 54626
rect 44658 54574 44670 54626
rect 41246 54562 41298 54574
rect 2606 54514 2658 54526
rect 2606 54450 2658 54462
rect 2942 54514 2994 54526
rect 4398 54514 4450 54526
rect 7086 54514 7138 54526
rect 3714 54462 3726 54514
rect 3778 54462 3790 54514
rect 6626 54462 6638 54514
rect 6690 54462 6702 54514
rect 2942 54450 2994 54462
rect 4398 54450 4450 54462
rect 7086 54450 7138 54462
rect 7422 54514 7474 54526
rect 7422 54450 7474 54462
rect 11902 54514 11954 54526
rect 18286 54514 18338 54526
rect 27246 54514 27298 54526
rect 12226 54462 12238 54514
rect 12290 54462 12302 54514
rect 18498 54462 18510 54514
rect 18562 54462 18574 54514
rect 19618 54462 19630 54514
rect 19682 54462 19694 54514
rect 24546 54462 24558 54514
rect 24610 54462 24622 54514
rect 11902 54450 11954 54462
rect 18286 54450 18338 54462
rect 27246 54450 27298 54462
rect 28814 54514 28866 54526
rect 35298 54462 35310 54514
rect 35362 54462 35374 54514
rect 45378 54462 45390 54514
rect 45442 54462 45454 54514
rect 28814 54450 28866 54462
rect 4958 54402 5010 54414
rect 9886 54402 9938 54414
rect 15150 54402 15202 54414
rect 32286 54402 32338 54414
rect 3602 54350 3614 54402
rect 3666 54350 3678 54402
rect 6850 54350 6862 54402
rect 6914 54350 6926 54402
rect 7746 54350 7758 54402
rect 7810 54350 7822 54402
rect 13010 54350 13022 54402
rect 13074 54350 13086 54402
rect 18386 54350 18398 54402
rect 18450 54350 18462 54402
rect 20402 54350 20414 54402
rect 20466 54350 20478 54402
rect 22530 54350 22542 54402
rect 22594 54350 22606 54402
rect 4958 54338 5010 54350
rect 9886 54338 9938 54350
rect 15150 54338 15202 54350
rect 32286 54338 32338 54350
rect 33182 54402 33234 54414
rect 33182 54338 33234 54350
rect 34302 54402 34354 54414
rect 34302 54338 34354 54350
rect 34862 54402 34914 54414
rect 42142 54402 42194 54414
rect 45838 54402 45890 54414
rect 35970 54350 35982 54402
rect 36034 54350 36046 54402
rect 38098 54350 38110 54402
rect 38162 54350 38174 54402
rect 42466 54350 42478 54402
rect 42530 54350 42542 54402
rect 34862 54338 34914 54350
rect 42142 54338 42194 54350
rect 45838 54338 45890 54350
rect 48078 54402 48130 54414
rect 48078 54338 48130 54350
rect 16942 54290 16994 54302
rect 18834 54238 18846 54290
rect 18898 54238 18910 54290
rect 16942 54226 16994 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 17502 53954 17554 53966
rect 18958 53954 19010 53966
rect 17826 53902 17838 53954
rect 17890 53902 17902 53954
rect 17502 53890 17554 53902
rect 18958 53890 19010 53902
rect 24670 53954 24722 53966
rect 24670 53890 24722 53902
rect 5070 53842 5122 53854
rect 18398 53842 18450 53854
rect 4610 53790 4622 53842
rect 4674 53790 4686 53842
rect 9650 53790 9662 53842
rect 9714 53790 9726 53842
rect 12898 53790 12910 53842
rect 12962 53790 12974 53842
rect 5070 53778 5122 53790
rect 18398 53778 18450 53790
rect 22990 53842 23042 53854
rect 42926 53842 42978 53854
rect 34066 53790 34078 53842
rect 34130 53790 34142 53842
rect 35186 53790 35198 53842
rect 35250 53790 35262 53842
rect 38658 53790 38670 53842
rect 38722 53790 38734 53842
rect 43250 53790 43262 53842
rect 43314 53790 43326 53842
rect 47730 53790 47742 53842
rect 47794 53790 47806 53842
rect 51314 53790 51326 53842
rect 51378 53790 51390 53842
rect 22990 53778 23042 53790
rect 42926 53778 42978 53790
rect 13470 53730 13522 53742
rect 1810 53678 1822 53730
rect 1874 53678 1886 53730
rect 6738 53678 6750 53730
rect 6802 53678 6814 53730
rect 9986 53678 9998 53730
rect 10050 53678 10062 53730
rect 13470 53666 13522 53678
rect 17278 53730 17330 53742
rect 17278 53666 17330 53678
rect 18622 53730 18674 53742
rect 18622 53666 18674 53678
rect 19182 53730 19234 53742
rect 19182 53666 19234 53678
rect 20302 53730 20354 53742
rect 20302 53666 20354 53678
rect 21870 53730 21922 53742
rect 21870 53666 21922 53678
rect 23662 53730 23714 53742
rect 39902 53730 39954 53742
rect 24658 53678 24670 53730
rect 24722 53678 24734 53730
rect 31154 53678 31166 53730
rect 31218 53678 31230 53730
rect 38882 53678 38894 53730
rect 38946 53678 38958 53730
rect 39218 53678 39230 53730
rect 39282 53678 39294 53730
rect 43474 53678 43486 53730
rect 43538 53678 43550 53730
rect 44818 53678 44830 53730
rect 44882 53678 44894 53730
rect 48402 53678 48414 53730
rect 48466 53678 48478 53730
rect 23662 53666 23714 53678
rect 39902 53666 39954 53678
rect 19742 53618 19794 53630
rect 2482 53566 2494 53618
rect 2546 53566 2558 53618
rect 7522 53566 7534 53618
rect 7586 53566 7598 53618
rect 10770 53566 10782 53618
rect 10834 53566 10846 53618
rect 19742 53554 19794 53566
rect 23102 53618 23154 53630
rect 23102 53554 23154 53566
rect 23438 53618 23490 53630
rect 23438 53554 23490 53566
rect 23998 53618 24050 53630
rect 23998 53554 24050 53566
rect 24334 53618 24386 53630
rect 24334 53554 24386 53566
rect 25006 53618 25058 53630
rect 25006 53554 25058 53566
rect 27134 53618 27186 53630
rect 27134 53554 27186 53566
rect 30718 53618 30770 53630
rect 34638 53618 34690 53630
rect 31938 53566 31950 53618
rect 32002 53566 32014 53618
rect 30718 53554 30770 53566
rect 34638 53554 34690 53566
rect 35534 53618 35586 53630
rect 35534 53554 35586 53566
rect 35870 53618 35922 53630
rect 35870 53554 35922 53566
rect 36206 53618 36258 53630
rect 36206 53554 36258 53566
rect 38670 53618 38722 53630
rect 38670 53554 38722 53566
rect 40350 53618 40402 53630
rect 45602 53566 45614 53618
rect 45666 53566 45678 53618
rect 49186 53566 49198 53618
rect 49250 53566 49262 53618
rect 40350 53554 40402 53566
rect 19294 53506 19346 53518
rect 13794 53454 13806 53506
rect 13858 53454 13870 53506
rect 19294 53442 19346 53454
rect 19630 53506 19682 53518
rect 19630 53442 19682 53454
rect 19854 53506 19906 53518
rect 19854 53442 19906 53454
rect 20638 53506 20690 53518
rect 20638 53442 20690 53454
rect 21422 53506 21474 53518
rect 21422 53442 21474 53454
rect 22542 53506 22594 53518
rect 22542 53442 22594 53454
rect 22878 53506 22930 53518
rect 22878 53442 22930 53454
rect 23774 53506 23826 53518
rect 23774 53442 23826 53454
rect 25678 53506 25730 53518
rect 25678 53442 25730 53454
rect 29262 53506 29314 53518
rect 29262 53442 29314 53454
rect 30382 53506 30434 53518
rect 30382 53442 30434 53454
rect 34750 53506 34802 53518
rect 34750 53442 34802 53454
rect 34974 53506 35026 53518
rect 34974 53442 35026 53454
rect 35310 53506 35362 53518
rect 35310 53442 35362 53454
rect 38446 53506 38498 53518
rect 40238 53506 40290 53518
rect 39554 53454 39566 53506
rect 39618 53454 39630 53506
rect 38446 53442 38498 53454
rect 40238 53442 40290 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 2830 53170 2882 53182
rect 2830 53106 2882 53118
rect 3614 53170 3666 53182
rect 3614 53106 3666 53118
rect 14366 53170 14418 53182
rect 14366 53106 14418 53118
rect 24110 53170 24162 53182
rect 24110 53106 24162 53118
rect 31390 53170 31442 53182
rect 31390 53106 31442 53118
rect 32174 53170 32226 53182
rect 32174 53106 32226 53118
rect 33854 53170 33906 53182
rect 33854 53106 33906 53118
rect 34638 53170 34690 53182
rect 34638 53106 34690 53118
rect 36766 53170 36818 53182
rect 36766 53106 36818 53118
rect 39454 53170 39506 53182
rect 45614 53170 45666 53182
rect 39666 53118 39678 53170
rect 39730 53118 39742 53170
rect 39454 53106 39506 53118
rect 45614 53106 45666 53118
rect 47966 53170 48018 53182
rect 47966 53106 48018 53118
rect 48974 53170 49026 53182
rect 48974 53106 49026 53118
rect 2718 53058 2770 53070
rect 2718 52994 2770 53006
rect 3390 53058 3442 53070
rect 3390 52994 3442 53006
rect 4510 53058 4562 53070
rect 4510 52994 4562 53006
rect 9998 53058 10050 53070
rect 9998 52994 10050 53006
rect 11566 53058 11618 53070
rect 11566 52994 11618 53006
rect 14478 53058 14530 53070
rect 23998 53058 24050 53070
rect 20178 53006 20190 53058
rect 20242 53006 20254 53058
rect 14478 52994 14530 53006
rect 23998 52994 24050 53006
rect 25454 53058 25506 53070
rect 32510 53058 32562 53070
rect 28802 53006 28814 53058
rect 28866 53006 28878 53058
rect 25454 52994 25506 53006
rect 32510 52994 32562 53006
rect 33966 53058 34018 53070
rect 33966 52994 34018 53006
rect 37214 53058 37266 53070
rect 37214 52994 37266 53006
rect 38670 53058 38722 53070
rect 38670 52994 38722 53006
rect 41022 53058 41074 53070
rect 41022 52994 41074 53006
rect 41918 53058 41970 53070
rect 41918 52994 41970 53006
rect 42254 53058 42306 53070
rect 42254 52994 42306 53006
rect 42590 53058 42642 53070
rect 42590 52994 42642 53006
rect 45502 53058 45554 53070
rect 45502 52994 45554 53006
rect 3726 52946 3778 52958
rect 3042 52894 3054 52946
rect 3106 52894 3118 52946
rect 3726 52882 3778 52894
rect 3838 52946 3890 52958
rect 3838 52882 3890 52894
rect 4398 52946 4450 52958
rect 4398 52882 4450 52894
rect 4622 52946 4674 52958
rect 4622 52882 4674 52894
rect 6414 52946 6466 52958
rect 6414 52882 6466 52894
rect 6526 52946 6578 52958
rect 6974 52946 7026 52958
rect 6738 52894 6750 52946
rect 6802 52894 6814 52946
rect 6526 52882 6578 52894
rect 6974 52882 7026 52894
rect 7422 52946 7474 52958
rect 7422 52882 7474 52894
rect 7534 52946 7586 52958
rect 7534 52882 7586 52894
rect 10334 52946 10386 52958
rect 12910 52946 12962 52958
rect 12450 52894 12462 52946
rect 12514 52894 12526 52946
rect 10334 52882 10386 52894
rect 12910 52882 12962 52894
rect 13358 52946 13410 52958
rect 13358 52882 13410 52894
rect 13694 52946 13746 52958
rect 13694 52882 13746 52894
rect 13918 52946 13970 52958
rect 23774 52946 23826 52958
rect 19394 52894 19406 52946
rect 19458 52894 19470 52946
rect 23538 52894 23550 52946
rect 23602 52894 23614 52946
rect 13918 52882 13970 52894
rect 23774 52882 23826 52894
rect 26014 52946 26066 52958
rect 35534 52946 35586 52958
rect 28018 52894 28030 52946
rect 28082 52894 28094 52946
rect 34178 52894 34190 52946
rect 34242 52894 34254 52946
rect 34402 52894 34414 52946
rect 34466 52894 34478 52946
rect 26014 52882 26066 52894
rect 35534 52882 35586 52894
rect 35870 52946 35922 52958
rect 35870 52882 35922 52894
rect 36094 52946 36146 52958
rect 36094 52882 36146 52894
rect 38110 52946 38162 52958
rect 38110 52882 38162 52894
rect 38446 52946 38498 52958
rect 38446 52882 38498 52894
rect 38782 52946 38834 52958
rect 38782 52882 38834 52894
rect 39230 52946 39282 52958
rect 39230 52882 39282 52894
rect 40238 52946 40290 52958
rect 40238 52882 40290 52894
rect 40910 52946 40962 52958
rect 40910 52882 40962 52894
rect 46062 52946 46114 52958
rect 46062 52882 46114 52894
rect 46622 52946 46674 52958
rect 48738 52894 48750 52946
rect 48802 52894 48814 52946
rect 50082 52894 50094 52946
rect 50146 52894 50158 52946
rect 46622 52882 46674 52894
rect 7198 52834 7250 52846
rect 7198 52770 7250 52782
rect 9662 52834 9714 52846
rect 9662 52770 9714 52782
rect 13022 52834 13074 52846
rect 13022 52770 13074 52782
rect 13470 52834 13522 52846
rect 13470 52770 13522 52782
rect 14254 52834 14306 52846
rect 14254 52770 14306 52782
rect 16606 52834 16658 52846
rect 16606 52770 16658 52782
rect 19070 52834 19122 52846
rect 35086 52834 35138 52846
rect 49086 52834 49138 52846
rect 22306 52782 22318 52834
rect 22370 52782 22382 52834
rect 24098 52782 24110 52834
rect 24162 52782 24174 52834
rect 30930 52782 30942 52834
rect 30994 52782 31006 52834
rect 43026 52782 43038 52834
rect 43090 52782 43102 52834
rect 19070 52770 19122 52782
rect 35086 52770 35138 52782
rect 49086 52770 49138 52782
rect 49422 52834 49474 52846
rect 50306 52782 50318 52834
rect 50370 52782 50382 52834
rect 49422 52770 49474 52782
rect 10110 52722 10162 52734
rect 5058 52670 5070 52722
rect 5122 52670 5134 52722
rect 5954 52670 5966 52722
rect 6018 52670 6030 52722
rect 10110 52658 10162 52670
rect 10446 52722 10498 52734
rect 10446 52658 10498 52670
rect 11678 52722 11730 52734
rect 11678 52658 11730 52670
rect 16494 52722 16546 52734
rect 16494 52658 16546 52670
rect 25230 52722 25282 52734
rect 25230 52658 25282 52670
rect 25566 52722 25618 52734
rect 25566 52658 25618 52670
rect 35310 52722 35362 52734
rect 35310 52658 35362 52670
rect 36318 52722 36370 52734
rect 36318 52658 36370 52670
rect 37662 52722 37714 52734
rect 37662 52658 37714 52670
rect 37886 52722 37938 52734
rect 37886 52658 37938 52670
rect 40014 52722 40066 52734
rect 40014 52658 40066 52670
rect 41022 52722 41074 52734
rect 41022 52658 41074 52670
rect 45726 52722 45778 52734
rect 45726 52658 45778 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 20302 52386 20354 52398
rect 39118 52386 39170 52398
rect 10882 52334 10894 52386
rect 10946 52334 10958 52386
rect 33842 52334 33854 52386
rect 33906 52383 33918 52386
rect 34290 52383 34302 52386
rect 33906 52337 34302 52383
rect 33906 52334 33918 52337
rect 34290 52334 34302 52337
rect 34354 52334 34366 52386
rect 20302 52322 20354 52334
rect 39118 52322 39170 52334
rect 45838 52386 45890 52398
rect 45838 52322 45890 52334
rect 4610 52248 4622 52300
rect 4674 52248 4686 52300
rect 5070 52274 5122 52286
rect 5070 52210 5122 52222
rect 11342 52274 11394 52286
rect 22766 52274 22818 52286
rect 28590 52274 28642 52286
rect 35870 52274 35922 52286
rect 18274 52222 18286 52274
rect 18338 52222 18350 52274
rect 24434 52222 24446 52274
rect 24498 52222 24510 52274
rect 25218 52222 25230 52274
rect 25282 52222 25294 52274
rect 27346 52222 27358 52274
rect 27410 52222 27422 52274
rect 33394 52222 33406 52274
rect 33458 52222 33470 52274
rect 34514 52222 34526 52274
rect 34578 52222 34590 52274
rect 11342 52210 11394 52222
rect 22766 52210 22818 52222
rect 28590 52210 28642 52222
rect 35870 52210 35922 52222
rect 38558 52274 38610 52286
rect 38558 52210 38610 52222
rect 39566 52274 39618 52286
rect 46622 52274 46674 52286
rect 41346 52222 41358 52274
rect 41410 52222 41422 52274
rect 39566 52210 39618 52222
rect 46622 52210 46674 52222
rect 7758 52162 7810 52174
rect 1810 52110 1822 52162
rect 1874 52110 1886 52162
rect 5618 52110 5630 52162
rect 5682 52110 5694 52162
rect 7758 52098 7810 52110
rect 10334 52162 10386 52174
rect 10334 52098 10386 52110
rect 10558 52162 10610 52174
rect 12574 52162 12626 52174
rect 12910 52162 12962 52174
rect 11554 52110 11566 52162
rect 11618 52110 11630 52162
rect 12786 52110 12798 52162
rect 12850 52110 12862 52162
rect 10558 52098 10610 52110
rect 12574 52098 12626 52110
rect 12910 52098 12962 52110
rect 13582 52162 13634 52174
rect 13582 52098 13634 52110
rect 13694 52162 13746 52174
rect 13694 52098 13746 52110
rect 13806 52162 13858 52174
rect 13806 52098 13858 52110
rect 14590 52162 14642 52174
rect 18734 52162 18786 52174
rect 15474 52110 15486 52162
rect 15538 52110 15550 52162
rect 14590 52098 14642 52110
rect 18734 52098 18786 52110
rect 19854 52162 19906 52174
rect 19854 52098 19906 52110
rect 23326 52162 23378 52174
rect 33854 52162 33906 52174
rect 23986 52110 23998 52162
rect 24050 52110 24062 52162
rect 28018 52110 28030 52162
rect 28082 52110 28094 52162
rect 30482 52110 30494 52162
rect 30546 52110 30558 52162
rect 23326 52098 23378 52110
rect 33854 52098 33906 52110
rect 34862 52162 34914 52174
rect 34862 52098 34914 52110
rect 37662 52162 37714 52174
rect 37662 52098 37714 52110
rect 38894 52162 38946 52174
rect 38894 52098 38946 52110
rect 39454 52162 39506 52174
rect 40686 52162 40738 52174
rect 39454 52098 39506 52110
rect 39678 52106 39730 52118
rect 40226 52110 40238 52162
rect 40290 52110 40302 52162
rect 8318 52050 8370 52062
rect 2482 51998 2494 52050
rect 2546 51998 2558 52050
rect 5730 51998 5742 52050
rect 5794 51998 5806 52050
rect 8318 51986 8370 51998
rect 11230 52050 11282 52062
rect 19182 52050 19234 52062
rect 16146 51998 16158 52050
rect 16210 51998 16222 52050
rect 11230 51986 11282 51998
rect 19182 51986 19234 51998
rect 20302 52050 20354 52062
rect 24446 52050 24498 52062
rect 35982 52050 36034 52062
rect 20302 51986 20354 51998
rect 20414 51994 20466 52006
rect 6974 51938 7026 51950
rect 19070 51938 19122 51950
rect 14242 51886 14254 51938
rect 14306 51886 14318 51938
rect 14914 51886 14926 51938
rect 14978 51886 14990 51938
rect 31266 51998 31278 52050
rect 31330 51998 31342 52050
rect 24446 51986 24498 51998
rect 35982 51986 36034 51998
rect 37998 52050 38050 52062
rect 40686 52098 40738 52110
rect 41022 52162 41074 52174
rect 41022 52098 41074 52110
rect 42030 52162 42082 52174
rect 42030 52098 42082 52110
rect 45614 52162 45666 52174
rect 45614 52098 45666 52110
rect 46510 52162 46562 52174
rect 46510 52098 46562 52110
rect 46734 52162 46786 52174
rect 46734 52098 46786 52110
rect 47742 52162 47794 52174
rect 47742 52098 47794 52110
rect 48078 52162 48130 52174
rect 48078 52098 48130 52110
rect 48190 52162 48242 52174
rect 48190 52098 48242 52110
rect 50318 52162 50370 52174
rect 50318 52098 50370 52110
rect 50542 52162 50594 52174
rect 50542 52098 50594 52110
rect 50878 52162 50930 52174
rect 50878 52098 50930 52110
rect 39678 52042 39730 52054
rect 39790 52050 39842 52062
rect 37998 51986 38050 51998
rect 39790 51986 39842 51998
rect 41470 52050 41522 52062
rect 41470 51986 41522 51998
rect 41694 52050 41746 52062
rect 43598 52050 43650 52062
rect 42466 51998 42478 52050
rect 42530 51998 42542 52050
rect 42802 51998 42814 52050
rect 42866 51998 42878 52050
rect 41694 51986 41746 51998
rect 43598 51986 43650 51998
rect 43710 52050 43762 52062
rect 43710 51986 43762 51998
rect 47070 52050 47122 52062
rect 47070 51986 47122 51998
rect 50094 52050 50146 52062
rect 50094 51986 50146 51998
rect 51102 52050 51154 52062
rect 51102 51986 51154 51998
rect 51214 52050 51266 52062
rect 51214 51986 51266 51998
rect 20414 51930 20466 51942
rect 24222 51938 24274 51950
rect 6974 51874 7026 51886
rect 19070 51874 19122 51886
rect 24222 51874 24274 51886
rect 24558 51938 24610 51950
rect 24558 51874 24610 51886
rect 34638 51938 34690 51950
rect 34638 51874 34690 51886
rect 35534 51938 35586 51950
rect 35534 51874 35586 51886
rect 35758 51938 35810 51950
rect 35758 51874 35810 51886
rect 37886 51938 37938 51950
rect 37886 51874 37938 51886
rect 38446 51938 38498 51950
rect 38446 51874 38498 51886
rect 38670 51938 38722 51950
rect 38670 51874 38722 51886
rect 40910 51938 40962 51950
rect 43374 51938 43426 51950
rect 49422 51938 49474 51950
rect 50318 51938 50370 51950
rect 42130 51886 42142 51938
rect 42194 51886 42206 51938
rect 46162 51886 46174 51938
rect 46226 51886 46238 51938
rect 47394 51886 47406 51938
rect 47458 51886 47470 51938
rect 49746 51886 49758 51938
rect 49810 51886 49822 51938
rect 40910 51874 40962 51886
rect 43374 51874 43426 51886
rect 49422 51874 49474 51886
rect 50318 51874 50370 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 4510 51602 4562 51614
rect 16270 51602 16322 51614
rect 10098 51550 10110 51602
rect 10162 51550 10174 51602
rect 4510 51538 4562 51550
rect 16270 51538 16322 51550
rect 17726 51602 17778 51614
rect 17726 51538 17778 51550
rect 21870 51602 21922 51614
rect 21870 51538 21922 51550
rect 22542 51602 22594 51614
rect 22542 51538 22594 51550
rect 34862 51602 34914 51614
rect 34862 51538 34914 51550
rect 35982 51602 36034 51614
rect 35982 51538 36034 51550
rect 36094 51602 36146 51614
rect 36094 51538 36146 51550
rect 38110 51602 38162 51614
rect 38110 51538 38162 51550
rect 38782 51602 38834 51614
rect 38782 51538 38834 51550
rect 44942 51602 44994 51614
rect 49646 51602 49698 51614
rect 46610 51550 46622 51602
rect 46674 51550 46686 51602
rect 44942 51538 44994 51550
rect 49646 51538 49698 51550
rect 11006 51490 11058 51502
rect 11006 51426 11058 51438
rect 13246 51490 13298 51502
rect 13246 51426 13298 51438
rect 15374 51490 15426 51502
rect 15374 51426 15426 51438
rect 15822 51490 15874 51502
rect 15822 51426 15874 51438
rect 17614 51490 17666 51502
rect 17614 51426 17666 51438
rect 18174 51490 18226 51502
rect 18174 51426 18226 51438
rect 19070 51490 19122 51502
rect 19070 51426 19122 51438
rect 22654 51490 22706 51502
rect 23774 51490 23826 51502
rect 23426 51438 23438 51490
rect 23490 51438 23502 51490
rect 22654 51426 22706 51438
rect 23774 51426 23826 51438
rect 24558 51490 24610 51502
rect 24558 51426 24610 51438
rect 33854 51490 33906 51502
rect 33854 51426 33906 51438
rect 34526 51490 34578 51502
rect 34526 51426 34578 51438
rect 35534 51490 35586 51502
rect 35534 51426 35586 51438
rect 35758 51490 35810 51502
rect 35758 51426 35810 51438
rect 37326 51490 37378 51502
rect 37326 51426 37378 51438
rect 39230 51490 39282 51502
rect 39230 51426 39282 51438
rect 40126 51490 40178 51502
rect 40126 51426 40178 51438
rect 42142 51490 42194 51502
rect 43822 51490 43874 51502
rect 48078 51490 48130 51502
rect 42802 51438 42814 51490
rect 42866 51438 42878 51490
rect 43026 51438 43038 51490
rect 43090 51438 43102 51490
rect 45602 51438 45614 51490
rect 45666 51438 45678 51490
rect 46050 51438 46062 51490
rect 46114 51438 46126 51490
rect 47170 51438 47182 51490
rect 47234 51438 47246 51490
rect 42142 51426 42194 51438
rect 43822 51426 43874 51438
rect 48078 51426 48130 51438
rect 48862 51490 48914 51502
rect 48862 51426 48914 51438
rect 50654 51490 50706 51502
rect 53218 51438 53230 51490
rect 53282 51438 53294 51490
rect 50654 51426 50706 51438
rect 4622 51378 4674 51390
rect 10446 51378 10498 51390
rect 11790 51378 11842 51390
rect 4386 51326 4398 51378
rect 4450 51326 4462 51378
rect 5394 51326 5406 51378
rect 5458 51326 5470 51378
rect 11330 51326 11342 51378
rect 11394 51326 11406 51378
rect 4622 51314 4674 51326
rect 10446 51314 10498 51326
rect 11790 51314 11842 51326
rect 13582 51378 13634 51390
rect 15262 51378 15314 51390
rect 13794 51326 13806 51378
rect 13858 51326 13870 51378
rect 13582 51314 13634 51326
rect 15262 51314 15314 51326
rect 15598 51378 15650 51390
rect 16830 51378 16882 51390
rect 16482 51326 16494 51378
rect 16546 51326 16558 51378
rect 15598 51314 15650 51326
rect 16830 51314 16882 51326
rect 17950 51378 18002 51390
rect 17950 51314 18002 51326
rect 18398 51378 18450 51390
rect 19854 51378 19906 51390
rect 19282 51326 19294 51378
rect 19346 51326 19358 51378
rect 18398 51314 18450 51326
rect 19854 51314 19906 51326
rect 20190 51378 20242 51390
rect 20190 51314 20242 51326
rect 20414 51378 20466 51390
rect 23102 51378 23154 51390
rect 34078 51378 34130 51390
rect 22082 51326 22094 51378
rect 22146 51326 22158 51378
rect 23986 51326 23998 51378
rect 24050 51326 24062 51378
rect 20414 51314 20466 51326
rect 23102 51314 23154 51326
rect 34078 51314 34130 51326
rect 34302 51378 34354 51390
rect 36766 51378 36818 51390
rect 37998 51378 38050 51390
rect 39566 51378 39618 51390
rect 36306 51326 36318 51378
rect 36370 51326 36382 51378
rect 36530 51326 36542 51378
rect 36594 51326 36606 51378
rect 37090 51326 37102 51378
rect 37154 51326 37166 51378
rect 38546 51326 38558 51378
rect 38610 51326 38622 51378
rect 38882 51326 38894 51378
rect 38946 51326 38958 51378
rect 34302 51314 34354 51326
rect 36766 51314 36818 51326
rect 37998 51314 38050 51326
rect 39566 51314 39618 51326
rect 41358 51378 41410 51390
rect 41358 51314 41410 51326
rect 41582 51378 41634 51390
rect 43710 51378 43762 51390
rect 43362 51326 43374 51378
rect 43426 51326 43438 51378
rect 41582 51314 41634 51326
rect 43710 51314 43762 51326
rect 45278 51378 45330 51390
rect 47966 51378 48018 51390
rect 50318 51378 50370 51390
rect 46498 51326 46510 51378
rect 46562 51326 46574 51378
rect 47058 51326 47070 51378
rect 47122 51326 47134 51378
rect 49186 51326 49198 51378
rect 49250 51326 49262 51378
rect 49410 51326 49422 51378
rect 49474 51326 49486 51378
rect 49970 51326 49982 51378
rect 50034 51326 50046 51378
rect 45278 51314 45330 51326
rect 47966 51314 48018 51326
rect 50318 51314 50370 51326
rect 50430 51378 50482 51390
rect 50430 51314 50482 51326
rect 50766 51378 50818 51390
rect 53890 51326 53902 51378
rect 53954 51326 53966 51378
rect 50766 51314 50818 51326
rect 8766 51266 8818 51278
rect 6178 51214 6190 51266
rect 6242 51214 6254 51266
rect 8306 51214 8318 51266
rect 8370 51214 8382 51266
rect 8766 51202 8818 51214
rect 10670 51266 10722 51278
rect 10670 51202 10722 51214
rect 16046 51266 16098 51278
rect 16046 51202 16098 51214
rect 18734 51266 18786 51278
rect 18734 51202 18786 51214
rect 20078 51266 20130 51278
rect 20078 51202 20130 51214
rect 21758 51266 21810 51278
rect 21758 51202 21810 51214
rect 33742 51266 33794 51278
rect 33742 51202 33794 51214
rect 36990 51266 37042 51278
rect 40226 51214 40238 51266
rect 40290 51214 40302 51266
rect 51090 51214 51102 51266
rect 51154 51214 51166 51266
rect 36990 51202 37042 51214
rect 4846 51154 4898 51166
rect 4846 51090 4898 51102
rect 11342 51154 11394 51166
rect 11342 51090 11394 51102
rect 13358 51154 13410 51166
rect 13358 51090 13410 51102
rect 16270 51154 16322 51166
rect 16270 51090 16322 51102
rect 22430 51154 22482 51166
rect 22430 51090 22482 51102
rect 24446 51154 24498 51166
rect 24446 51090 24498 51102
rect 34974 51154 35026 51166
rect 34974 51090 35026 51102
rect 35198 51154 35250 51166
rect 35198 51090 35250 51102
rect 38110 51154 38162 51166
rect 38110 51090 38162 51102
rect 39454 51154 39506 51166
rect 39454 51090 39506 51102
rect 39902 51154 39954 51166
rect 43822 51154 43874 51166
rect 41906 51102 41918 51154
rect 41970 51102 41982 51154
rect 39902 51090 39954 51102
rect 43822 51090 43874 51102
rect 48078 51154 48130 51166
rect 48078 51090 48130 51102
rect 48750 51154 48802 51166
rect 48750 51090 48802 51102
rect 49758 51154 49810 51166
rect 49758 51090 49810 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 5742 50818 5794 50830
rect 5742 50754 5794 50766
rect 6526 50818 6578 50830
rect 6526 50754 6578 50766
rect 6638 50818 6690 50830
rect 6638 50754 6690 50766
rect 11566 50818 11618 50830
rect 11566 50754 11618 50766
rect 11790 50818 11842 50830
rect 33630 50818 33682 50830
rect 12114 50766 12126 50818
rect 12178 50815 12190 50818
rect 12562 50815 12574 50818
rect 12178 50769 12574 50815
rect 12178 50766 12190 50769
rect 12562 50766 12574 50769
rect 12626 50766 12638 50818
rect 11790 50754 11842 50766
rect 33630 50754 33682 50766
rect 36318 50818 36370 50830
rect 36318 50754 36370 50766
rect 38222 50818 38274 50830
rect 38222 50754 38274 50766
rect 42590 50818 42642 50830
rect 42590 50754 42642 50766
rect 7534 50706 7586 50718
rect 12350 50706 12402 50718
rect 19966 50706 20018 50718
rect 23550 50706 23602 50718
rect 27470 50706 27522 50718
rect 36430 50706 36482 50718
rect 42478 50706 42530 50718
rect 48302 50706 48354 50718
rect 51662 50706 51714 50718
rect 10994 50654 11006 50706
rect 11058 50654 11070 50706
rect 14690 50654 14702 50706
rect 14754 50654 14766 50706
rect 18946 50654 18958 50706
rect 19010 50654 19022 50706
rect 22530 50654 22542 50706
rect 22594 50654 22606 50706
rect 24098 50654 24110 50706
rect 24162 50654 24174 50706
rect 32050 50654 32062 50706
rect 32114 50654 32126 50706
rect 40786 50654 40798 50706
rect 40850 50654 40862 50706
rect 45490 50654 45502 50706
rect 45554 50654 45566 50706
rect 50306 50654 50318 50706
rect 50370 50654 50382 50706
rect 7534 50642 7586 50654
rect 12350 50642 12402 50654
rect 19966 50642 20018 50654
rect 23550 50642 23602 50654
rect 27470 50642 27522 50654
rect 36430 50642 36482 50654
rect 42478 50642 42530 50654
rect 48302 50642 48354 50654
rect 51662 50642 51714 50654
rect 52110 50706 52162 50718
rect 55570 50654 55582 50706
rect 55634 50654 55646 50706
rect 52110 50642 52162 50654
rect 5966 50594 6018 50606
rect 6862 50594 6914 50606
rect 12798 50594 12850 50606
rect 19294 50594 19346 50606
rect 6178 50542 6190 50594
rect 6242 50542 6254 50594
rect 7074 50542 7086 50594
rect 7138 50542 7150 50594
rect 8082 50542 8094 50594
rect 8146 50542 8158 50594
rect 11330 50542 11342 50594
rect 11394 50542 11406 50594
rect 13458 50542 13470 50594
rect 13522 50542 13534 50594
rect 15362 50542 15374 50594
rect 15426 50542 15438 50594
rect 18162 50542 18174 50594
rect 18226 50542 18238 50594
rect 5966 50530 6018 50542
rect 6862 50530 6914 50542
rect 12798 50530 12850 50542
rect 19294 50530 19346 50542
rect 19742 50594 19794 50606
rect 19742 50530 19794 50542
rect 20190 50594 20242 50606
rect 20190 50530 20242 50542
rect 20414 50594 20466 50606
rect 23326 50594 23378 50606
rect 23090 50542 23102 50594
rect 23154 50542 23166 50594
rect 20414 50530 20466 50542
rect 23326 50530 23378 50542
rect 23774 50594 23826 50606
rect 33518 50594 33570 50606
rect 27010 50542 27022 50594
rect 27074 50542 27086 50594
rect 29138 50542 29150 50594
rect 29202 50542 29214 50594
rect 23774 50530 23826 50542
rect 33518 50530 33570 50542
rect 33742 50594 33794 50606
rect 33742 50530 33794 50542
rect 34190 50594 34242 50606
rect 36990 50594 37042 50606
rect 38670 50594 38722 50606
rect 34738 50542 34750 50594
rect 34802 50542 34814 50594
rect 35186 50542 35198 50594
rect 35250 50542 35262 50594
rect 35746 50542 35758 50594
rect 35810 50542 35822 50594
rect 37538 50542 37550 50594
rect 37602 50542 37614 50594
rect 38322 50542 38334 50594
rect 38386 50542 38398 50594
rect 34190 50530 34242 50542
rect 36990 50530 37042 50542
rect 38670 50530 38722 50542
rect 39006 50594 39058 50606
rect 43262 50594 43314 50606
rect 48190 50594 48242 50606
rect 40450 50542 40462 50594
rect 40514 50542 40526 50594
rect 41122 50542 41134 50594
rect 41186 50542 41198 50594
rect 42242 50542 42254 50594
rect 42306 50542 42318 50594
rect 47282 50542 47294 50594
rect 47346 50542 47358 50594
rect 39006 50530 39058 50542
rect 43262 50530 43314 50542
rect 48190 50530 48242 50542
rect 48414 50594 48466 50606
rect 48414 50530 48466 50542
rect 48862 50594 48914 50606
rect 50754 50542 50766 50594
rect 50818 50542 50830 50594
rect 52658 50542 52670 50594
rect 52722 50542 52734 50594
rect 48862 50530 48914 50542
rect 5630 50482 5682 50494
rect 11902 50482 11954 50494
rect 8866 50430 8878 50482
rect 8930 50430 8942 50482
rect 5630 50418 5682 50430
rect 11902 50418 11954 50430
rect 12910 50482 12962 50494
rect 19070 50482 19122 50494
rect 14914 50430 14926 50482
rect 14978 50430 14990 50482
rect 15922 50430 15934 50482
rect 15986 50430 15998 50482
rect 18386 50430 18398 50482
rect 18450 50430 18462 50482
rect 12910 50418 12962 50430
rect 19070 50418 19122 50430
rect 22206 50482 22258 50494
rect 22206 50418 22258 50430
rect 22878 50482 22930 50494
rect 27806 50482 27858 50494
rect 26226 50430 26238 50482
rect 26290 50430 26302 50482
rect 22878 50418 22930 50430
rect 27806 50418 27858 50430
rect 27918 50482 27970 50494
rect 27918 50418 27970 50430
rect 28478 50482 28530 50494
rect 28478 50418 28530 50430
rect 28590 50482 28642 50494
rect 33966 50482 34018 50494
rect 29922 50430 29934 50482
rect 29986 50430 29998 50482
rect 28590 50418 28642 50430
rect 33966 50418 34018 50430
rect 34414 50482 34466 50494
rect 38894 50482 38946 50494
rect 41582 50482 41634 50494
rect 43934 50482 43986 50494
rect 35858 50430 35870 50482
rect 35922 50430 35934 50482
rect 38434 50430 38446 50482
rect 38498 50430 38510 50482
rect 39890 50430 39902 50482
rect 39954 50430 39966 50482
rect 40114 50430 40126 50482
rect 40178 50430 40190 50482
rect 41010 50430 41022 50482
rect 41074 50430 41086 50482
rect 42914 50430 42926 50482
rect 42978 50430 42990 50482
rect 43586 50430 43598 50482
rect 43650 50430 43662 50482
rect 34414 50418 34466 50430
rect 38894 50418 38946 50430
rect 41582 50418 41634 50430
rect 43934 50418 43986 50430
rect 49646 50482 49698 50494
rect 49646 50418 49698 50430
rect 49870 50482 49922 50494
rect 49870 50418 49922 50430
rect 51214 50482 51266 50494
rect 53442 50430 53454 50482
rect 53506 50430 53518 50482
rect 51214 50418 51266 50430
rect 7422 50370 7474 50382
rect 22430 50370 22482 50382
rect 18498 50318 18510 50370
rect 18562 50318 18574 50370
rect 7422 50306 7474 50318
rect 22430 50306 22482 50318
rect 23886 50370 23938 50382
rect 23886 50306 23938 50318
rect 28142 50370 28194 50382
rect 28142 50306 28194 50318
rect 28254 50370 28306 50382
rect 28254 50306 28306 50318
rect 32510 50370 32562 50382
rect 41358 50370 41410 50382
rect 39442 50318 39454 50370
rect 39506 50318 39518 50370
rect 32510 50306 32562 50318
rect 41358 50306 41410 50318
rect 44942 50370 44994 50382
rect 44942 50306 44994 50318
rect 49758 50370 49810 50382
rect 49758 50306 49810 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 7198 50034 7250 50046
rect 6066 49982 6078 50034
rect 6130 49982 6142 50034
rect 7198 49970 7250 49982
rect 16158 50034 16210 50046
rect 18286 50034 18338 50046
rect 24110 50034 24162 50046
rect 17938 49982 17950 50034
rect 18002 49982 18014 50034
rect 23202 49982 23214 50034
rect 23266 49982 23278 50034
rect 16158 49970 16210 49982
rect 18286 49970 18338 49982
rect 24110 49970 24162 49982
rect 35982 50034 36034 50046
rect 35982 49970 36034 49982
rect 36094 50034 36146 50046
rect 36094 49970 36146 49982
rect 36318 50034 36370 50046
rect 42478 50034 42530 50046
rect 37650 49982 37662 50034
rect 37714 49982 37726 50034
rect 36318 49970 36370 49982
rect 42478 49970 42530 49982
rect 43598 50034 43650 50046
rect 43598 49970 43650 49982
rect 51550 50034 51602 50046
rect 51550 49970 51602 49982
rect 51998 50034 52050 50046
rect 51998 49970 52050 49982
rect 52222 50034 52274 50046
rect 52222 49970 52274 49982
rect 6414 49922 6466 49934
rect 2482 49870 2494 49922
rect 2546 49870 2558 49922
rect 6414 49858 6466 49870
rect 6638 49922 6690 49934
rect 6638 49858 6690 49870
rect 7310 49922 7362 49934
rect 7310 49858 7362 49870
rect 11902 49922 11954 49934
rect 11902 49858 11954 49870
rect 15934 49922 15986 49934
rect 15934 49858 15986 49870
rect 17390 49922 17442 49934
rect 17390 49858 17442 49870
rect 18734 49922 18786 49934
rect 18734 49858 18786 49870
rect 20750 49922 20802 49934
rect 20750 49858 20802 49870
rect 31166 49922 31218 49934
rect 31166 49858 31218 49870
rect 31502 49922 31554 49934
rect 31502 49858 31554 49870
rect 31838 49922 31890 49934
rect 36542 49922 36594 49934
rect 35410 49870 35422 49922
rect 35474 49870 35486 49922
rect 31838 49858 31890 49870
rect 36542 49858 36594 49870
rect 36878 49922 36930 49934
rect 36878 49858 36930 49870
rect 37102 49922 37154 49934
rect 37102 49858 37154 49870
rect 37998 49922 38050 49934
rect 43038 49922 43090 49934
rect 40002 49870 40014 49922
rect 40066 49870 40078 49922
rect 37998 49858 38050 49870
rect 43038 49858 43090 49870
rect 43822 49922 43874 49934
rect 43822 49858 43874 49870
rect 43934 49922 43986 49934
rect 43934 49858 43986 49870
rect 48750 49922 48802 49934
rect 48750 49858 48802 49870
rect 50766 49922 50818 49934
rect 50766 49858 50818 49870
rect 51886 49922 51938 49934
rect 51886 49858 51938 49870
rect 5742 49810 5794 49822
rect 1810 49758 1822 49810
rect 1874 49758 1886 49810
rect 5742 49746 5794 49758
rect 7086 49810 7138 49822
rect 12126 49810 12178 49822
rect 14142 49810 14194 49822
rect 10882 49758 10894 49810
rect 10946 49758 10958 49810
rect 13346 49758 13358 49810
rect 13410 49758 13422 49810
rect 13682 49758 13694 49810
rect 13746 49758 13758 49810
rect 7086 49746 7138 49758
rect 12126 49746 12178 49758
rect 14142 49746 14194 49758
rect 14366 49810 14418 49822
rect 14366 49746 14418 49758
rect 15038 49810 15090 49822
rect 17614 49810 17666 49822
rect 19182 49810 19234 49822
rect 16370 49758 16382 49810
rect 16434 49758 16446 49810
rect 18498 49758 18510 49810
rect 18562 49758 18574 49810
rect 15038 49746 15090 49758
rect 17614 49746 17666 49758
rect 19182 49746 19234 49758
rect 19518 49810 19570 49822
rect 19518 49746 19570 49758
rect 19854 49810 19906 49822
rect 19854 49746 19906 49758
rect 20302 49810 20354 49822
rect 20302 49746 20354 49758
rect 20862 49810 20914 49822
rect 20862 49746 20914 49758
rect 22878 49810 22930 49822
rect 22878 49746 22930 49758
rect 23214 49810 23266 49822
rect 23998 49810 24050 49822
rect 23538 49758 23550 49810
rect 23602 49758 23614 49810
rect 23214 49746 23266 49758
rect 23998 49746 24050 49758
rect 24222 49810 24274 49822
rect 30942 49810 30994 49822
rect 37438 49810 37490 49822
rect 41470 49810 41522 49822
rect 42590 49810 42642 49822
rect 24546 49758 24558 49810
rect 24610 49758 24622 49810
rect 27458 49758 27470 49810
rect 27522 49758 27534 49810
rect 35634 49758 35646 49810
rect 35698 49758 35710 49810
rect 38770 49758 38782 49810
rect 38834 49758 38846 49810
rect 39218 49758 39230 49810
rect 39282 49758 39294 49810
rect 39890 49758 39902 49810
rect 39954 49758 39966 49810
rect 42354 49758 42366 49810
rect 42418 49758 42430 49810
rect 24222 49746 24274 49758
rect 30942 49746 30994 49758
rect 37438 49746 37490 49758
rect 41470 49746 41522 49758
rect 42590 49746 42642 49758
rect 43150 49810 43202 49822
rect 51214 49810 51266 49822
rect 43362 49758 43374 49810
rect 43426 49758 43438 49810
rect 47058 49758 47070 49810
rect 47122 49758 47134 49810
rect 48962 49758 48974 49810
rect 49026 49758 49038 49810
rect 49858 49758 49870 49810
rect 49922 49758 49934 49810
rect 50978 49758 50990 49810
rect 51042 49758 51054 49810
rect 51314 49758 51326 49810
rect 51378 49758 51390 49810
rect 43150 49746 43202 49758
rect 51214 49746 51266 49758
rect 5070 49698 5122 49710
rect 4610 49646 4622 49698
rect 4674 49646 4686 49698
rect 5070 49634 5122 49646
rect 5518 49698 5570 49710
rect 5518 49634 5570 49646
rect 6526 49698 6578 49710
rect 6526 49634 6578 49646
rect 11342 49698 11394 49710
rect 11342 49634 11394 49646
rect 12462 49698 12514 49710
rect 19406 49698 19458 49710
rect 13794 49646 13806 49698
rect 13858 49646 13870 49698
rect 12462 49634 12514 49646
rect 19406 49634 19458 49646
rect 23326 49698 23378 49710
rect 23326 49634 23378 49646
rect 27022 49698 27074 49710
rect 32286 49698 32338 49710
rect 28130 49646 28142 49698
rect 28194 49646 28206 49698
rect 30258 49646 30270 49698
rect 30322 49646 30334 49698
rect 27022 49634 27074 49646
rect 32286 49634 32338 49646
rect 33182 49698 33234 49710
rect 33182 49634 33234 49646
rect 37214 49698 37266 49710
rect 37214 49634 37266 49646
rect 40910 49698 40962 49710
rect 40910 49634 40962 49646
rect 44606 49698 44658 49710
rect 45378 49646 45390 49698
rect 45442 49646 45454 49698
rect 49074 49646 49086 49698
rect 49138 49646 49150 49698
rect 49970 49646 49982 49698
rect 50034 49646 50046 49698
rect 44606 49634 44658 49646
rect 14590 49586 14642 49598
rect 14590 49522 14642 49534
rect 14814 49586 14866 49598
rect 14814 49522 14866 49534
rect 15486 49586 15538 49598
rect 15486 49522 15538 49534
rect 15822 49586 15874 49598
rect 15822 49522 15874 49534
rect 18174 49586 18226 49598
rect 18174 49522 18226 49534
rect 20526 49586 20578 49598
rect 20526 49522 20578 49534
rect 21086 49586 21138 49598
rect 21086 49522 21138 49534
rect 30606 49586 30658 49598
rect 39778 49534 39790 49586
rect 39842 49534 39854 49586
rect 30606 49522 30658 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 6302 49250 6354 49262
rect 35982 49250 36034 49262
rect 21858 49198 21870 49250
rect 21922 49198 21934 49250
rect 6302 49186 6354 49198
rect 35982 49186 36034 49198
rect 42142 49250 42194 49262
rect 42142 49186 42194 49198
rect 42926 49250 42978 49262
rect 42926 49186 42978 49198
rect 7870 49138 7922 49150
rect 7870 49074 7922 49086
rect 11342 49138 11394 49150
rect 23774 49138 23826 49150
rect 16706 49086 16718 49138
rect 16770 49086 16782 49138
rect 19954 49086 19966 49138
rect 20018 49086 20030 49138
rect 22754 49086 22766 49138
rect 22818 49086 22830 49138
rect 11342 49074 11394 49086
rect 23774 49074 23826 49086
rect 24334 49138 24386 49150
rect 24334 49074 24386 49086
rect 26014 49138 26066 49150
rect 26014 49074 26066 49086
rect 26798 49138 26850 49150
rect 26798 49074 26850 49086
rect 29598 49138 29650 49150
rect 39566 49138 39618 49150
rect 48302 49138 48354 49150
rect 31154 49086 31166 49138
rect 31218 49086 31230 49138
rect 47730 49086 47742 49138
rect 47794 49086 47806 49138
rect 50978 49086 50990 49138
rect 51042 49086 51054 49138
rect 29598 49074 29650 49086
rect 39566 49074 39618 49086
rect 48302 49074 48354 49086
rect 6078 49026 6130 49038
rect 12686 49026 12738 49038
rect 16606 49026 16658 49038
rect 21310 49026 21362 49038
rect 7186 48974 7198 49026
rect 7250 48974 7262 49026
rect 13458 48974 13470 49026
rect 13522 48974 13534 49026
rect 17154 48974 17166 49026
rect 17218 48974 17230 49026
rect 6078 48962 6130 48974
rect 12686 48962 12738 48974
rect 16606 48962 16658 48974
rect 21310 48962 21362 48974
rect 21534 49026 21586 49038
rect 21534 48962 21586 48974
rect 23102 49026 23154 49038
rect 23102 48962 23154 48974
rect 23214 49026 23266 49038
rect 23214 48962 23266 48974
rect 23886 49026 23938 49038
rect 29038 49026 29090 49038
rect 27346 48974 27358 49026
rect 27410 48974 27422 49026
rect 27570 48974 27582 49026
rect 27634 48974 27646 49026
rect 28466 48974 28478 49026
rect 28530 48974 28542 49026
rect 23886 48962 23938 48974
rect 29038 48962 29090 48974
rect 29486 49026 29538 49038
rect 36094 49026 36146 49038
rect 34066 48974 34078 49026
rect 34130 48974 34142 49026
rect 29486 48962 29538 48974
rect 36094 48962 36146 48974
rect 39342 49026 39394 49038
rect 41470 49026 41522 49038
rect 40786 48974 40798 49026
rect 40850 48974 40862 49026
rect 39342 48962 39394 48974
rect 41470 48962 41522 48974
rect 43262 49026 43314 49038
rect 49310 49026 49362 49038
rect 43698 48974 43710 49026
rect 43762 48974 43774 49026
rect 44930 48974 44942 49026
rect 44994 48974 45006 49026
rect 43262 48962 43314 48974
rect 49310 48962 49362 48974
rect 50654 49026 50706 49038
rect 50654 48962 50706 48974
rect 12798 48914 12850 48926
rect 20302 48914 20354 48926
rect 14130 48862 14142 48914
rect 14194 48862 14206 48914
rect 15138 48862 15150 48914
rect 15202 48862 15214 48914
rect 17826 48862 17838 48914
rect 17890 48862 17902 48914
rect 12798 48850 12850 48862
rect 20302 48850 20354 48862
rect 20638 48914 20690 48926
rect 20638 48850 20690 48862
rect 22766 48914 22818 48926
rect 22766 48850 22818 48862
rect 26686 48914 26738 48926
rect 30830 48914 30882 48926
rect 35982 48914 36034 48926
rect 41806 48914 41858 48926
rect 50878 48914 50930 48926
rect 27234 48862 27246 48914
rect 27298 48862 27310 48914
rect 30034 48862 30046 48914
rect 30098 48862 30110 48914
rect 33282 48862 33294 48914
rect 33346 48862 33358 48914
rect 40114 48862 40126 48914
rect 40178 48862 40190 48914
rect 40674 48862 40686 48914
rect 40738 48862 40750 48914
rect 41122 48862 41134 48914
rect 41186 48862 41198 48914
rect 44034 48862 44046 48914
rect 44098 48862 44110 48914
rect 45602 48862 45614 48914
rect 45666 48862 45678 48914
rect 50306 48862 50318 48914
rect 50370 48862 50382 48914
rect 26686 48850 26738 48862
rect 30830 48850 30882 48862
rect 35982 48850 36034 48862
rect 41806 48850 41858 48862
rect 50878 48850 50930 48862
rect 13022 48802 13074 48814
rect 6626 48750 6638 48802
rect 6690 48750 6702 48802
rect 6962 48750 6974 48802
rect 7026 48750 7038 48802
rect 13022 48738 13074 48750
rect 22542 48802 22594 48814
rect 22542 48738 22594 48750
rect 23662 48802 23714 48814
rect 23662 48738 23714 48750
rect 25566 48802 25618 48814
rect 25566 48738 25618 48750
rect 26462 48802 26514 48814
rect 26462 48738 26514 48750
rect 26910 48802 26962 48814
rect 26910 48738 26962 48750
rect 29710 48802 29762 48814
rect 29710 48738 29762 48750
rect 30382 48802 30434 48814
rect 30382 48738 30434 48750
rect 30718 48802 30770 48814
rect 30718 48738 30770 48750
rect 34526 48802 34578 48814
rect 42030 48802 42082 48814
rect 38994 48750 39006 48802
rect 39058 48750 39070 48802
rect 34526 48738 34578 48750
rect 42030 48738 42082 48750
rect 49086 48802 49138 48814
rect 49982 48802 50034 48814
rect 49634 48750 49646 48802
rect 49698 48750 49710 48802
rect 49086 48738 49138 48750
rect 49982 48738 50034 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 2830 48466 2882 48478
rect 2830 48402 2882 48414
rect 17614 48466 17666 48478
rect 19966 48466 20018 48478
rect 19506 48414 19518 48466
rect 19570 48414 19582 48466
rect 17614 48402 17666 48414
rect 19966 48402 20018 48414
rect 20190 48466 20242 48478
rect 20190 48402 20242 48414
rect 20974 48466 21026 48478
rect 23214 48466 23266 48478
rect 22978 48414 22990 48466
rect 23042 48414 23054 48466
rect 20974 48402 21026 48414
rect 23214 48402 23266 48414
rect 26350 48466 26402 48478
rect 26350 48402 26402 48414
rect 27470 48466 27522 48478
rect 27470 48402 27522 48414
rect 27582 48466 27634 48478
rect 27582 48402 27634 48414
rect 28702 48466 28754 48478
rect 28702 48402 28754 48414
rect 28814 48466 28866 48478
rect 28814 48402 28866 48414
rect 39230 48466 39282 48478
rect 40014 48466 40066 48478
rect 39666 48414 39678 48466
rect 39730 48414 39742 48466
rect 39230 48402 39282 48414
rect 40014 48402 40066 48414
rect 45838 48466 45890 48478
rect 49522 48414 49534 48466
rect 49586 48414 49598 48466
rect 45838 48402 45890 48414
rect 12126 48354 12178 48366
rect 12126 48290 12178 48302
rect 14142 48354 14194 48366
rect 14142 48290 14194 48302
rect 15598 48354 15650 48366
rect 15598 48290 15650 48302
rect 17726 48354 17778 48366
rect 19182 48354 19234 48366
rect 18834 48302 18846 48354
rect 18898 48302 18910 48354
rect 17726 48290 17778 48302
rect 19182 48290 19234 48302
rect 20414 48354 20466 48366
rect 20414 48290 20466 48302
rect 20526 48354 20578 48366
rect 20526 48290 20578 48302
rect 23438 48354 23490 48366
rect 23438 48290 23490 48302
rect 24670 48354 24722 48366
rect 27134 48354 27186 48366
rect 26674 48302 26686 48354
rect 26738 48302 26750 48354
rect 24670 48290 24722 48302
rect 27134 48290 27186 48302
rect 30606 48354 30658 48366
rect 39342 48354 39394 48366
rect 31826 48302 31838 48354
rect 31890 48302 31902 48354
rect 30606 48290 30658 48302
rect 39342 48290 39394 48302
rect 44494 48354 44546 48366
rect 47854 48354 47906 48366
rect 46386 48302 46398 48354
rect 46450 48302 46462 48354
rect 44494 48290 44546 48302
rect 47854 48290 47906 48302
rect 8318 48242 8370 48254
rect 7634 48190 7646 48242
rect 7698 48190 7710 48242
rect 8318 48178 8370 48190
rect 8430 48242 8482 48254
rect 12350 48242 12402 48254
rect 10210 48190 10222 48242
rect 10274 48190 10286 48242
rect 10882 48190 10894 48242
rect 10946 48190 10958 48242
rect 11330 48190 11342 48242
rect 11394 48190 11406 48242
rect 8430 48178 8482 48190
rect 12350 48178 12402 48190
rect 14702 48242 14754 48254
rect 17278 48242 17330 48254
rect 16818 48190 16830 48242
rect 16882 48190 16894 48242
rect 14702 48178 14754 48190
rect 17278 48178 17330 48190
rect 17950 48242 18002 48254
rect 19854 48242 19906 48254
rect 18610 48190 18622 48242
rect 18674 48190 18686 48242
rect 17950 48178 18002 48190
rect 19854 48178 19906 48190
rect 23550 48242 23602 48254
rect 25790 48242 25842 48254
rect 24322 48190 24334 48242
rect 24386 48190 24398 48242
rect 23550 48178 23602 48190
rect 25790 48178 25842 48190
rect 26014 48242 26066 48254
rect 26014 48178 26066 48190
rect 27358 48242 27410 48254
rect 27358 48178 27410 48190
rect 27694 48242 27746 48254
rect 27694 48178 27746 48190
rect 28926 48242 28978 48254
rect 29374 48242 29426 48254
rect 29026 48190 29038 48242
rect 29090 48190 29102 48242
rect 28926 48178 28978 48190
rect 29374 48178 29426 48190
rect 30046 48242 30098 48254
rect 46622 48242 46674 48254
rect 30370 48190 30382 48242
rect 30434 48190 30446 48242
rect 31378 48190 31390 48242
rect 31442 48190 31454 48242
rect 32050 48190 32062 48242
rect 32114 48190 32126 48242
rect 33394 48190 33406 48242
rect 33458 48190 33470 48242
rect 46050 48190 46062 48242
rect 46114 48190 46126 48242
rect 30046 48178 30098 48190
rect 46622 48178 46674 48190
rect 47070 48242 47122 48254
rect 47070 48178 47122 48190
rect 47182 48242 47234 48254
rect 47182 48178 47234 48190
rect 47630 48242 47682 48254
rect 50094 48242 50146 48254
rect 48066 48190 48078 48242
rect 48130 48190 48142 48242
rect 50530 48190 50542 48242
rect 50594 48190 50606 48242
rect 47630 48178 47682 48190
rect 50094 48178 50146 48190
rect 2942 48130 2994 48142
rect 8094 48130 8146 48142
rect 4722 48078 4734 48130
rect 4786 48078 4798 48130
rect 6850 48078 6862 48130
rect 6914 48078 6926 48130
rect 2942 48066 2994 48078
rect 8094 48066 8146 48078
rect 10670 48130 10722 48142
rect 22430 48130 22482 48142
rect 11666 48078 11678 48130
rect 11730 48078 11742 48130
rect 15474 48078 15486 48130
rect 15538 48078 15550 48130
rect 10670 48066 10722 48078
rect 22430 48066 22482 48078
rect 28142 48130 28194 48142
rect 28142 48066 28194 48078
rect 28254 48130 28306 48142
rect 28254 48066 28306 48078
rect 30942 48130 30994 48142
rect 46174 48130 46226 48142
rect 34178 48078 34190 48130
rect 34242 48078 34254 48130
rect 36306 48078 36318 48130
rect 36370 48078 36382 48130
rect 30942 48066 30994 48078
rect 46174 48066 46226 48078
rect 47406 48130 47458 48142
rect 47406 48066 47458 48078
rect 49198 48130 49250 48142
rect 51314 48078 51326 48130
rect 51378 48078 51390 48130
rect 53442 48078 53454 48130
rect 53506 48078 53518 48130
rect 49198 48066 49250 48078
rect 3054 48018 3106 48030
rect 3054 47954 3106 47966
rect 7982 48018 8034 48030
rect 7982 47954 8034 47966
rect 9662 48018 9714 48030
rect 9662 47954 9714 47966
rect 9774 48018 9826 48030
rect 9774 47954 9826 47966
rect 9998 48018 10050 48030
rect 9998 47954 10050 47966
rect 10558 48018 10610 48030
rect 10558 47954 10610 47966
rect 12686 48018 12738 48030
rect 12686 47954 12738 47966
rect 22654 48018 22706 48030
rect 22654 47954 22706 47966
rect 24334 48018 24386 48030
rect 24334 47954 24386 47966
rect 25454 48018 25506 48030
rect 25454 47954 25506 47966
rect 29598 48018 29650 48030
rect 29598 47954 29650 47966
rect 30270 48018 30322 48030
rect 49870 48018 49922 48030
rect 49074 47966 49086 48018
rect 49138 48015 49150 48018
rect 49298 48015 49310 48018
rect 49138 47969 49310 48015
rect 49138 47966 49150 47969
rect 49298 47966 49310 47969
rect 49362 47966 49374 48018
rect 30270 47954 30322 47966
rect 49870 47954 49922 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 19966 47682 20018 47694
rect 19966 47618 20018 47630
rect 29262 47682 29314 47694
rect 29262 47618 29314 47630
rect 50430 47682 50482 47694
rect 50430 47618 50482 47630
rect 50542 47682 50594 47694
rect 50542 47618 50594 47630
rect 50878 47682 50930 47694
rect 50878 47618 50930 47630
rect 12238 47570 12290 47582
rect 23886 47570 23938 47582
rect 33966 47570 34018 47582
rect 1698 47518 1710 47570
rect 1762 47518 1774 47570
rect 3826 47518 3838 47570
rect 3890 47518 3902 47570
rect 8978 47518 8990 47570
rect 9042 47518 9054 47570
rect 11106 47518 11118 47570
rect 11170 47518 11182 47570
rect 18610 47518 18622 47570
rect 18674 47518 18686 47570
rect 32386 47518 32398 47570
rect 32450 47518 32462 47570
rect 12238 47506 12290 47518
rect 23886 47506 23938 47518
rect 33966 47506 34018 47518
rect 34750 47570 34802 47582
rect 34750 47506 34802 47518
rect 34862 47570 34914 47582
rect 44830 47570 44882 47582
rect 48526 47570 48578 47582
rect 44258 47518 44270 47570
rect 44322 47518 44334 47570
rect 45154 47518 45166 47570
rect 45218 47518 45230 47570
rect 47954 47518 47966 47570
rect 48018 47518 48030 47570
rect 34862 47506 34914 47518
rect 44830 47506 44882 47518
rect 48526 47506 48578 47518
rect 48862 47570 48914 47582
rect 48862 47506 48914 47518
rect 49086 47570 49138 47582
rect 49086 47506 49138 47518
rect 12686 47458 12738 47470
rect 15934 47458 15986 47470
rect 4610 47406 4622 47458
rect 4674 47406 4686 47458
rect 6066 47406 6078 47458
rect 6130 47406 6142 47458
rect 7074 47406 7086 47458
rect 7138 47406 7150 47458
rect 8194 47406 8206 47458
rect 8258 47406 8270 47458
rect 11666 47406 11678 47458
rect 11730 47406 11742 47458
rect 13794 47406 13806 47458
rect 13858 47406 13870 47458
rect 12686 47394 12738 47406
rect 15934 47394 15986 47406
rect 18174 47458 18226 47470
rect 18174 47394 18226 47406
rect 20190 47458 20242 47470
rect 22318 47458 22370 47470
rect 20190 47394 20242 47406
rect 20526 47402 20578 47414
rect 16382 47346 16434 47358
rect 6178 47294 6190 47346
rect 6242 47294 6254 47346
rect 7634 47294 7646 47346
rect 7698 47294 7710 47346
rect 13906 47294 13918 47346
rect 13970 47294 13982 47346
rect 22318 47394 22370 47406
rect 22654 47458 22706 47470
rect 22654 47394 22706 47406
rect 24110 47458 24162 47470
rect 24110 47394 24162 47406
rect 27582 47458 27634 47470
rect 27582 47394 27634 47406
rect 27918 47458 27970 47470
rect 27918 47394 27970 47406
rect 28254 47458 28306 47470
rect 33742 47458 33794 47470
rect 45502 47458 45554 47470
rect 33170 47406 33182 47458
rect 33234 47406 33246 47458
rect 35074 47406 35086 47458
rect 35138 47406 35150 47458
rect 41346 47406 41358 47458
rect 41410 47406 41422 47458
rect 28254 47394 28306 47406
rect 33742 47394 33794 47406
rect 45502 47394 45554 47406
rect 45838 47458 45890 47470
rect 45838 47394 45890 47406
rect 46174 47458 46226 47470
rect 46174 47394 46226 47406
rect 46398 47458 46450 47470
rect 50766 47458 50818 47470
rect 47282 47406 47294 47458
rect 47346 47406 47358 47458
rect 47506 47406 47518 47458
rect 47570 47406 47582 47458
rect 46398 47394 46450 47406
rect 50766 47394 50818 47406
rect 20526 47338 20578 47350
rect 22094 47346 22146 47358
rect 16382 47282 16434 47294
rect 22094 47282 22146 47294
rect 29150 47346 29202 47358
rect 29150 47282 29202 47294
rect 29262 47346 29314 47358
rect 29262 47282 29314 47294
rect 34190 47346 34242 47358
rect 34190 47282 34242 47294
rect 34414 47346 34466 47358
rect 46622 47346 46674 47358
rect 42130 47294 42142 47346
rect 42194 47294 42206 47346
rect 34414 47282 34466 47294
rect 46622 47282 46674 47294
rect 48302 47346 48354 47358
rect 48302 47282 48354 47294
rect 5070 47234 5122 47246
rect 11454 47234 11506 47246
rect 6290 47182 6302 47234
rect 6354 47182 6366 47234
rect 5070 47170 5122 47182
rect 11454 47170 11506 47182
rect 12350 47234 12402 47246
rect 12350 47170 12402 47182
rect 12798 47234 12850 47246
rect 12798 47170 12850 47182
rect 13022 47234 13074 47246
rect 19182 47234 19234 47246
rect 20638 47234 20690 47246
rect 15250 47182 15262 47234
rect 15314 47182 15326 47234
rect 19618 47182 19630 47234
rect 19682 47182 19694 47234
rect 13022 47170 13074 47182
rect 19182 47170 19234 47182
rect 20638 47170 20690 47182
rect 20862 47234 20914 47246
rect 20862 47170 20914 47182
rect 22318 47234 22370 47246
rect 22318 47170 22370 47182
rect 24446 47234 24498 47246
rect 24446 47170 24498 47182
rect 24670 47234 24722 47246
rect 24670 47170 24722 47182
rect 24782 47234 24834 47246
rect 24782 47170 24834 47182
rect 25006 47234 25058 47246
rect 25790 47234 25842 47246
rect 26574 47234 26626 47246
rect 25330 47182 25342 47234
rect 25394 47182 25406 47234
rect 26114 47182 26126 47234
rect 26178 47182 26190 47234
rect 25006 47170 25058 47182
rect 25790 47170 25842 47182
rect 26574 47170 26626 47182
rect 27134 47234 27186 47246
rect 27134 47170 27186 47182
rect 27806 47234 27858 47246
rect 27806 47170 27858 47182
rect 35646 47234 35698 47246
rect 35646 47170 35698 47182
rect 45054 47234 45106 47246
rect 45054 47170 45106 47182
rect 45614 47234 45666 47246
rect 45614 47170 45666 47182
rect 46510 47234 46562 47246
rect 46510 47170 46562 47182
rect 49646 47234 49698 47246
rect 51326 47234 51378 47246
rect 49970 47182 49982 47234
rect 50034 47182 50046 47234
rect 49646 47170 49698 47182
rect 51326 47170 51378 47182
rect 51774 47234 51826 47246
rect 51774 47170 51826 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 4286 46898 4338 46910
rect 16382 46898 16434 46910
rect 9874 46846 9886 46898
rect 9938 46846 9950 46898
rect 4286 46834 4338 46846
rect 16382 46834 16434 46846
rect 26798 46898 26850 46910
rect 26798 46834 26850 46846
rect 27582 46898 27634 46910
rect 27582 46834 27634 46846
rect 28254 46898 28306 46910
rect 28254 46834 28306 46846
rect 28702 46898 28754 46910
rect 28702 46834 28754 46846
rect 30830 46898 30882 46910
rect 30830 46834 30882 46846
rect 31390 46898 31442 46910
rect 31390 46834 31442 46846
rect 48078 46898 48130 46910
rect 48078 46834 48130 46846
rect 50206 46898 50258 46910
rect 50206 46834 50258 46846
rect 2158 46786 2210 46798
rect 2158 46722 2210 46734
rect 2270 46786 2322 46798
rect 2270 46722 2322 46734
rect 2606 46786 2658 46798
rect 2606 46722 2658 46734
rect 4510 46786 4562 46798
rect 12910 46786 12962 46798
rect 6290 46734 6302 46786
rect 6354 46734 6366 46786
rect 4510 46722 4562 46734
rect 12910 46722 12962 46734
rect 14366 46786 14418 46798
rect 14366 46722 14418 46734
rect 15710 46786 15762 46798
rect 22542 46786 22594 46798
rect 18722 46734 18734 46786
rect 18786 46734 18798 46786
rect 15710 46722 15762 46734
rect 22542 46722 22594 46734
rect 23886 46786 23938 46798
rect 23886 46722 23938 46734
rect 27022 46786 27074 46798
rect 27022 46722 27074 46734
rect 28814 46786 28866 46798
rect 30046 46786 30098 46798
rect 29474 46734 29486 46786
rect 29538 46734 29550 46786
rect 28814 46722 28866 46734
rect 30046 46722 30098 46734
rect 30718 46786 30770 46798
rect 32062 46786 32114 46798
rect 31714 46734 31726 46786
rect 31778 46734 31790 46786
rect 30718 46722 30770 46734
rect 32062 46722 32114 46734
rect 41134 46786 41186 46798
rect 41134 46722 41186 46734
rect 46734 46786 46786 46798
rect 46734 46722 46786 46734
rect 2718 46674 2770 46686
rect 3950 46674 4002 46686
rect 3042 46622 3054 46674
rect 3106 46622 3118 46674
rect 2718 46610 2770 46622
rect 3950 46610 4002 46622
rect 4174 46674 4226 46686
rect 4174 46610 4226 46622
rect 6638 46674 6690 46686
rect 6638 46610 6690 46622
rect 10222 46674 10274 46686
rect 10222 46610 10274 46622
rect 11678 46674 11730 46686
rect 11678 46610 11730 46622
rect 12014 46674 12066 46686
rect 14478 46674 14530 46686
rect 16270 46674 16322 46686
rect 21198 46674 21250 46686
rect 26462 46674 26514 46686
rect 28478 46674 28530 46686
rect 30606 46674 30658 46686
rect 12674 46622 12686 46674
rect 12738 46622 12750 46674
rect 13458 46622 13470 46674
rect 13522 46622 13534 46674
rect 14018 46622 14030 46674
rect 14082 46622 14094 46674
rect 15026 46622 15038 46674
rect 15090 46622 15102 46674
rect 15810 46622 15822 46674
rect 15874 46622 15886 46674
rect 19394 46622 19406 46674
rect 19458 46622 19470 46674
rect 20066 46622 20078 46674
rect 20130 46622 20142 46674
rect 20738 46622 20750 46674
rect 20802 46622 20814 46674
rect 22306 46622 22318 46674
rect 22370 46622 22382 46674
rect 23202 46622 23214 46674
rect 23266 46622 23278 46674
rect 25666 46622 25678 46674
rect 25730 46622 25742 46674
rect 27346 46622 27358 46674
rect 27410 46622 27422 46674
rect 29250 46622 29262 46674
rect 29314 46622 29326 46674
rect 12014 46610 12066 46622
rect 14478 46610 14530 46622
rect 16270 46610 16322 46622
rect 21198 46610 21250 46622
rect 26462 46610 26514 46622
rect 28478 46610 28530 46622
rect 30606 46610 30658 46622
rect 31166 46674 31218 46686
rect 31166 46610 31218 46622
rect 32174 46674 32226 46686
rect 32174 46610 32226 46622
rect 33070 46674 33122 46686
rect 40350 46674 40402 46686
rect 45614 46674 45666 46686
rect 35858 46622 35870 46674
rect 35922 46622 35934 46674
rect 44930 46622 44942 46674
rect 44994 46622 45006 46674
rect 33070 46610 33122 46622
rect 40350 46610 40402 46622
rect 45614 46610 45666 46622
rect 46622 46674 46674 46686
rect 46622 46610 46674 46622
rect 46846 46674 46898 46686
rect 47966 46674 48018 46686
rect 47282 46622 47294 46674
rect 47346 46622 47358 46674
rect 46846 46610 46898 46622
rect 47966 46610 48018 46622
rect 48078 46674 48130 46686
rect 48078 46610 48130 46622
rect 48862 46674 48914 46686
rect 49758 46674 49810 46686
rect 50542 46674 50594 46686
rect 49074 46622 49086 46674
rect 49138 46622 49150 46674
rect 50082 46622 50094 46674
rect 50146 46622 50158 46674
rect 48862 46610 48914 46622
rect 49758 46610 49810 46622
rect 50542 46610 50594 46622
rect 51774 46674 51826 46686
rect 51774 46610 51826 46622
rect 51886 46674 51938 46686
rect 51886 46610 51938 46622
rect 10446 46562 10498 46574
rect 10446 46498 10498 46510
rect 11230 46562 11282 46574
rect 11230 46498 11282 46510
rect 11902 46562 11954 46574
rect 11902 46498 11954 46510
rect 14254 46562 14306 46574
rect 14254 46498 14306 46510
rect 17390 46562 17442 46574
rect 17390 46498 17442 46510
rect 17614 46562 17666 46574
rect 24446 46562 24498 46574
rect 26238 46562 26290 46574
rect 19506 46510 19518 46562
rect 19570 46510 19582 46562
rect 22530 46510 22542 46562
rect 22594 46510 22606 46562
rect 22978 46510 22990 46562
rect 23042 46510 23054 46562
rect 25330 46510 25342 46562
rect 25394 46510 25406 46562
rect 17614 46498 17666 46510
rect 24446 46498 24498 46510
rect 26238 46498 26290 46510
rect 28142 46562 28194 46574
rect 28142 46498 28194 46510
rect 29822 46562 29874 46574
rect 34078 46562 34130 46574
rect 33506 46510 33518 46562
rect 33570 46510 33582 46562
rect 29822 46498 29874 46510
rect 34078 46498 34130 46510
rect 34526 46562 34578 46574
rect 34526 46498 34578 46510
rect 35646 46562 35698 46574
rect 44382 46562 44434 46574
rect 36642 46510 36654 46562
rect 36706 46510 36718 46562
rect 38770 46510 38782 46562
rect 38834 46510 38846 46562
rect 35646 46498 35698 46510
rect 44382 46498 44434 46510
rect 45278 46562 45330 46574
rect 45278 46498 45330 46510
rect 2158 46450 2210 46462
rect 2158 46386 2210 46398
rect 11566 46450 11618 46462
rect 11566 46386 11618 46398
rect 16382 46450 16434 46462
rect 16382 46386 16434 46398
rect 17950 46450 18002 46462
rect 17950 46386 18002 46398
rect 27134 46450 27186 46462
rect 27134 46386 27186 46398
rect 27694 46450 27746 46462
rect 27694 46386 27746 46398
rect 30158 46450 30210 46462
rect 30158 46386 30210 46398
rect 40910 46450 40962 46462
rect 40910 46386 40962 46398
rect 41246 46450 41298 46462
rect 41246 46386 41298 46398
rect 44606 46450 44658 46462
rect 44606 46386 44658 46398
rect 45390 46450 45442 46462
rect 45390 46386 45442 46398
rect 45726 46450 45778 46462
rect 45726 46386 45778 46398
rect 47742 46450 47794 46462
rect 47742 46386 47794 46398
rect 50318 46450 50370 46462
rect 50318 46386 50370 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 7758 46114 7810 46126
rect 7758 46050 7810 46062
rect 15150 46114 15202 46126
rect 15150 46050 15202 46062
rect 26126 46114 26178 46126
rect 26126 46050 26178 46062
rect 31278 46114 31330 46126
rect 31278 46050 31330 46062
rect 11902 46002 11954 46014
rect 1698 45950 1710 46002
rect 1762 45950 1774 46002
rect 3826 45950 3838 46002
rect 3890 45950 3902 46002
rect 11902 45938 11954 45950
rect 14254 46002 14306 46014
rect 18386 45950 18398 46002
rect 18450 45950 18462 46002
rect 19394 45950 19406 46002
rect 19458 45950 19470 46002
rect 22194 45950 22206 46002
rect 22258 45950 22270 46002
rect 24322 45950 24334 46002
rect 24386 45950 24398 46002
rect 26450 45950 26462 46002
rect 26514 45950 26526 46002
rect 29362 45950 29374 46002
rect 29426 45950 29438 46002
rect 31602 45950 31614 46002
rect 31666 45950 31678 46002
rect 34738 45950 34750 46002
rect 34802 45950 34814 46002
rect 38882 45950 38894 46002
rect 38946 45950 38958 46002
rect 39666 45950 39678 46002
rect 39730 45950 39742 46002
rect 41794 45950 41806 46002
rect 41858 45950 41870 46002
rect 46162 45950 46174 46002
rect 46226 45950 46238 46002
rect 48290 45950 48302 46002
rect 48354 45950 48366 46002
rect 14254 45938 14306 45950
rect 12574 45890 12626 45902
rect 4610 45838 4622 45890
rect 4674 45838 4686 45890
rect 5730 45838 5742 45890
rect 5794 45838 5806 45890
rect 6514 45838 6526 45890
rect 6578 45838 6590 45890
rect 6962 45838 6974 45890
rect 7026 45838 7038 45890
rect 12574 45826 12626 45838
rect 13694 45890 13746 45902
rect 20190 45890 20242 45902
rect 14578 45838 14590 45890
rect 14642 45838 14654 45890
rect 14802 45838 14814 45890
rect 14866 45838 14878 45890
rect 18162 45838 18174 45890
rect 18226 45838 18238 45890
rect 19058 45838 19070 45890
rect 19122 45838 19134 45890
rect 13694 45826 13746 45838
rect 20190 45826 20242 45838
rect 20750 45890 20802 45902
rect 26686 45890 26738 45902
rect 22418 45838 22430 45890
rect 22482 45838 22494 45890
rect 23538 45838 23550 45890
rect 23602 45838 23614 45890
rect 24098 45838 24110 45890
rect 24162 45838 24174 45890
rect 24546 45838 24558 45890
rect 24610 45838 24622 45890
rect 20750 45826 20802 45838
rect 26686 45826 26738 45838
rect 27134 45890 27186 45902
rect 27134 45826 27186 45838
rect 27358 45890 27410 45902
rect 27358 45826 27410 45838
rect 27806 45890 27858 45902
rect 35534 45890 35586 45902
rect 43038 45890 43090 45902
rect 29474 45838 29486 45890
rect 29538 45838 29550 45890
rect 30034 45838 30046 45890
rect 30098 45838 30110 45890
rect 30370 45838 30382 45890
rect 30434 45838 30446 45890
rect 33058 45838 33070 45890
rect 33122 45838 33134 45890
rect 38658 45838 38670 45890
rect 38722 45838 38734 45890
rect 42578 45838 42590 45890
rect 42642 45838 42654 45890
rect 45490 45838 45502 45890
rect 45554 45838 45566 45890
rect 49074 45838 49086 45890
rect 49138 45838 49150 45890
rect 27806 45826 27858 45838
rect 35534 45826 35586 45838
rect 43038 45826 43090 45838
rect 7198 45778 7250 45790
rect 5618 45726 5630 45778
rect 5682 45726 5694 45778
rect 7198 45714 7250 45726
rect 7534 45778 7586 45790
rect 7534 45714 7586 45726
rect 9774 45778 9826 45790
rect 9774 45714 9826 45726
rect 11454 45778 11506 45790
rect 15710 45778 15762 45790
rect 12898 45726 12910 45778
rect 12962 45726 12974 45778
rect 11454 45714 11506 45726
rect 15710 45714 15762 45726
rect 26350 45778 26402 45790
rect 26350 45714 26402 45726
rect 31502 45778 31554 45790
rect 31502 45714 31554 45726
rect 39342 45778 39394 45790
rect 39342 45714 39394 45726
rect 45726 45778 45778 45790
rect 45726 45714 45778 45726
rect 5070 45666 5122 45678
rect 5070 45602 5122 45614
rect 7646 45666 7698 45678
rect 7646 45602 7698 45614
rect 10110 45666 10162 45678
rect 10110 45602 10162 45614
rect 11118 45666 11170 45678
rect 11118 45602 11170 45614
rect 11342 45666 11394 45678
rect 11342 45602 11394 45614
rect 11790 45666 11842 45678
rect 11790 45602 11842 45614
rect 15038 45666 15090 45678
rect 15038 45602 15090 45614
rect 15822 45666 15874 45678
rect 15822 45602 15874 45614
rect 16046 45666 16098 45678
rect 16046 45602 16098 45614
rect 27246 45666 27298 45678
rect 27246 45602 27298 45614
rect 27694 45666 27746 45678
rect 27694 45602 27746 45614
rect 28366 45666 28418 45678
rect 28366 45602 28418 45614
rect 45054 45666 45106 45678
rect 45054 45602 45106 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 9662 45330 9714 45342
rect 13918 45330 13970 45342
rect 5394 45278 5406 45330
rect 5458 45278 5470 45330
rect 12338 45278 12350 45330
rect 12402 45278 12414 45330
rect 9662 45266 9714 45278
rect 13918 45266 13970 45278
rect 14254 45330 14306 45342
rect 14254 45266 14306 45278
rect 14478 45330 14530 45342
rect 14478 45266 14530 45278
rect 14814 45330 14866 45342
rect 14814 45266 14866 45278
rect 28366 45330 28418 45342
rect 28366 45266 28418 45278
rect 38334 45330 38386 45342
rect 38334 45266 38386 45278
rect 44942 45330 44994 45342
rect 44942 45266 44994 45278
rect 49198 45330 49250 45342
rect 49198 45266 49250 45278
rect 2830 45218 2882 45230
rect 2830 45154 2882 45166
rect 4286 45218 4338 45230
rect 4286 45154 4338 45166
rect 14702 45218 14754 45230
rect 18958 45218 19010 45230
rect 24558 45218 24610 45230
rect 26798 45218 26850 45230
rect 31950 45218 32002 45230
rect 16482 45166 16494 45218
rect 16546 45166 16558 45218
rect 17602 45166 17614 45218
rect 17666 45166 17678 45218
rect 19394 45166 19406 45218
rect 19458 45166 19470 45218
rect 21746 45166 21758 45218
rect 21810 45166 21822 45218
rect 22754 45166 22766 45218
rect 22818 45166 22830 45218
rect 25218 45166 25230 45218
rect 25282 45166 25294 45218
rect 29586 45166 29598 45218
rect 29650 45166 29662 45218
rect 30594 45166 30606 45218
rect 30658 45166 30670 45218
rect 14702 45154 14754 45166
rect 18958 45154 19010 45166
rect 24558 45154 24610 45166
rect 26798 45154 26850 45166
rect 31950 45154 32002 45166
rect 33966 45218 34018 45230
rect 40350 45218 40402 45230
rect 35186 45166 35198 45218
rect 35250 45166 35262 45218
rect 37986 45166 37998 45218
rect 38050 45166 38062 45218
rect 50306 45166 50318 45218
rect 50370 45166 50382 45218
rect 33966 45154 34018 45166
rect 40350 45154 40402 45166
rect 12014 45106 12066 45118
rect 1698 45054 1710 45106
rect 1762 45054 1774 45106
rect 3714 45054 3726 45106
rect 3778 45054 3790 45106
rect 5954 45054 5966 45106
rect 6018 45054 6030 45106
rect 10434 45054 10446 45106
rect 10498 45054 10510 45106
rect 10770 45054 10782 45106
rect 10834 45054 10846 45106
rect 12014 45042 12066 45054
rect 14142 45106 14194 45118
rect 19070 45106 19122 45118
rect 16706 45054 16718 45106
rect 16770 45054 16782 45106
rect 17378 45054 17390 45106
rect 17442 45054 17454 45106
rect 14142 45042 14194 45054
rect 19070 45042 19122 45054
rect 19742 45106 19794 45118
rect 19742 45042 19794 45054
rect 20078 45106 20130 45118
rect 20078 45042 20130 45054
rect 20302 45106 20354 45118
rect 20302 45042 20354 45054
rect 20974 45106 21026 45118
rect 24334 45106 24386 45118
rect 21186 45054 21198 45106
rect 21250 45054 21262 45106
rect 20974 45042 21026 45054
rect 24334 45042 24386 45054
rect 25566 45106 25618 45118
rect 27134 45106 27186 45118
rect 26002 45054 26014 45106
rect 26066 45054 26078 45106
rect 25566 45042 25618 45054
rect 27134 45042 27186 45054
rect 27470 45106 27522 45118
rect 27470 45042 27522 45054
rect 27694 45106 27746 45118
rect 27694 45042 27746 45054
rect 27918 45106 27970 45118
rect 27918 45042 27970 45054
rect 28590 45106 28642 45118
rect 33182 45106 33234 45118
rect 29250 45054 29262 45106
rect 29314 45054 29326 45106
rect 31042 45054 31054 45106
rect 31106 45054 31118 45106
rect 31378 45054 31390 45106
rect 31442 45054 31454 45106
rect 32274 45054 32286 45106
rect 32338 45054 32350 45106
rect 28590 45042 28642 45054
rect 33182 45042 33234 45054
rect 33518 45106 33570 45118
rect 33518 45042 33570 45054
rect 33742 45106 33794 45118
rect 33742 45042 33794 45054
rect 34190 45106 34242 45118
rect 34514 45054 34526 45106
rect 34578 45054 34590 45106
rect 39666 45054 39678 45106
rect 39730 45054 39742 45106
rect 41458 45054 41470 45106
rect 41522 45054 41534 45106
rect 49522 45054 49534 45106
rect 49586 45054 49598 45106
rect 34190 45042 34242 45054
rect 11790 44994 11842 45006
rect 6626 44942 6638 44994
rect 6690 44942 6702 44994
rect 8754 44942 8766 44994
rect 8818 44942 8830 44994
rect 10546 44942 10558 44994
rect 10610 44942 10622 44994
rect 11790 44930 11842 44942
rect 15374 44994 15426 45006
rect 15374 44930 15426 44942
rect 15934 44994 15986 45006
rect 27246 44994 27298 45006
rect 18050 44942 18062 44994
rect 18114 44942 18126 44994
rect 26338 44942 26350 44994
rect 26402 44942 26414 44994
rect 15934 44930 15986 44942
rect 27246 44930 27298 44942
rect 28142 44994 28194 45006
rect 32062 44994 32114 45006
rect 41134 44994 41186 45006
rect 28466 44942 28478 44994
rect 28530 44942 28542 44994
rect 29362 44942 29374 44994
rect 29426 44942 29438 44994
rect 31154 44942 31166 44994
rect 31218 44942 31230 44994
rect 37314 44942 37326 44994
rect 37378 44942 37390 44994
rect 40002 44942 40014 44994
rect 40066 44942 40078 44994
rect 42130 44942 42142 44994
rect 42194 44942 42206 44994
rect 44370 44942 44382 44994
rect 44434 44942 44446 44994
rect 52434 44942 52446 44994
rect 52498 44942 52510 44994
rect 28142 44930 28194 44942
rect 32062 44930 32114 44942
rect 41134 44930 41186 44942
rect 18958 44882 19010 44894
rect 10210 44830 10222 44882
rect 10274 44830 10286 44882
rect 15362 44830 15374 44882
rect 15426 44879 15438 44882
rect 15922 44879 15934 44882
rect 15426 44833 15934 44879
rect 15426 44830 15438 44833
rect 15922 44830 15934 44833
rect 15986 44830 15998 44882
rect 18958 44818 19010 44830
rect 20526 44882 20578 44894
rect 20526 44818 20578 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 2046 44546 2098 44558
rect 6190 44546 6242 44558
rect 3266 44494 3278 44546
rect 3330 44494 3342 44546
rect 2046 44482 2098 44494
rect 6190 44482 6242 44494
rect 6526 44546 6578 44558
rect 6526 44482 6578 44494
rect 17278 44546 17330 44558
rect 17278 44482 17330 44494
rect 23102 44546 23154 44558
rect 23102 44482 23154 44494
rect 23326 44546 23378 44558
rect 23326 44482 23378 44494
rect 30046 44546 30098 44558
rect 30046 44482 30098 44494
rect 34414 44546 34466 44558
rect 34414 44482 34466 44494
rect 2494 44434 2546 44446
rect 2494 44370 2546 44382
rect 4622 44434 4674 44446
rect 4622 44370 4674 44382
rect 7646 44434 7698 44446
rect 14030 44434 14082 44446
rect 10994 44382 11006 44434
rect 11058 44382 11070 44434
rect 12674 44382 12686 44434
rect 12738 44382 12750 44434
rect 7646 44370 7698 44382
rect 14030 44370 14082 44382
rect 17390 44434 17442 44446
rect 17390 44370 17442 44382
rect 23550 44434 23602 44446
rect 42366 44434 42418 44446
rect 48190 44434 48242 44446
rect 23874 44382 23886 44434
rect 23938 44382 23950 44434
rect 30930 44382 30942 44434
rect 30994 44382 31006 44434
rect 32610 44382 32622 44434
rect 32674 44382 32686 44434
rect 33618 44382 33630 44434
rect 33682 44382 33694 44434
rect 44818 44382 44830 44434
rect 44882 44382 44894 44434
rect 23550 44370 23602 44382
rect 42366 44370 42418 44382
rect 48190 44370 48242 44382
rect 2382 44322 2434 44334
rect 2382 44258 2434 44270
rect 2606 44322 2658 44334
rect 2606 44258 2658 44270
rect 3054 44322 3106 44334
rect 3054 44258 3106 44270
rect 3614 44322 3666 44334
rect 3614 44258 3666 44270
rect 3838 44322 3890 44334
rect 4398 44322 4450 44334
rect 4162 44270 4174 44322
rect 4226 44270 4238 44322
rect 3838 44258 3890 44270
rect 4398 44258 4450 44270
rect 6302 44322 6354 44334
rect 7422 44322 7474 44334
rect 11902 44322 11954 44334
rect 6738 44270 6750 44322
rect 6802 44270 6814 44322
rect 7074 44270 7086 44322
rect 7138 44270 7150 44322
rect 8194 44270 8206 44322
rect 8258 44270 8270 44322
rect 6302 44258 6354 44270
rect 7422 44258 7474 44270
rect 11902 44258 11954 44270
rect 13582 44322 13634 44334
rect 13582 44258 13634 44270
rect 13806 44322 13858 44334
rect 13806 44258 13858 44270
rect 14254 44322 14306 44334
rect 14254 44258 14306 44270
rect 14478 44322 14530 44334
rect 14478 44258 14530 44270
rect 15038 44322 15090 44334
rect 15038 44258 15090 44270
rect 15262 44322 15314 44334
rect 15262 44258 15314 44270
rect 16382 44322 16434 44334
rect 16382 44258 16434 44270
rect 16606 44322 16658 44334
rect 16606 44258 16658 44270
rect 16830 44322 16882 44334
rect 16830 44258 16882 44270
rect 17502 44322 17554 44334
rect 19294 44322 19346 44334
rect 18050 44270 18062 44322
rect 18114 44270 18126 44322
rect 18722 44270 18734 44322
rect 18786 44270 18798 44322
rect 17502 44258 17554 44270
rect 19294 44258 19346 44270
rect 19518 44322 19570 44334
rect 19518 44258 19570 44270
rect 19630 44322 19682 44334
rect 19630 44258 19682 44270
rect 20414 44322 20466 44334
rect 20414 44258 20466 44270
rect 21534 44322 21586 44334
rect 21534 44258 21586 44270
rect 22094 44322 22146 44334
rect 23998 44322 24050 44334
rect 25006 44322 25058 44334
rect 29710 44322 29762 44334
rect 22530 44270 22542 44322
rect 22594 44270 22606 44322
rect 24434 44270 24446 44322
rect 24498 44270 24510 44322
rect 25778 44270 25790 44322
rect 25842 44270 25854 44322
rect 26562 44270 26574 44322
rect 26626 44270 26638 44322
rect 26898 44270 26910 44322
rect 26962 44270 26974 44322
rect 29362 44270 29374 44322
rect 29426 44270 29438 44322
rect 22094 44258 22146 44270
rect 23998 44258 24050 44270
rect 25006 44258 25058 44270
rect 29710 44258 29762 44270
rect 29934 44322 29986 44334
rect 30830 44322 30882 44334
rect 30594 44270 30606 44322
rect 30658 44270 30670 44322
rect 29934 44258 29986 44270
rect 30830 44258 30882 44270
rect 31166 44322 31218 44334
rect 31166 44258 31218 44270
rect 31838 44322 31890 44334
rect 31838 44258 31890 44270
rect 33406 44322 33458 44334
rect 40126 44322 40178 44334
rect 40798 44322 40850 44334
rect 41694 44322 41746 44334
rect 38546 44270 38558 44322
rect 38610 44270 38622 44322
rect 39442 44270 39454 44322
rect 39506 44270 39518 44322
rect 39890 44270 39902 44322
rect 39954 44270 39966 44322
rect 40450 44270 40462 44322
rect 40514 44270 40526 44322
rect 41346 44270 41358 44322
rect 41410 44270 41422 44322
rect 33406 44258 33458 44270
rect 40126 44258 40178 44270
rect 40798 44258 40850 44270
rect 41694 44258 41746 44270
rect 42142 44322 42194 44334
rect 42142 44258 42194 44270
rect 42478 44322 42530 44334
rect 42478 44258 42530 44270
rect 42702 44322 42754 44334
rect 47618 44270 47630 44322
rect 47682 44270 47694 44322
rect 42702 44258 42754 44270
rect 1934 44210 1986 44222
rect 1934 44146 1986 44158
rect 4734 44210 4786 44222
rect 4734 44146 4786 44158
rect 5742 44210 5794 44222
rect 5742 44146 5794 44158
rect 5854 44210 5906 44222
rect 12350 44210 12402 44222
rect 8866 44158 8878 44210
rect 8930 44158 8942 44210
rect 5854 44146 5906 44158
rect 12350 44146 12402 44158
rect 12574 44210 12626 44222
rect 12574 44146 12626 44158
rect 15598 44210 15650 44222
rect 15598 44146 15650 44158
rect 16158 44210 16210 44222
rect 31614 44210 31666 44222
rect 17714 44158 17726 44210
rect 17778 44158 17790 44210
rect 25442 44158 25454 44210
rect 25506 44158 25518 44210
rect 27346 44158 27358 44210
rect 27410 44158 27422 44210
rect 16158 44146 16210 44158
rect 31614 44146 31666 44158
rect 32286 44210 32338 44222
rect 32286 44146 32338 44158
rect 33182 44210 33234 44222
rect 33182 44146 33234 44158
rect 33630 44210 33682 44222
rect 33630 44146 33682 44158
rect 34638 44210 34690 44222
rect 41806 44210 41858 44222
rect 38322 44158 38334 44210
rect 38386 44158 38398 44210
rect 46946 44158 46958 44210
rect 47010 44158 47022 44210
rect 34638 44146 34690 44158
rect 41806 44146 41858 44158
rect 11566 44098 11618 44110
rect 11566 44034 11618 44046
rect 13694 44098 13746 44110
rect 13694 44034 13746 44046
rect 14702 44098 14754 44110
rect 14702 44034 14754 44046
rect 14926 44098 14978 44110
rect 14926 44034 14978 44046
rect 15486 44098 15538 44110
rect 15486 44034 15538 44046
rect 20750 44098 20802 44110
rect 23774 44098 23826 44110
rect 22754 44046 22766 44098
rect 22818 44046 22830 44098
rect 20750 44034 20802 44046
rect 23774 44034 23826 44046
rect 24782 44098 24834 44110
rect 24782 44034 24834 44046
rect 24894 44098 24946 44110
rect 27806 44098 27858 44110
rect 27122 44046 27134 44098
rect 27186 44046 27198 44098
rect 24894 44034 24946 44046
rect 27806 44034 27858 44046
rect 28590 44098 28642 44110
rect 28590 44034 28642 44046
rect 29038 44098 29090 44110
rect 29038 44034 29090 44046
rect 29150 44098 29202 44110
rect 29150 44034 29202 44046
rect 30382 44098 30434 44110
rect 30382 44034 30434 44046
rect 31390 44098 31442 44110
rect 31390 44034 31442 44046
rect 32510 44098 32562 44110
rect 32510 44034 32562 44046
rect 33742 44098 33794 44110
rect 33742 44034 33794 44046
rect 34526 44098 34578 44110
rect 34526 44034 34578 44046
rect 37550 44098 37602 44110
rect 37550 44034 37602 44046
rect 40910 44098 40962 44110
rect 40910 44034 40962 44046
rect 41022 44098 41074 44110
rect 41022 44034 41074 44046
rect 41918 44098 41970 44110
rect 41918 44034 41970 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 12126 43762 12178 43774
rect 12126 43698 12178 43710
rect 15710 43762 15762 43774
rect 24334 43762 24386 43774
rect 21746 43710 21758 43762
rect 21810 43710 21822 43762
rect 15710 43698 15762 43710
rect 24334 43698 24386 43710
rect 27582 43762 27634 43774
rect 27582 43698 27634 43710
rect 29262 43762 29314 43774
rect 29262 43698 29314 43710
rect 34190 43762 34242 43774
rect 34190 43698 34242 43710
rect 48190 43762 48242 43774
rect 48190 43698 48242 43710
rect 5070 43650 5122 43662
rect 3826 43598 3838 43650
rect 3890 43598 3902 43650
rect 5070 43586 5122 43598
rect 5182 43650 5234 43662
rect 10110 43650 10162 43662
rect 5618 43598 5630 43650
rect 5682 43598 5694 43650
rect 5182 43586 5234 43598
rect 10110 43586 10162 43598
rect 11118 43650 11170 43662
rect 11118 43586 11170 43598
rect 11678 43650 11730 43662
rect 11678 43586 11730 43598
rect 12350 43650 12402 43662
rect 17614 43650 17666 43662
rect 14802 43598 14814 43650
rect 14866 43598 14878 43650
rect 12350 43586 12402 43598
rect 17614 43586 17666 43598
rect 17726 43650 17778 43662
rect 17726 43586 17778 43598
rect 20862 43650 20914 43662
rect 24222 43650 24274 43662
rect 28030 43650 28082 43662
rect 23090 43598 23102 43650
rect 23154 43598 23166 43650
rect 25330 43598 25342 43650
rect 25394 43598 25406 43650
rect 26338 43598 26350 43650
rect 26402 43598 26414 43650
rect 20862 43586 20914 43598
rect 24222 43586 24274 43598
rect 28030 43586 28082 43598
rect 28254 43650 28306 43662
rect 33966 43650 34018 43662
rect 39006 43650 39058 43662
rect 29586 43598 29598 43650
rect 29650 43598 29662 43650
rect 33394 43598 33406 43650
rect 33458 43598 33470 43650
rect 35634 43598 35646 43650
rect 35698 43598 35710 43650
rect 28254 43586 28306 43598
rect 33966 43586 34018 43598
rect 39006 43586 39058 43598
rect 39230 43650 39282 43662
rect 39230 43586 39282 43598
rect 39678 43650 39730 43662
rect 39678 43586 39730 43598
rect 40238 43650 40290 43662
rect 40238 43586 40290 43598
rect 46510 43650 46562 43662
rect 46510 43586 46562 43598
rect 47070 43650 47122 43662
rect 47070 43586 47122 43598
rect 52110 43650 52162 43662
rect 52110 43586 52162 43598
rect 5966 43538 6018 43550
rect 10446 43538 10498 43550
rect 11230 43538 11282 43550
rect 4610 43486 4622 43538
rect 4674 43486 4686 43538
rect 6850 43486 6862 43538
rect 6914 43486 6926 43538
rect 10658 43486 10670 43538
rect 10722 43486 10734 43538
rect 5966 43474 6018 43486
rect 10446 43474 10498 43486
rect 11230 43474 11282 43486
rect 12798 43538 12850 43550
rect 12798 43474 12850 43486
rect 13022 43538 13074 43550
rect 14030 43538 14082 43550
rect 13794 43486 13806 43538
rect 13858 43486 13870 43538
rect 13022 43474 13074 43486
rect 14030 43474 14082 43486
rect 14254 43538 14306 43550
rect 14254 43474 14306 43486
rect 15150 43538 15202 43550
rect 15150 43474 15202 43486
rect 16158 43538 16210 43550
rect 16158 43474 16210 43486
rect 16606 43538 16658 43550
rect 18286 43538 18338 43550
rect 21646 43538 21698 43550
rect 23774 43538 23826 43550
rect 17938 43486 17950 43538
rect 18002 43486 18014 43538
rect 19058 43486 19070 43538
rect 19122 43486 19134 43538
rect 19842 43486 19854 43538
rect 19906 43486 19918 43538
rect 23426 43486 23438 43538
rect 23490 43486 23502 43538
rect 16606 43474 16658 43486
rect 18286 43474 18338 43486
rect 21646 43474 21698 43486
rect 23774 43474 23826 43486
rect 24446 43538 24498 43550
rect 27806 43538 27858 43550
rect 25666 43486 25678 43538
rect 25730 43486 25742 43538
rect 26114 43486 26126 43538
rect 26178 43486 26190 43538
rect 27010 43486 27022 43538
rect 27074 43486 27086 43538
rect 24446 43474 24498 43486
rect 27806 43474 27858 43486
rect 28478 43538 28530 43550
rect 31726 43538 31778 43550
rect 29810 43486 29822 43538
rect 29874 43486 29886 43538
rect 30594 43486 30606 43538
rect 30658 43486 30670 43538
rect 31266 43486 31278 43538
rect 31330 43486 31342 43538
rect 28478 43474 28530 43486
rect 31726 43474 31778 43486
rect 33070 43538 33122 43550
rect 33070 43474 33122 43486
rect 33854 43538 33906 43550
rect 38894 43538 38946 43550
rect 40350 43538 40402 43550
rect 45614 43538 45666 43550
rect 51998 43538 52050 43550
rect 34850 43486 34862 43538
rect 34914 43486 34926 43538
rect 39442 43486 39454 43538
rect 39506 43486 39518 43538
rect 40786 43486 40798 43538
rect 40850 43486 40862 43538
rect 41570 43486 41582 43538
rect 41634 43486 41646 43538
rect 44930 43486 44942 43538
rect 44994 43486 45006 43538
rect 45938 43486 45950 43538
rect 46002 43486 46014 43538
rect 48850 43486 48862 43538
rect 48914 43486 48926 43538
rect 33854 43474 33906 43486
rect 38894 43474 38946 43486
rect 40350 43474 40402 43486
rect 45614 43474 45666 43486
rect 51998 43474 52050 43486
rect 4958 43426 5010 43438
rect 9886 43426 9938 43438
rect 1698 43374 1710 43426
rect 1762 43374 1774 43426
rect 8194 43374 8206 43426
rect 8258 43374 8270 43426
rect 4958 43362 5010 43374
rect 9886 43362 9938 43374
rect 12238 43426 12290 43438
rect 12238 43362 12290 43374
rect 12910 43426 12962 43438
rect 12910 43362 12962 43374
rect 13246 43426 13298 43438
rect 13246 43362 13298 43374
rect 16830 43426 16882 43438
rect 16830 43362 16882 43374
rect 19518 43426 19570 43438
rect 34526 43426 34578 43438
rect 47518 43426 47570 43438
rect 23314 43374 23326 43426
rect 23378 43374 23390 43426
rect 37762 43374 37774 43426
rect 37826 43374 37838 43426
rect 41794 43374 41806 43426
rect 41858 43374 41870 43426
rect 44706 43374 44718 43426
rect 44770 43374 44782 43426
rect 49522 43374 49534 43426
rect 49586 43374 49598 43426
rect 51650 43374 51662 43426
rect 51714 43374 51726 43426
rect 19518 43362 19570 43374
rect 34526 43362 34578 43374
rect 47518 43362 47570 43374
rect 10222 43314 10274 43326
rect 10222 43250 10274 43262
rect 11118 43314 11170 43326
rect 11118 43250 11170 43262
rect 13470 43314 13522 43326
rect 13470 43250 13522 43262
rect 14366 43314 14418 43326
rect 14366 43250 14418 43262
rect 16382 43314 16434 43326
rect 16382 43250 16434 43262
rect 28366 43314 28418 43326
rect 39790 43314 39842 43326
rect 30930 43262 30942 43314
rect 30994 43262 31006 43314
rect 28366 43250 28418 43262
rect 39790 43250 39842 43262
rect 40238 43314 40290 43326
rect 46174 43314 46226 43326
rect 41906 43262 41918 43314
rect 41970 43262 41982 43314
rect 40238 43250 40290 43262
rect 46174 43250 46226 43262
rect 46398 43314 46450 43326
rect 46398 43250 46450 43262
rect 52110 43314 52162 43326
rect 52110 43250 52162 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 11790 42978 11842 42990
rect 16382 42978 16434 42990
rect 3602 42926 3614 42978
rect 3666 42926 3678 42978
rect 14354 42926 14366 42978
rect 14418 42975 14430 42978
rect 15026 42975 15038 42978
rect 14418 42929 15038 42975
rect 14418 42926 14430 42929
rect 15026 42926 15038 42929
rect 15090 42926 15102 42978
rect 11790 42914 11842 42926
rect 16382 42914 16434 42926
rect 18174 42978 18226 42990
rect 18174 42914 18226 42926
rect 18510 42978 18562 42990
rect 18510 42914 18562 42926
rect 19182 42978 19234 42990
rect 19182 42914 19234 42926
rect 27806 42978 27858 42990
rect 27806 42914 27858 42926
rect 34302 42978 34354 42990
rect 34302 42914 34354 42926
rect 52782 42978 52834 42990
rect 52782 42914 52834 42926
rect 4174 42866 4226 42878
rect 4174 42802 4226 42814
rect 5742 42866 5794 42878
rect 11566 42866 11618 42878
rect 8866 42814 8878 42866
rect 8930 42814 8942 42866
rect 10994 42814 11006 42866
rect 11058 42814 11070 42866
rect 5742 42802 5794 42814
rect 11566 42802 11618 42814
rect 13694 42866 13746 42878
rect 13694 42802 13746 42814
rect 15038 42866 15090 42878
rect 15038 42802 15090 42814
rect 15710 42866 15762 42878
rect 15710 42802 15762 42814
rect 18622 42866 18674 42878
rect 18622 42802 18674 42814
rect 22990 42866 23042 42878
rect 22990 42802 23042 42814
rect 27358 42866 27410 42878
rect 27358 42802 27410 42814
rect 29598 42866 29650 42878
rect 29598 42802 29650 42814
rect 35422 42866 35474 42878
rect 35422 42802 35474 42814
rect 50542 42866 50594 42878
rect 50542 42802 50594 42814
rect 3950 42754 4002 42766
rect 12798 42754 12850 42766
rect 8194 42702 8206 42754
rect 8258 42702 8270 42754
rect 3950 42690 4002 42702
rect 12798 42690 12850 42702
rect 13582 42754 13634 42766
rect 13582 42690 13634 42702
rect 14254 42754 14306 42766
rect 14254 42690 14306 42702
rect 21310 42754 21362 42766
rect 21310 42690 21362 42702
rect 21870 42754 21922 42766
rect 21870 42690 21922 42702
rect 22878 42754 22930 42766
rect 22878 42690 22930 42702
rect 23102 42754 23154 42766
rect 24334 42754 24386 42766
rect 23874 42702 23886 42754
rect 23938 42702 23950 42754
rect 23102 42690 23154 42702
rect 24334 42690 24386 42702
rect 25566 42754 25618 42766
rect 25566 42690 25618 42702
rect 27918 42754 27970 42766
rect 29710 42754 29762 42766
rect 29138 42702 29150 42754
rect 29202 42702 29214 42754
rect 27918 42690 27970 42702
rect 29710 42690 29762 42702
rect 30382 42754 30434 42766
rect 30382 42690 30434 42702
rect 30718 42754 30770 42766
rect 30718 42690 30770 42702
rect 34526 42754 34578 42766
rect 40238 42754 40290 42766
rect 35858 42702 35870 42754
rect 35922 42702 35934 42754
rect 34526 42690 34578 42702
rect 40238 42690 40290 42702
rect 40574 42754 40626 42766
rect 40574 42690 40626 42702
rect 40798 42754 40850 42766
rect 42254 42754 42306 42766
rect 41906 42702 41918 42754
rect 41970 42702 41982 42754
rect 40798 42690 40850 42702
rect 42254 42690 42306 42702
rect 43038 42754 43090 42766
rect 49870 42754 49922 42766
rect 48850 42702 48862 42754
rect 48914 42702 48926 42754
rect 49074 42702 49086 42754
rect 49138 42702 49150 42754
rect 43038 42690 43090 42702
rect 49870 42690 49922 42702
rect 50766 42754 50818 42766
rect 50766 42690 50818 42702
rect 52670 42754 52722 42766
rect 52670 42690 52722 42702
rect 12462 42642 12514 42654
rect 12462 42578 12514 42590
rect 16494 42642 16546 42654
rect 16494 42578 16546 42590
rect 16942 42642 16994 42654
rect 16942 42578 16994 42590
rect 17838 42642 17890 42654
rect 17838 42578 17890 42590
rect 18062 42642 18114 42654
rect 18062 42578 18114 42590
rect 19294 42642 19346 42654
rect 19294 42578 19346 42590
rect 24446 42642 24498 42654
rect 24446 42578 24498 42590
rect 25230 42642 25282 42654
rect 25230 42578 25282 42590
rect 25342 42642 25394 42654
rect 25342 42578 25394 42590
rect 25790 42642 25842 42654
rect 25790 42578 25842 42590
rect 27806 42642 27858 42654
rect 27806 42578 27858 42590
rect 30494 42642 30546 42654
rect 30494 42578 30546 42590
rect 34862 42642 34914 42654
rect 34862 42578 34914 42590
rect 36990 42642 37042 42654
rect 36990 42578 37042 42590
rect 40350 42642 40402 42654
rect 40350 42578 40402 42590
rect 40910 42642 40962 42654
rect 40910 42578 40962 42590
rect 42814 42642 42866 42654
rect 42814 42578 42866 42590
rect 46062 42642 46114 42654
rect 46062 42578 46114 42590
rect 49310 42642 49362 42654
rect 51438 42642 51490 42654
rect 51090 42590 51102 42642
rect 51154 42590 51166 42642
rect 49310 42578 49362 42590
rect 51438 42578 51490 42590
rect 51662 42642 51714 42654
rect 51662 42578 51714 42590
rect 51998 42642 52050 42654
rect 51998 42578 52050 42590
rect 4958 42530 5010 42542
rect 12574 42530 12626 42542
rect 12114 42478 12126 42530
rect 12178 42478 12190 42530
rect 4958 42466 5010 42478
rect 12574 42466 12626 42478
rect 13806 42530 13858 42542
rect 13806 42466 13858 42478
rect 14702 42530 14754 42542
rect 14702 42466 14754 42478
rect 16270 42530 16322 42542
rect 16270 42466 16322 42478
rect 16718 42530 16770 42542
rect 16718 42466 16770 42478
rect 17502 42530 17554 42542
rect 17502 42466 17554 42478
rect 18734 42530 18786 42542
rect 18734 42466 18786 42478
rect 22654 42530 22706 42542
rect 22654 42466 22706 42478
rect 25902 42530 25954 42542
rect 25902 42466 25954 42478
rect 29486 42530 29538 42542
rect 29486 42466 29538 42478
rect 32622 42530 32674 42542
rect 32622 42466 32674 42478
rect 33966 42530 34018 42542
rect 33966 42466 34018 42478
rect 34750 42530 34802 42542
rect 34750 42466 34802 42478
rect 34974 42530 35026 42542
rect 34974 42466 35026 42478
rect 36430 42530 36482 42542
rect 36430 42466 36482 42478
rect 37102 42530 37154 42542
rect 37102 42466 37154 42478
rect 37214 42530 37266 42542
rect 37214 42466 37266 42478
rect 41134 42530 41186 42542
rect 41134 42466 41186 42478
rect 42366 42530 42418 42542
rect 42366 42466 42418 42478
rect 42478 42530 42530 42542
rect 45614 42530 45666 42542
rect 43362 42478 43374 42530
rect 43426 42478 43438 42530
rect 42478 42466 42530 42478
rect 45614 42466 45666 42478
rect 47406 42530 47458 42542
rect 51774 42530 51826 42542
rect 47730 42478 47742 42530
rect 47794 42478 47806 42530
rect 50194 42478 50206 42530
rect 50258 42478 50270 42530
rect 47406 42466 47458 42478
rect 51774 42466 51826 42478
rect 52782 42530 52834 42542
rect 52782 42466 52834 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 14590 42194 14642 42206
rect 11554 42142 11566 42194
rect 11618 42142 11630 42194
rect 12898 42142 12910 42194
rect 12962 42142 12974 42194
rect 14590 42130 14642 42142
rect 16270 42194 16322 42206
rect 16270 42130 16322 42142
rect 16718 42194 16770 42206
rect 16718 42130 16770 42142
rect 17614 42194 17666 42206
rect 17614 42130 17666 42142
rect 20750 42194 20802 42206
rect 22990 42194 23042 42206
rect 22194 42142 22206 42194
rect 22258 42142 22270 42194
rect 20750 42130 20802 42142
rect 22990 42130 23042 42142
rect 23998 42194 24050 42206
rect 23998 42130 24050 42142
rect 24110 42194 24162 42206
rect 24110 42130 24162 42142
rect 26910 42194 26962 42206
rect 26910 42130 26962 42142
rect 27134 42194 27186 42206
rect 27134 42130 27186 42142
rect 27918 42194 27970 42206
rect 27918 42130 27970 42142
rect 28142 42194 28194 42206
rect 31950 42194 32002 42206
rect 31154 42142 31166 42194
rect 31218 42142 31230 42194
rect 28142 42130 28194 42142
rect 31950 42130 32002 42142
rect 32174 42194 32226 42206
rect 32174 42130 32226 42142
rect 35422 42194 35474 42206
rect 35422 42130 35474 42142
rect 41806 42194 41858 42206
rect 53106 42142 53118 42194
rect 53170 42142 53182 42194
rect 41806 42130 41858 42142
rect 16830 42082 16882 42094
rect 19742 42082 19794 42094
rect 12786 42030 12798 42082
rect 12850 42030 12862 42082
rect 18386 42030 18398 42082
rect 18450 42030 18462 42082
rect 16830 42018 16882 42030
rect 19742 42018 19794 42030
rect 20638 42082 20690 42094
rect 20638 42018 20690 42030
rect 25118 42082 25170 42094
rect 25118 42018 25170 42030
rect 25342 42082 25394 42094
rect 25342 42018 25394 42030
rect 25454 42082 25506 42094
rect 25454 42018 25506 42030
rect 25902 42082 25954 42094
rect 25902 42018 25954 42030
rect 26350 42082 26402 42094
rect 26350 42018 26402 42030
rect 26798 42082 26850 42094
rect 29822 42082 29874 42094
rect 28914 42030 28926 42082
rect 28978 42030 28990 42082
rect 26798 42018 26850 42030
rect 29822 42018 29874 42030
rect 33294 42082 33346 42094
rect 33294 42018 33346 42030
rect 39790 42082 39842 42094
rect 39790 42018 39842 42030
rect 40126 42082 40178 42094
rect 40126 42018 40178 42030
rect 40238 42082 40290 42094
rect 40238 42018 40290 42030
rect 53006 42082 53058 42094
rect 53778 42030 53790 42082
rect 53842 42030 53854 42082
rect 53006 42018 53058 42030
rect 8878 41970 8930 41982
rect 1810 41918 1822 41970
rect 1874 41918 1886 41970
rect 8418 41918 8430 41970
rect 8482 41918 8494 41970
rect 8878 41906 8930 41918
rect 9662 41970 9714 41982
rect 9662 41906 9714 41918
rect 11006 41970 11058 41982
rect 11006 41906 11058 41918
rect 11230 41970 11282 41982
rect 11230 41906 11282 41918
rect 12462 41970 12514 41982
rect 12462 41906 12514 41918
rect 13246 41970 13298 41982
rect 13246 41906 13298 41918
rect 13470 41970 13522 41982
rect 13470 41906 13522 41918
rect 14142 41970 14194 41982
rect 14142 41906 14194 41918
rect 15486 41970 15538 41982
rect 15486 41906 15538 41918
rect 15934 41970 15986 41982
rect 15934 41906 15986 41918
rect 16158 41970 16210 41982
rect 16158 41906 16210 41918
rect 16494 41970 16546 41982
rect 16494 41906 16546 41918
rect 17390 41970 17442 41982
rect 17390 41906 17442 41918
rect 17502 41970 17554 41982
rect 20302 41970 20354 41982
rect 17938 41918 17950 41970
rect 18002 41918 18014 41970
rect 18834 41918 18846 41970
rect 18898 41918 18910 41970
rect 19954 41918 19966 41970
rect 20018 41918 20030 41970
rect 17502 41906 17554 41918
rect 20302 41906 20354 41918
rect 21646 41970 21698 41982
rect 21646 41906 21698 41918
rect 22430 41970 22482 41982
rect 23886 41970 23938 41982
rect 22754 41918 22766 41970
rect 22818 41918 22830 41970
rect 22430 41906 22482 41918
rect 23886 41906 23938 41918
rect 24558 41970 24610 41982
rect 24558 41906 24610 41918
rect 25790 41970 25842 41982
rect 25790 41906 25842 41918
rect 26462 41970 26514 41982
rect 26462 41906 26514 41918
rect 27694 41970 27746 41982
rect 27694 41906 27746 41918
rect 28366 41970 28418 41982
rect 28366 41906 28418 41918
rect 29262 41970 29314 41982
rect 29262 41906 29314 41918
rect 30830 41970 30882 41982
rect 30830 41906 30882 41918
rect 31502 41970 31554 41982
rect 31502 41906 31554 41918
rect 31726 41970 31778 41982
rect 31726 41906 31778 41918
rect 32062 41970 32114 41982
rect 32062 41906 32114 41918
rect 34190 41970 34242 41982
rect 34190 41906 34242 41918
rect 34750 41970 34802 41982
rect 34750 41906 34802 41918
rect 35198 41970 35250 41982
rect 39230 41970 39282 41982
rect 35746 41918 35758 41970
rect 35810 41918 35822 41970
rect 36530 41918 36542 41970
rect 36594 41918 36606 41970
rect 38994 41918 39006 41970
rect 39058 41918 39070 41970
rect 35198 41906 35250 41918
rect 39230 41906 39282 41918
rect 39678 41970 39730 41982
rect 39678 41906 39730 41918
rect 40462 41970 40514 41982
rect 40462 41906 40514 41918
rect 41694 41970 41746 41982
rect 42242 41918 42254 41970
rect 42306 41918 42318 41970
rect 43362 41918 43374 41970
rect 43426 41918 43438 41970
rect 44146 41918 44158 41970
rect 44210 41918 44222 41970
rect 45042 41918 45054 41970
rect 45106 41918 45118 41970
rect 45490 41918 45502 41970
rect 45554 41918 45566 41970
rect 49410 41918 49422 41970
rect 49474 41918 49486 41970
rect 49746 41918 49758 41970
rect 49810 41918 49822 41970
rect 51762 41918 51774 41970
rect 51826 41918 51838 41970
rect 52322 41918 52334 41970
rect 52386 41918 52398 41970
rect 52770 41918 52782 41970
rect 52834 41918 52846 41970
rect 53666 41918 53678 41970
rect 53730 41918 53742 41970
rect 41694 41906 41746 41918
rect 5518 41858 5570 41870
rect 12238 41858 12290 41870
rect 2482 41806 2494 41858
rect 2546 41806 2558 41858
rect 4610 41806 4622 41858
rect 4674 41806 4686 41858
rect 4946 41806 4958 41858
rect 5010 41806 5022 41858
rect 6066 41806 6078 41858
rect 6130 41806 6142 41858
rect 5518 41794 5570 41806
rect 12238 41794 12290 41806
rect 14702 41858 14754 41870
rect 19406 41858 19458 41870
rect 18946 41806 18958 41858
rect 19010 41806 19022 41858
rect 14702 41794 14754 41806
rect 19406 41794 19458 41806
rect 20078 41858 20130 41870
rect 33182 41858 33234 41870
rect 29922 41806 29934 41858
rect 29986 41806 29998 41858
rect 20078 41794 20130 41806
rect 33182 41794 33234 41806
rect 34526 41858 34578 41870
rect 34526 41794 34578 41806
rect 35310 41858 35362 41870
rect 47182 41858 47234 41870
rect 38658 41806 38670 41858
rect 38722 41806 38734 41858
rect 46722 41806 46734 41858
rect 46786 41806 46798 41858
rect 48738 41806 48750 41858
rect 48802 41806 48814 41858
rect 50754 41806 50766 41858
rect 50818 41806 50830 41858
rect 35310 41794 35362 41806
rect 47182 41794 47234 41806
rect 5294 41746 5346 41758
rect 5294 41682 5346 41694
rect 13022 41746 13074 41758
rect 13022 41682 13074 41694
rect 14254 41746 14306 41758
rect 14254 41682 14306 41694
rect 15374 41746 15426 41758
rect 15374 41682 15426 41694
rect 20862 41746 20914 41758
rect 20862 41682 20914 41694
rect 21870 41746 21922 41758
rect 21870 41682 21922 41694
rect 23102 41746 23154 41758
rect 23102 41682 23154 41694
rect 26350 41746 26402 41758
rect 26350 41682 26402 41694
rect 27806 41746 27858 41758
rect 27806 41682 27858 41694
rect 29598 41746 29650 41758
rect 29598 41682 29650 41694
rect 33070 41746 33122 41758
rect 39454 41746 39506 41758
rect 34178 41694 34190 41746
rect 34242 41743 34254 41746
rect 34626 41743 34638 41746
rect 34242 41697 34638 41743
rect 34242 41694 34254 41697
rect 34626 41694 34638 41697
rect 34690 41694 34702 41746
rect 33070 41682 33122 41694
rect 39454 41682 39506 41694
rect 41806 41746 41858 41758
rect 41806 41682 41858 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 2942 41410 2994 41422
rect 2942 41346 2994 41358
rect 6862 41410 6914 41422
rect 18286 41410 18338 41422
rect 17938 41358 17950 41410
rect 18002 41358 18014 41410
rect 6862 41346 6914 41358
rect 18286 41346 18338 41358
rect 18622 41410 18674 41422
rect 18622 41346 18674 41358
rect 19294 41410 19346 41422
rect 19294 41346 19346 41358
rect 19966 41410 20018 41422
rect 19966 41346 20018 41358
rect 22094 41410 22146 41422
rect 39566 41410 39618 41422
rect 23314 41358 23326 41410
rect 23378 41358 23390 41410
rect 26786 41358 26798 41410
rect 26850 41358 26862 41410
rect 22094 41346 22146 41358
rect 39566 41346 39618 41358
rect 39902 41410 39954 41422
rect 39902 41346 39954 41358
rect 49870 41410 49922 41422
rect 52782 41410 52834 41422
rect 51986 41358 51998 41410
rect 52050 41358 52062 41410
rect 49870 41346 49922 41358
rect 52782 41346 52834 41358
rect 4958 41298 5010 41310
rect 23774 41298 23826 41310
rect 8978 41246 8990 41298
rect 9042 41246 9054 41298
rect 11106 41246 11118 41298
rect 11170 41246 11182 41298
rect 4958 41234 5010 41246
rect 23774 41234 23826 41246
rect 24558 41298 24610 41310
rect 39230 41298 39282 41310
rect 48638 41298 48690 41310
rect 25890 41246 25902 41298
rect 25954 41246 25966 41298
rect 29922 41246 29934 41298
rect 29986 41246 29998 41298
rect 32722 41246 32734 41298
rect 32786 41246 32798 41298
rect 34850 41246 34862 41298
rect 34914 41246 34926 41298
rect 45154 41246 45166 41298
rect 45218 41246 45230 41298
rect 24558 41234 24610 41246
rect 39230 41234 39282 41246
rect 48638 41234 48690 41246
rect 3278 41186 3330 41198
rect 3278 41122 3330 41134
rect 3726 41186 3778 41198
rect 3726 41122 3778 41134
rect 3838 41186 3890 41198
rect 3838 41122 3890 41134
rect 4286 41186 4338 41198
rect 6190 41186 6242 41198
rect 5954 41134 5966 41186
rect 6018 41134 6030 41186
rect 4286 41122 4338 41134
rect 6190 41122 6242 41134
rect 6414 41186 6466 41198
rect 6414 41122 6466 41134
rect 6974 41186 7026 41198
rect 14142 41186 14194 41198
rect 8306 41134 8318 41186
rect 8370 41134 8382 41186
rect 6974 41122 7026 41134
rect 14142 41122 14194 41134
rect 14478 41186 14530 41198
rect 14478 41122 14530 41134
rect 15038 41186 15090 41198
rect 15038 41122 15090 41134
rect 16046 41186 16098 41198
rect 16046 41122 16098 41134
rect 16270 41186 16322 41198
rect 16270 41122 16322 41134
rect 16494 41186 16546 41198
rect 16494 41122 16546 41134
rect 16942 41186 16994 41198
rect 16942 41122 16994 41134
rect 17390 41186 17442 41198
rect 22766 41186 22818 41198
rect 18274 41134 18286 41186
rect 18338 41134 18350 41186
rect 19954 41134 19966 41186
rect 20018 41134 20030 41186
rect 20402 41134 20414 41186
rect 20466 41134 20478 41186
rect 17390 41122 17442 41134
rect 22766 41122 22818 41134
rect 22878 41186 22930 41198
rect 22878 41122 22930 41134
rect 23998 41186 24050 41198
rect 23998 41122 24050 41134
rect 24110 41186 24162 41198
rect 24110 41122 24162 41134
rect 24670 41186 24722 41198
rect 26574 41186 26626 41198
rect 27918 41186 27970 41198
rect 25442 41134 25454 41186
rect 25506 41134 25518 41186
rect 25666 41134 25678 41186
rect 25730 41134 25742 41186
rect 26898 41134 26910 41186
rect 26962 41134 26974 41186
rect 24670 41122 24722 41134
rect 26574 41122 26626 41134
rect 27918 41122 27970 41134
rect 28590 41186 28642 41198
rect 28590 41122 28642 41134
rect 29150 41186 29202 41198
rect 30270 41186 30322 41198
rect 35198 41186 35250 41198
rect 29810 41134 29822 41186
rect 29874 41134 29886 41186
rect 31938 41134 31950 41186
rect 32002 41134 32014 41186
rect 29150 41122 29202 41134
rect 30270 41122 30322 41134
rect 35198 41122 35250 41134
rect 35534 41186 35586 41198
rect 35534 41122 35586 41134
rect 36990 41186 37042 41198
rect 48974 41186 49026 41198
rect 42914 41134 42926 41186
rect 42978 41134 42990 41186
rect 43250 41134 43262 41186
rect 43314 41134 43326 41186
rect 48066 41134 48078 41186
rect 48130 41134 48142 41186
rect 36990 41122 37042 41134
rect 48974 41122 49026 41134
rect 50318 41186 50370 41198
rect 50318 41122 50370 41134
rect 50542 41186 50594 41198
rect 51438 41186 51490 41198
rect 51202 41134 51214 41186
rect 51266 41134 51278 41186
rect 50542 41122 50594 41134
rect 51438 41122 51490 41134
rect 51550 41186 51602 41198
rect 51550 41122 51602 41134
rect 3054 41074 3106 41086
rect 3054 41010 3106 41022
rect 4846 41074 4898 41086
rect 4846 41010 4898 41022
rect 5070 41074 5122 41086
rect 5070 41010 5122 41022
rect 6526 41074 6578 41086
rect 6526 41010 6578 41022
rect 7086 41074 7138 41086
rect 7086 41010 7138 41022
rect 15150 41074 15202 41086
rect 15150 41010 15202 41022
rect 17278 41074 17330 41086
rect 17278 41010 17330 41022
rect 17502 41074 17554 41086
rect 17502 41010 17554 41022
rect 18958 41074 19010 41086
rect 18958 41010 19010 41022
rect 19630 41074 19682 41086
rect 19630 41010 19682 41022
rect 20638 41074 20690 41086
rect 20638 41010 20690 41022
rect 22094 41074 22146 41086
rect 22094 41010 22146 41022
rect 22206 41074 22258 41086
rect 22206 41010 22258 41022
rect 22654 41074 22706 41086
rect 22654 41010 22706 41022
rect 23662 41074 23714 41086
rect 23662 41010 23714 41022
rect 28478 41074 28530 41086
rect 28478 41010 28530 41022
rect 29486 41074 29538 41086
rect 35758 41074 35810 41086
rect 30594 41022 30606 41074
rect 30658 41022 30670 41074
rect 29486 41010 29538 41022
rect 35758 41010 35810 41022
rect 36430 41074 36482 41086
rect 36430 41010 36482 41022
rect 37102 41074 37154 41086
rect 39790 41074 39842 41086
rect 38434 41022 38446 41074
rect 38498 41022 38510 41074
rect 37102 41010 37154 41022
rect 39790 41010 39842 41022
rect 41582 41074 41634 41086
rect 44270 41074 44322 41086
rect 49870 41074 49922 41086
rect 42578 41022 42590 41074
rect 42642 41022 42654 41074
rect 47282 41022 47294 41074
rect 47346 41022 47358 41074
rect 41582 41010 41634 41022
rect 44270 41010 44322 41022
rect 49870 41010 49922 41022
rect 49982 41074 50034 41086
rect 49982 41010 50034 41022
rect 52894 41074 52946 41086
rect 52894 41010 52946 41022
rect 3614 40962 3666 40974
rect 3614 40898 3666 40910
rect 7870 40962 7922 40974
rect 7870 40898 7922 40910
rect 14030 40962 14082 40974
rect 14030 40898 14082 40910
rect 14590 40962 14642 40974
rect 14590 40898 14642 40910
rect 14814 40962 14866 40974
rect 14814 40898 14866 40910
rect 15374 40962 15426 40974
rect 15374 40898 15426 40910
rect 16382 40962 16434 40974
rect 16382 40898 16434 40910
rect 19182 40962 19234 40974
rect 19182 40898 19234 40910
rect 28366 40962 28418 40974
rect 28366 40898 28418 40910
rect 29374 40962 29426 40974
rect 29374 40898 29426 40910
rect 35646 40962 35698 40974
rect 35646 40898 35698 40910
rect 36206 40962 36258 40974
rect 36206 40898 36258 40910
rect 36318 40962 36370 40974
rect 36318 40898 36370 40910
rect 37214 40962 37266 40974
rect 37214 40898 37266 40910
rect 37438 40962 37490 40974
rect 37438 40898 37490 40910
rect 38110 40962 38162 40974
rect 38110 40898 38162 40910
rect 38782 40962 38834 40974
rect 38782 40898 38834 40910
rect 41470 40962 41522 40974
rect 41470 40898 41522 40910
rect 41694 40962 41746 40974
rect 41694 40898 41746 40910
rect 41918 40962 41970 40974
rect 44158 40962 44210 40974
rect 43474 40910 43486 40962
rect 43538 40910 43550 40962
rect 43698 40910 43710 40962
rect 43762 40910 43774 40962
rect 41918 40898 41970 40910
rect 44158 40898 44210 40910
rect 49534 40962 49586 40974
rect 52782 40962 52834 40974
rect 50866 40910 50878 40962
rect 50930 40910 50942 40962
rect 49534 40898 49586 40910
rect 52782 40898 52834 40910
rect 53342 40962 53394 40974
rect 53342 40898 53394 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 4510 40626 4562 40638
rect 4510 40562 4562 40574
rect 11342 40626 11394 40638
rect 11342 40562 11394 40574
rect 11678 40626 11730 40638
rect 17614 40626 17666 40638
rect 15474 40574 15486 40626
rect 15538 40574 15550 40626
rect 11678 40562 11730 40574
rect 17614 40562 17666 40574
rect 21198 40626 21250 40638
rect 21198 40562 21250 40574
rect 22318 40626 22370 40638
rect 22318 40562 22370 40574
rect 22654 40626 22706 40638
rect 22654 40562 22706 40574
rect 24110 40626 24162 40638
rect 24110 40562 24162 40574
rect 25790 40626 25842 40638
rect 25790 40562 25842 40574
rect 28366 40626 28418 40638
rect 28366 40562 28418 40574
rect 28926 40626 28978 40638
rect 28926 40562 28978 40574
rect 29150 40626 29202 40638
rect 29150 40562 29202 40574
rect 29822 40626 29874 40638
rect 34526 40626 34578 40638
rect 31826 40574 31838 40626
rect 31890 40574 31902 40626
rect 29822 40562 29874 40574
rect 34526 40562 34578 40574
rect 45278 40626 45330 40638
rect 45278 40562 45330 40574
rect 46510 40626 46562 40638
rect 46510 40562 46562 40574
rect 46846 40626 46898 40638
rect 46846 40562 46898 40574
rect 47630 40626 47682 40638
rect 47630 40562 47682 40574
rect 49198 40626 49250 40638
rect 49198 40562 49250 40574
rect 51438 40626 51490 40638
rect 51438 40562 51490 40574
rect 53790 40626 53842 40638
rect 53790 40562 53842 40574
rect 13246 40514 13298 40526
rect 7634 40462 7646 40514
rect 7698 40462 7710 40514
rect 12002 40462 12014 40514
rect 12066 40462 12078 40514
rect 12674 40462 12686 40514
rect 12738 40462 12750 40514
rect 13246 40450 13298 40462
rect 13470 40514 13522 40526
rect 18510 40514 18562 40526
rect 16146 40462 16158 40514
rect 16210 40462 16222 40514
rect 13470 40450 13522 40462
rect 18510 40450 18562 40462
rect 22094 40514 22146 40526
rect 22094 40450 22146 40462
rect 25566 40514 25618 40526
rect 25566 40450 25618 40462
rect 26014 40514 26066 40526
rect 26014 40450 26066 40462
rect 27358 40514 27410 40526
rect 27358 40450 27410 40462
rect 27582 40514 27634 40526
rect 27582 40450 27634 40462
rect 27918 40514 27970 40526
rect 42142 40514 42194 40526
rect 30146 40462 30158 40514
rect 30210 40462 30222 40514
rect 30930 40462 30942 40514
rect 30994 40462 31006 40514
rect 32498 40462 32510 40514
rect 32562 40462 32574 40514
rect 35634 40462 35646 40514
rect 35698 40462 35710 40514
rect 40002 40462 40014 40514
rect 40066 40462 40078 40514
rect 27918 40450 27970 40462
rect 42142 40450 42194 40462
rect 44942 40514 44994 40526
rect 51886 40514 51938 40526
rect 46162 40462 46174 40514
rect 46226 40462 46238 40514
rect 47170 40462 47182 40514
rect 47234 40462 47246 40514
rect 44942 40450 44994 40462
rect 51886 40450 51938 40462
rect 52446 40514 52498 40526
rect 52446 40450 52498 40462
rect 4846 40402 4898 40414
rect 12350 40402 12402 40414
rect 8306 40350 8318 40402
rect 8370 40350 8382 40402
rect 4846 40338 4898 40350
rect 12350 40338 12402 40350
rect 13582 40402 13634 40414
rect 13582 40338 13634 40350
rect 13806 40402 13858 40414
rect 13806 40338 13858 40350
rect 14030 40402 14082 40414
rect 14030 40338 14082 40350
rect 14590 40402 14642 40414
rect 14590 40338 14642 40350
rect 14926 40402 14978 40414
rect 17950 40402 18002 40414
rect 15922 40350 15934 40402
rect 15986 40350 15998 40402
rect 14926 40338 14978 40350
rect 17950 40338 18002 40350
rect 19294 40402 19346 40414
rect 19294 40338 19346 40350
rect 19966 40402 20018 40414
rect 19966 40338 20018 40350
rect 21422 40402 21474 40414
rect 21422 40338 21474 40350
rect 21534 40402 21586 40414
rect 21534 40338 21586 40350
rect 21646 40402 21698 40414
rect 21646 40338 21698 40350
rect 21982 40402 22034 40414
rect 21982 40338 22034 40350
rect 22542 40402 22594 40414
rect 25454 40402 25506 40414
rect 24322 40350 24334 40402
rect 24386 40350 24398 40402
rect 22542 40338 22594 40350
rect 25454 40338 25506 40350
rect 26350 40402 26402 40414
rect 28702 40402 28754 40414
rect 31950 40402 32002 40414
rect 40350 40402 40402 40414
rect 44270 40402 44322 40414
rect 28130 40350 28142 40402
rect 28194 40350 28206 40402
rect 31378 40350 31390 40402
rect 31442 40350 31454 40402
rect 34850 40350 34862 40402
rect 34914 40350 34926 40402
rect 41458 40350 41470 40402
rect 41522 40350 41534 40402
rect 41906 40350 41918 40402
rect 41970 40350 41982 40402
rect 42690 40350 42702 40402
rect 42754 40350 42766 40402
rect 26350 40338 26402 40350
rect 28702 40338 28754 40350
rect 31950 40338 32002 40350
rect 40350 40338 40402 40350
rect 44270 40338 44322 40350
rect 44718 40402 44770 40414
rect 44718 40338 44770 40350
rect 45838 40402 45890 40414
rect 45838 40338 45890 40350
rect 48078 40402 48130 40414
rect 48078 40338 48130 40350
rect 48974 40402 49026 40414
rect 48974 40338 49026 40350
rect 49198 40402 49250 40414
rect 49198 40338 49250 40350
rect 49534 40402 49586 40414
rect 49534 40338 49586 40350
rect 50766 40402 50818 40414
rect 50766 40338 50818 40350
rect 50878 40402 50930 40414
rect 50878 40338 50930 40350
rect 51326 40402 51378 40414
rect 51326 40338 51378 40350
rect 51550 40402 51602 40414
rect 51550 40338 51602 40350
rect 52110 40402 52162 40414
rect 52110 40338 52162 40350
rect 53454 40402 53506 40414
rect 53454 40338 53506 40350
rect 8878 40290 8930 40302
rect 5506 40238 5518 40290
rect 5570 40238 5582 40290
rect 8878 40226 8930 40238
rect 19406 40290 19458 40302
rect 19406 40226 19458 40238
rect 26238 40290 26290 40302
rect 26238 40226 26290 40238
rect 27470 40290 27522 40302
rect 27470 40226 27522 40238
rect 28814 40290 28866 40302
rect 44494 40290 44546 40302
rect 37762 40238 37774 40290
rect 37826 40238 37838 40290
rect 43138 40238 43150 40290
rect 43202 40238 43214 40290
rect 28814 40226 28866 40238
rect 44494 40226 44546 40238
rect 49982 40290 50034 40302
rect 49982 40226 50034 40238
rect 52334 40290 52386 40302
rect 52334 40226 52386 40238
rect 52894 40290 52946 40302
rect 52894 40226 52946 40238
rect 4510 40178 4562 40190
rect 4510 40114 4562 40126
rect 4622 40178 4674 40190
rect 4622 40114 4674 40126
rect 15150 40178 15202 40190
rect 15150 40114 15202 40126
rect 19630 40178 19682 40190
rect 19630 40114 19682 40126
rect 19854 40178 19906 40190
rect 19854 40114 19906 40126
rect 23998 40178 24050 40190
rect 23998 40114 24050 40126
rect 28478 40178 28530 40190
rect 28478 40114 28530 40126
rect 43934 40178 43986 40190
rect 43934 40114 43986 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 5742 39842 5794 39854
rect 5742 39778 5794 39790
rect 27022 39842 27074 39854
rect 27022 39778 27074 39790
rect 14366 39730 14418 39742
rect 2482 39678 2494 39730
rect 2546 39678 2558 39730
rect 4610 39678 4622 39730
rect 4674 39678 4686 39730
rect 6514 39678 6526 39730
rect 6578 39678 6590 39730
rect 9426 39678 9438 39730
rect 9490 39678 9502 39730
rect 11554 39678 11566 39730
rect 11618 39678 11630 39730
rect 14366 39666 14418 39678
rect 17390 39730 17442 39742
rect 17390 39666 17442 39678
rect 19070 39730 19122 39742
rect 26350 39730 26402 39742
rect 34750 39730 34802 39742
rect 21746 39678 21758 39730
rect 21810 39678 21822 39730
rect 34290 39678 34302 39730
rect 34354 39678 34366 39730
rect 19070 39666 19122 39678
rect 26350 39666 26402 39678
rect 34750 39666 34802 39678
rect 36430 39730 36482 39742
rect 48974 39730 49026 39742
rect 50542 39730 50594 39742
rect 37762 39678 37774 39730
rect 37826 39678 37838 39730
rect 39890 39678 39902 39730
rect 39954 39678 39966 39730
rect 41682 39678 41694 39730
rect 41746 39678 41758 39730
rect 42802 39678 42814 39730
rect 42866 39678 42878 39730
rect 45602 39678 45614 39730
rect 45666 39678 45678 39730
rect 48178 39678 48190 39730
rect 48242 39678 48254 39730
rect 50194 39678 50206 39730
rect 50258 39678 50270 39730
rect 52658 39678 52670 39730
rect 52722 39678 52734 39730
rect 54786 39678 54798 39730
rect 54850 39678 54862 39730
rect 36430 39666 36482 39678
rect 48974 39666 49026 39678
rect 50542 39666 50594 39678
rect 5518 39618 5570 39630
rect 14254 39618 14306 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 8642 39566 8654 39618
rect 8706 39566 8718 39618
rect 5518 39554 5570 39566
rect 14254 39554 14306 39566
rect 14926 39618 14978 39630
rect 26910 39618 26962 39630
rect 16930 39566 16942 39618
rect 16994 39566 17006 39618
rect 19394 39566 19406 39618
rect 19458 39566 19470 39618
rect 25218 39566 25230 39618
rect 25282 39566 25294 39618
rect 14926 39554 14978 39566
rect 26910 39554 26962 39566
rect 27582 39618 27634 39630
rect 27582 39554 27634 39566
rect 27918 39618 27970 39630
rect 46062 39618 46114 39630
rect 28242 39566 28254 39618
rect 28306 39566 28318 39618
rect 31490 39566 31502 39618
rect 31554 39566 31566 39618
rect 37090 39566 37102 39618
rect 37154 39566 37166 39618
rect 41346 39566 41358 39618
rect 41410 39566 41422 39618
rect 42578 39566 42590 39618
rect 42642 39566 42654 39618
rect 45378 39566 45390 39618
rect 45442 39566 45454 39618
rect 27918 39554 27970 39566
rect 46062 39554 46114 39566
rect 46286 39618 46338 39630
rect 46286 39554 46338 39566
rect 46734 39618 46786 39630
rect 46734 39554 46786 39566
rect 46846 39618 46898 39630
rect 50878 39618 50930 39630
rect 48514 39566 48526 39618
rect 48578 39566 48590 39618
rect 49858 39566 49870 39618
rect 49922 39566 49934 39618
rect 55458 39566 55470 39618
rect 55522 39566 55534 39618
rect 46846 39554 46898 39566
rect 50878 39554 50930 39566
rect 6638 39506 6690 39518
rect 6638 39442 6690 39454
rect 6862 39506 6914 39518
rect 7534 39506 7586 39518
rect 7186 39454 7198 39506
rect 7250 39454 7262 39506
rect 6862 39442 6914 39454
rect 7534 39442 7586 39454
rect 15150 39506 15202 39518
rect 15150 39442 15202 39454
rect 15486 39506 15538 39518
rect 15486 39442 15538 39454
rect 16606 39506 16658 39518
rect 16606 39442 16658 39454
rect 19966 39506 20018 39518
rect 19966 39442 20018 39454
rect 21534 39506 21586 39518
rect 26798 39506 26850 39518
rect 22530 39454 22542 39506
rect 22594 39454 22606 39506
rect 25442 39454 25454 39506
rect 25506 39454 25518 39506
rect 21534 39442 21586 39454
rect 26798 39442 26850 39454
rect 27694 39506 27746 39518
rect 42030 39506 42082 39518
rect 28466 39454 28478 39506
rect 28530 39454 28542 39506
rect 32162 39454 32174 39506
rect 32226 39454 32238 39506
rect 27694 39442 27746 39454
rect 42030 39442 42082 39454
rect 43486 39506 43538 39518
rect 51090 39454 51102 39506
rect 51154 39454 51166 39506
rect 51874 39454 51886 39506
rect 51938 39454 51950 39506
rect 43486 39442 43538 39454
rect 5070 39394 5122 39406
rect 5070 39330 5122 39342
rect 5854 39394 5906 39406
rect 5854 39330 5906 39342
rect 6078 39394 6130 39406
rect 6078 39330 6130 39342
rect 8318 39394 8370 39406
rect 8318 39330 8370 39342
rect 14478 39394 14530 39406
rect 14478 39330 14530 39342
rect 16158 39394 16210 39406
rect 16158 39330 16210 39342
rect 16718 39394 16770 39406
rect 16718 39330 16770 39342
rect 17278 39394 17330 39406
rect 17278 39330 17330 39342
rect 18062 39394 18114 39406
rect 18062 39330 18114 39342
rect 19518 39394 19570 39406
rect 19518 39330 19570 39342
rect 20078 39394 20130 39406
rect 20078 39330 20130 39342
rect 20750 39394 20802 39406
rect 20750 39330 20802 39342
rect 22206 39394 22258 39406
rect 22206 39330 22258 39342
rect 23438 39394 23490 39406
rect 23438 39330 23490 39342
rect 25902 39394 25954 39406
rect 25902 39330 25954 39342
rect 44270 39394 44322 39406
rect 44270 39330 44322 39342
rect 46622 39394 46674 39406
rect 46622 39330 46674 39342
rect 47518 39394 47570 39406
rect 51426 39342 51438 39394
rect 51490 39342 51502 39394
rect 47518 39330 47570 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 4398 39058 4450 39070
rect 7646 39058 7698 39070
rect 5954 39006 5966 39058
rect 6018 39006 6030 39058
rect 6290 39006 6302 39058
rect 6354 39006 6366 39058
rect 4398 38994 4450 39006
rect 7646 38994 7698 39006
rect 7758 39058 7810 39070
rect 7758 38994 7810 39006
rect 11678 39058 11730 39070
rect 11678 38994 11730 39006
rect 15150 39058 15202 39070
rect 15150 38994 15202 39006
rect 15710 39058 15762 39070
rect 15710 38994 15762 39006
rect 21758 39058 21810 39070
rect 26126 39058 26178 39070
rect 23986 39006 23998 39058
rect 24050 39006 24062 39058
rect 25554 39006 25566 39058
rect 25618 39006 25630 39058
rect 21758 38994 21810 39006
rect 26126 38994 26178 39006
rect 26910 39058 26962 39070
rect 26910 38994 26962 39006
rect 28366 39058 28418 39070
rect 29150 39058 29202 39070
rect 28690 39006 28702 39058
rect 28754 39006 28766 39058
rect 28366 38994 28418 39006
rect 29150 38994 29202 39006
rect 31614 39058 31666 39070
rect 31614 38994 31666 39006
rect 32286 39058 32338 39070
rect 32286 38994 32338 39006
rect 33182 39058 33234 39070
rect 33182 38994 33234 39006
rect 42142 39058 42194 39070
rect 43822 39058 43874 39070
rect 43026 39006 43038 39058
rect 43090 39006 43102 39058
rect 42142 38994 42194 39006
rect 43822 38994 43874 39006
rect 44046 39058 44098 39070
rect 44046 38994 44098 39006
rect 45614 39058 45666 39070
rect 45614 38994 45666 39006
rect 45726 39058 45778 39070
rect 45726 38994 45778 39006
rect 46286 39058 46338 39070
rect 46286 38994 46338 39006
rect 48302 39058 48354 39070
rect 48302 38994 48354 39006
rect 49870 39058 49922 39070
rect 49870 38994 49922 39006
rect 49982 39058 50034 39070
rect 49982 38994 50034 39006
rect 50094 39058 50146 39070
rect 50094 38994 50146 39006
rect 3726 38946 3778 38958
rect 3042 38894 3054 38946
rect 3106 38894 3118 38946
rect 3726 38882 3778 38894
rect 3950 38946 4002 38958
rect 3950 38882 4002 38894
rect 4510 38946 4562 38958
rect 4510 38882 4562 38894
rect 5406 38946 5458 38958
rect 5406 38882 5458 38894
rect 5518 38946 5570 38958
rect 5518 38882 5570 38894
rect 14814 38946 14866 38958
rect 14814 38882 14866 38894
rect 15934 38946 15986 38958
rect 15934 38882 15986 38894
rect 17390 38946 17442 38958
rect 17390 38882 17442 38894
rect 17726 38946 17778 38958
rect 17726 38882 17778 38894
rect 17950 38946 18002 38958
rect 26014 38946 26066 38958
rect 18834 38894 18846 38946
rect 18898 38894 18910 38946
rect 19842 38894 19854 38946
rect 19906 38894 19918 38946
rect 17950 38882 18002 38894
rect 26014 38882 26066 38894
rect 33294 38946 33346 38958
rect 33294 38882 33346 38894
rect 37102 38946 37154 38958
rect 37102 38882 37154 38894
rect 37886 38946 37938 38958
rect 37886 38882 37938 38894
rect 38446 38946 38498 38958
rect 38446 38882 38498 38894
rect 43710 38946 43762 38958
rect 43710 38882 43762 38894
rect 44270 38946 44322 38958
rect 44270 38882 44322 38894
rect 46510 38946 46562 38958
rect 46510 38882 46562 38894
rect 48078 38946 48130 38958
rect 48078 38882 48130 38894
rect 49198 38946 49250 38958
rect 49198 38882 49250 38894
rect 3390 38834 3442 38846
rect 2818 38782 2830 38834
rect 2882 38782 2894 38834
rect 3390 38770 3442 38782
rect 3502 38834 3554 38846
rect 3502 38770 3554 38782
rect 4286 38834 4338 38846
rect 6638 38834 6690 38846
rect 4834 38782 4846 38834
rect 4898 38782 4910 38834
rect 5170 38782 5182 38834
rect 5234 38782 5246 38834
rect 4286 38770 4338 38782
rect 6638 38770 6690 38782
rect 6862 38834 6914 38846
rect 6862 38770 6914 38782
rect 7086 38834 7138 38846
rect 7086 38770 7138 38782
rect 7534 38834 7586 38846
rect 13358 38834 13410 38846
rect 12338 38782 12350 38834
rect 12402 38782 12414 38834
rect 12562 38782 12574 38834
rect 12626 38782 12638 38834
rect 7534 38770 7586 38782
rect 13358 38770 13410 38782
rect 15038 38834 15090 38846
rect 15038 38770 15090 38782
rect 16606 38834 16658 38846
rect 16606 38770 16658 38782
rect 16830 38834 16882 38846
rect 21422 38834 21474 38846
rect 19506 38782 19518 38834
rect 19570 38782 19582 38834
rect 16830 38770 16882 38782
rect 21422 38770 21474 38782
rect 22094 38834 22146 38846
rect 23662 38834 23714 38846
rect 22418 38782 22430 38834
rect 22482 38782 22494 38834
rect 22978 38782 22990 38834
rect 23042 38782 23054 38834
rect 22094 38770 22146 38782
rect 23662 38770 23714 38782
rect 24446 38834 24498 38846
rect 24446 38770 24498 38782
rect 25230 38834 25282 38846
rect 25230 38770 25282 38782
rect 27246 38834 27298 38846
rect 32062 38834 32114 38846
rect 27682 38782 27694 38834
rect 27746 38782 27758 38834
rect 30818 38782 30830 38834
rect 30882 38782 30894 38834
rect 27246 38770 27298 38782
rect 32062 38770 32114 38782
rect 32174 38834 32226 38846
rect 32174 38770 32226 38782
rect 32622 38834 32674 38846
rect 32622 38770 32674 38782
rect 32958 38834 33010 38846
rect 32958 38770 33010 38782
rect 37774 38834 37826 38846
rect 37774 38770 37826 38782
rect 38334 38834 38386 38846
rect 38334 38770 38386 38782
rect 38670 38834 38722 38846
rect 38670 38770 38722 38782
rect 42478 38834 42530 38846
rect 42478 38770 42530 38782
rect 42702 38834 42754 38846
rect 42702 38770 42754 38782
rect 45166 38834 45218 38846
rect 45166 38770 45218 38782
rect 45838 38834 45890 38846
rect 45838 38770 45890 38782
rect 46846 38834 46898 38846
rect 46846 38770 46898 38782
rect 47406 38834 47458 38846
rect 47406 38770 47458 38782
rect 47966 38834 48018 38846
rect 47966 38770 48018 38782
rect 49310 38834 49362 38846
rect 49522 38782 49534 38834
rect 49586 38782 49598 38834
rect 50418 38782 50430 38834
rect 50482 38782 50494 38834
rect 54002 38782 54014 38834
rect 54066 38782 54078 38834
rect 49310 38770 49362 38782
rect 17502 38722 17554 38734
rect 37214 38722 37266 38734
rect 13010 38670 13022 38722
rect 13074 38670 13086 38722
rect 15586 38670 15598 38722
rect 15650 38670 15662 38722
rect 30482 38670 30494 38722
rect 30546 38670 30558 38722
rect 17502 38658 17554 38670
rect 37214 38658 37266 38670
rect 37326 38722 37378 38734
rect 47070 38722 47122 38734
rect 44594 38670 44606 38722
rect 44658 38670 44670 38722
rect 37326 38658 37378 38670
rect 47070 38658 47122 38670
rect 47630 38722 47682 38734
rect 51090 38670 51102 38722
rect 51154 38670 51166 38722
rect 53218 38670 53230 38722
rect 53282 38670 53294 38722
rect 47630 38658 47682 38670
rect 15150 38610 15202 38622
rect 20526 38610 20578 38622
rect 16258 38558 16270 38610
rect 16322 38558 16334 38610
rect 15150 38546 15202 38558
rect 20526 38546 20578 38558
rect 26126 38610 26178 38622
rect 26126 38546 26178 38558
rect 37886 38610 37938 38622
rect 37886 38546 37938 38558
rect 46622 38610 46674 38622
rect 48738 38558 48750 38610
rect 48802 38558 48814 38610
rect 46622 38546 46674 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 31614 38274 31666 38286
rect 50866 38222 50878 38274
rect 50930 38222 50942 38274
rect 31614 38210 31666 38222
rect 5070 38162 5122 38174
rect 13694 38162 13746 38174
rect 18734 38162 18786 38174
rect 2482 38110 2494 38162
rect 2546 38110 2558 38162
rect 4610 38110 4622 38162
rect 4674 38110 4686 38162
rect 6066 38110 6078 38162
rect 6130 38110 6142 38162
rect 8194 38110 8206 38162
rect 8258 38110 8270 38162
rect 10770 38110 10782 38162
rect 10834 38110 10846 38162
rect 12898 38110 12910 38162
rect 12962 38110 12974 38162
rect 17154 38110 17166 38162
rect 17218 38110 17230 38162
rect 5070 38098 5122 38110
rect 13694 38098 13746 38110
rect 18734 38098 18786 38110
rect 21310 38162 21362 38174
rect 21310 38098 21362 38110
rect 23886 38162 23938 38174
rect 36206 38162 36258 38174
rect 44270 38162 44322 38174
rect 25330 38110 25342 38162
rect 25394 38110 25406 38162
rect 27458 38110 27470 38162
rect 27522 38110 27534 38162
rect 38882 38110 38894 38162
rect 38946 38110 38958 38162
rect 40114 38110 40126 38162
rect 40178 38110 40190 38162
rect 23886 38098 23938 38110
rect 36206 38098 36258 38110
rect 44270 38098 44322 38110
rect 45054 38162 45106 38174
rect 45054 38098 45106 38110
rect 14366 38050 14418 38062
rect 1810 37998 1822 38050
rect 1874 37998 1886 38050
rect 8866 37998 8878 38050
rect 8930 37998 8942 38050
rect 10098 37998 10110 38050
rect 10162 37998 10174 38050
rect 14366 37986 14418 37998
rect 14814 38050 14866 38062
rect 14814 37986 14866 37998
rect 15038 38050 15090 38062
rect 19854 38050 19906 38062
rect 15250 37998 15262 38050
rect 15314 37998 15326 38050
rect 15810 37998 15822 38050
rect 15874 37998 15886 38050
rect 15038 37986 15090 37998
rect 19854 37986 19906 37998
rect 22654 38050 22706 38062
rect 29486 38050 29538 38062
rect 23202 37998 23214 38050
rect 23266 37998 23278 38050
rect 23650 37998 23662 38050
rect 23714 37998 23726 38050
rect 28130 37998 28142 38050
rect 28194 37998 28206 38050
rect 22654 37986 22706 37998
rect 29486 37986 29538 37998
rect 31054 38050 31106 38062
rect 31054 37986 31106 37998
rect 31278 38050 31330 38062
rect 31278 37986 31330 37998
rect 34078 38050 34130 38062
rect 34078 37986 34130 37998
rect 34526 38050 34578 38062
rect 43374 38050 43426 38062
rect 38322 37998 38334 38050
rect 38386 37998 38398 38050
rect 39218 37998 39230 38050
rect 39282 37998 39294 38050
rect 42914 37998 42926 38050
rect 42978 37998 42990 38050
rect 34526 37986 34578 37998
rect 43374 37986 43426 37998
rect 44158 38050 44210 38062
rect 44158 37986 44210 37998
rect 44830 38050 44882 38062
rect 44830 37986 44882 37998
rect 45278 38050 45330 38062
rect 45278 37986 45330 37998
rect 45390 38050 45442 38062
rect 45390 37986 45442 37998
rect 45838 38050 45890 38062
rect 45838 37986 45890 37998
rect 46622 38050 46674 38062
rect 49534 38050 49586 38062
rect 51326 38050 51378 38062
rect 52670 38050 52722 38062
rect 47618 37998 47630 38050
rect 47682 37998 47694 38050
rect 48850 37998 48862 38050
rect 48914 37998 48926 38050
rect 50194 37998 50206 38050
rect 50258 37998 50270 38050
rect 51762 37998 51774 38050
rect 51826 37998 51838 38050
rect 53106 37998 53118 38050
rect 53170 37998 53182 38050
rect 46622 37986 46674 37998
rect 49534 37986 49586 37998
rect 51326 37986 51378 37998
rect 52670 37986 52722 37998
rect 13582 37938 13634 37950
rect 13582 37874 13634 37886
rect 14030 37938 14082 37950
rect 14030 37874 14082 37886
rect 14590 37938 14642 37950
rect 14590 37874 14642 37886
rect 18622 37938 18674 37950
rect 18622 37874 18674 37886
rect 19182 37938 19234 37950
rect 19182 37874 19234 37886
rect 24222 37938 24274 37950
rect 24222 37874 24274 37886
rect 24334 37938 24386 37950
rect 24334 37874 24386 37886
rect 24446 37938 24498 37950
rect 24446 37874 24498 37886
rect 29822 37938 29874 37950
rect 29822 37874 29874 37886
rect 30382 37938 30434 37950
rect 30382 37874 30434 37886
rect 30718 37938 30770 37950
rect 30718 37874 30770 37886
rect 33742 37938 33794 37950
rect 43710 37938 43762 37950
rect 37650 37886 37662 37938
rect 37714 37886 37726 37938
rect 42242 37886 42254 37938
rect 42306 37886 42318 37938
rect 33742 37874 33794 37886
rect 43710 37874 43762 37886
rect 44942 37938 44994 37950
rect 44942 37874 44994 37886
rect 9438 37826 9490 37838
rect 9438 37762 9490 37774
rect 14142 37826 14194 37838
rect 14142 37762 14194 37774
rect 14926 37826 14978 37838
rect 14926 37762 14978 37774
rect 19294 37826 19346 37838
rect 19294 37762 19346 37774
rect 19518 37826 19570 37838
rect 19518 37762 19570 37774
rect 19742 37826 19794 37838
rect 19742 37762 19794 37774
rect 20302 37826 20354 37838
rect 20302 37762 20354 37774
rect 21870 37826 21922 37838
rect 21870 37762 21922 37774
rect 25118 37826 25170 37838
rect 25118 37762 25170 37774
rect 33966 37826 34018 37838
rect 33966 37762 34018 37774
rect 34190 37826 34242 37838
rect 34190 37762 34242 37774
rect 34638 37826 34690 37838
rect 34638 37762 34690 37774
rect 34750 37826 34802 37838
rect 34750 37762 34802 37774
rect 46174 37826 46226 37838
rect 46174 37762 46226 37774
rect 47070 37826 47122 37838
rect 47070 37762 47122 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 4398 37490 4450 37502
rect 4398 37426 4450 37438
rect 15822 37490 15874 37502
rect 15822 37426 15874 37438
rect 16158 37490 16210 37502
rect 16158 37426 16210 37438
rect 16382 37490 16434 37502
rect 16382 37426 16434 37438
rect 21422 37490 21474 37502
rect 25342 37490 25394 37502
rect 24434 37438 24446 37490
rect 24498 37438 24510 37490
rect 21422 37426 21474 37438
rect 25342 37426 25394 37438
rect 25790 37490 25842 37502
rect 25790 37426 25842 37438
rect 27022 37490 27074 37502
rect 27022 37426 27074 37438
rect 30830 37490 30882 37502
rect 36430 37490 36482 37502
rect 39678 37490 39730 37502
rect 31490 37438 31502 37490
rect 31554 37438 31566 37490
rect 37650 37438 37662 37490
rect 37714 37438 37726 37490
rect 30830 37426 30882 37438
rect 36430 37426 36482 37438
rect 39678 37426 39730 37438
rect 41022 37490 41074 37502
rect 47630 37490 47682 37502
rect 44594 37438 44606 37490
rect 44658 37438 44670 37490
rect 41022 37426 41074 37438
rect 47630 37426 47682 37438
rect 53790 37490 53842 37502
rect 53790 37426 53842 37438
rect 4622 37378 4674 37390
rect 4622 37314 4674 37326
rect 4846 37378 4898 37390
rect 4846 37314 4898 37326
rect 14702 37378 14754 37390
rect 14702 37314 14754 37326
rect 15038 37378 15090 37390
rect 15038 37314 15090 37326
rect 15598 37378 15650 37390
rect 15598 37314 15650 37326
rect 20078 37378 20130 37390
rect 20078 37314 20130 37326
rect 23774 37378 23826 37390
rect 23774 37314 23826 37326
rect 26798 37378 26850 37390
rect 26798 37314 26850 37326
rect 32174 37378 32226 37390
rect 37102 37378 37154 37390
rect 33842 37326 33854 37378
rect 33906 37326 33918 37378
rect 32174 37314 32226 37326
rect 37102 37314 37154 37326
rect 37214 37378 37266 37390
rect 37214 37314 37266 37326
rect 40238 37378 40290 37390
rect 40238 37314 40290 37326
rect 40350 37378 40402 37390
rect 45726 37378 45778 37390
rect 43250 37326 43262 37378
rect 43314 37326 43326 37378
rect 44818 37326 44830 37378
rect 44882 37326 44894 37378
rect 40350 37314 40402 37326
rect 45726 37314 45778 37326
rect 55694 37378 55746 37390
rect 55694 37314 55746 37326
rect 4174 37266 4226 37278
rect 15262 37266 15314 37278
rect 9650 37214 9662 37266
rect 9714 37214 9726 37266
rect 4174 37202 4226 37214
rect 15262 37202 15314 37214
rect 16494 37266 16546 37278
rect 16494 37202 16546 37214
rect 18062 37266 18114 37278
rect 18062 37202 18114 37214
rect 18286 37266 18338 37278
rect 20862 37266 20914 37278
rect 24110 37266 24162 37278
rect 19058 37214 19070 37266
rect 19122 37214 19134 37266
rect 23314 37214 23326 37266
rect 23378 37214 23390 37266
rect 18286 37202 18338 37214
rect 20862 37202 20914 37214
rect 24110 37202 24162 37214
rect 25566 37266 25618 37278
rect 31166 37266 31218 37278
rect 36206 37266 36258 37278
rect 27570 37214 27582 37266
rect 27634 37214 27646 37266
rect 31938 37214 31950 37266
rect 32002 37214 32014 37266
rect 33058 37214 33070 37266
rect 33122 37214 33134 37266
rect 25566 37202 25618 37214
rect 31166 37202 31218 37214
rect 36206 37202 36258 37214
rect 36542 37266 36594 37278
rect 38894 37266 38946 37278
rect 36866 37214 36878 37266
rect 36930 37214 36942 37266
rect 38434 37214 38446 37266
rect 38498 37214 38510 37266
rect 36542 37202 36594 37214
rect 38894 37202 38946 37214
rect 40014 37266 40066 37278
rect 44270 37266 44322 37278
rect 43138 37214 43150 37266
rect 43202 37214 43214 37266
rect 40014 37202 40066 37214
rect 44270 37202 44322 37214
rect 45166 37266 45218 37278
rect 45166 37202 45218 37214
rect 45390 37266 45442 37278
rect 54686 37266 54738 37278
rect 48178 37214 48190 37266
rect 48242 37214 48254 37266
rect 50082 37214 50094 37266
rect 50146 37214 50158 37266
rect 51202 37214 51214 37266
rect 51266 37214 51278 37266
rect 51762 37214 51774 37266
rect 51826 37214 51838 37266
rect 52210 37214 52222 37266
rect 52274 37214 52286 37266
rect 45390 37202 45442 37214
rect 54686 37202 54738 37214
rect 54910 37266 54962 37278
rect 54910 37202 54962 37214
rect 55358 37266 55410 37278
rect 55358 37202 55410 37214
rect 55806 37266 55858 37278
rect 55806 37202 55858 37214
rect 12910 37154 12962 37166
rect 10322 37102 10334 37154
rect 10386 37102 10398 37154
rect 12450 37102 12462 37154
rect 12514 37102 12526 37154
rect 12910 37090 12962 37102
rect 13358 37154 13410 37166
rect 13358 37090 13410 37102
rect 14478 37154 14530 37166
rect 14478 37090 14530 37102
rect 14814 37154 14866 37166
rect 14814 37090 14866 37102
rect 17614 37154 17666 37166
rect 17614 37090 17666 37102
rect 22094 37154 22146 37166
rect 25678 37154 25730 37166
rect 22866 37102 22878 37154
rect 22930 37102 22942 37154
rect 22094 37090 22146 37102
rect 25678 37090 25730 37102
rect 26462 37154 26514 37166
rect 39006 37154 39058 37166
rect 27122 37102 27134 37154
rect 27186 37102 27198 37154
rect 28242 37102 28254 37154
rect 28306 37102 28318 37154
rect 30370 37102 30382 37154
rect 30434 37102 30446 37154
rect 35970 37102 35982 37154
rect 36034 37102 36046 37154
rect 26462 37090 26514 37102
rect 39006 37090 39058 37102
rect 39454 37154 39506 37166
rect 39454 37090 39506 37102
rect 42814 37154 42866 37166
rect 42814 37090 42866 37102
rect 45614 37154 45666 37166
rect 45614 37090 45666 37102
rect 47070 37154 47122 37166
rect 55134 37154 55186 37166
rect 49970 37102 49982 37154
rect 50034 37102 50046 37154
rect 53442 37102 53454 37154
rect 53506 37102 53518 37154
rect 54226 37102 54238 37154
rect 54290 37102 54302 37154
rect 47070 37090 47122 37102
rect 55134 37090 55186 37102
rect 15934 37042 15986 37054
rect 15934 36978 15986 36990
rect 17838 37042 17890 37054
rect 17838 36978 17890 36990
rect 18734 37042 18786 37054
rect 18734 36978 18786 36990
rect 21982 37042 22034 37054
rect 39790 37042 39842 37054
rect 47854 37042 47906 37054
rect 30594 36990 30606 37042
rect 30658 37039 30670 37042
rect 30930 37039 30942 37042
rect 30658 36993 30942 37039
rect 30658 36990 30670 36993
rect 30930 36990 30942 36993
rect 30994 36990 31006 37042
rect 47058 36990 47070 37042
rect 47122 37039 47134 37042
rect 47506 37039 47518 37042
rect 47122 36993 47518 37039
rect 47122 36990 47134 36993
rect 47506 36990 47518 36993
rect 47570 36990 47582 37042
rect 21982 36978 22034 36990
rect 39790 36978 39842 36990
rect 47854 36978 47906 36990
rect 48190 37042 48242 37054
rect 48190 36978 48242 36990
rect 55694 37042 55746 37054
rect 55694 36978 55746 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 18958 36706 19010 36718
rect 18958 36642 19010 36654
rect 19854 36706 19906 36718
rect 19854 36642 19906 36654
rect 20750 36706 20802 36718
rect 20750 36642 20802 36654
rect 31502 36706 31554 36718
rect 31502 36642 31554 36654
rect 37550 36706 37602 36718
rect 37550 36642 37602 36654
rect 38894 36706 38946 36718
rect 38894 36642 38946 36654
rect 45502 36706 45554 36718
rect 53006 36706 53058 36718
rect 47730 36654 47742 36706
rect 47794 36654 47806 36706
rect 56354 36654 56366 36706
rect 56418 36654 56430 36706
rect 45502 36642 45554 36654
rect 53006 36642 53058 36654
rect 19070 36594 19122 36606
rect 19070 36530 19122 36542
rect 19630 36594 19682 36606
rect 27582 36594 27634 36606
rect 23650 36542 23662 36594
rect 23714 36542 23726 36594
rect 24098 36542 24110 36594
rect 24162 36542 24174 36594
rect 26226 36542 26238 36594
rect 26290 36542 26302 36594
rect 19630 36530 19682 36542
rect 27582 36530 27634 36542
rect 28590 36594 28642 36606
rect 37998 36594 38050 36606
rect 47630 36594 47682 36606
rect 33394 36542 33406 36594
rect 33458 36542 33470 36594
rect 40450 36542 40462 36594
rect 40514 36542 40526 36594
rect 42578 36542 42590 36594
rect 42642 36542 42654 36594
rect 28590 36530 28642 36542
rect 37998 36530 38050 36542
rect 47630 36530 47682 36542
rect 50878 36594 50930 36606
rect 54674 36542 54686 36594
rect 54738 36542 54750 36594
rect 50878 36530 50930 36542
rect 18622 36482 18674 36494
rect 20078 36482 20130 36494
rect 17490 36430 17502 36482
rect 17554 36430 17566 36482
rect 19282 36430 19294 36482
rect 19346 36430 19358 36482
rect 18622 36418 18674 36430
rect 20078 36418 20130 36430
rect 20302 36482 20354 36494
rect 22206 36482 22258 36494
rect 36990 36482 37042 36494
rect 21522 36430 21534 36482
rect 21586 36430 21598 36482
rect 23314 36430 23326 36482
rect 23378 36430 23390 36482
rect 27010 36430 27022 36482
rect 27074 36430 27086 36482
rect 30706 36430 30718 36482
rect 30770 36430 30782 36482
rect 32050 36430 32062 36482
rect 32114 36430 32126 36482
rect 33730 36430 33742 36482
rect 33794 36430 33806 36482
rect 36082 36430 36094 36482
rect 36146 36430 36158 36482
rect 20302 36418 20354 36430
rect 22206 36418 22258 36430
rect 36990 36418 37042 36430
rect 37214 36482 37266 36494
rect 37214 36418 37266 36430
rect 37886 36482 37938 36494
rect 37886 36418 37938 36430
rect 38110 36482 38162 36494
rect 38110 36418 38162 36430
rect 38558 36482 38610 36494
rect 46174 36482 46226 36494
rect 48078 36482 48130 36494
rect 39666 36430 39678 36482
rect 39730 36430 39742 36482
rect 45826 36430 45838 36482
rect 45890 36430 45902 36482
rect 47282 36430 47294 36482
rect 47346 36430 47358 36482
rect 38558 36418 38610 36430
rect 46174 36418 46226 36430
rect 48078 36418 48130 36430
rect 48526 36482 48578 36494
rect 50542 36482 50594 36494
rect 49634 36430 49646 36482
rect 49698 36430 49710 36482
rect 50306 36430 50318 36482
rect 50370 36430 50382 36482
rect 48526 36418 48578 36430
rect 50542 36418 50594 36430
rect 50654 36482 50706 36494
rect 53230 36482 53282 36494
rect 51314 36430 51326 36482
rect 51378 36430 51390 36482
rect 50654 36418 50706 36430
rect 53230 36418 53282 36430
rect 53454 36482 53506 36494
rect 57038 36482 57090 36494
rect 55010 36430 55022 36482
rect 55074 36430 55086 36482
rect 56354 36430 56366 36482
rect 56418 36430 56430 36482
rect 53454 36418 53506 36430
rect 57038 36418 57090 36430
rect 22654 36370 22706 36382
rect 14578 36318 14590 36370
rect 14642 36318 14654 36370
rect 16034 36318 16046 36370
rect 16098 36318 16110 36370
rect 21298 36318 21310 36370
rect 21362 36318 21374 36370
rect 22654 36306 22706 36318
rect 30158 36370 30210 36382
rect 30158 36306 30210 36318
rect 31166 36370 31218 36382
rect 39006 36370 39058 36382
rect 35858 36318 35870 36370
rect 35922 36318 35934 36370
rect 31166 36306 31218 36318
rect 39006 36306 39058 36318
rect 44830 36370 44882 36382
rect 49086 36370 49138 36382
rect 46498 36318 46510 36370
rect 46562 36318 46574 36370
rect 44830 36306 44882 36318
rect 49086 36306 49138 36318
rect 50990 36370 51042 36382
rect 55470 36370 55522 36382
rect 51650 36318 51662 36370
rect 51714 36318 51726 36370
rect 51986 36318 51998 36370
rect 52050 36318 52062 36370
rect 50990 36306 51042 36318
rect 55470 36306 55522 36318
rect 55806 36370 55858 36382
rect 56018 36318 56030 36370
rect 56082 36318 56094 36370
rect 55806 36306 55858 36318
rect 14926 36258 14978 36270
rect 22766 36258 22818 36270
rect 18274 36206 18286 36258
rect 18338 36206 18350 36258
rect 14926 36194 14978 36206
rect 22766 36194 22818 36206
rect 22878 36258 22930 36270
rect 31390 36258 31442 36270
rect 30482 36206 30494 36258
rect 30546 36206 30558 36258
rect 22878 36194 22930 36206
rect 31390 36194 31442 36206
rect 31838 36258 31890 36270
rect 31838 36194 31890 36206
rect 38894 36258 38946 36270
rect 38894 36194 38946 36206
rect 43038 36258 43090 36270
rect 43038 36194 43090 36206
rect 44270 36258 44322 36270
rect 45614 36258 45666 36270
rect 45154 36206 45166 36258
rect 45218 36206 45230 36258
rect 44270 36194 44322 36206
rect 45614 36194 45666 36206
rect 48638 36258 48690 36270
rect 48638 36194 48690 36206
rect 48750 36258 48802 36270
rect 48750 36194 48802 36206
rect 49198 36258 49250 36270
rect 49198 36194 49250 36206
rect 49310 36258 49362 36270
rect 49310 36194 49362 36206
rect 52558 36258 52610 36270
rect 52558 36194 52610 36206
rect 53902 36258 53954 36270
rect 57486 36258 57538 36270
rect 56242 36206 56254 36258
rect 56306 36206 56318 36258
rect 53902 36194 53954 36206
rect 57486 36194 57538 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 16830 35922 16882 35934
rect 18286 35922 18338 35934
rect 17378 35870 17390 35922
rect 17442 35870 17454 35922
rect 16830 35858 16882 35870
rect 18286 35858 18338 35870
rect 21422 35922 21474 35934
rect 21422 35858 21474 35870
rect 21870 35922 21922 35934
rect 21870 35858 21922 35870
rect 24782 35922 24834 35934
rect 30494 35922 30546 35934
rect 25442 35870 25454 35922
rect 25506 35870 25518 35922
rect 24782 35858 24834 35870
rect 30494 35858 30546 35870
rect 31166 35922 31218 35934
rect 31166 35858 31218 35870
rect 31614 35922 31666 35934
rect 31614 35858 31666 35870
rect 40126 35922 40178 35934
rect 40126 35858 40178 35870
rect 45166 35922 45218 35934
rect 45166 35858 45218 35870
rect 48078 35922 48130 35934
rect 48078 35858 48130 35870
rect 57374 35922 57426 35934
rect 57374 35858 57426 35870
rect 20526 35810 20578 35822
rect 25790 35810 25842 35822
rect 26462 35810 26514 35822
rect 16146 35758 16158 35810
rect 16210 35758 16222 35810
rect 22866 35758 22878 35810
rect 22930 35758 22942 35810
rect 26114 35758 26126 35810
rect 26178 35758 26190 35810
rect 20526 35746 20578 35758
rect 25790 35746 25842 35758
rect 26462 35746 26514 35758
rect 34414 35810 34466 35822
rect 34414 35746 34466 35758
rect 37550 35810 37602 35822
rect 37550 35746 37602 35758
rect 44718 35810 44770 35822
rect 44718 35746 44770 35758
rect 47854 35810 47906 35822
rect 47854 35746 47906 35758
rect 48190 35810 48242 35822
rect 56590 35810 56642 35822
rect 54002 35758 54014 35810
rect 54066 35758 54078 35810
rect 48190 35746 48242 35758
rect 56590 35746 56642 35758
rect 15486 35698 15538 35710
rect 12002 35646 12014 35698
rect 12066 35646 12078 35698
rect 15486 35634 15538 35646
rect 15710 35698 15762 35710
rect 15710 35634 15762 35646
rect 15934 35698 15986 35710
rect 15934 35634 15986 35646
rect 16494 35698 16546 35710
rect 16494 35634 16546 35646
rect 17726 35698 17778 35710
rect 17726 35634 17778 35646
rect 17950 35698 18002 35710
rect 17950 35634 18002 35646
rect 18622 35698 18674 35710
rect 18622 35634 18674 35646
rect 20078 35698 20130 35710
rect 20078 35634 20130 35646
rect 22430 35698 22482 35710
rect 27246 35698 27298 35710
rect 30270 35698 30322 35710
rect 23426 35646 23438 35698
rect 23490 35646 23502 35698
rect 23874 35646 23886 35698
rect 23938 35646 23950 35698
rect 29922 35646 29934 35698
rect 29986 35646 29998 35698
rect 22430 35634 22482 35646
rect 27246 35634 27298 35646
rect 30270 35634 30322 35646
rect 31390 35698 31442 35710
rect 31390 35634 31442 35646
rect 34638 35698 34690 35710
rect 39006 35698 39058 35710
rect 36978 35646 36990 35698
rect 37042 35646 37054 35698
rect 38546 35646 38558 35698
rect 38610 35646 38622 35698
rect 34638 35634 34690 35646
rect 39006 35634 39058 35646
rect 39342 35698 39394 35710
rect 44942 35698 44994 35710
rect 47742 35698 47794 35710
rect 39666 35646 39678 35698
rect 39730 35646 39742 35698
rect 46722 35646 46734 35698
rect 46786 35646 46798 35698
rect 47058 35646 47070 35698
rect 47122 35646 47134 35698
rect 48738 35646 48750 35698
rect 48802 35646 48814 35698
rect 49522 35646 49534 35698
rect 49586 35646 49598 35698
rect 50642 35646 50654 35698
rect 50706 35646 50718 35698
rect 52098 35646 52110 35698
rect 52162 35646 52174 35698
rect 53218 35646 53230 35698
rect 53282 35646 53294 35698
rect 54338 35646 54350 35698
rect 54402 35646 54414 35698
rect 55122 35646 55134 35698
rect 55186 35646 55198 35698
rect 56914 35646 56926 35698
rect 56978 35646 56990 35698
rect 39342 35634 39394 35646
rect 44942 35634 44994 35646
rect 47742 35634 47794 35646
rect 15598 35586 15650 35598
rect 12674 35534 12686 35586
rect 12738 35534 12750 35586
rect 14802 35534 14814 35586
rect 14866 35534 14878 35586
rect 15598 35522 15650 35534
rect 19742 35586 19794 35598
rect 30382 35586 30434 35598
rect 23538 35534 23550 35586
rect 23602 35534 23614 35586
rect 19742 35522 19794 35534
rect 30382 35522 30434 35534
rect 31502 35586 31554 35598
rect 43150 35586 43202 35598
rect 36754 35534 36766 35586
rect 36818 35534 36830 35586
rect 38098 35534 38110 35586
rect 38162 35534 38174 35586
rect 31502 35522 31554 35534
rect 43150 35522 43202 35534
rect 44270 35586 44322 35598
rect 44270 35522 44322 35534
rect 45054 35586 45106 35598
rect 55806 35586 55858 35598
rect 45602 35534 45614 35586
rect 45666 35534 45678 35586
rect 51426 35534 51438 35586
rect 51490 35534 51502 35586
rect 45054 35522 45106 35534
rect 55806 35522 55858 35534
rect 56702 35586 56754 35598
rect 56702 35522 56754 35534
rect 57822 35586 57874 35598
rect 57822 35522 57874 35534
rect 34862 35474 34914 35486
rect 34862 35410 34914 35422
rect 35086 35474 35138 35486
rect 35086 35410 35138 35422
rect 35534 35474 35586 35486
rect 35534 35410 35586 35422
rect 39678 35474 39730 35486
rect 57362 35422 57374 35474
rect 57426 35471 57438 35474
rect 58034 35471 58046 35474
rect 57426 35425 58046 35471
rect 57426 35422 57438 35425
rect 58034 35422 58046 35425
rect 58098 35422 58110 35474
rect 39678 35410 39730 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 13470 35138 13522 35150
rect 13470 35074 13522 35086
rect 13806 35138 13858 35150
rect 13806 35074 13858 35086
rect 15038 35138 15090 35150
rect 15038 35074 15090 35086
rect 30382 35138 30434 35150
rect 30382 35074 30434 35086
rect 31390 35138 31442 35150
rect 31390 35074 31442 35086
rect 44046 35138 44098 35150
rect 44046 35074 44098 35086
rect 44158 35138 44210 35150
rect 44158 35074 44210 35086
rect 46174 35138 46226 35150
rect 54574 35138 54626 35150
rect 53106 35086 53118 35138
rect 53170 35086 53182 35138
rect 46174 35074 46226 35086
rect 54574 35074 54626 35086
rect 14590 35026 14642 35038
rect 14590 34962 14642 34974
rect 14814 35026 14866 35038
rect 19070 35026 19122 35038
rect 18610 34974 18622 35026
rect 18674 34974 18686 35026
rect 14814 34962 14866 34974
rect 19070 34962 19122 34974
rect 21534 35026 21586 35038
rect 25902 35026 25954 35038
rect 22418 34974 22430 35026
rect 22482 34974 22494 35026
rect 21534 34962 21586 34974
rect 25902 34962 25954 34974
rect 26238 35026 26290 35038
rect 29710 35026 29762 35038
rect 45278 35026 45330 35038
rect 49758 35026 49810 35038
rect 27122 34974 27134 35026
rect 27186 34974 27198 35026
rect 30034 34974 30046 35026
rect 30098 34974 30110 35026
rect 37538 34974 37550 35026
rect 37602 34974 37614 35026
rect 40002 34974 40014 35026
rect 40066 34974 40078 35026
rect 42130 34974 42142 35026
rect 42194 34974 42206 35026
rect 49410 34974 49422 35026
rect 49474 34974 49486 35026
rect 26238 34962 26290 34974
rect 29710 34962 29762 34974
rect 45278 34962 45330 34974
rect 49758 34962 49810 34974
rect 52894 35026 52946 35038
rect 52894 34962 52946 34974
rect 54462 35026 54514 35038
rect 55234 34974 55246 35026
rect 55298 34974 55310 35026
rect 57362 34974 57374 35026
rect 57426 34974 57438 35026
rect 54462 34962 54514 34974
rect 19518 34914 19570 34926
rect 15810 34862 15822 34914
rect 15874 34862 15886 34914
rect 19518 34850 19570 34862
rect 19966 34914 20018 34926
rect 19966 34850 20018 34862
rect 20750 34914 20802 34926
rect 27582 34914 27634 34926
rect 21970 34862 21982 34914
rect 22034 34862 22046 34914
rect 22642 34862 22654 34914
rect 22706 34862 22718 34914
rect 26786 34862 26798 34914
rect 26850 34862 26862 34914
rect 20750 34850 20802 34862
rect 27582 34850 27634 34862
rect 28142 34914 28194 34926
rect 33518 34914 33570 34926
rect 31042 34862 31054 34914
rect 31106 34862 31118 34914
rect 28142 34850 28194 34862
rect 33518 34850 33570 34862
rect 34078 34914 34130 34926
rect 34078 34850 34130 34862
rect 34414 34914 34466 34926
rect 34414 34850 34466 34862
rect 34862 34914 34914 34926
rect 34862 34850 34914 34862
rect 34974 34914 35026 34926
rect 43822 34914 43874 34926
rect 45502 34914 45554 34926
rect 35298 34862 35310 34914
rect 35362 34862 35374 34914
rect 37202 34862 37214 34914
rect 37266 34862 37278 34914
rect 39330 34862 39342 34914
rect 39394 34862 39406 34914
rect 45042 34862 45054 34914
rect 45106 34862 45118 34914
rect 34974 34850 35026 34862
rect 43822 34850 43874 34862
rect 45502 34850 45554 34862
rect 45726 34914 45778 34926
rect 45726 34850 45778 34862
rect 46062 34914 46114 34926
rect 54798 34914 54850 34926
rect 47842 34862 47854 34914
rect 47906 34862 47918 34914
rect 48402 34862 48414 34914
rect 48466 34862 48478 34914
rect 50194 34862 50206 34914
rect 50258 34862 50270 34914
rect 50642 34862 50654 34914
rect 50706 34862 50718 34914
rect 52098 34862 52110 34914
rect 52162 34862 52174 34914
rect 53330 34862 53342 34914
rect 53394 34862 53406 34914
rect 53778 34862 53790 34914
rect 53842 34862 53854 34914
rect 58034 34862 58046 34914
rect 58098 34862 58110 34914
rect 46062 34850 46114 34862
rect 54798 34850 54850 34862
rect 20190 34802 20242 34814
rect 16482 34750 16494 34802
rect 16546 34750 16558 34802
rect 20190 34738 20242 34750
rect 33854 34802 33906 34814
rect 33854 34738 33906 34750
rect 43710 34802 43762 34814
rect 43710 34738 43762 34750
rect 44830 34802 44882 34814
rect 44830 34738 44882 34750
rect 46622 34802 46674 34814
rect 51090 34750 51102 34802
rect 51154 34750 51166 34802
rect 46622 34738 46674 34750
rect 13582 34690 13634 34702
rect 18958 34690 19010 34702
rect 15362 34638 15374 34690
rect 15426 34638 15438 34690
rect 13582 34626 13634 34638
rect 18958 34626 19010 34638
rect 19854 34690 19906 34702
rect 23550 34690 23602 34702
rect 23202 34638 23214 34690
rect 23266 34638 23278 34690
rect 19854 34626 19906 34638
rect 23550 34626 23602 34638
rect 23998 34690 24050 34702
rect 23998 34626 24050 34638
rect 26350 34690 26402 34702
rect 26350 34626 26402 34638
rect 28590 34690 28642 34702
rect 28590 34626 28642 34638
rect 29150 34690 29202 34702
rect 29150 34626 29202 34638
rect 30158 34690 30210 34702
rect 30158 34626 30210 34638
rect 31278 34690 31330 34702
rect 31278 34626 31330 34638
rect 33966 34690 34018 34702
rect 33966 34626 34018 34638
rect 34750 34690 34802 34702
rect 34750 34626 34802 34638
rect 38446 34690 38498 34702
rect 42926 34690 42978 34702
rect 42578 34638 42590 34690
rect 42642 34638 42654 34690
rect 38446 34626 38498 34638
rect 42926 34626 42978 34638
rect 43374 34690 43426 34702
rect 43374 34626 43426 34638
rect 45614 34690 45666 34702
rect 54462 34690 54514 34702
rect 50978 34638 50990 34690
rect 51042 34638 51054 34690
rect 51986 34638 51998 34690
rect 52050 34638 52062 34690
rect 45614 34626 45666 34638
rect 54462 34626 54514 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 15598 34354 15650 34366
rect 15598 34290 15650 34302
rect 15934 34354 15986 34366
rect 15934 34290 15986 34302
rect 17502 34354 17554 34366
rect 17502 34290 17554 34302
rect 22654 34354 22706 34366
rect 22654 34290 22706 34302
rect 25454 34354 25506 34366
rect 25454 34290 25506 34302
rect 27582 34354 27634 34366
rect 27582 34290 27634 34302
rect 36654 34354 36706 34366
rect 36654 34290 36706 34302
rect 46958 34354 47010 34366
rect 46958 34290 47010 34302
rect 47966 34354 48018 34366
rect 47966 34290 48018 34302
rect 54014 34354 54066 34366
rect 54014 34290 54066 34302
rect 56030 34354 56082 34366
rect 56030 34290 56082 34302
rect 57374 34354 57426 34366
rect 57374 34290 57426 34302
rect 58046 34354 58098 34366
rect 58046 34290 58098 34302
rect 14030 34242 14082 34254
rect 14030 34178 14082 34190
rect 14702 34242 14754 34254
rect 14702 34178 14754 34190
rect 17390 34242 17442 34254
rect 17390 34178 17442 34190
rect 17726 34242 17778 34254
rect 17726 34178 17778 34190
rect 18846 34242 18898 34254
rect 23214 34242 23266 34254
rect 47854 34242 47906 34254
rect 21410 34190 21422 34242
rect 21474 34190 21486 34242
rect 29362 34190 29374 34242
rect 29426 34190 29438 34242
rect 33842 34190 33854 34242
rect 33906 34190 33918 34242
rect 43362 34190 43374 34242
rect 43426 34190 43438 34242
rect 18846 34178 18898 34190
rect 23214 34178 23266 34190
rect 47854 34178 47906 34190
rect 48078 34242 48130 34254
rect 48078 34178 48130 34190
rect 54238 34242 54290 34254
rect 54238 34178 54290 34190
rect 54798 34242 54850 34254
rect 55918 34242 55970 34254
rect 57262 34242 57314 34254
rect 55010 34190 55022 34242
rect 55074 34190 55086 34242
rect 56578 34190 56590 34242
rect 56642 34190 56654 34242
rect 54798 34178 54850 34190
rect 55918 34178 55970 34190
rect 57262 34178 57314 34190
rect 57486 34242 57538 34254
rect 57486 34178 57538 34190
rect 16382 34130 16434 34142
rect 16382 34066 16434 34078
rect 17950 34130 18002 34142
rect 36766 34130 36818 34142
rect 46734 34130 46786 34142
rect 55246 34130 55298 34142
rect 22082 34078 22094 34130
rect 22146 34078 22158 34130
rect 23538 34078 23550 34130
rect 23602 34078 23614 34130
rect 24434 34078 24446 34130
rect 24498 34078 24510 34130
rect 28690 34078 28702 34130
rect 28754 34078 28766 34130
rect 33058 34078 33070 34130
rect 33122 34078 33134 34130
rect 37090 34078 37102 34130
rect 37154 34078 37166 34130
rect 38210 34078 38222 34130
rect 38274 34078 38286 34130
rect 39330 34078 39342 34130
rect 39394 34078 39406 34130
rect 42690 34078 42702 34130
rect 42754 34078 42766 34130
rect 47170 34078 47182 34130
rect 47234 34078 47246 34130
rect 47506 34078 47518 34130
rect 47570 34078 47582 34130
rect 50306 34078 50318 34130
rect 50370 34078 50382 34130
rect 50978 34078 50990 34130
rect 51042 34078 51054 34130
rect 53218 34078 53230 34130
rect 53282 34078 53294 34130
rect 53442 34078 53454 34130
rect 53506 34078 53518 34130
rect 55458 34078 55470 34130
rect 55522 34078 55534 34130
rect 56802 34078 56814 34130
rect 56866 34078 56878 34130
rect 17950 34066 18002 34078
rect 36766 34066 36818 34078
rect 46734 34066 46786 34078
rect 55246 34066 55298 34078
rect 14142 34018 14194 34030
rect 14142 33954 14194 33966
rect 16942 34018 16994 34030
rect 32062 34018 32114 34030
rect 45950 34018 46002 34030
rect 54910 34018 54962 34030
rect 18498 33966 18510 34018
rect 18562 33966 18574 34018
rect 19282 33966 19294 34018
rect 19346 33966 19358 34018
rect 23426 33966 23438 34018
rect 23490 33966 23502 34018
rect 31490 33966 31502 34018
rect 31554 33966 31566 34018
rect 35970 33966 35982 34018
rect 36034 33966 36046 34018
rect 45490 33966 45502 34018
rect 45554 33966 45566 34018
rect 47058 33966 47070 34018
rect 47122 33966 47134 34018
rect 49858 33966 49870 34018
rect 49922 33966 49934 34018
rect 53890 33966 53902 34018
rect 53954 33966 53966 34018
rect 16942 33954 16994 33966
rect 32062 33954 32114 33966
rect 45950 33954 46002 33966
rect 54910 33954 54962 33966
rect 14254 33906 14306 33918
rect 14254 33842 14306 33854
rect 24110 33906 24162 33918
rect 24110 33842 24162 33854
rect 24446 33906 24498 33918
rect 24446 33842 24498 33854
rect 36654 33906 36706 33918
rect 38546 33854 38558 33906
rect 38610 33854 38622 33906
rect 50194 33854 50206 33906
rect 50258 33854 50270 33906
rect 36654 33842 36706 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 17278 33570 17330 33582
rect 17278 33506 17330 33518
rect 43822 33570 43874 33582
rect 43822 33506 43874 33518
rect 48974 33570 49026 33582
rect 48974 33506 49026 33518
rect 49310 33570 49362 33582
rect 49310 33506 49362 33518
rect 50206 33570 50258 33582
rect 50206 33506 50258 33518
rect 54798 33570 54850 33582
rect 54798 33506 54850 33518
rect 20750 33458 20802 33470
rect 49982 33458 50034 33470
rect 14242 33406 14254 33458
rect 14306 33406 14318 33458
rect 16370 33406 16382 33458
rect 16434 33406 16446 33458
rect 16930 33406 16942 33458
rect 16994 33406 17006 33458
rect 24546 33406 24558 33458
rect 24610 33406 24622 33458
rect 26674 33406 26686 33458
rect 26738 33406 26750 33458
rect 31714 33406 31726 33458
rect 31778 33406 31790 33458
rect 33842 33406 33854 33458
rect 33906 33406 33918 33458
rect 40338 33406 40350 33458
rect 40402 33406 40414 33458
rect 43586 33406 43598 33458
rect 43650 33406 43662 33458
rect 55234 33406 55246 33458
rect 55298 33406 55310 33458
rect 57362 33406 57374 33458
rect 57426 33406 57438 33458
rect 20750 33394 20802 33406
rect 49982 33394 50034 33406
rect 18398 33346 18450 33358
rect 13570 33294 13582 33346
rect 13634 33294 13646 33346
rect 18398 33282 18450 33294
rect 18958 33346 19010 33358
rect 18958 33282 19010 33294
rect 19630 33346 19682 33358
rect 19630 33282 19682 33294
rect 21310 33346 21362 33358
rect 21310 33282 21362 33294
rect 21646 33346 21698 33358
rect 21646 33282 21698 33294
rect 21982 33346 22034 33358
rect 21982 33282 22034 33294
rect 22766 33346 22818 33358
rect 27470 33346 27522 33358
rect 46846 33346 46898 33358
rect 23762 33294 23774 33346
rect 23826 33294 23838 33346
rect 27570 33294 27582 33346
rect 27634 33294 27646 33346
rect 31042 33294 31054 33346
rect 31106 33294 31118 33346
rect 35522 33294 35534 33346
rect 35586 33294 35598 33346
rect 37426 33294 37438 33346
rect 37490 33294 37502 33346
rect 40898 33294 40910 33346
rect 40962 33294 40974 33346
rect 42018 33294 42030 33346
rect 42082 33294 42094 33346
rect 43474 33294 43486 33346
rect 43538 33294 43550 33346
rect 22766 33282 22818 33294
rect 27470 33282 27522 33294
rect 46846 33282 46898 33294
rect 50318 33346 50370 33358
rect 53330 33294 53342 33346
rect 53394 33294 53406 33346
rect 54338 33294 54350 33346
rect 54402 33294 54414 33346
rect 58146 33294 58158 33346
rect 58210 33294 58222 33346
rect 50318 33282 50370 33294
rect 17054 33234 17106 33246
rect 17054 33170 17106 33182
rect 27022 33234 27074 33246
rect 45838 33234 45890 33246
rect 27234 33182 27246 33234
rect 27298 33182 27310 33234
rect 35074 33182 35086 33234
rect 35138 33182 35150 33234
rect 35634 33182 35646 33234
rect 35698 33182 35710 33234
rect 38210 33182 38222 33234
rect 38274 33182 38286 33234
rect 41010 33182 41022 33234
rect 41074 33182 41086 33234
rect 42578 33182 42590 33234
rect 42642 33182 42654 33234
rect 27022 33170 27074 33182
rect 45838 33170 45890 33182
rect 46062 33234 46114 33246
rect 46062 33170 46114 33182
rect 46510 33234 46562 33246
rect 46510 33170 46562 33182
rect 49086 33234 49138 33246
rect 54686 33234 54738 33246
rect 52770 33182 52782 33234
rect 52834 33182 52846 33234
rect 54226 33182 54238 33234
rect 54290 33182 54302 33234
rect 49086 33170 49138 33182
rect 54686 33170 54738 33182
rect 17726 33122 17778 33134
rect 17726 33058 17778 33070
rect 17838 33122 17890 33134
rect 17838 33058 17890 33070
rect 17950 33122 18002 33134
rect 17950 33058 18002 33070
rect 20190 33122 20242 33134
rect 20190 33058 20242 33070
rect 21758 33122 21810 33134
rect 23438 33122 23490 33134
rect 23090 33070 23102 33122
rect 23154 33070 23166 33122
rect 21758 33058 21810 33070
rect 23438 33058 23490 33070
rect 27806 33122 27858 33134
rect 27806 33058 27858 33070
rect 34302 33122 34354 33134
rect 34302 33058 34354 33070
rect 36206 33122 36258 33134
rect 36206 33058 36258 33070
rect 37102 33122 37154 33134
rect 43262 33122 43314 33134
rect 41906 33070 41918 33122
rect 41970 33070 41982 33122
rect 37102 33058 37154 33070
rect 43262 33058 43314 33070
rect 45950 33122 46002 33134
rect 45950 33058 46002 33070
rect 46622 33122 46674 33134
rect 46622 33058 46674 33070
rect 51102 33122 51154 33134
rect 51102 33058 51154 33070
rect 52110 33122 52162 33134
rect 53218 33070 53230 33122
rect 53282 33070 53294 33122
rect 52110 33058 52162 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 15598 32786 15650 32798
rect 15598 32722 15650 32734
rect 18510 32786 18562 32798
rect 18510 32722 18562 32734
rect 19294 32786 19346 32798
rect 19294 32722 19346 32734
rect 30046 32786 30098 32798
rect 30046 32722 30098 32734
rect 32174 32786 32226 32798
rect 34190 32786 34242 32798
rect 36990 32786 37042 32798
rect 32498 32734 32510 32786
rect 32562 32734 32574 32786
rect 35074 32734 35086 32786
rect 35138 32734 35150 32786
rect 32174 32722 32226 32734
rect 34190 32722 34242 32734
rect 36990 32722 37042 32734
rect 37662 32786 37714 32798
rect 37662 32722 37714 32734
rect 38110 32786 38162 32798
rect 38110 32722 38162 32734
rect 38558 32786 38610 32798
rect 38558 32722 38610 32734
rect 41246 32786 41298 32798
rect 41246 32722 41298 32734
rect 45054 32786 45106 32798
rect 45054 32722 45106 32734
rect 45390 32786 45442 32798
rect 45390 32722 45442 32734
rect 45726 32786 45778 32798
rect 49870 32786 49922 32798
rect 56702 32786 56754 32798
rect 49074 32734 49086 32786
rect 49138 32734 49150 32786
rect 52210 32734 52222 32786
rect 52274 32734 52286 32786
rect 45726 32722 45778 32734
rect 49870 32722 49922 32734
rect 56702 32722 56754 32734
rect 18846 32674 18898 32686
rect 25566 32674 25618 32686
rect 19618 32622 19630 32674
rect 19682 32622 19694 32674
rect 18846 32610 18898 32622
rect 25566 32610 25618 32622
rect 26014 32674 26066 32686
rect 37438 32674 37490 32686
rect 28802 32622 28814 32674
rect 28866 32622 28878 32674
rect 30818 32622 30830 32674
rect 30882 32622 30894 32674
rect 26014 32610 26066 32622
rect 37438 32610 37490 32622
rect 43262 32674 43314 32686
rect 43262 32610 43314 32622
rect 43486 32674 43538 32686
rect 43486 32610 43538 32622
rect 45278 32674 45330 32686
rect 45278 32610 45330 32622
rect 47406 32674 47458 32686
rect 47406 32610 47458 32622
rect 49534 32674 49586 32686
rect 49534 32610 49586 32622
rect 50318 32674 50370 32686
rect 50318 32610 50370 32622
rect 53342 32674 53394 32686
rect 53342 32610 53394 32622
rect 54798 32674 54850 32686
rect 54798 32610 54850 32622
rect 16270 32562 16322 32574
rect 12338 32510 12350 32562
rect 12402 32510 12414 32562
rect 16270 32498 16322 32510
rect 16382 32562 16434 32574
rect 16382 32498 16434 32510
rect 16606 32562 16658 32574
rect 17502 32562 17554 32574
rect 16818 32510 16830 32562
rect 16882 32510 16894 32562
rect 16606 32498 16658 32510
rect 17502 32498 17554 32510
rect 17614 32562 17666 32574
rect 17614 32498 17666 32510
rect 17726 32562 17778 32574
rect 17726 32498 17778 32510
rect 17838 32562 17890 32574
rect 18398 32562 18450 32574
rect 18050 32510 18062 32562
rect 18114 32510 18126 32562
rect 17838 32498 17890 32510
rect 18398 32498 18450 32510
rect 18622 32562 18674 32574
rect 23550 32562 23602 32574
rect 20066 32510 20078 32562
rect 20130 32510 20142 32562
rect 23314 32510 23326 32562
rect 23378 32510 23390 32562
rect 18622 32498 18674 32510
rect 23550 32498 23602 32510
rect 23774 32562 23826 32574
rect 24334 32562 24386 32574
rect 23986 32510 23998 32562
rect 24050 32510 24062 32562
rect 23774 32498 23826 32510
rect 24334 32498 24386 32510
rect 26126 32562 26178 32574
rect 37326 32562 37378 32574
rect 26338 32510 26350 32562
rect 26402 32510 26414 32562
rect 29586 32510 29598 32562
rect 29650 32510 29662 32562
rect 30594 32510 30606 32562
rect 30658 32510 30670 32562
rect 33506 32510 33518 32562
rect 33570 32510 33582 32562
rect 35298 32510 35310 32562
rect 35362 32510 35374 32562
rect 26126 32498 26178 32510
rect 37326 32498 37378 32510
rect 37886 32562 37938 32574
rect 37886 32498 37938 32510
rect 38334 32562 38386 32574
rect 43038 32562 43090 32574
rect 47630 32562 47682 32574
rect 49758 32562 49810 32574
rect 41570 32510 41582 32562
rect 41634 32510 41646 32562
rect 44818 32510 44830 32562
rect 44882 32510 44894 32562
rect 45602 32510 45614 32562
rect 45666 32510 45678 32562
rect 47058 32510 47070 32562
rect 47122 32510 47134 32562
rect 48850 32510 48862 32562
rect 48914 32510 48926 32562
rect 38334 32498 38386 32510
rect 43038 32498 43090 32510
rect 47630 32498 47682 32510
rect 49758 32498 49810 32510
rect 49982 32562 50034 32574
rect 49982 32498 50034 32510
rect 50542 32562 50594 32574
rect 50542 32498 50594 32510
rect 50878 32562 50930 32574
rect 50878 32498 50930 32510
rect 51662 32562 51714 32574
rect 51662 32498 51714 32510
rect 51774 32562 51826 32574
rect 52098 32510 52110 32562
rect 52162 32510 52174 32562
rect 55906 32510 55918 32562
rect 55970 32510 55982 32562
rect 51774 32498 51826 32510
rect 16494 32450 16546 32462
rect 23662 32450 23714 32462
rect 13010 32398 13022 32450
rect 13074 32398 13086 32450
rect 15138 32398 15150 32450
rect 15202 32398 15214 32450
rect 20738 32398 20750 32450
rect 20802 32398 20814 32450
rect 22866 32398 22878 32450
rect 22930 32398 22942 32450
rect 16494 32386 16546 32398
rect 23662 32386 23714 32398
rect 24446 32450 24498 32462
rect 24446 32386 24498 32398
rect 25678 32450 25730 32462
rect 34750 32450 34802 32462
rect 26674 32398 26686 32450
rect 26738 32398 26750 32450
rect 33170 32398 33182 32450
rect 33234 32398 33246 32450
rect 25678 32386 25730 32398
rect 34750 32386 34802 32398
rect 38222 32450 38274 32462
rect 38222 32386 38274 32398
rect 41806 32450 41858 32462
rect 41806 32386 41858 32398
rect 41918 32450 41970 32462
rect 41918 32386 41970 32398
rect 42702 32450 42754 32462
rect 42702 32386 42754 32398
rect 43150 32450 43202 32462
rect 43150 32386 43202 32398
rect 47518 32450 47570 32462
rect 47518 32386 47570 32398
rect 48190 32450 48242 32462
rect 48190 32386 48242 32398
rect 50766 32450 50818 32462
rect 50766 32386 50818 32398
rect 51438 32450 51490 32462
rect 51438 32386 51490 32398
rect 57150 32450 57202 32462
rect 57150 32386 57202 32398
rect 45838 32338 45890 32350
rect 45838 32274 45890 32286
rect 46062 32338 46114 32350
rect 46062 32274 46114 32286
rect 46286 32338 46338 32350
rect 46286 32274 46338 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 27470 32002 27522 32014
rect 18722 31950 18734 32002
rect 18786 31950 18798 32002
rect 23538 31950 23550 32002
rect 23602 31950 23614 32002
rect 27470 31938 27522 31950
rect 37550 32002 37602 32014
rect 37550 31938 37602 31950
rect 48974 32002 49026 32014
rect 51538 31950 51550 32002
rect 51602 31950 51614 32002
rect 48974 31938 49026 31950
rect 15598 31890 15650 31902
rect 28366 31890 28418 31902
rect 13682 31838 13694 31890
rect 13746 31838 13758 31890
rect 21858 31838 21870 31890
rect 21922 31838 21934 31890
rect 24546 31838 24558 31890
rect 24610 31838 24622 31890
rect 15598 31826 15650 31838
rect 28366 31826 28418 31838
rect 33518 31890 33570 31902
rect 33518 31826 33570 31838
rect 38782 31890 38834 31902
rect 53230 31890 53282 31902
rect 40674 31838 40686 31890
rect 40738 31838 40750 31890
rect 41906 31838 41918 31890
rect 41970 31838 41982 31890
rect 44034 31838 44046 31890
rect 44098 31838 44110 31890
rect 46946 31838 46958 31890
rect 47010 31838 47022 31890
rect 53890 31838 53902 31890
rect 53954 31838 53966 31890
rect 38782 31826 38834 31838
rect 53230 31826 53282 31838
rect 16158 31778 16210 31790
rect 22206 31778 22258 31790
rect 23662 31778 23714 31790
rect 13794 31726 13806 31778
rect 13858 31726 13870 31778
rect 16594 31726 16606 31778
rect 16658 31726 16670 31778
rect 17378 31726 17390 31778
rect 17442 31726 17454 31778
rect 18834 31726 18846 31778
rect 18898 31726 18910 31778
rect 19506 31726 19518 31778
rect 19570 31726 19582 31778
rect 23090 31726 23102 31778
rect 23154 31726 23166 31778
rect 16158 31714 16210 31726
rect 22206 31714 22258 31726
rect 23662 31714 23714 31726
rect 27022 31778 27074 31790
rect 30270 31778 30322 31790
rect 27234 31726 27246 31778
rect 27298 31726 27310 31778
rect 27794 31726 27806 31778
rect 27858 31726 27870 31778
rect 27022 31714 27074 31726
rect 30270 31714 30322 31726
rect 31502 31778 31554 31790
rect 31502 31714 31554 31726
rect 32062 31778 32114 31790
rect 32062 31714 32114 31726
rect 34190 31778 34242 31790
rect 34190 31714 34242 31726
rect 34302 31778 34354 31790
rect 34302 31714 34354 31726
rect 34526 31778 34578 31790
rect 34526 31714 34578 31726
rect 37438 31778 37490 31790
rect 49422 31778 49474 31790
rect 37650 31726 37662 31778
rect 37714 31726 37726 31778
rect 41234 31726 41246 31778
rect 41298 31726 41310 31778
rect 46274 31726 46286 31778
rect 46338 31726 46350 31778
rect 48066 31726 48078 31778
rect 48130 31726 48142 31778
rect 37438 31714 37490 31726
rect 49422 31714 49474 31726
rect 49646 31778 49698 31790
rect 49646 31714 49698 31726
rect 50654 31778 50706 31790
rect 50654 31714 50706 31726
rect 50878 31778 50930 31790
rect 52110 31778 52162 31790
rect 51538 31726 51550 31778
rect 51602 31726 51614 31778
rect 51874 31726 51886 31778
rect 51938 31726 51950 31778
rect 50878 31714 50930 31726
rect 52110 31714 52162 31726
rect 52670 31778 52722 31790
rect 56690 31726 56702 31778
rect 56754 31726 56766 31778
rect 52670 31714 52722 31726
rect 13470 31666 13522 31678
rect 13470 31602 13522 31614
rect 15710 31666 15762 31678
rect 15710 31602 15762 31614
rect 17054 31666 17106 31678
rect 21870 31666 21922 31678
rect 20066 31614 20078 31666
rect 20130 31614 20142 31666
rect 17054 31602 17106 31614
rect 21870 31602 21922 31614
rect 22430 31666 22482 31678
rect 26350 31666 26402 31678
rect 33854 31666 33906 31678
rect 24882 31614 24894 31666
rect 24946 31614 24958 31666
rect 29922 31614 29934 31666
rect 29986 31614 29998 31666
rect 22430 31602 22482 31614
rect 26350 31602 26402 31614
rect 33854 31602 33906 31614
rect 34750 31666 34802 31678
rect 34750 31602 34802 31614
rect 37102 31666 37154 31678
rect 37102 31602 37154 31614
rect 38894 31666 38946 31678
rect 38894 31602 38946 31614
rect 40350 31666 40402 31678
rect 40350 31602 40402 31614
rect 40574 31666 40626 31678
rect 40574 31602 40626 31614
rect 45838 31666 45890 31678
rect 45838 31602 45890 31614
rect 47182 31666 47234 31678
rect 48862 31666 48914 31678
rect 48290 31614 48302 31666
rect 48354 31614 48366 31666
rect 47182 31602 47234 31614
rect 48862 31602 48914 31614
rect 49982 31666 50034 31678
rect 49982 31602 50034 31614
rect 51998 31666 52050 31678
rect 56018 31614 56030 31666
rect 56082 31614 56094 31666
rect 51998 31602 52050 31614
rect 14254 31554 14306 31566
rect 14254 31490 14306 31502
rect 15486 31554 15538 31566
rect 15486 31490 15538 31502
rect 21982 31554 22034 31566
rect 21982 31490 22034 31502
rect 25678 31554 25730 31566
rect 27806 31554 27858 31566
rect 26674 31502 26686 31554
rect 26738 31502 26750 31554
rect 25678 31490 25730 31502
rect 27806 31490 27858 31502
rect 34302 31554 34354 31566
rect 34302 31490 34354 31502
rect 35198 31554 35250 31566
rect 35198 31490 35250 31502
rect 35982 31554 36034 31566
rect 35982 31490 36034 31502
rect 36430 31554 36482 31566
rect 38334 31554 38386 31566
rect 37538 31502 37550 31554
rect 37602 31502 37614 31554
rect 36430 31490 36482 31502
rect 38334 31490 38386 31502
rect 44942 31554 44994 31566
rect 44942 31490 44994 31502
rect 46958 31554 47010 31566
rect 46958 31490 47010 31502
rect 48974 31554 49026 31566
rect 48974 31490 49026 31502
rect 49758 31554 49810 31566
rect 50306 31502 50318 31554
rect 50370 31502 50382 31554
rect 49758 31490 49810 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 13470 31218 13522 31230
rect 13470 31154 13522 31166
rect 14030 31218 14082 31230
rect 14030 31154 14082 31166
rect 17390 31218 17442 31230
rect 24222 31218 24274 31230
rect 19170 31166 19182 31218
rect 19234 31166 19246 31218
rect 22978 31166 22990 31218
rect 23042 31166 23054 31218
rect 17390 31154 17442 31166
rect 24222 31154 24274 31166
rect 47070 31218 47122 31230
rect 47070 31154 47122 31166
rect 47518 31218 47570 31230
rect 53666 31166 53678 31218
rect 53730 31166 53742 31218
rect 47518 31154 47570 31166
rect 13246 31106 13298 31118
rect 13246 31042 13298 31054
rect 16830 31106 16882 31118
rect 16830 31042 16882 31054
rect 17502 31106 17554 31118
rect 24446 31106 24498 31118
rect 41918 31106 41970 31118
rect 18274 31054 18286 31106
rect 18338 31054 18350 31106
rect 23090 31054 23102 31106
rect 23154 31054 23166 31106
rect 23874 31054 23886 31106
rect 23938 31054 23950 31106
rect 34402 31054 34414 31106
rect 34466 31054 34478 31106
rect 37650 31054 37662 31106
rect 37714 31054 37726 31106
rect 17502 31042 17554 31054
rect 24446 31042 24498 31054
rect 41918 31042 41970 31054
rect 43486 31106 43538 31118
rect 43934 31106 43986 31118
rect 43586 31054 43598 31106
rect 43650 31054 43662 31106
rect 43486 31042 43538 31054
rect 43934 31042 43986 31054
rect 44718 31106 44770 31118
rect 44718 31042 44770 31054
rect 45838 31106 45890 31118
rect 45838 31042 45890 31054
rect 48750 31106 48802 31118
rect 48750 31042 48802 31054
rect 54462 31106 54514 31118
rect 54462 31042 54514 31054
rect 24558 30994 24610 31006
rect 32510 30994 32562 31006
rect 41470 30994 41522 31006
rect 9538 30942 9550 30994
rect 9602 30942 9614 30994
rect 16146 30942 16158 30994
rect 16210 30942 16222 30994
rect 18162 30942 18174 30994
rect 18226 30942 18238 30994
rect 19058 30942 19070 30994
rect 19122 30942 19134 30994
rect 19618 30942 19630 30994
rect 19682 30942 19694 30994
rect 23986 30942 23998 30994
rect 24050 30942 24062 30994
rect 32050 30942 32062 30994
rect 32114 30942 32126 30994
rect 33730 30942 33742 30994
rect 33794 30942 33806 30994
rect 36866 30942 36878 30994
rect 36930 30942 36942 30994
rect 24558 30930 24610 30942
rect 32510 30930 32562 30942
rect 41470 30930 41522 30942
rect 42142 30994 42194 31006
rect 44158 30994 44210 31006
rect 43250 30942 43262 30994
rect 43314 30942 43326 30994
rect 42142 30930 42194 30942
rect 44158 30930 44210 30942
rect 44270 30994 44322 31006
rect 44270 30930 44322 30942
rect 44830 30994 44882 31006
rect 44830 30930 44882 30942
rect 45502 30994 45554 31006
rect 45502 30930 45554 30942
rect 46398 30994 46450 31006
rect 46398 30930 46450 30942
rect 48078 30994 48130 31006
rect 48078 30930 48130 30942
rect 48862 30994 48914 31006
rect 48862 30930 48914 30942
rect 49086 30994 49138 31006
rect 49086 30930 49138 30942
rect 49198 30994 49250 31006
rect 52446 30994 52498 31006
rect 51090 30942 51102 30994
rect 51154 30942 51166 30994
rect 51426 30942 51438 30994
rect 51490 30942 51502 30994
rect 49198 30930 49250 30942
rect 52446 30930 52498 30942
rect 52782 30994 52834 31006
rect 52782 30930 52834 30942
rect 53006 30994 53058 31006
rect 53890 30942 53902 30994
rect 53954 30942 53966 30994
rect 53006 30930 53058 30942
rect 12910 30882 12962 30894
rect 10322 30830 10334 30882
rect 10386 30830 10398 30882
rect 12450 30830 12462 30882
rect 12514 30830 12526 30882
rect 16370 30830 16382 30882
rect 16434 30830 16446 30882
rect 20402 30830 20414 30882
rect 20466 30830 20478 30882
rect 22530 30830 22542 30882
rect 22594 30830 22606 30882
rect 29138 30830 29150 30882
rect 29202 30830 29214 30882
rect 31266 30830 31278 30882
rect 31330 30830 31342 30882
rect 36530 30830 36542 30882
rect 36594 30830 36606 30882
rect 39778 30830 39790 30882
rect 39842 30830 39854 30882
rect 41010 30830 41022 30882
rect 41074 30830 41086 30882
rect 49858 30830 49870 30882
rect 49922 30830 49934 30882
rect 51986 30830 51998 30882
rect 52050 30830 52062 30882
rect 12910 30818 12962 30830
rect 13582 30770 13634 30782
rect 13582 30706 13634 30718
rect 13918 30770 13970 30782
rect 13918 30706 13970 30718
rect 14254 30770 14306 30782
rect 14254 30706 14306 30718
rect 42478 30770 42530 30782
rect 42478 30706 42530 30718
rect 44718 30770 44770 30782
rect 44718 30706 44770 30718
rect 45390 30770 45442 30782
rect 45390 30706 45442 30718
rect 45726 30770 45778 30782
rect 45726 30706 45778 30718
rect 46286 30770 46338 30782
rect 46286 30706 46338 30718
rect 46622 30770 46674 30782
rect 53330 30718 53342 30770
rect 53394 30718 53406 30770
rect 46622 30706 46674 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 20414 30434 20466 30446
rect 20414 30370 20466 30382
rect 20750 30434 20802 30446
rect 20750 30370 20802 30382
rect 21310 30434 21362 30446
rect 21310 30370 21362 30382
rect 21646 30434 21698 30446
rect 21646 30370 21698 30382
rect 29822 30434 29874 30446
rect 29822 30370 29874 30382
rect 36094 30434 36146 30446
rect 36094 30370 36146 30382
rect 39566 30434 39618 30446
rect 39566 30370 39618 30382
rect 19294 30322 19346 30334
rect 35758 30322 35810 30334
rect 14242 30270 14254 30322
rect 14306 30270 14318 30322
rect 16370 30270 16382 30322
rect 16434 30270 16446 30322
rect 25218 30270 25230 30322
rect 25282 30270 25294 30322
rect 19294 30258 19346 30270
rect 35758 30258 35810 30270
rect 16830 30210 16882 30222
rect 19742 30210 19794 30222
rect 26574 30210 26626 30222
rect 28254 30210 28306 30222
rect 36990 30210 37042 30222
rect 39454 30210 39506 30222
rect 13458 30158 13470 30210
rect 13522 30158 13534 30210
rect 17490 30158 17502 30210
rect 17554 30158 17566 30210
rect 18610 30158 18622 30210
rect 18674 30158 18686 30210
rect 21298 30158 21310 30210
rect 21362 30158 21374 30210
rect 22978 30158 22990 30210
rect 23042 30158 23054 30210
rect 24322 30158 24334 30210
rect 24386 30158 24398 30210
rect 25442 30158 25454 30210
rect 25506 30158 25518 30210
rect 27010 30158 27022 30210
rect 27074 30158 27086 30210
rect 29810 30158 29822 30210
rect 29874 30158 29886 30210
rect 30258 30158 30270 30210
rect 30322 30158 30334 30210
rect 33618 30158 33630 30210
rect 33682 30158 33694 30210
rect 37314 30158 37326 30210
rect 37378 30158 37390 30210
rect 38098 30158 38110 30210
rect 38162 30158 38174 30210
rect 38770 30158 38782 30210
rect 38834 30158 38846 30210
rect 16830 30146 16882 30158
rect 19742 30146 19794 30158
rect 26574 30146 26626 30158
rect 28254 30146 28306 30158
rect 36990 30146 37042 30158
rect 39454 30146 39506 30158
rect 40126 30210 40178 30222
rect 40126 30146 40178 30158
rect 40798 30210 40850 30222
rect 40798 30146 40850 30158
rect 41134 30210 41186 30222
rect 41134 30146 41186 30158
rect 41806 30210 41858 30222
rect 41806 30146 41858 30158
rect 42478 30210 42530 30222
rect 42478 30146 42530 30158
rect 43150 30210 43202 30222
rect 43150 30146 43202 30158
rect 45054 30210 45106 30222
rect 45054 30146 45106 30158
rect 45614 30210 45666 30222
rect 46274 30158 46286 30210
rect 46338 30158 46350 30210
rect 46834 30158 46846 30210
rect 46898 30158 46910 30210
rect 47618 30158 47630 30210
rect 47682 30158 47694 30210
rect 48962 30158 48974 30210
rect 49026 30158 49038 30210
rect 50194 30158 50206 30210
rect 50258 30158 50270 30210
rect 50530 30158 50542 30210
rect 50594 30158 50606 30210
rect 53106 30158 53118 30210
rect 53170 30158 53182 30210
rect 53778 30158 53790 30210
rect 53842 30158 53854 30210
rect 45614 30146 45666 30158
rect 9550 30098 9602 30110
rect 9550 30034 9602 30046
rect 9886 30098 9938 30110
rect 20526 30098 20578 30110
rect 26462 30098 26514 30110
rect 17938 30046 17950 30098
rect 18002 30046 18014 30098
rect 25778 30046 25790 30098
rect 25842 30046 25854 30098
rect 9886 30034 9938 30046
rect 20526 30034 20578 30046
rect 26462 30034 26514 30046
rect 28590 30098 28642 30110
rect 28590 30034 28642 30046
rect 29486 30098 29538 30110
rect 41470 30098 41522 30110
rect 39218 30046 39230 30098
rect 39282 30046 39294 30098
rect 40450 30046 40462 30098
rect 40514 30046 40526 30098
rect 29486 30034 29538 30046
rect 41470 30034 41522 30046
rect 45166 30098 45218 30110
rect 46946 30046 46958 30098
rect 47010 30046 47022 30098
rect 47954 30046 47966 30098
rect 48018 30046 48030 30098
rect 51538 30046 51550 30098
rect 51602 30046 51614 30098
rect 53554 30046 53566 30098
rect 53618 30046 53630 30098
rect 45166 30034 45218 30046
rect 22094 29986 22146 29998
rect 18386 29934 18398 29986
rect 18450 29934 18462 29986
rect 22094 29922 22146 29934
rect 28478 29986 28530 29998
rect 28478 29922 28530 29934
rect 35982 29986 36034 29998
rect 35982 29922 36034 29934
rect 39790 29986 39842 29998
rect 45278 29986 45330 29998
rect 42130 29934 42142 29986
rect 42194 29934 42206 29986
rect 42802 29934 42814 29986
rect 42866 29934 42878 29986
rect 43474 29934 43486 29986
rect 43538 29934 43550 29986
rect 39790 29922 39842 29934
rect 45278 29922 45330 29934
rect 45726 29986 45778 29998
rect 50866 29934 50878 29986
rect 50930 29934 50942 29986
rect 52882 29934 52894 29986
rect 52946 29934 52958 29986
rect 45726 29922 45778 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 10334 29650 10386 29662
rect 10334 29586 10386 29598
rect 16270 29650 16322 29662
rect 16270 29586 16322 29598
rect 18174 29650 18226 29662
rect 18174 29586 18226 29598
rect 19518 29650 19570 29662
rect 19518 29586 19570 29598
rect 29038 29650 29090 29662
rect 29038 29586 29090 29598
rect 31278 29650 31330 29662
rect 31278 29586 31330 29598
rect 32398 29650 32450 29662
rect 32398 29586 32450 29598
rect 33182 29650 33234 29662
rect 48862 29650 48914 29662
rect 34850 29598 34862 29650
rect 34914 29598 34926 29650
rect 47506 29598 47518 29650
rect 47570 29598 47582 29650
rect 51650 29598 51662 29650
rect 51714 29598 51726 29650
rect 33182 29586 33234 29598
rect 48862 29586 48914 29598
rect 28814 29538 28866 29550
rect 11218 29486 11230 29538
rect 11282 29486 11294 29538
rect 13682 29486 13694 29538
rect 13746 29486 13758 29538
rect 25330 29486 25342 29538
rect 25394 29486 25406 29538
rect 28814 29474 28866 29486
rect 29486 29538 29538 29550
rect 29486 29474 29538 29486
rect 30158 29538 30210 29550
rect 30158 29474 30210 29486
rect 30270 29538 30322 29550
rect 30270 29474 30322 29486
rect 30830 29538 30882 29550
rect 30830 29474 30882 29486
rect 35422 29538 35474 29550
rect 48078 29538 48130 29550
rect 52110 29538 52162 29550
rect 41234 29486 41246 29538
rect 41298 29486 41310 29538
rect 45826 29486 45838 29538
rect 45890 29486 45902 29538
rect 46498 29486 46510 29538
rect 46562 29486 46574 29538
rect 49634 29486 49646 29538
rect 49698 29486 49710 29538
rect 35422 29474 35474 29486
rect 48078 29474 48130 29486
rect 52110 29474 52162 29486
rect 52222 29538 52274 29550
rect 52222 29474 52274 29486
rect 53342 29538 53394 29550
rect 53342 29474 53394 29486
rect 8542 29426 8594 29438
rect 28702 29426 28754 29438
rect 5282 29374 5294 29426
rect 5346 29374 5358 29426
rect 11442 29374 11454 29426
rect 11506 29374 11518 29426
rect 12898 29374 12910 29426
rect 12962 29374 12974 29426
rect 21298 29374 21310 29426
rect 21362 29374 21374 29426
rect 25442 29374 25454 29426
rect 25506 29374 25518 29426
rect 25666 29374 25678 29426
rect 25730 29374 25742 29426
rect 26450 29374 26462 29426
rect 26514 29374 26526 29426
rect 8542 29362 8594 29374
rect 28702 29362 28754 29374
rect 29374 29426 29426 29438
rect 29374 29362 29426 29374
rect 29934 29426 29986 29438
rect 29934 29362 29986 29374
rect 31950 29426 32002 29438
rect 31950 29362 32002 29374
rect 32174 29426 32226 29438
rect 32174 29362 32226 29374
rect 32622 29426 32674 29438
rect 44158 29426 44210 29438
rect 50430 29426 50482 29438
rect 53454 29426 53506 29438
rect 34178 29374 34190 29426
rect 34242 29374 34254 29426
rect 41010 29374 41022 29426
rect 41074 29374 41086 29426
rect 45154 29374 45166 29426
rect 45218 29374 45230 29426
rect 46050 29374 46062 29426
rect 46114 29374 46126 29426
rect 46610 29374 46622 29426
rect 46674 29374 46686 29426
rect 49746 29374 49758 29426
rect 49810 29374 49822 29426
rect 50530 29374 50542 29426
rect 50594 29374 50606 29426
rect 52434 29374 52446 29426
rect 52498 29374 52510 29426
rect 53106 29374 53118 29426
rect 53170 29374 53182 29426
rect 32622 29362 32674 29374
rect 44158 29362 44210 29374
rect 50430 29362 50482 29374
rect 53454 29362 53506 29374
rect 53678 29426 53730 29438
rect 53678 29362 53730 29374
rect 54574 29426 54626 29438
rect 54574 29362 54626 29374
rect 18286 29314 18338 29326
rect 5954 29262 5966 29314
rect 6018 29262 6030 29314
rect 8082 29262 8094 29314
rect 8146 29262 8158 29314
rect 15810 29262 15822 29314
rect 15874 29262 15886 29314
rect 18286 29250 18338 29262
rect 18958 29314 19010 29326
rect 24670 29314 24722 29326
rect 21970 29262 21982 29314
rect 22034 29262 22046 29314
rect 24098 29262 24110 29314
rect 24162 29262 24174 29314
rect 18958 29250 19010 29262
rect 24670 29250 24722 29262
rect 29710 29314 29762 29326
rect 29710 29250 29762 29262
rect 33518 29314 33570 29326
rect 35198 29314 35250 29326
rect 34402 29262 34414 29314
rect 34466 29262 34478 29314
rect 33518 29250 33570 29262
rect 35198 29250 35250 29262
rect 43710 29314 43762 29326
rect 47854 29314 47906 29326
rect 54014 29314 54066 29326
rect 46946 29262 46958 29314
rect 47010 29262 47022 29314
rect 49970 29262 49982 29314
rect 50034 29262 50046 29314
rect 43710 29250 43762 29262
rect 47854 29250 47906 29262
rect 54014 29250 54066 29262
rect 55022 29314 55074 29326
rect 55022 29250 55074 29262
rect 10670 29202 10722 29214
rect 10670 29138 10722 29150
rect 30270 29202 30322 29214
rect 30270 29138 30322 29150
rect 30718 29202 30770 29214
rect 30718 29138 30770 29150
rect 52670 29202 52722 29214
rect 52670 29138 52722 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 21982 28866 22034 28878
rect 21982 28802 22034 28814
rect 27582 28866 27634 28878
rect 27582 28802 27634 28814
rect 28254 28866 28306 28878
rect 28254 28802 28306 28814
rect 33406 28866 33458 28878
rect 33406 28802 33458 28814
rect 35198 28866 35250 28878
rect 35198 28802 35250 28814
rect 46174 28866 46226 28878
rect 46174 28802 46226 28814
rect 46846 28866 46898 28878
rect 46846 28802 46898 28814
rect 19518 28754 19570 28766
rect 12002 28702 12014 28754
rect 12066 28702 12078 28754
rect 16706 28702 16718 28754
rect 16770 28702 16782 28754
rect 19518 28690 19570 28702
rect 23214 28754 23266 28766
rect 37102 28754 37154 28766
rect 23538 28702 23550 28754
rect 23602 28702 23614 28754
rect 27906 28702 27918 28754
rect 27970 28702 27982 28754
rect 28578 28702 28590 28754
rect 28642 28702 28654 28754
rect 29138 28702 29150 28754
rect 29202 28702 29214 28754
rect 31266 28702 31278 28754
rect 31330 28702 31342 28754
rect 23214 28690 23266 28702
rect 37102 28690 37154 28702
rect 37998 28754 38050 28766
rect 37998 28690 38050 28702
rect 39678 28754 39730 28766
rect 39678 28690 39730 28702
rect 45502 28754 45554 28766
rect 45502 28690 45554 28702
rect 45614 28754 45666 28766
rect 48626 28702 48638 28754
rect 48690 28702 48702 28754
rect 55234 28702 55246 28754
rect 55298 28702 55310 28754
rect 57362 28702 57374 28754
rect 57426 28702 57438 28754
rect 45614 28690 45666 28702
rect 7198 28642 7250 28654
rect 6514 28590 6526 28642
rect 6578 28590 6590 28642
rect 7198 28578 7250 28590
rect 7534 28642 7586 28654
rect 12462 28642 12514 28654
rect 26686 28642 26738 28654
rect 9202 28590 9214 28642
rect 9266 28590 9278 28642
rect 15922 28590 15934 28642
rect 15986 28590 15998 28642
rect 23650 28590 23662 28642
rect 23714 28590 23726 28642
rect 7534 28578 7586 28590
rect 12462 28578 12514 28590
rect 26686 28578 26738 28590
rect 26798 28642 26850 28654
rect 32622 28642 32674 28654
rect 27122 28590 27134 28642
rect 27186 28590 27198 28642
rect 32050 28590 32062 28642
rect 32114 28590 32126 28642
rect 26798 28578 26850 28590
rect 32622 28578 32674 28590
rect 32958 28642 33010 28654
rect 32958 28578 33010 28590
rect 33182 28642 33234 28654
rect 33966 28642 34018 28654
rect 33618 28590 33630 28642
rect 33682 28590 33694 28642
rect 33182 28578 33234 28590
rect 33966 28578 34018 28590
rect 34526 28642 34578 28654
rect 34526 28578 34578 28590
rect 34862 28642 34914 28654
rect 34862 28578 34914 28590
rect 36206 28642 36258 28654
rect 40014 28642 40066 28654
rect 42590 28642 42642 28654
rect 37538 28590 37550 28642
rect 37602 28590 37614 28642
rect 38322 28590 38334 28642
rect 38386 28590 38398 28642
rect 40674 28590 40686 28642
rect 40738 28590 40750 28642
rect 36206 28578 36258 28590
rect 40014 28578 40066 28590
rect 42590 28578 42642 28590
rect 43374 28642 43426 28654
rect 43374 28578 43426 28590
rect 43934 28642 43986 28654
rect 43934 28578 43986 28590
rect 45166 28642 45218 28654
rect 45166 28578 45218 28590
rect 45950 28642 46002 28654
rect 50318 28642 50370 28654
rect 52670 28642 52722 28654
rect 49298 28590 49310 28642
rect 49362 28590 49374 28642
rect 50978 28590 50990 28642
rect 51042 28590 51054 28642
rect 52098 28590 52110 28642
rect 52162 28590 52174 28642
rect 53218 28590 53230 28642
rect 53282 28590 53294 28642
rect 53890 28590 53902 28642
rect 53954 28590 53966 28642
rect 54562 28590 54574 28642
rect 54626 28590 54638 28642
rect 45950 28578 46002 28590
rect 50318 28578 50370 28590
rect 52670 28578 52722 28590
rect 6302 28530 6354 28542
rect 21310 28530 21362 28542
rect 7746 28478 7758 28530
rect 7810 28478 7822 28530
rect 8082 28478 8094 28530
rect 8146 28478 8158 28530
rect 9874 28478 9886 28530
rect 9938 28478 9950 28530
rect 6302 28466 6354 28478
rect 21310 28466 21362 28478
rect 22094 28530 22146 28542
rect 22094 28466 22146 28478
rect 22318 28530 22370 28542
rect 22318 28466 22370 28478
rect 26350 28530 26402 28542
rect 26350 28466 26402 28478
rect 27806 28530 27858 28542
rect 27806 28466 27858 28478
rect 28478 28530 28530 28542
rect 28478 28466 28530 28478
rect 32510 28530 32562 28542
rect 32510 28466 32562 28478
rect 35310 28530 35362 28542
rect 35310 28466 35362 28478
rect 38670 28530 38722 28542
rect 38670 28466 38722 28478
rect 41022 28530 41074 28542
rect 41022 28466 41074 28478
rect 46958 28530 47010 28542
rect 51986 28478 51998 28530
rect 52050 28478 52062 28530
rect 52882 28478 52894 28530
rect 52946 28478 52958 28530
rect 46958 28466 47010 28478
rect 27134 28418 27186 28430
rect 18946 28366 18958 28418
rect 19010 28366 19022 28418
rect 21634 28366 21646 28418
rect 21698 28366 21710 28418
rect 27134 28354 27186 28366
rect 32846 28418 32898 28430
rect 32846 28354 32898 28366
rect 34638 28418 34690 28430
rect 34638 28354 34690 28366
rect 35198 28418 35250 28430
rect 35198 28354 35250 28366
rect 35758 28418 35810 28430
rect 40910 28418 40962 28430
rect 52782 28418 52834 28430
rect 40338 28366 40350 28418
rect 40402 28366 40414 28418
rect 42914 28366 42926 28418
rect 42978 28366 42990 28418
rect 46498 28366 46510 28418
rect 46562 28366 46574 28418
rect 51090 28366 51102 28418
rect 51154 28366 51166 28418
rect 35758 28354 35810 28366
rect 40910 28354 40962 28366
rect 52782 28354 52834 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 9774 28082 9826 28094
rect 9774 28018 9826 28030
rect 19742 28082 19794 28094
rect 19742 28018 19794 28030
rect 19854 28082 19906 28094
rect 19854 28018 19906 28030
rect 25454 28082 25506 28094
rect 41694 28082 41746 28094
rect 47630 28082 47682 28094
rect 39330 28030 39342 28082
rect 39394 28030 39406 28082
rect 46274 28030 46286 28082
rect 46338 28030 46350 28082
rect 25454 28018 25506 28030
rect 41694 28018 41746 28030
rect 47630 28018 47682 28030
rect 47854 28082 47906 28094
rect 47854 28018 47906 28030
rect 52110 28082 52162 28094
rect 52110 28018 52162 28030
rect 55134 28082 55186 28094
rect 55134 28018 55186 28030
rect 55582 28082 55634 28094
rect 55582 28018 55634 28030
rect 55694 28082 55746 28094
rect 55694 28018 55746 28030
rect 56590 28082 56642 28094
rect 56590 28018 56642 28030
rect 8430 27970 8482 27982
rect 20526 27970 20578 27982
rect 7858 27918 7870 27970
rect 7922 27918 7934 27970
rect 11442 27918 11454 27970
rect 11506 27918 11518 27970
rect 19282 27918 19294 27970
rect 19346 27918 19358 27970
rect 8430 27906 8482 27918
rect 20526 27906 20578 27918
rect 22318 27970 22370 27982
rect 25342 27970 25394 27982
rect 22642 27918 22654 27970
rect 22706 27918 22718 27970
rect 22318 27906 22370 27918
rect 25342 27906 25394 27918
rect 25566 27970 25618 27982
rect 34526 27970 34578 27982
rect 36206 27970 36258 27982
rect 39230 27970 39282 27982
rect 28130 27918 28142 27970
rect 28194 27918 28206 27970
rect 30146 27918 30158 27970
rect 30210 27918 30222 27970
rect 35970 27918 35982 27970
rect 36034 27918 36046 27970
rect 36642 27918 36654 27970
rect 36706 27918 36718 27970
rect 25566 27906 25618 27918
rect 34526 27906 34578 27918
rect 36206 27906 36258 27918
rect 39230 27906 39282 27918
rect 46734 27970 46786 27982
rect 52658 27918 52670 27970
rect 52722 27918 52734 27970
rect 52994 27918 53006 27970
rect 53058 27918 53070 27970
rect 46734 27906 46786 27918
rect 10110 27858 10162 27870
rect 3490 27806 3502 27858
rect 3554 27806 3566 27858
rect 7746 27806 7758 27858
rect 7810 27806 7822 27858
rect 10110 27794 10162 27806
rect 10558 27858 10610 27870
rect 21086 27858 21138 27870
rect 23998 27858 24050 27870
rect 11330 27806 11342 27858
rect 11394 27806 11406 27858
rect 19058 27806 19070 27858
rect 19122 27806 19134 27858
rect 20738 27806 20750 27858
rect 20802 27806 20814 27858
rect 21634 27806 21646 27858
rect 21698 27806 21710 27858
rect 22866 27806 22878 27858
rect 22930 27806 22942 27858
rect 10558 27794 10610 27806
rect 21086 27794 21138 27806
rect 23998 27794 24050 27806
rect 24446 27858 24498 27870
rect 24446 27794 24498 27806
rect 24558 27858 24610 27870
rect 34078 27858 34130 27870
rect 28802 27806 28814 27858
rect 28866 27806 28878 27858
rect 29362 27806 29374 27858
rect 29426 27806 29438 27858
rect 33394 27806 33406 27858
rect 33458 27806 33470 27858
rect 24558 27794 24610 27806
rect 34078 27794 34130 27806
rect 34302 27858 34354 27870
rect 34302 27794 34354 27806
rect 34750 27858 34802 27870
rect 34750 27794 34802 27806
rect 34862 27858 34914 27870
rect 38670 27858 38722 27870
rect 35522 27806 35534 27858
rect 35586 27806 35598 27858
rect 36530 27806 36542 27858
rect 36594 27806 36606 27858
rect 34862 27794 34914 27806
rect 38670 27794 38722 27806
rect 41806 27858 41858 27870
rect 41806 27794 41858 27806
rect 41918 27858 41970 27870
rect 46846 27858 46898 27870
rect 43026 27806 43038 27858
rect 43090 27806 43102 27858
rect 41918 27794 41970 27806
rect 46846 27794 46898 27806
rect 46958 27858 47010 27870
rect 46958 27794 47010 27806
rect 47406 27858 47458 27870
rect 51662 27858 51714 27870
rect 49186 27806 49198 27858
rect 49250 27806 49262 27858
rect 47406 27794 47458 27806
rect 51662 27794 51714 27806
rect 51886 27858 51938 27870
rect 54350 27858 54402 27870
rect 56702 27858 56754 27870
rect 52770 27806 52782 27858
rect 52834 27806 52846 27858
rect 54674 27806 54686 27858
rect 54738 27806 54750 27858
rect 54898 27806 54910 27858
rect 54962 27806 54974 27858
rect 51886 27794 51938 27806
rect 54350 27794 54402 27806
rect 56702 27794 56754 27806
rect 7086 27746 7138 27758
rect 4162 27694 4174 27746
rect 4226 27694 4238 27746
rect 6290 27694 6302 27746
rect 6354 27694 6366 27746
rect 7086 27682 7138 27694
rect 18734 27746 18786 27758
rect 24222 27746 24274 27758
rect 36094 27746 36146 27758
rect 21410 27694 21422 27746
rect 21474 27694 21486 27746
rect 26002 27694 26014 27746
rect 26066 27694 26078 27746
rect 32386 27694 32398 27746
rect 32450 27694 32462 27746
rect 33282 27694 33294 27746
rect 33346 27694 33358 27746
rect 18734 27682 18786 27694
rect 24222 27682 24274 27694
rect 36094 27682 36146 27694
rect 42142 27746 42194 27758
rect 47518 27746 47570 27758
rect 51774 27746 51826 27758
rect 43698 27694 43710 27746
rect 43762 27694 43774 27746
rect 45826 27694 45838 27746
rect 45890 27694 45902 27746
rect 50418 27694 50430 27746
rect 50482 27694 50494 27746
rect 42142 27682 42194 27694
rect 47518 27682 47570 27694
rect 51774 27682 51826 27694
rect 53790 27746 53842 27758
rect 53790 27682 53842 27694
rect 55470 27746 55522 27758
rect 55470 27682 55522 27694
rect 6750 27634 6802 27646
rect 6750 27570 6802 27582
rect 8318 27634 8370 27646
rect 8318 27570 8370 27582
rect 10894 27634 10946 27646
rect 10894 27570 10946 27582
rect 19966 27634 20018 27646
rect 19966 27570 20018 27582
rect 20414 27634 20466 27646
rect 20414 27570 20466 27582
rect 35758 27634 35810 27646
rect 35758 27570 35810 27582
rect 42366 27634 42418 27646
rect 42366 27570 42418 27582
rect 54798 27634 54850 27646
rect 54798 27570 54850 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 34526 27298 34578 27310
rect 34526 27234 34578 27246
rect 37438 27298 37490 27310
rect 37438 27234 37490 27246
rect 7086 27186 7138 27198
rect 19406 27186 19458 27198
rect 16258 27134 16270 27186
rect 16322 27134 16334 27186
rect 18386 27134 18398 27186
rect 18450 27134 18462 27186
rect 18722 27134 18734 27186
rect 18786 27134 18798 27186
rect 20290 27134 20302 27186
rect 20354 27134 20366 27186
rect 26562 27160 26574 27212
rect 26626 27160 26638 27212
rect 42366 27186 42418 27198
rect 49422 27186 49474 27198
rect 33506 27134 33518 27186
rect 33570 27134 33582 27186
rect 38770 27134 38782 27186
rect 38834 27134 38846 27186
rect 40898 27134 40910 27186
rect 40962 27134 40974 27186
rect 46722 27134 46734 27186
rect 46786 27134 46798 27186
rect 7086 27122 7138 27134
rect 19406 27122 19458 27134
rect 42366 27122 42418 27134
rect 49422 27122 49474 27134
rect 49646 27186 49698 27198
rect 49646 27122 49698 27134
rect 50206 27186 50258 27198
rect 53006 27186 53058 27198
rect 50530 27134 50542 27186
rect 50594 27134 50606 27186
rect 51986 27134 51998 27186
rect 52050 27134 52062 27186
rect 57026 27134 57038 27186
rect 57090 27134 57102 27186
rect 50206 27122 50258 27134
rect 53006 27122 53058 27134
rect 4958 27074 5010 27086
rect 21310 27074 21362 27086
rect 27022 27074 27074 27086
rect 15474 27022 15486 27074
rect 15538 27022 15550 27074
rect 20066 27022 20078 27074
rect 20130 27022 20142 27074
rect 21858 27022 21870 27074
rect 21922 27022 21934 27074
rect 22530 27022 22542 27074
rect 22594 27022 22606 27074
rect 23762 27022 23774 27074
rect 23826 27022 23838 27074
rect 4958 27010 5010 27022
rect 21310 27010 21362 27022
rect 27022 27010 27074 27022
rect 29262 27074 29314 27086
rect 37214 27074 37266 27086
rect 33394 27022 33406 27074
rect 33458 27022 33470 27074
rect 34402 27022 34414 27074
rect 34466 27022 34478 27074
rect 34626 27022 34638 27074
rect 34690 27022 34702 27074
rect 36082 27022 36094 27074
rect 36146 27022 36158 27074
rect 29262 27010 29314 27022
rect 37214 27010 37266 27022
rect 37550 27074 37602 27086
rect 37550 27010 37602 27022
rect 37998 27074 38050 27086
rect 42254 27074 42306 27086
rect 41682 27022 41694 27074
rect 41746 27022 41758 27074
rect 37998 27010 38050 27022
rect 42254 27010 42306 27022
rect 42926 27074 42978 27086
rect 42926 27010 42978 27022
rect 43710 27074 43762 27086
rect 43710 27010 43762 27022
rect 44158 27074 44210 27086
rect 48526 27074 48578 27086
rect 44818 27022 44830 27074
rect 44882 27022 44894 27074
rect 44158 27010 44210 27022
rect 48526 27010 48578 27022
rect 48862 27074 48914 27086
rect 48862 27010 48914 27022
rect 49870 27074 49922 27086
rect 51550 27074 51602 27086
rect 50642 27022 50654 27074
rect 50706 27022 50718 27074
rect 52770 27022 52782 27074
rect 52834 27022 52846 27074
rect 53218 27022 53230 27074
rect 53282 27022 53294 27074
rect 54114 27022 54126 27074
rect 54178 27022 54190 27074
rect 49870 27010 49922 27022
rect 51550 27010 51602 27022
rect 4622 26962 4674 26974
rect 4622 26898 4674 26910
rect 5630 26962 5682 26974
rect 5630 26898 5682 26910
rect 5966 26962 6018 26974
rect 5966 26898 6018 26910
rect 13470 26962 13522 26974
rect 13470 26898 13522 26910
rect 13806 26962 13858 26974
rect 13806 26898 13858 26910
rect 18846 26962 18898 26974
rect 18846 26898 18898 26910
rect 19070 26962 19122 26974
rect 19070 26898 19122 26910
rect 21198 26962 21250 26974
rect 29710 26962 29762 26974
rect 21522 26910 21534 26962
rect 21586 26910 21598 26962
rect 24434 26910 24446 26962
rect 24498 26910 24510 26962
rect 21198 26898 21250 26910
rect 29710 26898 29762 26910
rect 33854 26962 33906 26974
rect 33854 26898 33906 26910
rect 34190 26962 34242 26974
rect 36990 26962 37042 26974
rect 35858 26910 35870 26962
rect 35922 26910 35934 26962
rect 34190 26898 34242 26910
rect 36990 26898 37042 26910
rect 42478 26962 42530 26974
rect 42478 26898 42530 26910
rect 43150 26962 43202 26974
rect 43150 26898 43202 26910
rect 43262 26962 43314 26974
rect 43262 26898 43314 26910
rect 43486 26962 43538 26974
rect 43486 26898 43538 26910
rect 44046 26962 44098 26974
rect 44046 26898 44098 26910
rect 45950 26962 46002 26974
rect 53342 26962 53394 26974
rect 48626 26910 48638 26962
rect 48690 26910 48702 26962
rect 49186 26910 49198 26962
rect 49250 26910 49262 26962
rect 45950 26898 46002 26910
rect 53342 26898 53394 26910
rect 53454 26962 53506 26974
rect 54898 26910 54910 26962
rect 54962 26910 54974 26962
rect 53454 26898 53506 26910
rect 6526 26850 6578 26862
rect 6526 26786 6578 26798
rect 6974 26850 7026 26862
rect 6974 26786 7026 26798
rect 15150 26850 15202 26862
rect 15150 26786 15202 26798
rect 23438 26850 23490 26862
rect 23438 26786 23490 26798
rect 35086 26850 35138 26862
rect 35086 26786 35138 26798
rect 35534 26850 35586 26862
rect 35534 26786 35586 26798
rect 37102 26850 37154 26862
rect 37102 26786 37154 26798
rect 38334 26850 38386 26862
rect 38334 26786 38386 26798
rect 49982 26850 50034 26862
rect 49982 26786 50034 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 16606 26514 16658 26526
rect 25566 26514 25618 26526
rect 15362 26462 15374 26514
rect 15426 26462 15438 26514
rect 24210 26462 24222 26514
rect 24274 26462 24286 26514
rect 16606 26450 16658 26462
rect 25566 26450 25618 26462
rect 32510 26514 32562 26526
rect 32510 26450 32562 26462
rect 34862 26514 34914 26526
rect 34862 26450 34914 26462
rect 41918 26514 41970 26526
rect 46398 26514 46450 26526
rect 55582 26514 55634 26526
rect 44706 26462 44718 26514
rect 44770 26462 44782 26514
rect 47170 26462 47182 26514
rect 47234 26462 47246 26514
rect 41918 26450 41970 26462
rect 46398 26450 46450 26462
rect 55582 26450 55634 26462
rect 7982 26402 8034 26414
rect 4834 26350 4846 26402
rect 4898 26350 4910 26402
rect 7982 26338 8034 26350
rect 10110 26402 10162 26414
rect 19518 26402 19570 26414
rect 11666 26350 11678 26402
rect 11730 26350 11742 26402
rect 12898 26350 12910 26402
rect 12962 26350 12974 26402
rect 10110 26338 10162 26350
rect 19518 26338 19570 26350
rect 21982 26402 22034 26414
rect 21982 26338 22034 26350
rect 24446 26402 24498 26414
rect 34750 26402 34802 26414
rect 25218 26350 25230 26402
rect 25282 26350 25294 26402
rect 26450 26350 26462 26402
rect 26514 26350 26526 26402
rect 24446 26338 24498 26350
rect 34750 26338 34802 26350
rect 35086 26402 35138 26414
rect 35086 26338 35138 26350
rect 35198 26402 35250 26414
rect 40126 26402 40178 26414
rect 46622 26402 46674 26414
rect 36418 26350 36430 26402
rect 36482 26350 36494 26402
rect 45378 26350 45390 26402
rect 45442 26350 45454 26402
rect 35198 26338 35250 26350
rect 40126 26338 40178 26350
rect 46622 26338 46674 26350
rect 46846 26402 46898 26414
rect 46846 26338 46898 26350
rect 47742 26402 47794 26414
rect 47742 26338 47794 26350
rect 48302 26402 48354 26414
rect 48302 26338 48354 26350
rect 48750 26402 48802 26414
rect 48750 26338 48802 26350
rect 8318 26290 8370 26302
rect 10558 26290 10610 26302
rect 4162 26238 4174 26290
rect 4226 26238 4238 26290
rect 9874 26238 9886 26290
rect 9938 26238 9950 26290
rect 8318 26226 8370 26238
rect 10558 26226 10610 26238
rect 10894 26290 10946 26302
rect 15710 26290 15762 26302
rect 11442 26238 11454 26290
rect 11506 26238 11518 26290
rect 12226 26238 12238 26290
rect 12290 26238 12302 26290
rect 10894 26226 10946 26238
rect 15710 26226 15762 26238
rect 18286 26290 18338 26302
rect 18286 26226 18338 26238
rect 18622 26290 18674 26302
rect 20414 26290 20466 26302
rect 23998 26290 24050 26302
rect 19954 26238 19966 26290
rect 20018 26238 20030 26290
rect 21522 26238 21534 26290
rect 21586 26238 21598 26290
rect 22194 26238 22206 26290
rect 22258 26238 22270 26290
rect 22418 26238 22430 26290
rect 22482 26238 22494 26290
rect 22866 26238 22878 26290
rect 22930 26238 22942 26290
rect 23650 26238 23662 26290
rect 23714 26238 23726 26290
rect 18622 26226 18674 26238
rect 20414 26226 20466 26238
rect 23998 26226 24050 26238
rect 24110 26290 24162 26302
rect 29598 26290 29650 26302
rect 26226 26238 26238 26290
rect 26290 26238 26302 26290
rect 24110 26226 24162 26238
rect 29598 26226 29650 26238
rect 33070 26290 33122 26302
rect 33070 26226 33122 26238
rect 33294 26290 33346 26302
rect 33294 26226 33346 26238
rect 33518 26290 33570 26302
rect 34190 26290 34242 26302
rect 39790 26290 39842 26302
rect 33730 26238 33742 26290
rect 33794 26238 33806 26290
rect 33954 26238 33966 26290
rect 34018 26238 34030 26290
rect 34514 26238 34526 26290
rect 34578 26238 34590 26290
rect 35746 26238 35758 26290
rect 35810 26238 35822 26290
rect 38882 26238 38894 26290
rect 38946 26238 38958 26290
rect 33518 26226 33570 26238
rect 34190 26226 34242 26238
rect 39790 26226 39842 26238
rect 40350 26290 40402 26302
rect 40350 26226 40402 26238
rect 40910 26290 40962 26302
rect 46286 26290 46338 26302
rect 42802 26238 42814 26290
rect 42866 26238 42878 26290
rect 44034 26238 44046 26290
rect 44098 26238 44110 26290
rect 44370 26238 44382 26290
rect 44434 26238 44446 26290
rect 40910 26226 40962 26238
rect 46286 26226 46338 26238
rect 49086 26290 49138 26302
rect 49758 26290 49810 26302
rect 51438 26290 51490 26302
rect 49410 26238 49422 26290
rect 49474 26238 49486 26290
rect 50754 26238 50766 26290
rect 50818 26238 50830 26290
rect 52322 26238 52334 26290
rect 52386 26238 52398 26290
rect 49086 26226 49138 26238
rect 49758 26226 49810 26238
rect 51438 26226 51490 26238
rect 7422 26178 7474 26190
rect 16158 26178 16210 26190
rect 19182 26178 19234 26190
rect 6962 26126 6974 26178
rect 7026 26126 7038 26178
rect 15026 26126 15038 26178
rect 15090 26126 15102 26178
rect 17826 26126 17838 26178
rect 17890 26126 17902 26178
rect 7422 26114 7474 26126
rect 16158 26114 16210 26126
rect 19182 26114 19234 26126
rect 21086 26178 21138 26190
rect 21086 26114 21138 26126
rect 23326 26178 23378 26190
rect 33182 26178 33234 26190
rect 39902 26178 39954 26190
rect 49646 26178 49698 26190
rect 29138 26126 29150 26178
rect 29202 26126 29214 26178
rect 38546 26126 38558 26178
rect 38610 26126 38622 26178
rect 41346 26126 41358 26178
rect 41410 26126 41422 26178
rect 23326 26114 23378 26126
rect 33182 26114 33234 26126
rect 39902 26114 39954 26126
rect 49646 26114 49698 26126
rect 50094 26178 50146 26190
rect 51550 26178 51602 26190
rect 50866 26126 50878 26178
rect 50930 26126 50942 26178
rect 52994 26126 53006 26178
rect 53058 26126 53070 26178
rect 55122 26126 55134 26178
rect 55186 26126 55198 26178
rect 50094 26114 50146 26126
rect 51550 26114 51602 26126
rect 21870 26066 21922 26078
rect 7186 26014 7198 26066
rect 7250 26063 7262 26066
rect 7746 26063 7758 26066
rect 7250 26017 7758 26063
rect 7250 26014 7262 26017
rect 7746 26014 7758 26017
rect 7810 26014 7822 26066
rect 21870 26002 21922 26014
rect 38894 26066 38946 26078
rect 38894 26002 38946 26014
rect 39230 26066 39282 26078
rect 39230 26002 39282 26014
rect 47518 26066 47570 26078
rect 47518 26002 47570 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 13582 25730 13634 25742
rect 13582 25666 13634 25678
rect 13918 25730 13970 25742
rect 49758 25730 49810 25742
rect 23426 25678 23438 25730
rect 23490 25678 23502 25730
rect 13918 25666 13970 25678
rect 49758 25666 49810 25678
rect 50094 25730 50146 25742
rect 50094 25666 50146 25678
rect 45838 25618 45890 25630
rect 6962 25566 6974 25618
rect 7026 25566 7038 25618
rect 9090 25566 9102 25618
rect 9154 25566 9166 25618
rect 10210 25566 10222 25618
rect 10274 25566 10286 25618
rect 12338 25566 12350 25618
rect 12402 25566 12414 25618
rect 16034 25566 16046 25618
rect 16098 25566 16110 25618
rect 18162 25566 18174 25618
rect 18226 25566 18238 25618
rect 24434 25566 24446 25618
rect 24498 25566 24510 25618
rect 30706 25566 30718 25618
rect 30770 25566 30782 25618
rect 32834 25566 32846 25618
rect 32898 25566 32910 25618
rect 33618 25566 33630 25618
rect 33682 25566 33694 25618
rect 38434 25566 38446 25618
rect 38498 25566 38510 25618
rect 40562 25566 40574 25618
rect 40626 25566 40638 25618
rect 42466 25566 42478 25618
rect 42530 25566 42542 25618
rect 43250 25566 43262 25618
rect 43314 25566 43326 25618
rect 45838 25554 45890 25566
rect 46734 25618 46786 25630
rect 46734 25554 46786 25566
rect 47742 25618 47794 25630
rect 54686 25618 54738 25630
rect 52882 25566 52894 25618
rect 52946 25566 52958 25618
rect 47742 25554 47794 25566
rect 54686 25554 54738 25566
rect 18734 25506 18786 25518
rect 6290 25454 6302 25506
rect 6354 25454 6366 25506
rect 9538 25454 9550 25506
rect 9602 25454 9614 25506
rect 15250 25454 15262 25506
rect 15314 25454 15326 25506
rect 18734 25442 18786 25454
rect 18846 25506 18898 25518
rect 18846 25442 18898 25454
rect 20750 25506 20802 25518
rect 22766 25506 22818 25518
rect 21410 25454 21422 25506
rect 21474 25454 21486 25506
rect 22082 25454 22094 25506
rect 22146 25454 22158 25506
rect 20750 25442 20802 25454
rect 22766 25442 22818 25454
rect 23102 25506 23154 25518
rect 23102 25442 23154 25454
rect 23774 25506 23826 25518
rect 23774 25442 23826 25454
rect 23998 25506 24050 25518
rect 23998 25442 24050 25454
rect 27918 25506 27970 25518
rect 27918 25442 27970 25454
rect 28254 25506 28306 25518
rect 41918 25506 41970 25518
rect 44830 25506 44882 25518
rect 29922 25454 29934 25506
rect 29986 25454 29998 25506
rect 34178 25454 34190 25506
rect 34242 25454 34254 25506
rect 36418 25454 36430 25506
rect 36482 25454 36494 25506
rect 36978 25454 36990 25506
rect 37042 25454 37054 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 42354 25454 42366 25506
rect 42418 25454 42430 25506
rect 43138 25454 43150 25506
rect 43202 25454 43214 25506
rect 28254 25442 28306 25454
rect 41918 25442 41970 25454
rect 44830 25442 44882 25454
rect 45278 25506 45330 25518
rect 45278 25442 45330 25454
rect 45502 25506 45554 25518
rect 45502 25442 45554 25454
rect 47518 25506 47570 25518
rect 47518 25442 47570 25454
rect 47966 25506 48018 25518
rect 47966 25442 48018 25454
rect 48078 25506 48130 25518
rect 48078 25442 48130 25454
rect 48862 25506 48914 25518
rect 48862 25442 48914 25454
rect 49982 25506 50034 25518
rect 49982 25442 50034 25454
rect 50430 25506 50482 25518
rect 50430 25442 50482 25454
rect 50878 25506 50930 25518
rect 50878 25442 50930 25454
rect 51102 25506 51154 25518
rect 52670 25506 52722 25518
rect 52098 25454 52110 25506
rect 52162 25454 52174 25506
rect 53554 25454 53566 25506
rect 53618 25454 53630 25506
rect 51102 25442 51154 25454
rect 52670 25442 52722 25454
rect 18510 25394 18562 25406
rect 14130 25342 14142 25394
rect 14194 25342 14206 25394
rect 14466 25342 14478 25394
rect 14530 25342 14542 25394
rect 18510 25330 18562 25342
rect 19742 25394 19794 25406
rect 19742 25330 19794 25342
rect 20190 25394 20242 25406
rect 20190 25330 20242 25342
rect 22542 25394 22594 25406
rect 22542 25330 22594 25342
rect 22990 25394 23042 25406
rect 37326 25394 37378 25406
rect 46398 25394 46450 25406
rect 33954 25342 33966 25394
rect 34018 25342 34030 25394
rect 34850 25342 34862 25394
rect 34914 25342 34926 25394
rect 41010 25342 41022 25394
rect 41074 25342 41086 25394
rect 41682 25342 41694 25394
rect 41746 25342 41758 25394
rect 51426 25342 51438 25394
rect 51490 25342 51502 25394
rect 51986 25342 51998 25394
rect 52050 25342 52062 25394
rect 22990 25330 23042 25342
rect 37326 25330 37378 25342
rect 46398 25330 46450 25342
rect 12798 25282 12850 25294
rect 12798 25218 12850 25230
rect 21534 25282 21586 25294
rect 21534 25218 21586 25230
rect 24894 25282 24946 25294
rect 29598 25282 29650 25294
rect 27570 25230 27582 25282
rect 27634 25230 27646 25282
rect 28578 25230 28590 25282
rect 28642 25230 28654 25282
rect 24894 25218 24946 25230
rect 29598 25218 29650 25230
rect 37214 25282 37266 25294
rect 45390 25282 45442 25294
rect 41906 25230 41918 25282
rect 41970 25230 41982 25282
rect 37214 25218 37266 25230
rect 45390 25218 45442 25230
rect 47294 25282 47346 25294
rect 47294 25218 47346 25230
rect 48638 25282 48690 25294
rect 48638 25218 48690 25230
rect 48974 25282 49026 25294
rect 48974 25218 49026 25230
rect 49086 25282 49138 25294
rect 49086 25218 49138 25230
rect 50094 25282 50146 25294
rect 50094 25218 50146 25230
rect 50766 25282 50818 25294
rect 50766 25218 50818 25230
rect 54238 25282 54290 25294
rect 54238 25218 54290 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 6078 24946 6130 24958
rect 6078 24882 6130 24894
rect 7758 24946 7810 24958
rect 7758 24882 7810 24894
rect 9662 24946 9714 24958
rect 18398 24946 18450 24958
rect 11666 24894 11678 24946
rect 11730 24894 11742 24946
rect 9662 24882 9714 24894
rect 18398 24882 18450 24894
rect 26238 24946 26290 24958
rect 26238 24882 26290 24894
rect 41022 24946 41074 24958
rect 41022 24882 41074 24894
rect 41134 24946 41186 24958
rect 53678 24946 53730 24958
rect 44706 24894 44718 24946
rect 44770 24894 44782 24946
rect 41134 24882 41186 24894
rect 53678 24882 53730 24894
rect 54126 24946 54178 24958
rect 54126 24882 54178 24894
rect 2718 24834 2770 24846
rect 2718 24770 2770 24782
rect 3390 24834 3442 24846
rect 14030 24834 14082 24846
rect 7186 24782 7198 24834
rect 7250 24782 7262 24834
rect 8866 24782 8878 24834
rect 8930 24782 8942 24834
rect 3390 24770 3442 24782
rect 14030 24770 14082 24782
rect 18846 24834 18898 24846
rect 24558 24834 24610 24846
rect 46622 24834 46674 24846
rect 22194 24782 22206 24834
rect 22258 24782 22270 24834
rect 28690 24782 28702 24834
rect 28754 24782 28766 24834
rect 30146 24782 30158 24834
rect 30210 24782 30222 24834
rect 37874 24782 37886 24834
rect 37938 24782 37950 24834
rect 39106 24782 39118 24834
rect 39170 24782 39182 24834
rect 45714 24782 45726 24834
rect 45778 24782 45790 24834
rect 18846 24770 18898 24782
rect 24558 24770 24610 24782
rect 46622 24770 46674 24782
rect 3726 24722 3778 24734
rect 2930 24670 2942 24722
rect 2994 24670 3006 24722
rect 3726 24658 3778 24670
rect 6414 24722 6466 24734
rect 8094 24722 8146 24734
rect 12014 24722 12066 24734
rect 17950 24722 18002 24734
rect 24446 24722 24498 24734
rect 6850 24670 6862 24722
rect 6914 24670 6926 24722
rect 8642 24670 8654 24722
rect 8706 24670 8718 24722
rect 13794 24670 13806 24722
rect 13858 24670 13870 24722
rect 19842 24670 19854 24722
rect 19906 24670 19918 24722
rect 22754 24670 22766 24722
rect 22818 24670 22830 24722
rect 23426 24670 23438 24722
rect 23490 24670 23502 24722
rect 6414 24658 6466 24670
rect 8094 24658 8146 24670
rect 12014 24658 12066 24670
rect 17950 24658 18002 24670
rect 24446 24658 24498 24670
rect 24782 24722 24834 24734
rect 40910 24722 40962 24734
rect 46846 24722 46898 24734
rect 25666 24670 25678 24722
rect 25730 24670 25742 24722
rect 29362 24670 29374 24722
rect 29426 24670 29438 24722
rect 29922 24670 29934 24722
rect 29986 24670 29998 24722
rect 36306 24670 36318 24722
rect 36370 24670 36382 24722
rect 37202 24670 37214 24722
rect 37266 24670 37278 24722
rect 38546 24670 38558 24722
rect 38610 24670 38622 24722
rect 41458 24670 41470 24722
rect 41522 24670 41534 24722
rect 42242 24670 42254 24722
rect 42306 24670 42318 24722
rect 42802 24670 42814 24722
rect 42866 24670 42878 24722
rect 44930 24670 44942 24722
rect 44994 24670 45006 24722
rect 24782 24658 24834 24670
rect 40910 24658 40962 24670
rect 46846 24658 46898 24670
rect 47294 24722 47346 24734
rect 47294 24658 47346 24670
rect 47518 24722 47570 24734
rect 47518 24658 47570 24670
rect 47742 24722 47794 24734
rect 48738 24670 48750 24722
rect 48802 24670 48814 24722
rect 49074 24670 49086 24722
rect 49138 24670 49150 24722
rect 50642 24670 50654 24722
rect 50706 24670 50718 24722
rect 52098 24670 52110 24722
rect 52162 24670 52174 24722
rect 47742 24658 47794 24670
rect 12462 24610 12514 24622
rect 12462 24546 12514 24558
rect 13134 24610 13186 24622
rect 13134 24546 13186 24558
rect 14926 24610 14978 24622
rect 20078 24610 20130 24622
rect 25230 24610 25282 24622
rect 33966 24610 34018 24622
rect 40014 24610 40066 24622
rect 17490 24558 17502 24610
rect 17554 24558 17566 24610
rect 22418 24558 22430 24610
rect 22482 24558 22494 24610
rect 26562 24558 26574 24610
rect 26626 24558 26638 24610
rect 35746 24558 35758 24610
rect 35810 24558 35822 24610
rect 14926 24546 14978 24558
rect 20078 24546 20130 24558
rect 25230 24546 25282 24558
rect 33966 24546 34018 24558
rect 40014 24546 40066 24558
rect 41918 24610 41970 24622
rect 41918 24546 41970 24558
rect 47070 24610 47122 24622
rect 48850 24558 48862 24610
rect 48914 24558 48926 24610
rect 52210 24558 52222 24610
rect 52274 24558 52286 24610
rect 47070 24546 47122 24558
rect 48066 24446 48078 24498
rect 48130 24446 48142 24498
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 45390 24162 45442 24174
rect 12338 24110 12350 24162
rect 12402 24110 12414 24162
rect 25554 24110 25566 24162
rect 25618 24110 25630 24162
rect 41794 24110 41806 24162
rect 41858 24110 41870 24162
rect 43250 24110 43262 24162
rect 43314 24110 43326 24162
rect 50306 24110 50318 24162
rect 50370 24110 50382 24162
rect 45390 24098 45442 24110
rect 5742 24050 5794 24062
rect 2930 23998 2942 24050
rect 2994 23998 3006 24050
rect 5058 23998 5070 24050
rect 5122 23998 5134 24050
rect 5742 23986 5794 23998
rect 7310 24050 7362 24062
rect 7310 23986 7362 23998
rect 9550 24050 9602 24062
rect 9550 23986 9602 23998
rect 12910 24050 12962 24062
rect 47182 24050 47234 24062
rect 14242 23998 14254 24050
rect 14306 23998 14318 24050
rect 16370 23998 16382 24050
rect 16434 23998 16446 24050
rect 18722 23998 18734 24050
rect 18786 23998 18798 24050
rect 24322 23998 24334 24050
rect 24386 23998 24398 24050
rect 33170 23998 33182 24050
rect 33234 23998 33246 24050
rect 36082 23998 36094 24050
rect 36146 23998 36158 24050
rect 42578 23998 42590 24050
rect 42642 23998 42654 24050
rect 46274 23998 46286 24050
rect 46338 23998 46350 24050
rect 12910 23986 12962 23998
rect 47182 23986 47234 23998
rect 47630 24050 47682 24062
rect 54350 24050 54402 24062
rect 48738 23998 48750 24050
rect 48802 23998 48814 24050
rect 47630 23986 47682 23998
rect 54350 23986 54402 23998
rect 7646 23938 7698 23950
rect 2258 23886 2270 23938
rect 2322 23886 2334 23938
rect 7646 23874 7698 23886
rect 7982 23938 8034 23950
rect 7982 23874 8034 23886
rect 12686 23938 12738 23950
rect 24894 23938 24946 23950
rect 13458 23886 13470 23938
rect 13522 23886 13534 23938
rect 18386 23886 18398 23938
rect 18450 23886 18462 23938
rect 20738 23886 20750 23938
rect 20802 23886 20814 23938
rect 22978 23886 22990 23938
rect 23042 23886 23054 23938
rect 23202 23886 23214 23938
rect 23266 23886 23278 23938
rect 12686 23874 12738 23886
rect 24894 23874 24946 23886
rect 25342 23938 25394 23950
rect 43822 23938 43874 23950
rect 26114 23886 26126 23938
rect 26178 23886 26190 23938
rect 29250 23886 29262 23938
rect 29314 23886 29326 23938
rect 34290 23886 34302 23938
rect 34354 23886 34366 23938
rect 34626 23886 34638 23938
rect 34690 23886 34702 23938
rect 35186 23886 35198 23938
rect 35250 23886 35262 23938
rect 35634 23886 35646 23938
rect 35698 23886 35710 23938
rect 36978 23886 36990 23938
rect 37042 23886 37054 23938
rect 40786 23886 40798 23938
rect 40850 23886 40862 23938
rect 41346 23886 41358 23938
rect 41410 23886 41422 23938
rect 41794 23886 41806 23938
rect 41858 23886 41870 23938
rect 42242 23886 42254 23938
rect 42306 23886 42318 23938
rect 25342 23874 25394 23886
rect 43822 23874 43874 23886
rect 43934 23938 43986 23950
rect 43934 23874 43986 23886
rect 44942 23938 44994 23950
rect 44942 23874 44994 23886
rect 45166 23938 45218 23950
rect 45166 23874 45218 23886
rect 45950 23938 46002 23950
rect 47518 23938 47570 23950
rect 51662 23938 51714 23950
rect 46498 23886 46510 23938
rect 46562 23886 46574 23938
rect 48290 23886 48302 23938
rect 48354 23886 48366 23938
rect 49074 23886 49086 23938
rect 49138 23886 49150 23938
rect 49522 23886 49534 23938
rect 49586 23886 49598 23938
rect 51090 23886 51102 23938
rect 51154 23886 51166 23938
rect 45950 23874 46002 23886
rect 47518 23874 47570 23886
rect 51662 23874 51714 23886
rect 53342 23938 53394 23950
rect 53890 23886 53902 23938
rect 53954 23886 53966 23938
rect 53342 23874 53394 23886
rect 43710 23826 43762 23838
rect 49758 23826 49810 23838
rect 18050 23774 18062 23826
rect 18114 23774 18126 23826
rect 19058 23774 19070 23826
rect 19122 23774 19134 23826
rect 22754 23774 22766 23826
rect 22818 23774 22830 23826
rect 23986 23774 23998 23826
rect 24050 23774 24062 23826
rect 36194 23774 36206 23826
rect 36258 23774 36270 23826
rect 37090 23774 37102 23826
rect 37154 23774 37166 23826
rect 40674 23774 40686 23826
rect 40738 23774 40750 23826
rect 45602 23774 45614 23826
rect 45666 23774 45678 23826
rect 49186 23774 49198 23826
rect 49250 23774 49262 23826
rect 43710 23762 43762 23774
rect 49758 23762 49810 23774
rect 49870 23826 49922 23838
rect 49870 23762 49922 23774
rect 51774 23826 51826 23838
rect 51774 23762 51826 23774
rect 52670 23826 52722 23838
rect 52670 23762 52722 23774
rect 52894 23826 52946 23838
rect 52894 23762 52946 23774
rect 53566 23826 53618 23838
rect 53566 23762 53618 23774
rect 7422 23714 7474 23726
rect 7422 23650 7474 23662
rect 7870 23714 7922 23726
rect 7870 23650 7922 23662
rect 8542 23714 8594 23726
rect 8542 23650 8594 23662
rect 9662 23714 9714 23726
rect 9662 23650 9714 23662
rect 26350 23714 26402 23726
rect 26350 23650 26402 23662
rect 27918 23714 27970 23726
rect 27918 23650 27970 23662
rect 28366 23714 28418 23726
rect 28366 23650 28418 23662
rect 29486 23714 29538 23726
rect 53006 23714 53058 23726
rect 37202 23662 37214 23714
rect 37266 23662 37278 23714
rect 45490 23662 45502 23714
rect 45554 23662 45566 23714
rect 29486 23650 29538 23662
rect 53006 23650 53058 23662
rect 53678 23714 53730 23726
rect 53678 23650 53730 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 5406 23378 5458 23390
rect 5406 23314 5458 23326
rect 13582 23378 13634 23390
rect 13582 23314 13634 23326
rect 21870 23378 21922 23390
rect 21870 23314 21922 23326
rect 23438 23378 23490 23390
rect 23438 23314 23490 23326
rect 33630 23378 33682 23390
rect 33630 23314 33682 23326
rect 34974 23378 35026 23390
rect 34974 23314 35026 23326
rect 38446 23378 38498 23390
rect 38446 23314 38498 23326
rect 39006 23378 39058 23390
rect 39006 23314 39058 23326
rect 41358 23378 41410 23390
rect 41358 23314 41410 23326
rect 42590 23378 42642 23390
rect 42590 23314 42642 23326
rect 47406 23378 47458 23390
rect 47406 23314 47458 23326
rect 48190 23378 48242 23390
rect 48190 23314 48242 23326
rect 7534 23266 7586 23278
rect 2594 23214 2606 23266
rect 2658 23214 2670 23266
rect 6402 23214 6414 23266
rect 6466 23214 6478 23266
rect 7534 23202 7586 23214
rect 7646 23266 7698 23278
rect 7646 23202 7698 23214
rect 8206 23266 8258 23278
rect 16382 23266 16434 23278
rect 17502 23266 17554 23278
rect 20974 23266 21026 23278
rect 15250 23214 15262 23266
rect 15314 23214 15326 23266
rect 16706 23214 16718 23266
rect 16770 23214 16782 23266
rect 19842 23214 19854 23266
rect 19906 23214 19918 23266
rect 8206 23202 8258 23214
rect 16382 23202 16434 23214
rect 17502 23202 17554 23214
rect 20974 23202 21026 23214
rect 23886 23266 23938 23278
rect 33854 23266 33906 23278
rect 27346 23214 27358 23266
rect 27410 23214 27422 23266
rect 30706 23214 30718 23266
rect 30770 23214 30782 23266
rect 23886 23202 23938 23214
rect 33854 23202 33906 23214
rect 38558 23266 38610 23278
rect 45726 23266 45778 23278
rect 42018 23214 42030 23266
rect 42082 23214 42094 23266
rect 42914 23214 42926 23266
rect 42978 23214 42990 23266
rect 44706 23214 44718 23266
rect 44770 23214 44782 23266
rect 50418 23214 50430 23266
rect 50482 23214 50494 23266
rect 38558 23202 38610 23214
rect 45726 23202 45778 23214
rect 7310 23154 7362 23166
rect 13694 23154 13746 23166
rect 1922 23102 1934 23154
rect 1986 23102 1998 23154
rect 6514 23102 6526 23154
rect 6578 23102 6590 23154
rect 9650 23102 9662 23154
rect 9714 23102 9726 23154
rect 7310 23090 7362 23102
rect 13694 23090 13746 23102
rect 14478 23154 14530 23166
rect 18062 23154 18114 23166
rect 15138 23102 15150 23154
rect 15202 23102 15214 23154
rect 14478 23090 14530 23102
rect 18062 23090 18114 23102
rect 20526 23154 20578 23166
rect 20526 23090 20578 23102
rect 23326 23154 23378 23166
rect 23326 23090 23378 23102
rect 23662 23154 23714 23166
rect 34078 23154 34130 23166
rect 28130 23102 28142 23154
rect 28194 23102 28206 23154
rect 31378 23102 31390 23154
rect 31442 23102 31454 23154
rect 23662 23090 23714 23102
rect 34078 23090 34130 23102
rect 34526 23154 34578 23166
rect 39902 23154 39954 23166
rect 37426 23102 37438 23154
rect 37490 23102 37502 23154
rect 39778 23102 39790 23154
rect 39842 23102 39854 23154
rect 34526 23090 34578 23102
rect 39902 23090 39954 23102
rect 41694 23154 41746 23166
rect 41694 23090 41746 23102
rect 41806 23154 41858 23166
rect 41806 23090 41858 23102
rect 42366 23154 42418 23166
rect 45950 23154 46002 23166
rect 43698 23102 43710 23154
rect 43762 23102 43774 23154
rect 45154 23102 45166 23154
rect 45218 23102 45230 23154
rect 42366 23090 42418 23102
rect 45950 23090 46002 23102
rect 46398 23154 46450 23166
rect 46398 23090 46450 23102
rect 47182 23154 47234 23166
rect 49646 23154 49698 23166
rect 47730 23102 47742 23154
rect 47794 23102 47806 23154
rect 49298 23102 49310 23154
rect 49362 23102 49374 23154
rect 47182 23090 47234 23102
rect 49646 23090 49698 23102
rect 50094 23154 50146 23166
rect 50866 23102 50878 23154
rect 50930 23102 50942 23154
rect 50094 23090 50146 23102
rect 8766 23042 8818 23054
rect 13134 23042 13186 23054
rect 4722 22990 4734 23042
rect 4786 22990 4798 23042
rect 10322 22990 10334 23042
rect 10386 22990 10398 23042
rect 12450 22990 12462 23042
rect 12514 22990 12526 23042
rect 8766 22978 8818 22990
rect 13134 22978 13186 22990
rect 15822 23042 15874 23054
rect 22206 23042 22258 23054
rect 19618 22990 19630 23042
rect 19682 22990 19694 23042
rect 15822 22978 15874 22990
rect 22206 22978 22258 22990
rect 24110 23042 24162 23054
rect 34302 23042 34354 23054
rect 46174 23042 46226 23054
rect 25218 22990 25230 23042
rect 25282 22990 25294 23042
rect 28578 22990 28590 23042
rect 28642 22990 28654 23042
rect 35074 22990 35086 23042
rect 35138 22990 35150 23042
rect 36306 22990 36318 23042
rect 36370 22990 36382 23042
rect 39554 22990 39566 23042
rect 39618 22990 39630 23042
rect 24110 22978 24162 22990
rect 34302 22978 34354 22990
rect 46174 22978 46226 22990
rect 46734 23042 46786 23054
rect 46734 22978 46786 22990
rect 47294 23042 47346 23054
rect 47294 22978 47346 22990
rect 48750 23042 48802 23054
rect 51538 22990 51550 23042
rect 51602 22990 51614 23042
rect 53666 22990 53678 23042
rect 53730 22990 53742 23042
rect 48750 22978 48802 22990
rect 5742 22930 5794 22942
rect 5742 22866 5794 22878
rect 7982 22930 8034 22942
rect 7982 22866 8034 22878
rect 8318 22930 8370 22942
rect 8318 22866 8370 22878
rect 13582 22930 13634 22942
rect 13582 22866 13634 22878
rect 14142 22930 14194 22942
rect 14142 22866 14194 22878
rect 18286 22930 18338 22942
rect 24446 22930 24498 22942
rect 19730 22878 19742 22930
rect 19794 22878 19806 22930
rect 18286 22866 18338 22878
rect 24446 22866 24498 22878
rect 34750 22930 34802 22942
rect 34750 22866 34802 22878
rect 38334 22930 38386 22942
rect 38334 22866 38386 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 6078 22594 6130 22606
rect 6078 22530 6130 22542
rect 7310 22594 7362 22606
rect 7310 22530 7362 22542
rect 11790 22594 11842 22606
rect 11790 22530 11842 22542
rect 14030 22594 14082 22606
rect 14030 22530 14082 22542
rect 14366 22594 14418 22606
rect 14366 22530 14418 22542
rect 20302 22594 20354 22606
rect 20302 22530 20354 22542
rect 20638 22594 20690 22606
rect 20638 22530 20690 22542
rect 21758 22594 21810 22606
rect 21758 22530 21810 22542
rect 22542 22594 22594 22606
rect 22542 22530 22594 22542
rect 26574 22594 26626 22606
rect 26574 22530 26626 22542
rect 26910 22594 26962 22606
rect 26910 22530 26962 22542
rect 29262 22594 29314 22606
rect 29262 22530 29314 22542
rect 46622 22594 46674 22606
rect 46622 22530 46674 22542
rect 46958 22594 47010 22606
rect 46958 22530 47010 22542
rect 47518 22594 47570 22606
rect 52670 22594 52722 22606
rect 51426 22542 51438 22594
rect 51490 22542 51502 22594
rect 47518 22530 47570 22542
rect 52670 22530 52722 22542
rect 5070 22482 5122 22494
rect 5070 22418 5122 22430
rect 13694 22482 13746 22494
rect 13694 22418 13746 22430
rect 18510 22482 18562 22494
rect 18510 22418 18562 22430
rect 21534 22482 21586 22494
rect 21534 22418 21586 22430
rect 25678 22482 25730 22494
rect 25678 22418 25730 22430
rect 28478 22482 28530 22494
rect 28478 22418 28530 22430
rect 29598 22482 29650 22494
rect 36206 22482 36258 22494
rect 42590 22482 42642 22494
rect 34066 22430 34078 22482
rect 34130 22430 34142 22482
rect 37090 22430 37102 22482
rect 37154 22430 37166 22482
rect 40338 22430 40350 22482
rect 40402 22430 40414 22482
rect 29598 22418 29650 22430
rect 36206 22418 36258 22430
rect 42590 22418 42642 22430
rect 44270 22482 44322 22494
rect 44270 22418 44322 22430
rect 44830 22482 44882 22494
rect 47182 22482 47234 22494
rect 45714 22430 45726 22482
rect 45778 22430 45790 22482
rect 44830 22418 44882 22430
rect 47182 22418 47234 22430
rect 47854 22482 47906 22494
rect 47854 22418 47906 22430
rect 48414 22482 48466 22494
rect 48414 22418 48466 22430
rect 49646 22482 49698 22494
rect 49646 22418 49698 22430
rect 50430 22482 50482 22494
rect 50430 22418 50482 22430
rect 50878 22482 50930 22494
rect 50878 22418 50930 22430
rect 5742 22370 5794 22382
rect 10670 22370 10722 22382
rect 6514 22318 6526 22370
rect 6578 22318 6590 22370
rect 5742 22306 5794 22318
rect 10670 22306 10722 22318
rect 11454 22370 11506 22382
rect 18846 22370 18898 22382
rect 12562 22318 12574 22370
rect 12626 22318 12638 22370
rect 17938 22318 17950 22370
rect 18002 22318 18014 22370
rect 11454 22306 11506 22318
rect 18846 22306 18898 22318
rect 19182 22370 19234 22382
rect 19182 22306 19234 22318
rect 20526 22370 20578 22382
rect 20526 22306 20578 22318
rect 22430 22370 22482 22382
rect 22430 22306 22482 22318
rect 22878 22370 22930 22382
rect 22878 22306 22930 22318
rect 23102 22370 23154 22382
rect 23102 22306 23154 22318
rect 23774 22370 23826 22382
rect 23774 22306 23826 22318
rect 24222 22370 24274 22382
rect 35982 22370 36034 22382
rect 43486 22370 43538 22382
rect 46062 22370 46114 22382
rect 27682 22318 27694 22370
rect 27746 22318 27758 22370
rect 31154 22318 31166 22370
rect 31218 22318 31230 22370
rect 34626 22318 34638 22370
rect 34690 22318 34702 22370
rect 35522 22318 35534 22370
rect 35586 22318 35598 22370
rect 35746 22318 35758 22370
rect 35810 22318 35822 22370
rect 37314 22318 37326 22370
rect 37378 22318 37390 22370
rect 37986 22318 37998 22370
rect 38050 22318 38062 22370
rect 38210 22318 38222 22370
rect 38274 22318 38286 22370
rect 40562 22318 40574 22370
rect 40626 22318 40638 22370
rect 40786 22318 40798 22370
rect 40850 22318 40862 22370
rect 43698 22318 43710 22370
rect 43762 22318 43774 22370
rect 45266 22318 45278 22370
rect 45330 22318 45342 22370
rect 24222 22306 24274 22318
rect 35982 22306 36034 22318
rect 43486 22306 43538 22318
rect 46062 22306 46114 22318
rect 48862 22370 48914 22382
rect 52782 22370 52834 22382
rect 51202 22318 51214 22370
rect 51266 22318 51278 22370
rect 51762 22318 51774 22370
rect 51826 22318 51838 22370
rect 48862 22306 48914 22318
rect 52782 22306 52834 22318
rect 3614 22258 3666 22270
rect 10334 22258 10386 22270
rect 16718 22258 16770 22270
rect 6850 22206 6862 22258
rect 6914 22206 6926 22258
rect 12450 22206 12462 22258
rect 12514 22206 12526 22258
rect 14578 22206 14590 22258
rect 14642 22206 14654 22258
rect 14914 22206 14926 22258
rect 14978 22206 14990 22258
rect 3614 22194 3666 22206
rect 10334 22194 10386 22206
rect 16718 22194 16770 22206
rect 17166 22258 17218 22270
rect 19070 22258 19122 22270
rect 23326 22258 23378 22270
rect 18050 22206 18062 22258
rect 18114 22206 18126 22258
rect 18386 22206 18398 22258
rect 18450 22206 18462 22258
rect 19730 22206 19742 22258
rect 19794 22206 19806 22258
rect 17166 22194 17218 22206
rect 19070 22194 19122 22206
rect 23326 22194 23378 22206
rect 24894 22258 24946 22270
rect 24894 22194 24946 22206
rect 25230 22258 25282 22270
rect 36430 22258 36482 22270
rect 43374 22258 43426 22270
rect 27458 22206 27470 22258
rect 27522 22206 27534 22258
rect 29810 22206 29822 22258
rect 29874 22206 29886 22258
rect 30370 22206 30382 22258
rect 30434 22206 30446 22258
rect 31938 22206 31950 22258
rect 32002 22206 32014 22258
rect 40338 22206 40350 22258
rect 40402 22206 40414 22258
rect 41570 22206 41582 22258
rect 41634 22206 41646 22258
rect 25230 22194 25282 22206
rect 36430 22194 36482 22206
rect 43374 22194 43426 22206
rect 45838 22258 45890 22270
rect 45838 22194 45890 22206
rect 47630 22258 47682 22270
rect 47630 22194 47682 22206
rect 48302 22258 48354 22270
rect 48302 22194 48354 22206
rect 48526 22258 48578 22270
rect 51998 22258 52050 22270
rect 49186 22206 49198 22258
rect 49250 22206 49262 22258
rect 48526 22194 48578 22206
rect 51998 22194 52050 22206
rect 3278 22146 3330 22158
rect 3278 22082 3330 22094
rect 7422 22146 7474 22158
rect 7422 22082 7474 22094
rect 7534 22146 7586 22158
rect 16046 22146 16098 22158
rect 17502 22146 17554 22158
rect 22990 22146 23042 22158
rect 15698 22094 15710 22146
rect 15762 22094 15774 22146
rect 16370 22094 16382 22146
rect 16434 22094 16446 22146
rect 22082 22094 22094 22146
rect 22146 22094 22158 22146
rect 7534 22082 7586 22094
rect 16046 22082 16098 22094
rect 17502 22082 17554 22094
rect 22990 22082 23042 22094
rect 23886 22146 23938 22158
rect 23886 22082 23938 22094
rect 25006 22146 25058 22158
rect 25006 22082 25058 22094
rect 25790 22146 25842 22158
rect 25790 22082 25842 22094
rect 28590 22146 28642 22158
rect 35198 22146 35250 22158
rect 34402 22094 34414 22146
rect 34466 22094 34478 22146
rect 28590 22082 28642 22094
rect 35198 22082 35250 22094
rect 36542 22146 36594 22158
rect 42914 22094 42926 22146
rect 42978 22094 42990 22146
rect 51650 22094 51662 22146
rect 51714 22094 51726 22146
rect 36542 22082 36594 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 7758 21810 7810 21822
rect 7758 21746 7810 21758
rect 8878 21810 8930 21822
rect 8878 21746 8930 21758
rect 14590 21810 14642 21822
rect 14590 21746 14642 21758
rect 20302 21810 20354 21822
rect 20302 21746 20354 21758
rect 20750 21810 20802 21822
rect 20750 21746 20802 21758
rect 21422 21810 21474 21822
rect 21422 21746 21474 21758
rect 22654 21810 22706 21822
rect 22654 21746 22706 21758
rect 27022 21810 27074 21822
rect 27022 21746 27074 21758
rect 27694 21810 27746 21822
rect 27694 21746 27746 21758
rect 28478 21810 28530 21822
rect 28478 21746 28530 21758
rect 30270 21810 30322 21822
rect 30270 21746 30322 21758
rect 32062 21810 32114 21822
rect 32062 21746 32114 21758
rect 34974 21810 35026 21822
rect 34974 21746 35026 21758
rect 35198 21810 35250 21822
rect 35198 21746 35250 21758
rect 35534 21810 35586 21822
rect 35534 21746 35586 21758
rect 35758 21810 35810 21822
rect 45166 21810 45218 21822
rect 39218 21758 39230 21810
rect 39282 21758 39294 21810
rect 35758 21746 35810 21758
rect 45166 21746 45218 21758
rect 46846 21810 46898 21822
rect 47854 21810 47906 21822
rect 47394 21758 47406 21810
rect 47458 21758 47470 21810
rect 46846 21746 46898 21758
rect 47854 21746 47906 21758
rect 6974 21698 7026 21710
rect 3042 21646 3054 21698
rect 3106 21646 3118 21698
rect 6974 21634 7026 21646
rect 8094 21698 8146 21710
rect 8094 21634 8146 21646
rect 10558 21698 10610 21710
rect 10558 21634 10610 21646
rect 10894 21698 10946 21710
rect 10894 21634 10946 21646
rect 11118 21698 11170 21710
rect 13806 21698 13858 21710
rect 11666 21646 11678 21698
rect 11730 21646 11742 21698
rect 12114 21646 12126 21698
rect 12178 21646 12190 21698
rect 11118 21634 11170 21646
rect 13806 21634 13858 21646
rect 15934 21698 15986 21710
rect 20190 21698 20242 21710
rect 19058 21646 19070 21698
rect 19122 21646 19134 21698
rect 15934 21634 15986 21646
rect 20190 21634 20242 21646
rect 20862 21698 20914 21710
rect 20862 21634 20914 21646
rect 21646 21698 21698 21710
rect 22990 21698 23042 21710
rect 22306 21646 22318 21698
rect 22370 21646 22382 21698
rect 21646 21634 21698 21646
rect 22990 21634 23042 21646
rect 24558 21698 24610 21710
rect 26238 21698 26290 21710
rect 35310 21698 35362 21710
rect 25554 21646 25566 21698
rect 25618 21646 25630 21698
rect 28018 21646 28030 21698
rect 28082 21646 28094 21698
rect 29810 21646 29822 21698
rect 29874 21646 29886 21698
rect 33730 21646 33742 21698
rect 33794 21646 33806 21698
rect 34066 21646 34078 21698
rect 34130 21646 34142 21698
rect 24558 21634 24610 21646
rect 26238 21634 26290 21646
rect 35310 21634 35362 21646
rect 35870 21698 35922 21710
rect 44382 21698 44434 21710
rect 36978 21646 36990 21698
rect 37042 21646 37054 21698
rect 40338 21646 40350 21698
rect 40402 21646 40414 21698
rect 40898 21646 40910 21698
rect 40962 21646 40974 21698
rect 35870 21634 35922 21646
rect 44382 21634 44434 21646
rect 47966 21698 48018 21710
rect 47966 21634 48018 21646
rect 7422 21586 7474 21598
rect 8542 21586 8594 21598
rect 12350 21586 12402 21598
rect 14254 21586 14306 21598
rect 16718 21586 16770 21598
rect 20526 21586 20578 21598
rect 2258 21534 2270 21586
rect 2322 21534 2334 21586
rect 7186 21534 7198 21586
rect 7250 21534 7262 21586
rect 7746 21534 7758 21586
rect 7810 21534 7822 21586
rect 8306 21534 8318 21586
rect 8370 21534 8382 21586
rect 8642 21534 8654 21586
rect 8706 21534 8718 21586
rect 14018 21534 14030 21586
rect 14082 21534 14094 21586
rect 14354 21534 14366 21586
rect 14418 21534 14430 21586
rect 16146 21534 16158 21586
rect 16210 21534 16222 21586
rect 19170 21534 19182 21586
rect 19234 21534 19246 21586
rect 7422 21522 7474 21534
rect 8542 21522 8594 21534
rect 12350 21522 12402 21534
rect 14254 21522 14306 21534
rect 16718 21522 16770 21534
rect 20526 21522 20578 21534
rect 24334 21586 24386 21598
rect 26574 21586 26626 21598
rect 32398 21586 32450 21598
rect 25218 21534 25230 21586
rect 25282 21534 25294 21586
rect 29586 21534 29598 21586
rect 29650 21534 29662 21586
rect 24334 21522 24386 21534
rect 26574 21522 26626 21534
rect 32398 21522 32450 21534
rect 33182 21586 33234 21598
rect 42926 21586 42978 21598
rect 43934 21586 43986 21598
rect 36306 21534 36318 21586
rect 36370 21534 36382 21586
rect 39778 21534 39790 21586
rect 39842 21534 39854 21586
rect 42130 21534 42142 21586
rect 42194 21534 42206 21586
rect 42466 21534 42478 21586
rect 42530 21534 42542 21586
rect 43138 21534 43150 21586
rect 43202 21534 43214 21586
rect 43698 21534 43710 21586
rect 43762 21534 43774 21586
rect 33182 21522 33234 21534
rect 42926 21522 42978 21534
rect 43934 21522 43986 21534
rect 44494 21586 44546 21598
rect 47630 21586 47682 21598
rect 47170 21534 47182 21586
rect 47234 21534 47246 21586
rect 44494 21522 44546 21534
rect 47630 21522 47682 21534
rect 5630 21474 5682 21486
rect 5170 21422 5182 21474
rect 5234 21422 5246 21474
rect 5630 21410 5682 21422
rect 13246 21474 13298 21486
rect 13246 21410 13298 21422
rect 21534 21474 21586 21486
rect 30830 21474 30882 21486
rect 43038 21474 43090 21486
rect 25890 21422 25902 21474
rect 25954 21422 25966 21474
rect 40226 21422 40238 21474
rect 40290 21422 40302 21474
rect 21534 21410 21586 21422
rect 30830 21410 30882 21422
rect 43038 21410 43090 21422
rect 43374 21474 43426 21486
rect 43374 21410 43426 21422
rect 44158 21474 44210 21486
rect 44158 21410 44210 21422
rect 45278 21474 45330 21486
rect 45278 21410 45330 21422
rect 50878 21474 50930 21486
rect 50878 21410 50930 21422
rect 10782 21362 10834 21374
rect 5394 21310 5406 21362
rect 5458 21359 5470 21362
rect 5730 21359 5742 21362
rect 5458 21313 5742 21359
rect 5458 21310 5470 21313
rect 5730 21310 5742 21313
rect 5794 21310 5806 21362
rect 10782 21298 10834 21310
rect 12686 21362 12738 21374
rect 12686 21298 12738 21310
rect 18174 21362 18226 21374
rect 18174 21298 18226 21310
rect 18510 21362 18562 21374
rect 18510 21298 18562 21310
rect 23102 21362 23154 21374
rect 23102 21298 23154 21310
rect 23998 21362 24050 21374
rect 23998 21298 24050 21310
rect 33518 21362 33570 21374
rect 33518 21298 33570 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 5742 21026 5794 21038
rect 5742 20962 5794 20974
rect 9102 21026 9154 21038
rect 9102 20962 9154 20974
rect 10110 21026 10162 21038
rect 10110 20962 10162 20974
rect 13918 21026 13970 21038
rect 13918 20962 13970 20974
rect 38222 21026 38274 21038
rect 38222 20962 38274 20974
rect 38446 21026 38498 21038
rect 38446 20962 38498 20974
rect 38558 21026 38610 21038
rect 43586 21023 43598 21026
rect 38558 20962 38610 20974
rect 42817 20977 43598 21023
rect 8094 20914 8146 20926
rect 22654 20914 22706 20926
rect 37662 20914 37714 20926
rect 42254 20914 42306 20926
rect 42817 20914 42863 20977
rect 43586 20974 43598 20977
rect 43650 20974 43662 21026
rect 43598 20914 43650 20926
rect 48190 20914 48242 20926
rect 4610 20862 4622 20914
rect 4674 20862 4686 20914
rect 11330 20862 11342 20914
rect 11394 20862 11406 20914
rect 19730 20862 19742 20914
rect 19794 20862 19806 20914
rect 23426 20862 23438 20914
rect 23490 20862 23502 20914
rect 25778 20862 25790 20914
rect 25842 20862 25854 20914
rect 27906 20862 27918 20914
rect 27970 20862 27982 20914
rect 37314 20862 37326 20914
rect 37378 20862 37390 20914
rect 39666 20862 39678 20914
rect 39730 20862 39742 20914
rect 41794 20862 41806 20914
rect 41858 20862 41870 20914
rect 42802 20862 42814 20914
rect 42866 20862 42878 20914
rect 45602 20862 45614 20914
rect 45666 20862 45678 20914
rect 47730 20862 47742 20914
rect 47794 20862 47806 20914
rect 8094 20850 8146 20862
rect 22654 20850 22706 20862
rect 37662 20850 37714 20862
rect 42254 20850 42306 20862
rect 43598 20850 43650 20862
rect 48190 20850 48242 20862
rect 6078 20802 6130 20814
rect 1810 20750 1822 20802
rect 1874 20750 1886 20802
rect 6078 20738 6130 20750
rect 7646 20802 7698 20814
rect 9662 20802 9714 20814
rect 11006 20802 11058 20814
rect 8194 20750 8206 20802
rect 8258 20750 8270 20802
rect 9090 20750 9102 20802
rect 9154 20750 9166 20802
rect 10210 20750 10222 20802
rect 10274 20750 10286 20802
rect 7646 20738 7698 20750
rect 9662 20738 9714 20750
rect 11006 20738 11058 20750
rect 13470 20802 13522 20814
rect 20638 20802 20690 20814
rect 32846 20802 32898 20814
rect 35198 20802 35250 20814
rect 13682 20750 13694 20802
rect 13746 20750 13758 20802
rect 14018 20750 14030 20802
rect 14082 20750 14094 20802
rect 15138 20750 15150 20802
rect 15202 20750 15214 20802
rect 15362 20750 15374 20802
rect 15426 20750 15438 20802
rect 15586 20750 15598 20802
rect 15650 20750 15662 20802
rect 16930 20750 16942 20802
rect 16994 20750 17006 20802
rect 22978 20750 22990 20802
rect 23042 20750 23054 20802
rect 24098 20750 24110 20802
rect 24162 20750 24174 20802
rect 25106 20750 25118 20802
rect 25170 20750 25182 20802
rect 29362 20750 29374 20802
rect 29426 20750 29438 20802
rect 34514 20750 34526 20802
rect 34578 20750 34590 20802
rect 13470 20738 13522 20750
rect 20638 20738 20690 20750
rect 32846 20738 32898 20750
rect 35198 20738 35250 20750
rect 35534 20802 35586 20814
rect 35534 20738 35586 20750
rect 38110 20802 38162 20814
rect 42142 20802 42194 20814
rect 38994 20750 39006 20802
rect 39058 20750 39070 20802
rect 38110 20738 38162 20750
rect 42142 20738 42194 20750
rect 42366 20802 42418 20814
rect 42366 20738 42418 20750
rect 42814 20802 42866 20814
rect 44930 20750 44942 20802
rect 44994 20750 45006 20802
rect 42814 20738 42866 20750
rect 8766 20690 8818 20702
rect 11230 20690 11282 20702
rect 20302 20690 20354 20702
rect 2482 20638 2494 20690
rect 2546 20638 2558 20690
rect 6290 20638 6302 20690
rect 6354 20638 6366 20690
rect 6738 20638 6750 20690
rect 6802 20638 6814 20690
rect 7858 20638 7870 20690
rect 7922 20638 7934 20690
rect 9874 20638 9886 20690
rect 9938 20638 9950 20690
rect 10546 20638 10558 20690
rect 10610 20687 10622 20690
rect 10882 20687 10894 20690
rect 10610 20641 10894 20687
rect 10610 20638 10622 20641
rect 10882 20638 10894 20641
rect 10946 20638 10958 20690
rect 17602 20638 17614 20690
rect 17666 20638 17678 20690
rect 23650 20638 23662 20690
rect 23714 20638 23726 20690
rect 33058 20638 33070 20690
rect 33122 20638 33134 20690
rect 33618 20638 33630 20690
rect 33682 20638 33694 20690
rect 35746 20638 35758 20690
rect 35810 20638 35822 20690
rect 36082 20638 36094 20690
rect 36146 20638 36158 20690
rect 8766 20626 8818 20638
rect 11230 20626 11282 20638
rect 20302 20626 20354 20638
rect 5070 20578 5122 20590
rect 13582 20578 13634 20590
rect 8082 20526 8094 20578
rect 8146 20526 8158 20578
rect 10098 20526 10110 20578
rect 10162 20526 10174 20578
rect 5070 20514 5122 20526
rect 13582 20514 13634 20526
rect 16382 20578 16434 20590
rect 16382 20514 16434 20526
rect 20526 20578 20578 20590
rect 20526 20514 20578 20526
rect 21422 20578 21474 20590
rect 21422 20514 21474 20526
rect 24558 20578 24610 20590
rect 24558 20514 24610 20526
rect 28366 20578 28418 20590
rect 28366 20514 28418 20526
rect 29150 20578 29202 20590
rect 29150 20514 29202 20526
rect 32510 20578 32562 20590
rect 32510 20514 32562 20526
rect 34750 20578 34802 20590
rect 34750 20514 34802 20526
rect 43262 20578 43314 20590
rect 43262 20514 43314 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 2494 20242 2546 20254
rect 17502 20242 17554 20254
rect 10994 20190 11006 20242
rect 11058 20190 11070 20242
rect 15922 20190 15934 20242
rect 15986 20190 15998 20242
rect 2494 20178 2546 20190
rect 17502 20178 17554 20190
rect 22206 20242 22258 20254
rect 22206 20178 22258 20190
rect 22766 20242 22818 20254
rect 22766 20178 22818 20190
rect 26798 20242 26850 20254
rect 26798 20178 26850 20190
rect 39118 20242 39170 20254
rect 39118 20178 39170 20190
rect 41246 20242 41298 20254
rect 41246 20178 41298 20190
rect 48190 20242 48242 20254
rect 48190 20178 48242 20190
rect 7086 20130 7138 20142
rect 5954 20078 5966 20130
rect 6018 20078 6030 20130
rect 7086 20066 7138 20078
rect 7310 20130 7362 20142
rect 7310 20066 7362 20078
rect 7982 20130 8034 20142
rect 7982 20066 8034 20078
rect 13806 20130 13858 20142
rect 13806 20066 13858 20078
rect 17838 20130 17890 20142
rect 21422 20130 21474 20142
rect 19282 20078 19294 20130
rect 19346 20078 19358 20130
rect 17838 20066 17890 20078
rect 21422 20066 21474 20078
rect 21534 20130 21586 20142
rect 21534 20066 21586 20078
rect 21646 20130 21698 20142
rect 21646 20066 21698 20078
rect 22094 20130 22146 20142
rect 22094 20066 22146 20078
rect 22430 20130 22482 20142
rect 24558 20130 24610 20142
rect 32062 20130 32114 20142
rect 24098 20078 24110 20130
rect 24162 20078 24174 20130
rect 25554 20078 25566 20130
rect 25618 20078 25630 20130
rect 27682 20078 27694 20130
rect 27746 20078 27758 20130
rect 29138 20078 29150 20130
rect 29202 20078 29214 20130
rect 22430 20066 22482 20078
rect 24558 20066 24610 20078
rect 32062 20066 32114 20078
rect 32398 20130 32450 20142
rect 40350 20130 40402 20142
rect 35298 20078 35310 20130
rect 35362 20078 35374 20130
rect 32398 20066 32450 20078
rect 40350 20066 40402 20078
rect 41134 20130 41186 20142
rect 45602 20078 45614 20130
rect 45666 20078 45678 20130
rect 41134 20066 41186 20078
rect 2830 20018 2882 20030
rect 2830 19954 2882 19966
rect 5070 20018 5122 20030
rect 5070 19954 5122 19966
rect 5406 20018 5458 20030
rect 10558 20018 10610 20030
rect 11006 20018 11058 20030
rect 14926 20018 14978 20030
rect 24670 20018 24722 20030
rect 27134 20018 27186 20030
rect 39790 20018 39842 20030
rect 6178 19966 6190 20018
rect 6242 19966 6254 20018
rect 10770 19966 10782 20018
rect 10834 19966 10846 20018
rect 11106 19966 11118 20018
rect 11170 19966 11182 20018
rect 14130 19966 14142 20018
rect 14194 19966 14206 20018
rect 14690 19966 14702 20018
rect 14754 19966 14766 20018
rect 15810 19966 15822 20018
rect 15874 19966 15886 20018
rect 16034 19966 16046 20018
rect 16098 19966 16110 20018
rect 19170 19966 19182 20018
rect 19234 19966 19246 20018
rect 23090 19966 23102 20018
rect 23154 19966 23166 20018
rect 24210 19966 24222 20018
rect 24274 19966 24286 20018
rect 25218 19966 25230 20018
rect 25282 19966 25294 20018
rect 27906 19966 27918 20018
rect 27970 19966 27982 20018
rect 28354 19966 28366 20018
rect 28418 19966 28430 20018
rect 34626 19966 34638 20018
rect 34690 19966 34702 20018
rect 44930 19966 44942 20018
rect 44994 19966 45006 20018
rect 5406 19954 5458 19966
rect 10558 19954 10610 19966
rect 11006 19954 11058 19966
rect 14926 19954 14978 19966
rect 24670 19954 24722 19966
rect 27134 19954 27186 19966
rect 39790 19954 39842 19966
rect 14814 19906 14866 19918
rect 18174 19906 18226 19918
rect 7410 19854 7422 19906
rect 7474 19854 7486 19906
rect 15586 19854 15598 19906
rect 15650 19854 15662 19906
rect 14814 19842 14866 19854
rect 18174 19842 18226 19854
rect 18734 19906 18786 19918
rect 18734 19842 18786 19854
rect 20862 19906 20914 19918
rect 34302 19906 34354 19918
rect 37886 19906 37938 19918
rect 23538 19854 23550 19906
rect 23602 19854 23614 19906
rect 25890 19854 25902 19906
rect 25954 19854 25966 19906
rect 31266 19854 31278 19906
rect 31330 19854 31342 19906
rect 37426 19854 37438 19906
rect 37490 19854 37502 19906
rect 20862 19842 20914 19854
rect 34302 19842 34354 19854
rect 37886 19842 37938 19854
rect 38558 19906 38610 19918
rect 38558 19842 38610 19854
rect 39454 19906 39506 19918
rect 47730 19854 47742 19906
rect 47794 19854 47806 19906
rect 39454 19842 39506 19854
rect 13358 19794 13410 19806
rect 7634 19742 7646 19794
rect 7698 19791 7710 19794
rect 8082 19791 8094 19794
rect 7698 19745 8094 19791
rect 7698 19742 7710 19745
rect 8082 19742 8094 19745
rect 8146 19742 8158 19794
rect 13358 19730 13410 19742
rect 13470 19794 13522 19806
rect 13470 19730 13522 19742
rect 13694 19794 13746 19806
rect 18510 19794 18562 19806
rect 14354 19742 14366 19794
rect 14418 19742 14430 19794
rect 13694 19730 13746 19742
rect 18510 19730 18562 19742
rect 19966 19794 20018 19806
rect 19966 19730 20018 19742
rect 20302 19794 20354 19806
rect 20302 19730 20354 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 11118 19458 11170 19470
rect 11118 19394 11170 19406
rect 12574 19458 12626 19470
rect 12574 19394 12626 19406
rect 14926 19458 14978 19470
rect 14926 19394 14978 19406
rect 15262 19458 15314 19470
rect 15262 19394 15314 19406
rect 23550 19458 23602 19470
rect 23550 19394 23602 19406
rect 27022 19458 27074 19470
rect 27022 19394 27074 19406
rect 29262 19458 29314 19470
rect 29262 19394 29314 19406
rect 29598 19458 29650 19470
rect 29598 19394 29650 19406
rect 23326 19346 23378 19358
rect 7186 19294 7198 19346
rect 7250 19294 7262 19346
rect 23326 19282 23378 19294
rect 24334 19346 24386 19358
rect 37214 19346 37266 19358
rect 26674 19294 26686 19346
rect 26738 19294 26750 19346
rect 31938 19294 31950 19346
rect 32002 19294 32014 19346
rect 34066 19294 34078 19346
rect 34130 19294 34142 19346
rect 24334 19282 24386 19294
rect 37214 19282 37266 19294
rect 11006 19234 11058 19246
rect 15150 19234 15202 19246
rect 8418 19182 8430 19234
rect 8482 19182 8494 19234
rect 9762 19182 9774 19234
rect 9826 19182 9838 19234
rect 11330 19182 11342 19234
rect 11394 19182 11406 19234
rect 12674 19182 12686 19234
rect 12738 19182 12750 19234
rect 14242 19182 14254 19234
rect 14306 19182 14318 19234
rect 14690 19182 14702 19234
rect 14754 19182 14766 19234
rect 11006 19170 11058 19182
rect 15150 19170 15202 19182
rect 16158 19234 16210 19246
rect 16158 19170 16210 19182
rect 16494 19234 16546 19246
rect 19854 19234 19906 19246
rect 19170 19182 19182 19234
rect 19234 19182 19246 19234
rect 16494 19170 16546 19182
rect 19854 19170 19906 19182
rect 21982 19234 22034 19246
rect 21982 19170 22034 19182
rect 22318 19234 22370 19246
rect 35534 19234 35586 19246
rect 31154 19182 31166 19234
rect 31218 19182 31230 19234
rect 22318 19170 22370 19182
rect 35534 19170 35586 19182
rect 4062 19122 4114 19134
rect 4062 19058 4114 19070
rect 6862 19122 6914 19134
rect 6862 19058 6914 19070
rect 7086 19122 7138 19134
rect 7086 19058 7138 19070
rect 7646 19122 7698 19134
rect 7646 19058 7698 19070
rect 7758 19122 7810 19134
rect 7758 19058 7810 19070
rect 8094 19122 8146 19134
rect 8094 19058 8146 19070
rect 8766 19122 8818 19134
rect 8766 19058 8818 19070
rect 9102 19122 9154 19134
rect 9102 19058 9154 19070
rect 9998 19122 10050 19134
rect 9998 19058 10050 19070
rect 10670 19122 10722 19134
rect 10670 19058 10722 19070
rect 12126 19122 12178 19134
rect 26798 19122 26850 19134
rect 12338 19070 12350 19122
rect 12402 19070 12414 19122
rect 14018 19070 14030 19122
rect 14082 19070 14094 19122
rect 22642 19070 22654 19122
rect 22706 19070 22718 19122
rect 29810 19070 29822 19122
rect 29874 19070 29886 19122
rect 30370 19070 30382 19122
rect 30434 19070 30446 19122
rect 35746 19070 35758 19122
rect 35810 19070 35822 19122
rect 36082 19070 36094 19122
rect 36146 19070 36158 19122
rect 12126 19058 12178 19070
rect 26798 19058 26850 19070
rect 3726 19010 3778 19022
rect 3726 18946 3778 18958
rect 5742 19010 5794 19022
rect 5742 18946 5794 18958
rect 7422 19010 7474 19022
rect 7422 18946 7474 18958
rect 8206 19010 8258 19022
rect 12910 19010 12962 19022
rect 16606 19010 16658 19022
rect 10882 18958 10894 19010
rect 10946 18958 10958 19010
rect 15810 18958 15822 19010
rect 15874 18958 15886 19010
rect 8206 18946 8258 18958
rect 12910 18946 12962 18958
rect 16606 18946 16658 18958
rect 19406 19010 19458 19022
rect 19406 18946 19458 18958
rect 21646 19010 21698 19022
rect 24894 19010 24946 19022
rect 23874 18958 23886 19010
rect 23938 18958 23950 19010
rect 21646 18946 21698 18958
rect 24894 18946 24946 18958
rect 28030 19010 28082 19022
rect 28030 18946 28082 18958
rect 35198 19010 35250 19022
rect 35198 18946 35250 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 8318 18674 8370 18686
rect 13022 18674 13074 18686
rect 9986 18622 9998 18674
rect 10050 18622 10062 18674
rect 11554 18622 11566 18674
rect 11618 18622 11630 18674
rect 8318 18610 8370 18622
rect 13022 18610 13074 18622
rect 14366 18674 14418 18686
rect 14366 18610 14418 18622
rect 23214 18674 23266 18686
rect 23214 18610 23266 18622
rect 25230 18674 25282 18686
rect 25230 18610 25282 18622
rect 30830 18674 30882 18686
rect 30830 18610 30882 18622
rect 2270 18562 2322 18574
rect 7534 18562 7586 18574
rect 9550 18562 9602 18574
rect 3378 18510 3390 18562
rect 3442 18510 3454 18562
rect 6850 18510 6862 18562
rect 6914 18510 6926 18562
rect 8978 18510 8990 18562
rect 9042 18510 9054 18562
rect 2270 18498 2322 18510
rect 7534 18498 7586 18510
rect 9550 18498 9602 18510
rect 14478 18562 14530 18574
rect 14478 18498 14530 18510
rect 15374 18562 15426 18574
rect 24222 18562 24274 18574
rect 19506 18510 19518 18562
rect 19570 18510 19582 18562
rect 23538 18510 23550 18562
rect 23602 18510 23614 18562
rect 15374 18498 15426 18510
rect 24222 18498 24274 18510
rect 26014 18562 26066 18574
rect 26014 18498 26066 18510
rect 29710 18562 29762 18574
rect 29710 18498 29762 18510
rect 29934 18562 29986 18574
rect 29934 18498 29986 18510
rect 34078 18562 34130 18574
rect 34078 18498 34130 18510
rect 35198 18562 35250 18574
rect 35198 18498 35250 18510
rect 5966 18450 6018 18462
rect 2034 18398 2046 18450
rect 2098 18398 2110 18450
rect 2706 18398 2718 18450
rect 2770 18398 2782 18450
rect 5966 18386 6018 18398
rect 6302 18450 6354 18462
rect 7982 18450 8034 18462
rect 11118 18450 11170 18462
rect 11566 18450 11618 18462
rect 12238 18450 12290 18462
rect 12686 18450 12738 18462
rect 14142 18450 14194 18462
rect 15038 18450 15090 18462
rect 22094 18450 22146 18462
rect 25566 18450 25618 18462
rect 7074 18398 7086 18450
rect 7138 18398 7150 18450
rect 7746 18398 7758 18450
rect 7810 18398 7822 18450
rect 8306 18398 8318 18450
rect 8370 18398 8382 18450
rect 8754 18398 8766 18450
rect 8818 18398 8830 18450
rect 9762 18398 9774 18450
rect 9826 18398 9838 18450
rect 10098 18398 10110 18450
rect 10162 18398 10174 18450
rect 11330 18398 11342 18450
rect 11394 18398 11406 18450
rect 11666 18398 11678 18450
rect 11730 18398 11742 18450
rect 12450 18398 12462 18450
rect 12514 18398 12526 18450
rect 12786 18398 12798 18450
rect 12850 18398 12862 18450
rect 13682 18398 13694 18450
rect 13746 18398 13758 18450
rect 14802 18398 14814 18450
rect 14866 18398 14878 18450
rect 18722 18398 18734 18450
rect 18786 18398 18798 18450
rect 23986 18398 23998 18450
rect 24050 18398 24062 18450
rect 25218 18398 25230 18450
rect 25282 18398 25294 18450
rect 6302 18386 6354 18398
rect 7982 18386 8034 18398
rect 11118 18386 11170 18398
rect 11566 18386 11618 18398
rect 12238 18386 12290 18398
rect 12686 18386 12738 18398
rect 14142 18386 14194 18398
rect 15038 18386 15090 18398
rect 22094 18386 22146 18398
rect 25566 18386 25618 18398
rect 25678 18450 25730 18462
rect 33742 18450 33794 18462
rect 28354 18398 28366 18450
rect 28418 18398 28430 18450
rect 34962 18398 34974 18450
rect 35026 18398 35038 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 38434 18398 38446 18450
rect 38498 18398 38510 18450
rect 25678 18386 25730 18398
rect 33742 18386 33794 18398
rect 38894 18338 38946 18350
rect 5506 18286 5518 18338
rect 5570 18286 5582 18338
rect 21634 18286 21646 18338
rect 21698 18286 21710 18338
rect 35522 18286 35534 18338
rect 35586 18286 35598 18338
rect 38894 18274 38946 18286
rect 15262 18226 15314 18238
rect 10098 18174 10110 18226
rect 10162 18174 10174 18226
rect 13906 18174 13918 18226
rect 13970 18174 13982 18226
rect 15262 18162 15314 18174
rect 28030 18226 28082 18238
rect 28030 18162 28082 18174
rect 28366 18226 28418 18238
rect 28366 18162 28418 18174
rect 29598 18226 29650 18238
rect 29598 18162 29650 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 5742 17890 5794 17902
rect 5742 17826 5794 17838
rect 6078 17890 6130 17902
rect 6078 17826 6130 17838
rect 12462 17890 12514 17902
rect 12462 17826 12514 17838
rect 14030 17890 14082 17902
rect 14030 17826 14082 17838
rect 14254 17890 14306 17902
rect 14254 17826 14306 17838
rect 24446 17890 24498 17902
rect 24446 17826 24498 17838
rect 25342 17890 25394 17902
rect 25342 17826 25394 17838
rect 26350 17890 26402 17902
rect 26350 17826 26402 17838
rect 29598 17890 29650 17902
rect 29598 17826 29650 17838
rect 9886 17778 9938 17790
rect 2482 17726 2494 17778
rect 2546 17726 2558 17778
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 9886 17714 9938 17726
rect 17166 17778 17218 17790
rect 17166 17714 17218 17726
rect 27694 17778 27746 17790
rect 33394 17726 33406 17778
rect 33458 17726 33470 17778
rect 35522 17726 35534 17778
rect 35586 17726 35598 17778
rect 27694 17714 27746 17726
rect 8766 17666 8818 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 6850 17614 6862 17666
rect 6914 17614 6926 17666
rect 8766 17602 8818 17614
rect 9438 17666 9490 17678
rect 9438 17602 9490 17614
rect 12350 17666 12402 17678
rect 21534 17666 21586 17678
rect 26462 17666 26514 17678
rect 12562 17614 12574 17666
rect 12626 17614 12638 17666
rect 13794 17614 13806 17666
rect 13858 17614 13870 17666
rect 16594 17614 16606 17666
rect 16658 17614 16670 17666
rect 22530 17614 22542 17666
rect 22594 17614 22606 17666
rect 24098 17614 24110 17666
rect 24162 17614 24174 17666
rect 26114 17614 26126 17666
rect 26178 17614 26190 17666
rect 12350 17602 12402 17614
rect 21534 17602 21586 17614
rect 26462 17602 26514 17614
rect 29150 17666 29202 17678
rect 32174 17666 32226 17678
rect 37102 17666 37154 17678
rect 29362 17614 29374 17666
rect 29426 17614 29438 17666
rect 29698 17614 29710 17666
rect 29762 17614 29774 17666
rect 36194 17614 36206 17666
rect 36258 17614 36270 17666
rect 29150 17602 29202 17614
rect 32174 17602 32226 17614
rect 37102 17602 37154 17614
rect 12014 17554 12066 17566
rect 6738 17502 6750 17554
rect 6802 17502 6814 17554
rect 8418 17502 8430 17554
rect 8482 17502 8494 17554
rect 9090 17502 9102 17554
rect 9154 17502 9166 17554
rect 11330 17502 11342 17554
rect 11394 17502 11406 17554
rect 12014 17490 12066 17502
rect 15598 17554 15650 17566
rect 15598 17490 15650 17502
rect 15934 17554 15986 17566
rect 15934 17490 15986 17502
rect 16382 17554 16434 17566
rect 16382 17490 16434 17502
rect 22990 17554 23042 17566
rect 24894 17554 24946 17566
rect 23314 17502 23326 17554
rect 23378 17502 23390 17554
rect 24658 17502 24670 17554
rect 24722 17502 24734 17554
rect 22990 17490 23042 17502
rect 24894 17490 24946 17502
rect 25454 17554 25506 17566
rect 25454 17490 25506 17502
rect 26798 17554 26850 17566
rect 26798 17490 26850 17502
rect 30382 17554 30434 17566
rect 30382 17490 30434 17502
rect 31838 17554 31890 17566
rect 32386 17502 32398 17554
rect 32450 17502 32462 17554
rect 32722 17502 32734 17554
rect 32786 17502 32798 17554
rect 31838 17490 31890 17502
rect 5070 17442 5122 17454
rect 5070 17378 5122 17390
rect 11678 17442 11730 17454
rect 11678 17378 11730 17390
rect 12798 17442 12850 17454
rect 12798 17378 12850 17390
rect 13918 17442 13970 17454
rect 13918 17378 13970 17390
rect 21198 17442 21250 17454
rect 21198 17378 21250 17390
rect 21422 17442 21474 17454
rect 21422 17378 21474 17390
rect 21982 17442 22034 17454
rect 24110 17442 24162 17454
rect 22306 17390 22318 17442
rect 22370 17390 22382 17442
rect 21982 17378 22034 17390
rect 24110 17378 24162 17390
rect 25342 17442 25394 17454
rect 25342 17378 25394 17390
rect 26686 17442 26738 17454
rect 26686 17378 26738 17390
rect 27134 17442 27186 17454
rect 27134 17378 27186 17390
rect 29262 17442 29314 17454
rect 29262 17378 29314 17390
rect 30718 17442 30770 17454
rect 30718 17378 30770 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 6302 17106 6354 17118
rect 6302 17042 6354 17054
rect 7086 17106 7138 17118
rect 7086 17042 7138 17054
rect 8094 17106 8146 17118
rect 8094 17042 8146 17054
rect 8542 17106 8594 17118
rect 8542 17042 8594 17054
rect 10334 17106 10386 17118
rect 10334 17042 10386 17054
rect 11006 17106 11058 17118
rect 13694 17106 13746 17118
rect 13346 17054 13358 17106
rect 13410 17054 13422 17106
rect 11006 17042 11058 17054
rect 13694 17042 13746 17054
rect 14814 17106 14866 17118
rect 14814 17042 14866 17054
rect 15374 17106 15426 17118
rect 15374 17042 15426 17054
rect 16494 17106 16546 17118
rect 16494 17042 16546 17054
rect 20750 17106 20802 17118
rect 20750 17042 20802 17054
rect 22878 17106 22930 17118
rect 23774 17106 23826 17118
rect 23202 17054 23214 17106
rect 23266 17054 23278 17106
rect 22878 17042 22930 17054
rect 23774 17042 23826 17054
rect 24782 17106 24834 17118
rect 24782 17042 24834 17054
rect 33630 17106 33682 17118
rect 33630 17042 33682 17054
rect 16158 16994 16210 17006
rect 23998 16994 24050 17006
rect 7746 16942 7758 16994
rect 7810 16942 7822 16994
rect 15026 16942 15038 16994
rect 15090 16942 15102 16994
rect 16818 16942 16830 16994
rect 16882 16942 16894 16994
rect 16158 16930 16210 16942
rect 23998 16930 24050 16942
rect 24558 16994 24610 17006
rect 28142 16994 28194 17006
rect 26002 16942 26014 16994
rect 26066 16942 26078 16994
rect 28354 16942 28366 16994
rect 28418 16942 28430 16994
rect 31714 16942 31726 16994
rect 31778 16942 31790 16994
rect 34178 16942 34190 16994
rect 34242 16942 34254 16994
rect 34514 16942 34526 16994
rect 34578 16942 34590 16994
rect 24558 16930 24610 16942
rect 28142 16930 28194 16942
rect 6974 16882 7026 16894
rect 23550 16882 23602 16894
rect 15922 16830 15934 16882
rect 15986 16830 15998 16882
rect 17490 16830 17502 16882
rect 17554 16830 17566 16882
rect 6974 16818 7026 16830
rect 23550 16818 23602 16830
rect 24446 16882 24498 16894
rect 28590 16882 28642 16894
rect 33182 16882 33234 16894
rect 27794 16830 27806 16882
rect 27858 16830 27870 16882
rect 28690 16830 28702 16882
rect 28754 16830 28766 16882
rect 32498 16830 32510 16882
rect 32562 16830 32574 16882
rect 24446 16818 24498 16830
rect 28590 16818 28642 16830
rect 33182 16818 33234 16830
rect 6190 16770 6242 16782
rect 6190 16706 6242 16718
rect 10222 16770 10274 16782
rect 10222 16706 10274 16718
rect 11118 16770 11170 16782
rect 23662 16770 23714 16782
rect 18162 16718 18174 16770
rect 18226 16718 18238 16770
rect 20290 16718 20302 16770
rect 20354 16718 20366 16770
rect 11118 16706 11170 16718
rect 23662 16706 23714 16718
rect 28254 16770 28306 16782
rect 29586 16718 29598 16770
rect 29650 16718 29662 16770
rect 28254 16706 28306 16718
rect 33966 16658 34018 16670
rect 33966 16594 34018 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 14926 16322 14978 16334
rect 14926 16258 14978 16270
rect 16158 16322 16210 16334
rect 16158 16258 16210 16270
rect 19518 16322 19570 16334
rect 19518 16258 19570 16270
rect 26350 16322 26402 16334
rect 26350 16258 26402 16270
rect 26686 16322 26738 16334
rect 26686 16258 26738 16270
rect 29486 16322 29538 16334
rect 29486 16258 29538 16270
rect 30382 16322 30434 16334
rect 30382 16258 30434 16270
rect 30718 16322 30770 16334
rect 30718 16258 30770 16270
rect 11790 16210 11842 16222
rect 11330 16158 11342 16210
rect 11394 16158 11406 16210
rect 11790 16146 11842 16158
rect 17502 16210 17554 16222
rect 17502 16146 17554 16158
rect 23998 16210 24050 16222
rect 23998 16146 24050 16158
rect 24894 16210 24946 16222
rect 24894 16146 24946 16158
rect 25790 16210 25842 16222
rect 25790 16146 25842 16158
rect 6078 16098 6130 16110
rect 7198 16098 7250 16110
rect 6850 16046 6862 16098
rect 6914 16046 6926 16098
rect 6078 16034 6130 16046
rect 7198 16034 7250 16046
rect 7534 16098 7586 16110
rect 7534 16034 7586 16046
rect 7870 16098 7922 16110
rect 12798 16098 12850 16110
rect 15150 16098 15202 16110
rect 8530 16046 8542 16098
rect 8594 16046 8606 16098
rect 14130 16046 14142 16098
rect 14194 16046 14206 16098
rect 7870 16034 7922 16046
rect 12798 16034 12850 16046
rect 15150 16034 15202 16046
rect 15822 16098 15874 16110
rect 15822 16034 15874 16046
rect 17054 16098 17106 16110
rect 22878 16098 22930 16110
rect 20290 16046 20302 16098
rect 20354 16046 20366 16098
rect 17054 16034 17106 16046
rect 22878 16034 22930 16046
rect 25230 16098 25282 16110
rect 25230 16034 25282 16046
rect 25678 16098 25730 16110
rect 35534 16098 35586 16110
rect 27346 16046 27358 16098
rect 27410 16046 27422 16098
rect 29138 16046 29150 16098
rect 29202 16046 29214 16098
rect 25678 16034 25730 16046
rect 35534 16034 35586 16046
rect 4062 15986 4114 15998
rect 7422 15986 7474 15998
rect 16270 15986 16322 15998
rect 18286 15986 18338 15998
rect 6738 15934 6750 15986
rect 6802 15934 6814 15986
rect 9202 15934 9214 15986
rect 9266 15934 9278 15986
rect 13794 15934 13806 15986
rect 13858 15934 13870 15986
rect 16706 15934 16718 15986
rect 16770 15934 16782 15986
rect 4062 15922 4114 15934
rect 7422 15922 7474 15934
rect 16270 15922 16322 15934
rect 18286 15922 18338 15934
rect 18622 15986 18674 15998
rect 18622 15922 18674 15934
rect 19182 15986 19234 15998
rect 23662 15986 23714 15998
rect 20066 15934 20078 15986
rect 20130 15934 20142 15986
rect 19182 15922 19234 15934
rect 23662 15922 23714 15934
rect 24558 15986 24610 15998
rect 29934 15986 29986 15998
rect 27458 15934 27470 15986
rect 27522 15934 27534 15986
rect 29698 15934 29710 15986
rect 29762 15934 29774 15986
rect 30930 15934 30942 15986
rect 30994 15934 31006 15986
rect 31266 15934 31278 15986
rect 31330 15934 31342 15986
rect 35746 15934 35758 15986
rect 35810 15934 35822 15986
rect 36306 15934 36318 15986
rect 36370 15934 36382 15986
rect 24558 15922 24610 15934
rect 29934 15922 29986 15934
rect 3726 15874 3778 15886
rect 3726 15810 3778 15822
rect 5742 15874 5794 15886
rect 5742 15810 5794 15822
rect 7982 15874 8034 15886
rect 7982 15810 8034 15822
rect 8206 15874 8258 15886
rect 8206 15810 8258 15822
rect 12238 15874 12290 15886
rect 12238 15810 12290 15822
rect 12462 15874 12514 15886
rect 12462 15810 12514 15822
rect 12686 15874 12738 15886
rect 22654 15874 22706 15886
rect 23886 15874 23938 15886
rect 13570 15822 13582 15874
rect 13634 15822 13646 15874
rect 14578 15822 14590 15874
rect 14642 15822 14654 15874
rect 15474 15822 15486 15874
rect 15538 15822 15550 15874
rect 23202 15822 23214 15874
rect 23266 15822 23278 15874
rect 12686 15810 12738 15822
rect 22654 15810 22706 15822
rect 23886 15810 23938 15822
rect 24110 15874 24162 15886
rect 24110 15810 24162 15822
rect 24782 15874 24834 15886
rect 24782 15810 24834 15822
rect 25006 15874 25058 15886
rect 25006 15810 25058 15822
rect 25902 15874 25954 15886
rect 25902 15810 25954 15822
rect 28030 15874 28082 15886
rect 28030 15810 28082 15822
rect 29150 15874 29202 15886
rect 29150 15810 29202 15822
rect 35198 15874 35250 15886
rect 35198 15810 35250 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 6078 15538 6130 15550
rect 6078 15474 6130 15486
rect 7870 15538 7922 15550
rect 7870 15474 7922 15486
rect 8990 15538 9042 15550
rect 8990 15474 9042 15486
rect 13582 15538 13634 15550
rect 13582 15474 13634 15486
rect 14478 15538 14530 15550
rect 14478 15474 14530 15486
rect 15486 15538 15538 15550
rect 15486 15474 15538 15486
rect 16158 15538 16210 15550
rect 16158 15474 16210 15486
rect 16494 15538 16546 15550
rect 16494 15474 16546 15486
rect 17390 15538 17442 15550
rect 17390 15474 17442 15486
rect 23774 15538 23826 15550
rect 23774 15474 23826 15486
rect 27246 15538 27298 15550
rect 27246 15474 27298 15486
rect 2382 15426 2434 15438
rect 8430 15426 8482 15438
rect 3490 15374 3502 15426
rect 3554 15374 3566 15426
rect 7186 15374 7198 15426
rect 7250 15374 7262 15426
rect 2382 15362 2434 15374
rect 8430 15362 8482 15374
rect 13694 15426 13746 15438
rect 13694 15362 13746 15374
rect 14926 15426 14978 15438
rect 26238 15426 26290 15438
rect 35422 15426 35474 15438
rect 16818 15374 16830 15426
rect 16882 15374 16894 15426
rect 17714 15374 17726 15426
rect 17778 15374 17790 15426
rect 28578 15374 28590 15426
rect 28642 15374 28654 15426
rect 29026 15374 29038 15426
rect 29090 15374 29102 15426
rect 31378 15374 31390 15426
rect 31442 15374 31454 15426
rect 31714 15374 31726 15426
rect 31778 15374 31790 15426
rect 37874 15374 37886 15426
rect 37938 15374 37950 15426
rect 14926 15362 14978 15374
rect 26238 15362 26290 15374
rect 35422 15362 35474 15374
rect 6414 15314 6466 15326
rect 27022 15314 27074 15326
rect 2146 15262 2158 15314
rect 2210 15262 2222 15314
rect 2818 15262 2830 15314
rect 2882 15262 2894 15314
rect 6850 15262 6862 15314
rect 6914 15262 6926 15314
rect 8754 15262 8766 15314
rect 8818 15262 8830 15314
rect 9986 15262 9998 15314
rect 10050 15262 10062 15314
rect 20178 15262 20190 15314
rect 20242 15262 20254 15314
rect 24210 15262 24222 15314
rect 24274 15262 24286 15314
rect 25666 15262 25678 15314
rect 25730 15262 25742 15314
rect 26562 15262 26574 15314
rect 26626 15262 26638 15314
rect 6414 15250 6466 15262
rect 27022 15250 27074 15262
rect 27358 15314 27410 15326
rect 27358 15250 27410 15262
rect 27918 15314 27970 15326
rect 27918 15250 27970 15262
rect 28254 15314 28306 15326
rect 28254 15250 28306 15262
rect 35086 15314 35138 15326
rect 39118 15314 39170 15326
rect 38658 15262 38670 15314
rect 38722 15262 38734 15314
rect 35086 15250 35138 15262
rect 39118 15250 39170 15262
rect 12574 15202 12626 15214
rect 5618 15150 5630 15202
rect 5682 15150 5694 15202
rect 11778 15150 11790 15202
rect 11842 15150 11854 15202
rect 20850 15150 20862 15202
rect 20914 15150 20926 15202
rect 22978 15150 22990 15202
rect 23042 15150 23054 15202
rect 24546 15150 24558 15202
rect 24610 15150 24622 15202
rect 25778 15150 25790 15202
rect 25842 15150 25854 15202
rect 35746 15150 35758 15202
rect 35810 15150 35822 15202
rect 12574 15138 12626 15150
rect 13582 15090 13634 15102
rect 30830 15090 30882 15102
rect 26786 15038 26798 15090
rect 26850 15038 26862 15090
rect 13582 15026 13634 15038
rect 30830 15026 30882 15038
rect 31166 15090 31218 15102
rect 31166 15026 31218 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 11118 14754 11170 14766
rect 11118 14690 11170 14702
rect 11454 14754 11506 14766
rect 11454 14690 11506 14702
rect 28030 14754 28082 14766
rect 28030 14690 28082 14702
rect 35198 14754 35250 14766
rect 35198 14690 35250 14702
rect 5070 14642 5122 14654
rect 2482 14590 2494 14642
rect 2546 14590 2558 14642
rect 4610 14590 4622 14642
rect 4674 14590 4686 14642
rect 5070 14578 5122 14590
rect 5854 14642 5906 14654
rect 22878 14642 22930 14654
rect 9762 14590 9774 14642
rect 9826 14590 9838 14642
rect 19842 14590 19854 14642
rect 19906 14590 19918 14642
rect 24434 14590 24446 14642
rect 24498 14590 24510 14642
rect 31154 14590 31166 14642
rect 31218 14590 31230 14642
rect 5854 14578 5906 14590
rect 22878 14578 22930 14590
rect 14030 14530 14082 14542
rect 16606 14530 16658 14542
rect 22542 14530 22594 14542
rect 26574 14530 26626 14542
rect 28478 14530 28530 14542
rect 34526 14530 34578 14542
rect 1810 14478 1822 14530
rect 1874 14478 1886 14530
rect 6962 14478 6974 14530
rect 7026 14478 7038 14530
rect 12226 14478 12238 14530
rect 12290 14478 12302 14530
rect 14466 14478 14478 14530
rect 14530 14478 14542 14530
rect 16930 14478 16942 14530
rect 16994 14478 17006 14530
rect 20402 14478 20414 14530
rect 20466 14478 20478 14530
rect 22194 14478 22206 14530
rect 22258 14478 22270 14530
rect 22754 14478 22766 14530
rect 22818 14478 22830 14530
rect 23538 14478 23550 14530
rect 23602 14478 23614 14530
rect 26226 14478 26238 14530
rect 26290 14478 26302 14530
rect 26786 14478 26798 14530
rect 26850 14478 26862 14530
rect 27682 14478 27694 14530
rect 27746 14478 27758 14530
rect 28242 14478 28254 14530
rect 28306 14478 28318 14530
rect 30594 14478 30606 14530
rect 30658 14478 30670 14530
rect 33954 14478 33966 14530
rect 34018 14478 34030 14530
rect 14030 14466 14082 14478
rect 16606 14466 16658 14478
rect 22542 14466 22594 14478
rect 26574 14466 26626 14478
rect 28478 14466 28530 14478
rect 34526 14466 34578 14478
rect 35534 14530 35586 14542
rect 35534 14466 35586 14478
rect 10446 14418 10498 14430
rect 13470 14418 13522 14430
rect 7634 14366 7646 14418
rect 7698 14366 7710 14418
rect 12002 14366 12014 14418
rect 12066 14366 12078 14418
rect 10446 14354 10498 14366
rect 13470 14354 13522 14366
rect 16046 14418 16098 14430
rect 20638 14418 20690 14430
rect 17714 14366 17726 14418
rect 17778 14366 17790 14418
rect 16046 14354 16098 14366
rect 20638 14354 20690 14366
rect 22990 14418 23042 14430
rect 22990 14354 23042 14366
rect 27022 14418 27074 14430
rect 27022 14354 27074 14366
rect 30830 14418 30882 14430
rect 33282 14366 33294 14418
rect 33346 14366 33358 14418
rect 35746 14366 35758 14418
rect 35810 14366 35822 14418
rect 36082 14366 36094 14418
rect 36146 14366 36158 14418
rect 30830 14354 30882 14366
rect 10110 14306 10162 14318
rect 10110 14242 10162 14254
rect 12910 14306 12962 14318
rect 12910 14242 12962 14254
rect 14702 14306 14754 14318
rect 14702 14242 14754 14254
rect 26238 14306 26290 14318
rect 26238 14242 26290 14254
rect 27694 14306 27746 14318
rect 27694 14242 27746 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 7982 13970 8034 13982
rect 7982 13906 8034 13918
rect 9102 13970 9154 13982
rect 9102 13906 9154 13918
rect 11454 13970 11506 13982
rect 11454 13906 11506 13918
rect 16718 13970 16770 13982
rect 16718 13906 16770 13918
rect 21422 13970 21474 13982
rect 21422 13906 21474 13918
rect 22654 13970 22706 13982
rect 25566 13970 25618 13982
rect 23986 13918 23998 13970
rect 24050 13918 24062 13970
rect 22654 13906 22706 13918
rect 25566 13906 25618 13918
rect 26686 13970 26738 13982
rect 26686 13906 26738 13918
rect 27022 13970 27074 13982
rect 27022 13906 27074 13918
rect 28814 13970 28866 13982
rect 28814 13906 28866 13918
rect 29150 13970 29202 13982
rect 33182 13970 33234 13982
rect 29474 13918 29486 13970
rect 29538 13918 29550 13970
rect 29150 13906 29202 13918
rect 33182 13906 33234 13918
rect 2606 13858 2658 13870
rect 6066 13806 6078 13858
rect 6130 13806 6142 13858
rect 10770 13806 10782 13858
rect 10834 13806 10846 13858
rect 12450 13806 12462 13858
rect 12514 13806 12526 13858
rect 15138 13806 15150 13858
rect 15202 13806 15214 13858
rect 19506 13806 19518 13858
rect 19570 13806 19582 13858
rect 20290 13806 20302 13858
rect 20354 13806 20366 13858
rect 26114 13806 26126 13858
rect 26178 13806 26190 13858
rect 33730 13806 33742 13858
rect 33794 13806 33806 13858
rect 34178 13806 34190 13858
rect 34242 13806 34254 13858
rect 36306 13806 36318 13858
rect 36370 13806 36382 13858
rect 36530 13806 36542 13858
rect 36594 13806 36606 13858
rect 2606 13794 2658 13806
rect 2942 13746 2994 13758
rect 8318 13746 8370 13758
rect 6178 13694 6190 13746
rect 6242 13694 6254 13746
rect 2942 13682 2994 13694
rect 8318 13682 8370 13694
rect 9774 13746 9826 13758
rect 9774 13682 9826 13694
rect 10110 13746 10162 13758
rect 21086 13746 21138 13758
rect 10882 13694 10894 13746
rect 10946 13694 10958 13746
rect 12562 13694 12574 13746
rect 12626 13694 12638 13746
rect 15810 13694 15822 13746
rect 15874 13694 15886 13746
rect 19730 13694 19742 13746
rect 19794 13694 19806 13746
rect 20514 13694 20526 13746
rect 20578 13694 20590 13746
rect 10110 13682 10162 13694
rect 21086 13682 21138 13694
rect 21870 13746 21922 13758
rect 21870 13682 21922 13694
rect 22206 13746 22258 13758
rect 23550 13746 23602 13758
rect 22642 13694 22654 13746
rect 22706 13694 22718 13746
rect 22206 13682 22258 13694
rect 23550 13682 23602 13694
rect 23886 13746 23938 13758
rect 25902 13746 25954 13758
rect 27470 13746 27522 13758
rect 24098 13694 24110 13746
rect 24162 13694 24174 13746
rect 26450 13694 26462 13746
rect 26514 13694 26526 13746
rect 27234 13694 27246 13746
rect 27298 13694 27310 13746
rect 23886 13682 23938 13694
rect 25902 13682 25954 13694
rect 27470 13682 27522 13694
rect 27806 13746 27858 13758
rect 27806 13682 27858 13694
rect 33518 13746 33570 13758
rect 33518 13682 33570 13694
rect 35646 13746 35698 13758
rect 35646 13682 35698 13694
rect 35982 13746 36034 13758
rect 35982 13682 36034 13694
rect 13010 13582 13022 13634
rect 13074 13582 13086 13634
rect 5070 13522 5122 13534
rect 5070 13458 5122 13470
rect 5406 13522 5458 13534
rect 5406 13458 5458 13470
rect 11790 13522 11842 13534
rect 11790 13458 11842 13470
rect 18622 13522 18674 13534
rect 18622 13458 18674 13470
rect 18958 13522 19010 13534
rect 18958 13458 19010 13470
rect 22318 13522 22370 13534
rect 22318 13458 22370 13470
rect 23998 13522 24050 13534
rect 27358 13522 27410 13534
rect 26450 13470 26462 13522
rect 26514 13470 26526 13522
rect 23998 13458 24050 13470
rect 27358 13458 27410 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 5742 13186 5794 13198
rect 5742 13122 5794 13134
rect 8654 13186 8706 13198
rect 8654 13122 8706 13134
rect 8990 13186 9042 13198
rect 8990 13122 9042 13134
rect 14366 13186 14418 13198
rect 14366 13122 14418 13134
rect 14702 13186 14754 13198
rect 14702 13122 14754 13134
rect 19070 13186 19122 13198
rect 19070 13122 19122 13134
rect 20302 13186 20354 13198
rect 20302 13122 20354 13134
rect 22206 13186 22258 13198
rect 22206 13122 22258 13134
rect 24334 13186 24386 13198
rect 24334 13122 24386 13134
rect 27022 13186 27074 13198
rect 27022 13122 27074 13134
rect 6078 13074 6130 13086
rect 21310 13074 21362 13086
rect 2482 13022 2494 13074
rect 2546 13022 2558 13074
rect 4610 13022 4622 13074
rect 4674 13022 4686 13074
rect 12562 13022 12574 13074
rect 12626 13022 12638 13074
rect 6078 13010 6130 13022
rect 21310 13010 21362 13022
rect 22318 13074 22370 13086
rect 25442 13022 25454 13074
rect 25506 13022 25518 13074
rect 26226 13022 26238 13074
rect 26290 13022 26302 13074
rect 29138 13022 29150 13074
rect 29202 13022 29214 13074
rect 22318 13010 22370 13022
rect 18286 12962 18338 12974
rect 21646 12962 21698 12974
rect 23662 12962 23714 12974
rect 26686 12962 26738 12974
rect 1810 12910 1822 12962
rect 1874 12910 1886 12962
rect 7522 12910 7534 12962
rect 7586 12910 7598 12962
rect 9538 12910 9550 12962
rect 9602 12910 9614 12962
rect 10770 12910 10782 12962
rect 10834 12910 10846 12962
rect 19730 12910 19742 12962
rect 19794 12910 19806 12962
rect 22530 12910 22542 12962
rect 22594 12910 22606 12962
rect 23426 12910 23438 12962
rect 23490 12910 23502 12962
rect 23762 12910 23774 12962
rect 23826 12910 23838 12962
rect 25218 12910 25230 12962
rect 25282 12910 25294 12962
rect 18286 12898 18338 12910
rect 21646 12898 21698 12910
rect 23662 12898 23714 12910
rect 26686 12898 26738 12910
rect 27358 12962 27410 12974
rect 32510 12962 32562 12974
rect 28354 12910 28366 12962
rect 28418 12910 28430 12962
rect 32050 12910 32062 12962
rect 32114 12910 32126 12962
rect 27358 12898 27410 12910
rect 32510 12898 32562 12910
rect 36318 12962 36370 12974
rect 36318 12898 36370 12910
rect 17950 12850 18002 12862
rect 6290 12798 6302 12850
rect 6354 12798 6366 12850
rect 6738 12798 6750 12850
rect 6802 12798 6814 12850
rect 9762 12798 9774 12850
rect 9826 12798 9838 12850
rect 13794 12798 13806 12850
rect 13858 12798 13870 12850
rect 14018 12798 14030 12850
rect 14082 12798 14094 12850
rect 17950 12786 18002 12798
rect 18958 12850 19010 12862
rect 21870 12850 21922 12862
rect 23214 12850 23266 12862
rect 19506 12798 19518 12850
rect 19570 12798 19582 12850
rect 22754 12798 22766 12850
rect 22818 12847 22830 12850
rect 22978 12847 22990 12850
rect 22818 12801 22990 12847
rect 22818 12798 22830 12801
rect 22978 12798 22990 12801
rect 23042 12798 23054 12850
rect 18958 12786 19010 12798
rect 21870 12786 21922 12798
rect 23214 12786 23266 12798
rect 25790 12850 25842 12862
rect 25790 12786 25842 12798
rect 27134 12850 27186 12862
rect 27134 12786 27186 12798
rect 28590 12850 28642 12862
rect 35534 12850 35586 12862
rect 31266 12798 31278 12850
rect 31330 12798 31342 12850
rect 28590 12786 28642 12798
rect 35534 12786 35586 12798
rect 5070 12738 5122 12750
rect 5070 12674 5122 12686
rect 7310 12738 7362 12750
rect 7310 12674 7362 12686
rect 20638 12738 20690 12750
rect 20638 12674 20690 12686
rect 23998 12738 24050 12750
rect 23998 12674 24050 12686
rect 24446 12738 24498 12750
rect 24446 12674 24498 12686
rect 24558 12738 24610 12750
rect 24558 12674 24610 12686
rect 35870 12738 35922 12750
rect 35870 12674 35922 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 13134 12402 13186 12414
rect 13134 12338 13186 12350
rect 15038 12402 15090 12414
rect 15038 12338 15090 12350
rect 19966 12402 20018 12414
rect 19966 12338 20018 12350
rect 23550 12402 23602 12414
rect 23550 12338 23602 12350
rect 25790 12402 25842 12414
rect 25790 12338 25842 12350
rect 28254 12402 28306 12414
rect 28254 12338 28306 12350
rect 29598 12402 29650 12414
rect 29598 12338 29650 12350
rect 39678 12402 39730 12414
rect 39678 12338 39730 12350
rect 32510 12290 32562 12302
rect 6850 12238 6862 12290
rect 6914 12238 6926 12290
rect 10322 12238 10334 12290
rect 10386 12238 10398 12290
rect 14018 12238 14030 12290
rect 14082 12238 14094 12290
rect 14466 12238 14478 12290
rect 14530 12238 14542 12290
rect 28802 12238 28814 12290
rect 28866 12238 28878 12290
rect 30258 12238 30270 12290
rect 30322 12238 30334 12290
rect 30482 12238 30494 12290
rect 30546 12238 30558 12290
rect 33842 12238 33854 12290
rect 33906 12238 33918 12290
rect 38434 12238 38446 12290
rect 38498 12238 38510 12290
rect 32510 12226 32562 12238
rect 5630 12178 5682 12190
rect 26126 12178 26178 12190
rect 29038 12178 29090 12190
rect 2370 12126 2382 12178
rect 2434 12126 2446 12178
rect 6178 12126 6190 12178
rect 6242 12126 6254 12178
rect 9538 12126 9550 12178
rect 9602 12126 9614 12178
rect 23090 12126 23102 12178
rect 23154 12126 23166 12178
rect 26338 12126 26350 12178
rect 26402 12126 26414 12178
rect 28242 12126 28254 12178
rect 28306 12126 28318 12178
rect 5630 12114 5682 12126
rect 26126 12114 26178 12126
rect 29038 12114 29090 12126
rect 29934 12178 29986 12190
rect 32274 12126 32286 12178
rect 32338 12126 32350 12178
rect 33058 12126 33070 12178
rect 33122 12126 33134 12178
rect 39106 12126 39118 12178
rect 39170 12126 39182 12178
rect 29934 12114 29986 12126
rect 13470 12066 13522 12078
rect 3042 12014 3054 12066
rect 3106 12014 3118 12066
rect 5170 12014 5182 12066
rect 5234 12014 5246 12066
rect 8978 12014 8990 12066
rect 9042 12014 9054 12066
rect 12450 12014 12462 12066
rect 12514 12014 12526 12066
rect 13470 12002 13522 12014
rect 15598 12066 15650 12078
rect 26910 12066 26962 12078
rect 20178 12014 20190 12066
rect 20242 12014 20254 12066
rect 22306 12014 22318 12066
rect 22370 12014 22382 12066
rect 35970 12014 35982 12066
rect 36034 12014 36046 12066
rect 36306 12014 36318 12066
rect 36370 12014 36382 12066
rect 15598 12002 15650 12014
rect 26910 12002 26962 12014
rect 14702 11954 14754 11966
rect 28466 11902 28478 11954
rect 28530 11902 28542 11954
rect 14702 11890 14754 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 7310 11618 7362 11630
rect 7310 11554 7362 11566
rect 7646 11618 7698 11630
rect 7646 11554 7698 11566
rect 11230 11618 11282 11630
rect 11230 11554 11282 11566
rect 11566 11618 11618 11630
rect 11566 11554 11618 11566
rect 23886 11618 23938 11630
rect 23886 11554 23938 11566
rect 31950 11618 32002 11630
rect 31950 11554 32002 11566
rect 33182 11618 33234 11630
rect 33182 11554 33234 11566
rect 33518 11618 33570 11630
rect 33518 11554 33570 11566
rect 35198 11618 35250 11630
rect 35198 11554 35250 11566
rect 9214 11506 9266 11518
rect 20750 11506 20802 11518
rect 18498 11454 18510 11506
rect 18562 11454 18574 11506
rect 19954 11454 19966 11506
rect 20018 11454 20030 11506
rect 9214 11442 9266 11454
rect 20750 11442 20802 11454
rect 21422 11506 21474 11518
rect 21422 11442 21474 11454
rect 25678 11506 25730 11518
rect 29262 11506 29314 11518
rect 26114 11454 26126 11506
rect 26178 11454 26190 11506
rect 25678 11442 25730 11454
rect 29262 11442 29314 11454
rect 29710 11506 29762 11518
rect 29710 11442 29762 11454
rect 3726 11394 3778 11406
rect 15262 11394 15314 11406
rect 22206 11394 22258 11406
rect 8082 11342 8094 11394
rect 8146 11342 8158 11394
rect 12002 11342 12014 11394
rect 12066 11342 12078 11394
rect 13682 11342 13694 11394
rect 13746 11342 13758 11394
rect 15586 11342 15598 11394
rect 15650 11342 15662 11394
rect 20066 11342 20078 11394
rect 20130 11342 20142 11394
rect 3726 11330 3778 11342
rect 15262 11330 15314 11342
rect 22206 11330 22258 11342
rect 24222 11394 24274 11406
rect 35534 11394 35586 11406
rect 24882 11342 24894 11394
rect 24946 11342 24958 11394
rect 26226 11342 26238 11394
rect 26290 11342 26302 11394
rect 34290 11342 34302 11394
rect 34354 11342 34366 11394
rect 24222 11330 24274 11342
rect 35534 11330 35586 11342
rect 3390 11282 3442 11294
rect 19182 11282 19234 11294
rect 8194 11230 8206 11282
rect 8258 11230 8270 11282
rect 12114 11230 12126 11282
rect 12178 11230 12190 11282
rect 16370 11230 16382 11282
rect 16434 11230 16446 11282
rect 3390 11218 3442 11230
rect 19182 11218 19234 11230
rect 19518 11282 19570 11294
rect 19518 11218 19570 11230
rect 22542 11282 22594 11294
rect 22542 11218 22594 11230
rect 22878 11282 22930 11294
rect 26798 11282 26850 11294
rect 24994 11230 25006 11282
rect 25058 11230 25070 11282
rect 22878 11218 22930 11230
rect 26798 11218 26850 11230
rect 32062 11282 32114 11294
rect 32062 11218 32114 11230
rect 32286 11282 32338 11294
rect 34178 11230 34190 11282
rect 34242 11230 34254 11282
rect 35746 11230 35758 11282
rect 35810 11230 35822 11282
rect 36306 11230 36318 11282
rect 36370 11230 36382 11282
rect 32286 11218 32338 11230
rect 13470 11170 13522 11182
rect 13470 11106 13522 11118
rect 18846 11170 18898 11182
rect 18846 11106 18898 11118
rect 22990 11170 23042 11182
rect 22990 11106 23042 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 11566 10834 11618 10846
rect 11566 10770 11618 10782
rect 12126 10834 12178 10846
rect 12126 10770 12178 10782
rect 16382 10834 16434 10846
rect 16382 10770 16434 10782
rect 19182 10834 19234 10846
rect 19182 10770 19234 10782
rect 24222 10834 24274 10846
rect 24222 10770 24274 10782
rect 27134 10834 27186 10846
rect 27134 10770 27186 10782
rect 29486 10834 29538 10846
rect 29486 10770 29538 10782
rect 22766 10722 22818 10734
rect 26798 10722 26850 10734
rect 30494 10722 30546 10734
rect 7970 10670 7982 10722
rect 8034 10670 8046 10722
rect 11778 10670 11790 10722
rect 11842 10670 11854 10722
rect 13234 10670 13246 10722
rect 13298 10670 13310 10722
rect 15698 10670 15710 10722
rect 15762 10670 15774 10722
rect 18386 10670 18398 10722
rect 18450 10670 18462 10722
rect 19730 10670 19742 10722
rect 19794 10670 19806 10722
rect 20290 10670 20302 10722
rect 20354 10670 20366 10722
rect 25330 10670 25342 10722
rect 25394 10670 25406 10722
rect 28578 10670 28590 10722
rect 28642 10670 28654 10722
rect 28914 10670 28926 10722
rect 28978 10670 28990 10722
rect 29810 10670 29822 10722
rect 29874 10670 29886 10722
rect 31490 10670 31502 10722
rect 31554 10670 31566 10722
rect 32050 10670 32062 10722
rect 32114 10670 32126 10722
rect 22766 10658 22818 10670
rect 26798 10658 26850 10670
rect 30494 10658 30546 10670
rect 16046 10610 16098 10622
rect 8082 10558 8094 10610
rect 8146 10558 8158 10610
rect 12450 10558 12462 10610
rect 12514 10558 12526 10610
rect 16046 10546 16098 10558
rect 16718 10610 16770 10622
rect 16718 10546 16770 10558
rect 17502 10610 17554 10622
rect 26014 10610 26066 10622
rect 18610 10558 18622 10610
rect 18674 10558 18686 10610
rect 22978 10558 22990 10610
rect 23042 10558 23054 10610
rect 25554 10558 25566 10610
rect 25618 10558 25630 10610
rect 17502 10546 17554 10558
rect 26014 10546 26066 10558
rect 26462 10610 26514 10622
rect 31278 10610 31330 10622
rect 30258 10558 30270 10610
rect 30322 10558 30334 10610
rect 26462 10546 26514 10558
rect 31278 10546 31330 10558
rect 11006 10498 11058 10510
rect 19518 10498 19570 10510
rect 15362 10446 15374 10498
rect 15426 10446 15438 10498
rect 11006 10434 11058 10446
rect 19518 10434 19570 10446
rect 20862 10498 20914 10510
rect 20862 10434 20914 10446
rect 24670 10498 24722 10510
rect 24670 10434 24722 10446
rect 27246 10498 27298 10510
rect 27246 10434 27298 10446
rect 30942 10498 30994 10510
rect 30942 10434 30994 10446
rect 7086 10386 7138 10398
rect 7086 10322 7138 10334
rect 7422 10386 7474 10398
rect 7422 10322 7474 10334
rect 17838 10386 17890 10398
rect 17838 10322 17890 10334
rect 27918 10386 27970 10398
rect 27918 10322 27970 10334
rect 28254 10386 28306 10398
rect 28254 10322 28306 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 11678 10050 11730 10062
rect 11678 9986 11730 9998
rect 13694 10050 13746 10062
rect 13694 9986 13746 9998
rect 29934 10050 29986 10062
rect 29934 9986 29986 9998
rect 12014 9938 12066 9950
rect 11218 9886 11230 9938
rect 11282 9886 11294 9938
rect 12014 9874 12066 9886
rect 16382 9938 16434 9950
rect 29822 9938 29874 9950
rect 18386 9886 18398 9938
rect 18450 9886 18462 9938
rect 20514 9886 20526 9938
rect 20578 9886 20590 9938
rect 22194 9886 22206 9938
rect 22258 9886 22270 9938
rect 24322 9886 24334 9938
rect 24386 9886 24398 9938
rect 27570 9886 27582 9938
rect 27634 9886 27646 9938
rect 31042 9886 31054 9938
rect 31106 9886 31118 9938
rect 33170 9886 33182 9938
rect 33234 9886 33246 9938
rect 16382 9874 16434 9886
rect 29822 9874 29874 9886
rect 6862 9826 6914 9838
rect 14030 9826 14082 9838
rect 28030 9826 28082 9838
rect 8418 9774 8430 9826
rect 8482 9774 8494 9826
rect 12786 9774 12798 9826
rect 12850 9774 12862 9826
rect 17714 9774 17726 9826
rect 17778 9774 17790 9826
rect 21522 9774 21534 9826
rect 21586 9774 21598 9826
rect 24770 9774 24782 9826
rect 24834 9774 24846 9826
rect 6862 9762 6914 9774
rect 14030 9762 14082 9774
rect 28030 9762 28082 9774
rect 29486 9826 29538 9838
rect 30258 9774 30270 9826
rect 30322 9774 30334 9826
rect 29486 9762 29538 9774
rect 9090 9662 9102 9714
rect 9154 9662 9166 9714
rect 12562 9662 12574 9714
rect 12626 9662 12638 9714
rect 14242 9662 14254 9714
rect 14306 9662 14318 9714
rect 14690 9662 14702 9714
rect 14754 9662 14766 9714
rect 25442 9662 25454 9714
rect 25506 9662 25518 9714
rect 6526 9602 6578 9614
rect 6526 9538 6578 9550
rect 28366 9602 28418 9614
rect 29138 9550 29150 9602
rect 29202 9550 29214 9602
rect 28366 9538 28418 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 9550 9266 9602 9278
rect 9550 9202 9602 9214
rect 12238 9266 12290 9278
rect 12238 9202 12290 9214
rect 19294 9266 19346 9278
rect 19294 9202 19346 9214
rect 22206 9266 22258 9278
rect 22206 9202 22258 9214
rect 25342 9266 25394 9278
rect 25342 9202 25394 9214
rect 6402 9102 6414 9154
rect 6466 9102 6478 9154
rect 11330 9102 11342 9154
rect 11394 9102 11406 9154
rect 12786 9102 12798 9154
rect 12850 9102 12862 9154
rect 13346 9102 13358 9154
rect 13410 9102 13422 9154
rect 21522 9102 21534 9154
rect 21586 9102 21598 9154
rect 23202 9102 23214 9154
rect 23266 9102 23278 9154
rect 26898 9102 26910 9154
rect 26962 9102 26974 9154
rect 28466 9102 28478 9154
rect 28530 9102 28542 9154
rect 8990 9042 9042 9054
rect 5730 8990 5742 9042
rect 5794 8990 5806 9042
rect 8990 8978 9042 8990
rect 9886 9042 9938 9054
rect 9886 8978 9938 8990
rect 10446 9042 10498 9054
rect 10446 8978 10498 8990
rect 10782 9042 10834 9054
rect 23774 9042 23826 9054
rect 11554 8990 11566 9042
rect 11618 8990 11630 9042
rect 18610 8990 18622 9042
rect 18674 8990 18686 9042
rect 21634 8990 21646 9042
rect 21698 8990 21710 9042
rect 23314 8990 23326 9042
rect 23378 8990 23390 9042
rect 10782 8978 10834 8990
rect 23774 8978 23826 8990
rect 24110 9042 24162 9054
rect 26786 8990 26798 9042
rect 26850 8990 26862 9042
rect 27794 8990 27806 9042
rect 27858 8990 27870 9042
rect 24110 8978 24162 8990
rect 18062 8930 18114 8942
rect 19742 8930 19794 8942
rect 8530 8878 8542 8930
rect 8594 8878 8606 8930
rect 18386 8878 18398 8930
rect 18450 8878 18462 8930
rect 18062 8866 18114 8878
rect 19742 8866 19794 8878
rect 23998 8930 24050 8942
rect 30594 8878 30606 8930
rect 30658 8878 30670 8930
rect 23998 8866 24050 8878
rect 12574 8818 12626 8830
rect 20526 8818 20578 8830
rect 19058 8766 19070 8818
rect 19122 8815 19134 8818
rect 19394 8815 19406 8818
rect 19122 8769 19406 8815
rect 19122 8766 19134 8769
rect 19394 8766 19406 8769
rect 19458 8815 19470 8818
rect 19730 8815 19742 8818
rect 19458 8769 19742 8815
rect 19458 8766 19470 8769
rect 19730 8766 19742 8769
rect 19794 8766 19806 8818
rect 12574 8754 12626 8766
rect 20526 8754 20578 8766
rect 20862 8818 20914 8830
rect 20862 8754 20914 8766
rect 22542 8818 22594 8830
rect 22542 8754 22594 8766
rect 25790 8818 25842 8830
rect 25790 8754 25842 8766
rect 26126 8818 26178 8830
rect 26126 8754 26178 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 22194 8430 22206 8482
rect 22258 8430 22270 8482
rect 11454 8370 11506 8382
rect 11454 8306 11506 8318
rect 15262 8370 15314 8382
rect 20750 8370 20802 8382
rect 22766 8370 22818 8382
rect 18498 8318 18510 8370
rect 18562 8318 18574 8370
rect 19506 8318 19518 8370
rect 19570 8318 19582 8370
rect 21634 8318 21646 8370
rect 21698 8318 21710 8370
rect 15262 8306 15314 8318
rect 20750 8306 20802 8318
rect 22766 8306 22818 8318
rect 23102 8370 23154 8382
rect 23102 8306 23154 8318
rect 24446 8370 24498 8382
rect 24446 8306 24498 8318
rect 21982 8258 22034 8270
rect 25790 8258 25842 8270
rect 15586 8206 15598 8258
rect 15650 8206 15662 8258
rect 19394 8206 19406 8258
rect 19458 8206 19470 8258
rect 23874 8206 23886 8258
rect 23938 8206 23950 8258
rect 21982 8194 22034 8206
rect 25790 8194 25842 8206
rect 29934 8258 29986 8270
rect 29934 8194 29986 8206
rect 18846 8146 18898 8158
rect 16370 8094 16382 8146
rect 16434 8094 16446 8146
rect 18846 8082 18898 8094
rect 20078 8146 20130 8158
rect 25454 8146 25506 8158
rect 23650 8094 23662 8146
rect 23714 8094 23726 8146
rect 20078 8082 20130 8094
rect 25454 8082 25506 8094
rect 27358 8034 27410 8046
rect 27358 7970 27410 7982
rect 27806 8034 27858 8046
rect 27806 7970 27858 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 14702 7698 14754 7710
rect 14702 7634 14754 7646
rect 16382 7698 16434 7710
rect 16382 7634 16434 7646
rect 22878 7698 22930 7710
rect 22878 7634 22930 7646
rect 23326 7698 23378 7710
rect 23326 7634 23378 7646
rect 26350 7698 26402 7710
rect 26350 7634 26402 7646
rect 29150 7698 29202 7710
rect 29150 7634 29202 7646
rect 10222 7586 10274 7598
rect 25342 7586 25394 7598
rect 12226 7534 12238 7586
rect 12290 7534 12302 7586
rect 14130 7534 14142 7586
rect 14194 7534 14206 7586
rect 15810 7534 15822 7586
rect 15874 7534 15886 7586
rect 18050 7534 18062 7586
rect 18114 7534 18126 7586
rect 18498 7534 18510 7586
rect 18562 7534 18574 7586
rect 28242 7534 28254 7586
rect 28306 7534 28318 7586
rect 28690 7534 28702 7586
rect 28754 7534 28766 7586
rect 10222 7522 10274 7534
rect 25342 7522 25394 7534
rect 10558 7474 10610 7486
rect 10558 7410 10610 7422
rect 11118 7474 11170 7486
rect 11118 7410 11170 7422
rect 11454 7474 11506 7486
rect 13358 7474 13410 7486
rect 16718 7474 16770 7486
rect 12114 7422 12126 7474
rect 12178 7422 12190 7474
rect 14018 7422 14030 7474
rect 14082 7422 14094 7474
rect 15698 7422 15710 7474
rect 15762 7422 15774 7474
rect 11454 7410 11506 7422
rect 13358 7410 13410 7422
rect 16718 7410 16770 7422
rect 17502 7474 17554 7486
rect 17502 7410 17554 7422
rect 17838 7474 17890 7486
rect 25678 7474 25730 7486
rect 19506 7422 19518 7474
rect 19570 7422 19582 7474
rect 17838 7410 17890 7422
rect 25678 7410 25730 7422
rect 27918 7474 27970 7486
rect 27918 7410 27970 7422
rect 26462 7362 26514 7374
rect 20178 7310 20190 7362
rect 20242 7310 20254 7362
rect 22306 7310 22318 7362
rect 22370 7310 22382 7362
rect 26462 7298 26514 7310
rect 29262 7362 29314 7374
rect 29262 7298 29314 7310
rect 13022 7250 13074 7262
rect 13022 7186 13074 7198
rect 15038 7250 15090 7262
rect 15038 7186 15090 7198
rect 27582 7250 27634 7262
rect 27582 7186 27634 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 17166 6914 17218 6926
rect 17166 6850 17218 6862
rect 19854 6802 19906 6814
rect 28590 6802 28642 6814
rect 10098 6750 10110 6802
rect 10162 6750 10174 6802
rect 12226 6750 12238 6802
rect 12290 6750 12302 6802
rect 25330 6750 25342 6802
rect 25394 6750 25406 6802
rect 27458 6750 27470 6802
rect 27522 6750 27534 6802
rect 19854 6738 19906 6750
rect 28590 6738 28642 6750
rect 12686 6690 12738 6702
rect 22542 6690 22594 6702
rect 27806 6690 27858 6702
rect 9314 6638 9326 6690
rect 9378 6638 9390 6690
rect 13682 6638 13694 6690
rect 13746 6638 13758 6690
rect 17938 6638 17950 6690
rect 18002 6638 18014 6690
rect 20626 6638 20638 6690
rect 20690 6638 20702 6690
rect 24658 6638 24670 6690
rect 24722 6638 24734 6690
rect 12686 6626 12738 6638
rect 22542 6626 22594 6638
rect 27806 6626 27858 6638
rect 20414 6578 20466 6590
rect 17714 6526 17726 6578
rect 17778 6526 17790 6578
rect 20414 6514 20466 6526
rect 13470 6466 13522 6478
rect 13470 6402 13522 6414
rect 16270 6466 16322 6478
rect 16270 6402 16322 6414
rect 16830 6466 16882 6478
rect 16830 6402 16882 6414
rect 28142 6466 28194 6478
rect 28142 6402 28194 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 11790 6130 11842 6142
rect 11790 6066 11842 6078
rect 25678 6130 25730 6142
rect 25678 6066 25730 6078
rect 16382 6018 16434 6030
rect 12898 5966 12910 6018
rect 12962 5966 12974 6018
rect 16382 5954 16434 5966
rect 16718 6018 16770 6030
rect 21970 5966 21982 6018
rect 22034 5966 22046 6018
rect 23314 5966 23326 6018
rect 23378 5966 23390 6018
rect 23874 5966 23886 6018
rect 23938 5966 23950 6018
rect 26562 5966 26574 6018
rect 26626 5966 26638 6018
rect 28018 5966 28030 6018
rect 28082 5966 28094 6018
rect 16718 5954 16770 5966
rect 21422 5906 21474 5918
rect 23102 5906 23154 5918
rect 12114 5854 12126 5906
rect 12178 5854 12190 5906
rect 22194 5854 22206 5906
rect 22258 5854 22270 5906
rect 21422 5842 21474 5854
rect 23102 5842 23154 5854
rect 26014 5906 26066 5918
rect 26674 5854 26686 5906
rect 26738 5854 26750 5906
rect 27234 5854 27246 5906
rect 27298 5854 27310 5906
rect 26014 5842 26066 5854
rect 15026 5742 15038 5794
rect 15090 5742 15102 5794
rect 30146 5742 30158 5794
rect 30210 5742 30222 5794
rect 21086 5682 21138 5694
rect 21086 5618 21138 5630
rect 22766 5682 22818 5694
rect 22766 5618 22818 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 15374 5234 15426 5246
rect 25342 5234 25394 5246
rect 16370 5182 16382 5234
rect 16434 5182 16446 5234
rect 18498 5182 18510 5234
rect 18562 5182 18574 5234
rect 24882 5182 24894 5234
rect 24946 5182 24958 5234
rect 15374 5170 15426 5182
rect 25342 5170 25394 5182
rect 26910 5234 26962 5246
rect 26910 5170 26962 5182
rect 20414 5122 20466 5134
rect 15586 5070 15598 5122
rect 15650 5070 15662 5122
rect 20414 5058 20466 5070
rect 21310 5122 21362 5134
rect 22082 5070 22094 5122
rect 22146 5070 22158 5122
rect 22754 5070 22766 5122
rect 22818 5070 22830 5122
rect 21310 5058 21362 5070
rect 21646 5010 21698 5022
rect 21646 4946 21698 4958
rect 20750 4898 20802 4910
rect 20750 4834 20802 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 23774 4562 23826 4574
rect 23774 4498 23826 4510
rect 21186 4398 21198 4450
rect 21250 4398 21262 4450
rect 20514 4286 20526 4338
rect 20578 4286 20590 4338
rect 23314 4174 23326 4226
rect 23378 4174 23390 4226
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 12574 57038 12626 57090
rect 13134 57038 13186 57090
rect 54238 56814 54290 56866
rect 55022 56814 55074 56866
rect 16046 56702 16098 56754
rect 17054 56702 17106 56754
rect 17166 56590 17218 56642
rect 17950 56590 18002 56642
rect 18510 56590 18562 56642
rect 18958 56590 19010 56642
rect 24222 56590 24274 56642
rect 25006 56590 25058 56642
rect 28702 56590 28754 56642
rect 29374 56590 29426 56642
rect 44382 56590 44434 56642
rect 44942 56590 44994 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4622 56254 4674 56306
rect 6190 56254 6242 56306
rect 7422 56254 7474 56306
rect 8654 56254 8706 56306
rect 10110 56254 10162 56306
rect 11454 56254 11506 56306
rect 13134 56254 13186 56306
rect 14030 56254 14082 56306
rect 15038 56254 15090 56306
rect 17166 56254 17218 56306
rect 19406 56254 19458 56306
rect 20750 56254 20802 56306
rect 23214 56254 23266 56306
rect 30718 56254 30770 56306
rect 35310 56254 35362 56306
rect 39118 56254 39170 56306
rect 44046 56254 44098 56306
rect 45390 56254 45442 56306
rect 46398 56254 46450 56306
rect 47854 56254 47906 56306
rect 49086 56254 49138 56306
rect 50430 56254 50482 56306
rect 51774 56254 51826 56306
rect 53118 56254 53170 56306
rect 55022 56254 55074 56306
rect 55918 56254 55970 56306
rect 5518 56142 5570 56194
rect 5854 56142 5906 56194
rect 15710 56142 15762 56194
rect 16046 56142 16098 56194
rect 16382 56142 16434 56194
rect 17614 56142 17666 56194
rect 18622 56142 18674 56194
rect 18958 56142 19010 56194
rect 19854 56142 19906 56194
rect 20190 56142 20242 56194
rect 21310 56142 21362 56194
rect 15486 56030 15538 56082
rect 22430 56030 22482 56082
rect 23998 56030 24050 56082
rect 27358 56030 27410 56082
rect 28702 56030 28754 56082
rect 31390 56030 31442 56082
rect 32174 56030 32226 56082
rect 33742 56030 33794 56082
rect 35982 56030 36034 56082
rect 37550 56030 37602 56082
rect 39790 56030 39842 56082
rect 42478 56030 42530 56082
rect 4958 55918 5010 55970
rect 6974 55918 7026 55970
rect 8206 55918 8258 55970
rect 9662 55918 9714 55970
rect 11006 55918 11058 55970
rect 12350 55918 12402 55970
rect 13582 55918 13634 55970
rect 14590 55918 14642 55970
rect 17726 55918 17778 55970
rect 21982 55918 22034 55970
rect 24558 55918 24610 55970
rect 26686 55918 26738 55970
rect 29374 55918 29426 55970
rect 30494 55918 30546 55970
rect 32622 55918 32674 55970
rect 34190 55918 34242 55970
rect 36430 55918 36482 55970
rect 37998 55918 38050 55970
rect 40350 55918 40402 55970
rect 42030 55918 42082 55970
rect 42926 55918 42978 55970
rect 43598 55918 43650 55970
rect 44494 55918 44546 55970
rect 44942 55918 44994 55970
rect 45950 55918 46002 55970
rect 47406 55918 47458 55970
rect 48638 55918 48690 55970
rect 49982 55918 50034 55970
rect 51326 55918 51378 55970
rect 52670 55918 52722 55970
rect 54014 55918 54066 55970
rect 55470 55918 55522 55970
rect 17838 55806 17890 55858
rect 18286 55806 18338 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 15934 55470 15986 55522
rect 17838 55470 17890 55522
rect 18510 55470 18562 55522
rect 19406 55470 19458 55522
rect 20414 55470 20466 55522
rect 4622 55358 4674 55410
rect 5966 55358 6018 55410
rect 15598 55358 15650 55410
rect 18846 55358 18898 55410
rect 25230 55358 25282 55410
rect 28590 55358 28642 55410
rect 32062 55358 32114 55410
rect 35758 55358 35810 55410
rect 37438 55358 37490 55410
rect 39342 55358 39394 55410
rect 1822 55246 1874 55298
rect 8878 55246 8930 55298
rect 16942 55246 16994 55298
rect 17502 55246 17554 55298
rect 18062 55246 18114 55298
rect 22318 55246 22370 55298
rect 25790 55246 25842 55298
rect 29150 55246 29202 55298
rect 32958 55246 33010 55298
rect 38110 55246 38162 55298
rect 42142 55246 42194 55298
rect 2494 55134 2546 55186
rect 8094 55134 8146 55186
rect 16382 55134 16434 55186
rect 16830 55134 16882 55186
rect 17278 55134 17330 55186
rect 17614 55134 17666 55186
rect 19070 55134 19122 55186
rect 21758 55134 21810 55186
rect 23102 55134 23154 55186
rect 26462 55134 26514 55186
rect 29934 55134 29986 55186
rect 32398 55134 32450 55186
rect 33630 55134 33682 55186
rect 36094 55134 36146 55186
rect 38558 55134 38610 55186
rect 41470 55134 41522 55186
rect 42590 55134 42642 55186
rect 42702 55134 42754 55186
rect 43262 55134 43314 55186
rect 43934 55134 43986 55186
rect 5070 55022 5122 55074
rect 9326 55022 9378 55074
rect 16606 55022 16658 55074
rect 19966 55022 20018 55074
rect 21422 55022 21474 55074
rect 43598 55022 43650 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 2494 54686 2546 54738
rect 15934 54686 15986 54738
rect 16606 54686 16658 54738
rect 16830 54686 16882 54738
rect 22990 54686 23042 54738
rect 23886 54686 23938 54738
rect 25566 54686 25618 54738
rect 26462 54686 26514 54738
rect 27694 54686 27746 54738
rect 28030 54686 28082 54738
rect 29150 54686 29202 54738
rect 29822 54686 29874 54738
rect 31166 54686 31218 54738
rect 39230 54686 39282 54738
rect 40462 54686 40514 54738
rect 41582 54686 41634 54738
rect 2382 54574 2434 54626
rect 7646 54574 7698 54626
rect 16382 54574 16434 54626
rect 40910 54574 40962 54626
rect 41246 54574 41298 54626
rect 44606 54574 44658 54626
rect 2606 54462 2658 54514
rect 2942 54462 2994 54514
rect 3726 54462 3778 54514
rect 4398 54462 4450 54514
rect 6638 54462 6690 54514
rect 7086 54462 7138 54514
rect 7422 54462 7474 54514
rect 11902 54462 11954 54514
rect 12238 54462 12290 54514
rect 18286 54462 18338 54514
rect 18510 54462 18562 54514
rect 19630 54462 19682 54514
rect 24558 54462 24610 54514
rect 27246 54462 27298 54514
rect 28814 54462 28866 54514
rect 35310 54462 35362 54514
rect 45390 54462 45442 54514
rect 3614 54350 3666 54402
rect 4958 54350 5010 54402
rect 6862 54350 6914 54402
rect 7758 54350 7810 54402
rect 9886 54350 9938 54402
rect 13022 54350 13074 54402
rect 15150 54350 15202 54402
rect 18398 54350 18450 54402
rect 20414 54350 20466 54402
rect 22542 54350 22594 54402
rect 32286 54350 32338 54402
rect 33182 54350 33234 54402
rect 34302 54350 34354 54402
rect 34862 54350 34914 54402
rect 35982 54350 36034 54402
rect 38110 54350 38162 54402
rect 42142 54350 42194 54402
rect 42478 54350 42530 54402
rect 45838 54350 45890 54402
rect 48078 54350 48130 54402
rect 16942 54238 16994 54290
rect 18846 54238 18898 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 17502 53902 17554 53954
rect 17838 53902 17890 53954
rect 18958 53902 19010 53954
rect 24670 53902 24722 53954
rect 4622 53790 4674 53842
rect 5070 53790 5122 53842
rect 9662 53790 9714 53842
rect 12910 53790 12962 53842
rect 18398 53790 18450 53842
rect 22990 53790 23042 53842
rect 34078 53790 34130 53842
rect 35198 53790 35250 53842
rect 38670 53790 38722 53842
rect 42926 53790 42978 53842
rect 43262 53790 43314 53842
rect 47742 53790 47794 53842
rect 51326 53790 51378 53842
rect 1822 53678 1874 53730
rect 6750 53678 6802 53730
rect 9998 53678 10050 53730
rect 13470 53678 13522 53730
rect 17278 53678 17330 53730
rect 18622 53678 18674 53730
rect 19182 53678 19234 53730
rect 20302 53678 20354 53730
rect 21870 53678 21922 53730
rect 23662 53678 23714 53730
rect 24670 53678 24722 53730
rect 31166 53678 31218 53730
rect 38894 53678 38946 53730
rect 39230 53678 39282 53730
rect 39902 53678 39954 53730
rect 43486 53678 43538 53730
rect 44830 53678 44882 53730
rect 48414 53678 48466 53730
rect 2494 53566 2546 53618
rect 7534 53566 7586 53618
rect 10782 53566 10834 53618
rect 19742 53566 19794 53618
rect 23102 53566 23154 53618
rect 23438 53566 23490 53618
rect 23998 53566 24050 53618
rect 24334 53566 24386 53618
rect 25006 53566 25058 53618
rect 27134 53566 27186 53618
rect 30718 53566 30770 53618
rect 31950 53566 32002 53618
rect 34638 53566 34690 53618
rect 35534 53566 35586 53618
rect 35870 53566 35922 53618
rect 36206 53566 36258 53618
rect 38670 53566 38722 53618
rect 40350 53566 40402 53618
rect 45614 53566 45666 53618
rect 49198 53566 49250 53618
rect 13806 53454 13858 53506
rect 19294 53454 19346 53506
rect 19630 53454 19682 53506
rect 19854 53454 19906 53506
rect 20638 53454 20690 53506
rect 21422 53454 21474 53506
rect 22542 53454 22594 53506
rect 22878 53454 22930 53506
rect 23774 53454 23826 53506
rect 25678 53454 25730 53506
rect 29262 53454 29314 53506
rect 30382 53454 30434 53506
rect 34750 53454 34802 53506
rect 34974 53454 35026 53506
rect 35310 53454 35362 53506
rect 38446 53454 38498 53506
rect 39566 53454 39618 53506
rect 40238 53454 40290 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 2830 53118 2882 53170
rect 3614 53118 3666 53170
rect 14366 53118 14418 53170
rect 24110 53118 24162 53170
rect 31390 53118 31442 53170
rect 32174 53118 32226 53170
rect 33854 53118 33906 53170
rect 34638 53118 34690 53170
rect 36766 53118 36818 53170
rect 39454 53118 39506 53170
rect 39678 53118 39730 53170
rect 45614 53118 45666 53170
rect 47966 53118 48018 53170
rect 48974 53118 49026 53170
rect 2718 53006 2770 53058
rect 3390 53006 3442 53058
rect 4510 53006 4562 53058
rect 9998 53006 10050 53058
rect 11566 53006 11618 53058
rect 14478 53006 14530 53058
rect 20190 53006 20242 53058
rect 23998 53006 24050 53058
rect 25454 53006 25506 53058
rect 28814 53006 28866 53058
rect 32510 53006 32562 53058
rect 33966 53006 34018 53058
rect 37214 53006 37266 53058
rect 38670 53006 38722 53058
rect 41022 53006 41074 53058
rect 41918 53006 41970 53058
rect 42254 53006 42306 53058
rect 42590 53006 42642 53058
rect 45502 53006 45554 53058
rect 3054 52894 3106 52946
rect 3726 52894 3778 52946
rect 3838 52894 3890 52946
rect 4398 52894 4450 52946
rect 4622 52894 4674 52946
rect 6414 52894 6466 52946
rect 6526 52894 6578 52946
rect 6750 52894 6802 52946
rect 6974 52894 7026 52946
rect 7422 52894 7474 52946
rect 7534 52894 7586 52946
rect 10334 52894 10386 52946
rect 12462 52894 12514 52946
rect 12910 52894 12962 52946
rect 13358 52894 13410 52946
rect 13694 52894 13746 52946
rect 13918 52894 13970 52946
rect 19406 52894 19458 52946
rect 23550 52894 23602 52946
rect 23774 52894 23826 52946
rect 26014 52894 26066 52946
rect 28030 52894 28082 52946
rect 34190 52894 34242 52946
rect 34414 52894 34466 52946
rect 35534 52894 35586 52946
rect 35870 52894 35922 52946
rect 36094 52894 36146 52946
rect 38110 52894 38162 52946
rect 38446 52894 38498 52946
rect 38782 52894 38834 52946
rect 39230 52894 39282 52946
rect 40238 52894 40290 52946
rect 40910 52894 40962 52946
rect 46062 52894 46114 52946
rect 46622 52894 46674 52946
rect 48750 52894 48802 52946
rect 50094 52894 50146 52946
rect 7198 52782 7250 52834
rect 9662 52782 9714 52834
rect 13022 52782 13074 52834
rect 13470 52782 13522 52834
rect 14254 52782 14306 52834
rect 16606 52782 16658 52834
rect 19070 52782 19122 52834
rect 22318 52782 22370 52834
rect 24110 52782 24162 52834
rect 30942 52782 30994 52834
rect 35086 52782 35138 52834
rect 43038 52782 43090 52834
rect 49086 52782 49138 52834
rect 49422 52782 49474 52834
rect 50318 52782 50370 52834
rect 5070 52670 5122 52722
rect 5966 52670 6018 52722
rect 10110 52670 10162 52722
rect 10446 52670 10498 52722
rect 11678 52670 11730 52722
rect 16494 52670 16546 52722
rect 25230 52670 25282 52722
rect 25566 52670 25618 52722
rect 35310 52670 35362 52722
rect 36318 52670 36370 52722
rect 37662 52670 37714 52722
rect 37886 52670 37938 52722
rect 40014 52670 40066 52722
rect 41022 52670 41074 52722
rect 45726 52670 45778 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 10894 52334 10946 52386
rect 20302 52334 20354 52386
rect 33854 52334 33906 52386
rect 34302 52334 34354 52386
rect 39118 52334 39170 52386
rect 45838 52334 45890 52386
rect 4622 52248 4674 52300
rect 5070 52222 5122 52274
rect 11342 52222 11394 52274
rect 18286 52222 18338 52274
rect 22766 52222 22818 52274
rect 24446 52222 24498 52274
rect 25230 52222 25282 52274
rect 27358 52222 27410 52274
rect 28590 52222 28642 52274
rect 33406 52222 33458 52274
rect 34526 52222 34578 52274
rect 35870 52222 35922 52274
rect 38558 52222 38610 52274
rect 39566 52222 39618 52274
rect 41358 52222 41410 52274
rect 46622 52222 46674 52274
rect 1822 52110 1874 52162
rect 5630 52110 5682 52162
rect 7758 52110 7810 52162
rect 10334 52110 10386 52162
rect 10558 52110 10610 52162
rect 11566 52110 11618 52162
rect 12574 52110 12626 52162
rect 12798 52110 12850 52162
rect 12910 52110 12962 52162
rect 13582 52110 13634 52162
rect 13694 52110 13746 52162
rect 13806 52110 13858 52162
rect 14590 52110 14642 52162
rect 15486 52110 15538 52162
rect 18734 52110 18786 52162
rect 19854 52110 19906 52162
rect 23326 52110 23378 52162
rect 23998 52110 24050 52162
rect 28030 52110 28082 52162
rect 30494 52110 30546 52162
rect 33854 52110 33906 52162
rect 34862 52110 34914 52162
rect 37662 52110 37714 52162
rect 38894 52110 38946 52162
rect 39454 52110 39506 52162
rect 40238 52110 40290 52162
rect 40686 52110 40738 52162
rect 2494 51998 2546 52050
rect 5742 51998 5794 52050
rect 8318 51998 8370 52050
rect 11230 51998 11282 52050
rect 16158 51998 16210 52050
rect 19182 51998 19234 52050
rect 20302 51998 20354 52050
rect 6974 51886 7026 51938
rect 14254 51886 14306 51938
rect 14926 51886 14978 51938
rect 19070 51886 19122 51938
rect 20414 51942 20466 51994
rect 24446 51998 24498 52050
rect 31278 51998 31330 52050
rect 35982 51998 36034 52050
rect 37998 51998 38050 52050
rect 39678 52054 39730 52106
rect 41022 52110 41074 52162
rect 42030 52110 42082 52162
rect 45614 52110 45666 52162
rect 46510 52110 46562 52162
rect 46734 52110 46786 52162
rect 47742 52110 47794 52162
rect 48078 52110 48130 52162
rect 48190 52110 48242 52162
rect 50318 52110 50370 52162
rect 50542 52110 50594 52162
rect 50878 52110 50930 52162
rect 39790 51998 39842 52050
rect 41470 51998 41522 52050
rect 41694 51998 41746 52050
rect 42478 51998 42530 52050
rect 42814 51998 42866 52050
rect 43598 51998 43650 52050
rect 43710 51998 43762 52050
rect 47070 51998 47122 52050
rect 50094 51998 50146 52050
rect 51102 51998 51154 52050
rect 51214 51998 51266 52050
rect 24222 51886 24274 51938
rect 24558 51886 24610 51938
rect 34638 51886 34690 51938
rect 35534 51886 35586 51938
rect 35758 51886 35810 51938
rect 37886 51886 37938 51938
rect 38446 51886 38498 51938
rect 38670 51886 38722 51938
rect 40910 51886 40962 51938
rect 42142 51886 42194 51938
rect 43374 51886 43426 51938
rect 46174 51886 46226 51938
rect 47406 51886 47458 51938
rect 49422 51886 49474 51938
rect 49758 51886 49810 51938
rect 50318 51886 50370 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 4510 51550 4562 51602
rect 10110 51550 10162 51602
rect 16270 51550 16322 51602
rect 17726 51550 17778 51602
rect 21870 51550 21922 51602
rect 22542 51550 22594 51602
rect 34862 51550 34914 51602
rect 35982 51550 36034 51602
rect 36094 51550 36146 51602
rect 38110 51550 38162 51602
rect 38782 51550 38834 51602
rect 44942 51550 44994 51602
rect 46622 51550 46674 51602
rect 49646 51550 49698 51602
rect 11006 51438 11058 51490
rect 13246 51438 13298 51490
rect 15374 51438 15426 51490
rect 15822 51438 15874 51490
rect 17614 51438 17666 51490
rect 18174 51438 18226 51490
rect 19070 51438 19122 51490
rect 22654 51438 22706 51490
rect 23438 51438 23490 51490
rect 23774 51438 23826 51490
rect 24558 51438 24610 51490
rect 33854 51438 33906 51490
rect 34526 51438 34578 51490
rect 35534 51438 35586 51490
rect 35758 51438 35810 51490
rect 37326 51438 37378 51490
rect 39230 51438 39282 51490
rect 40126 51438 40178 51490
rect 42142 51438 42194 51490
rect 42814 51438 42866 51490
rect 43038 51438 43090 51490
rect 43822 51438 43874 51490
rect 45614 51438 45666 51490
rect 46062 51438 46114 51490
rect 47182 51438 47234 51490
rect 48078 51438 48130 51490
rect 48862 51438 48914 51490
rect 50654 51438 50706 51490
rect 53230 51438 53282 51490
rect 4398 51326 4450 51378
rect 4622 51326 4674 51378
rect 5406 51326 5458 51378
rect 10446 51326 10498 51378
rect 11342 51326 11394 51378
rect 11790 51326 11842 51378
rect 13582 51326 13634 51378
rect 13806 51326 13858 51378
rect 15262 51326 15314 51378
rect 15598 51326 15650 51378
rect 16494 51326 16546 51378
rect 16830 51326 16882 51378
rect 17950 51326 18002 51378
rect 18398 51326 18450 51378
rect 19294 51326 19346 51378
rect 19854 51326 19906 51378
rect 20190 51326 20242 51378
rect 20414 51326 20466 51378
rect 22094 51326 22146 51378
rect 23102 51326 23154 51378
rect 23998 51326 24050 51378
rect 34078 51326 34130 51378
rect 34302 51326 34354 51378
rect 36318 51326 36370 51378
rect 36542 51326 36594 51378
rect 36766 51326 36818 51378
rect 37102 51326 37154 51378
rect 37998 51326 38050 51378
rect 38558 51326 38610 51378
rect 38894 51326 38946 51378
rect 39566 51326 39618 51378
rect 41358 51326 41410 51378
rect 41582 51326 41634 51378
rect 43374 51326 43426 51378
rect 43710 51326 43762 51378
rect 45278 51326 45330 51378
rect 46510 51326 46562 51378
rect 47070 51326 47122 51378
rect 47966 51326 48018 51378
rect 49198 51326 49250 51378
rect 49422 51326 49474 51378
rect 49982 51326 50034 51378
rect 50318 51326 50370 51378
rect 50430 51326 50482 51378
rect 50766 51326 50818 51378
rect 53902 51326 53954 51378
rect 6190 51214 6242 51266
rect 8318 51214 8370 51266
rect 8766 51214 8818 51266
rect 10670 51214 10722 51266
rect 16046 51214 16098 51266
rect 18734 51214 18786 51266
rect 20078 51214 20130 51266
rect 21758 51214 21810 51266
rect 33742 51214 33794 51266
rect 36990 51214 37042 51266
rect 40238 51214 40290 51266
rect 51102 51214 51154 51266
rect 4846 51102 4898 51154
rect 11342 51102 11394 51154
rect 13358 51102 13410 51154
rect 16270 51102 16322 51154
rect 22430 51102 22482 51154
rect 24446 51102 24498 51154
rect 34974 51102 35026 51154
rect 35198 51102 35250 51154
rect 38110 51102 38162 51154
rect 39454 51102 39506 51154
rect 39902 51102 39954 51154
rect 41918 51102 41970 51154
rect 43822 51102 43874 51154
rect 48078 51102 48130 51154
rect 48750 51102 48802 51154
rect 49758 51102 49810 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 5742 50766 5794 50818
rect 6526 50766 6578 50818
rect 6638 50766 6690 50818
rect 11566 50766 11618 50818
rect 11790 50766 11842 50818
rect 12126 50766 12178 50818
rect 12574 50766 12626 50818
rect 33630 50766 33682 50818
rect 36318 50766 36370 50818
rect 38222 50766 38274 50818
rect 42590 50766 42642 50818
rect 7534 50654 7586 50706
rect 11006 50654 11058 50706
rect 12350 50654 12402 50706
rect 14702 50654 14754 50706
rect 18958 50654 19010 50706
rect 19966 50654 20018 50706
rect 22542 50654 22594 50706
rect 23550 50654 23602 50706
rect 24110 50654 24162 50706
rect 27470 50654 27522 50706
rect 32062 50654 32114 50706
rect 36430 50654 36482 50706
rect 40798 50654 40850 50706
rect 42478 50654 42530 50706
rect 45502 50654 45554 50706
rect 48302 50654 48354 50706
rect 50318 50654 50370 50706
rect 51662 50654 51714 50706
rect 52110 50654 52162 50706
rect 55582 50654 55634 50706
rect 5966 50542 6018 50594
rect 6190 50542 6242 50594
rect 6862 50542 6914 50594
rect 7086 50542 7138 50594
rect 8094 50542 8146 50594
rect 11342 50542 11394 50594
rect 12798 50542 12850 50594
rect 13470 50542 13522 50594
rect 15374 50542 15426 50594
rect 18174 50542 18226 50594
rect 19294 50542 19346 50594
rect 19742 50542 19794 50594
rect 20190 50542 20242 50594
rect 20414 50542 20466 50594
rect 23102 50542 23154 50594
rect 23326 50542 23378 50594
rect 23774 50542 23826 50594
rect 27022 50542 27074 50594
rect 29150 50542 29202 50594
rect 33518 50542 33570 50594
rect 33742 50542 33794 50594
rect 34190 50542 34242 50594
rect 34750 50542 34802 50594
rect 35198 50542 35250 50594
rect 35758 50542 35810 50594
rect 36990 50542 37042 50594
rect 37550 50542 37602 50594
rect 38334 50542 38386 50594
rect 38670 50542 38722 50594
rect 39006 50542 39058 50594
rect 40462 50542 40514 50594
rect 41134 50542 41186 50594
rect 42254 50542 42306 50594
rect 43262 50542 43314 50594
rect 47294 50542 47346 50594
rect 48190 50542 48242 50594
rect 48414 50542 48466 50594
rect 48862 50542 48914 50594
rect 50766 50542 50818 50594
rect 52670 50542 52722 50594
rect 5630 50430 5682 50482
rect 8878 50430 8930 50482
rect 11902 50430 11954 50482
rect 12910 50430 12962 50482
rect 14926 50430 14978 50482
rect 15934 50430 15986 50482
rect 18398 50430 18450 50482
rect 19070 50430 19122 50482
rect 22206 50430 22258 50482
rect 22878 50430 22930 50482
rect 26238 50430 26290 50482
rect 27806 50430 27858 50482
rect 27918 50430 27970 50482
rect 28478 50430 28530 50482
rect 28590 50430 28642 50482
rect 29934 50430 29986 50482
rect 33966 50430 34018 50482
rect 34414 50430 34466 50482
rect 35870 50430 35922 50482
rect 38446 50430 38498 50482
rect 38894 50430 38946 50482
rect 39902 50430 39954 50482
rect 40126 50430 40178 50482
rect 41022 50430 41074 50482
rect 41582 50430 41634 50482
rect 42926 50430 42978 50482
rect 43598 50430 43650 50482
rect 43934 50430 43986 50482
rect 49646 50430 49698 50482
rect 49870 50430 49922 50482
rect 51214 50430 51266 50482
rect 53454 50430 53506 50482
rect 7422 50318 7474 50370
rect 18510 50318 18562 50370
rect 22430 50318 22482 50370
rect 23886 50318 23938 50370
rect 28142 50318 28194 50370
rect 28254 50318 28306 50370
rect 32510 50318 32562 50370
rect 39454 50318 39506 50370
rect 41358 50318 41410 50370
rect 44942 50318 44994 50370
rect 49758 50318 49810 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 6078 49982 6130 50034
rect 7198 49982 7250 50034
rect 16158 49982 16210 50034
rect 17950 49982 18002 50034
rect 18286 49982 18338 50034
rect 23214 49982 23266 50034
rect 24110 49982 24162 50034
rect 35982 49982 36034 50034
rect 36094 49982 36146 50034
rect 36318 49982 36370 50034
rect 37662 49982 37714 50034
rect 42478 49982 42530 50034
rect 43598 49982 43650 50034
rect 51550 49982 51602 50034
rect 51998 49982 52050 50034
rect 52222 49982 52274 50034
rect 2494 49870 2546 49922
rect 6414 49870 6466 49922
rect 6638 49870 6690 49922
rect 7310 49870 7362 49922
rect 11902 49870 11954 49922
rect 15934 49870 15986 49922
rect 17390 49870 17442 49922
rect 18734 49870 18786 49922
rect 20750 49870 20802 49922
rect 31166 49870 31218 49922
rect 31502 49870 31554 49922
rect 31838 49870 31890 49922
rect 35422 49870 35474 49922
rect 36542 49870 36594 49922
rect 36878 49870 36930 49922
rect 37102 49870 37154 49922
rect 37998 49870 38050 49922
rect 40014 49870 40066 49922
rect 43038 49870 43090 49922
rect 43822 49870 43874 49922
rect 43934 49870 43986 49922
rect 48750 49870 48802 49922
rect 50766 49870 50818 49922
rect 51886 49870 51938 49922
rect 1822 49758 1874 49810
rect 5742 49758 5794 49810
rect 7086 49758 7138 49810
rect 10894 49758 10946 49810
rect 12126 49758 12178 49810
rect 13358 49758 13410 49810
rect 13694 49758 13746 49810
rect 14142 49758 14194 49810
rect 14366 49758 14418 49810
rect 15038 49758 15090 49810
rect 16382 49758 16434 49810
rect 17614 49758 17666 49810
rect 18510 49758 18562 49810
rect 19182 49758 19234 49810
rect 19518 49758 19570 49810
rect 19854 49758 19906 49810
rect 20302 49758 20354 49810
rect 20862 49758 20914 49810
rect 22878 49758 22930 49810
rect 23214 49758 23266 49810
rect 23550 49758 23602 49810
rect 23998 49758 24050 49810
rect 24222 49758 24274 49810
rect 24558 49758 24610 49810
rect 27470 49758 27522 49810
rect 30942 49758 30994 49810
rect 35646 49758 35698 49810
rect 37438 49758 37490 49810
rect 38782 49758 38834 49810
rect 39230 49758 39282 49810
rect 39902 49758 39954 49810
rect 41470 49758 41522 49810
rect 42366 49758 42418 49810
rect 42590 49758 42642 49810
rect 43150 49758 43202 49810
rect 43374 49758 43426 49810
rect 47070 49758 47122 49810
rect 48974 49758 49026 49810
rect 49870 49758 49922 49810
rect 50990 49758 51042 49810
rect 51214 49758 51266 49810
rect 51326 49758 51378 49810
rect 4622 49646 4674 49698
rect 5070 49646 5122 49698
rect 5518 49646 5570 49698
rect 6526 49646 6578 49698
rect 11342 49646 11394 49698
rect 12462 49646 12514 49698
rect 13806 49646 13858 49698
rect 19406 49646 19458 49698
rect 23326 49646 23378 49698
rect 27022 49646 27074 49698
rect 28142 49646 28194 49698
rect 30270 49646 30322 49698
rect 32286 49646 32338 49698
rect 33182 49646 33234 49698
rect 37214 49646 37266 49698
rect 40910 49646 40962 49698
rect 44606 49646 44658 49698
rect 45390 49646 45442 49698
rect 49086 49646 49138 49698
rect 49982 49646 50034 49698
rect 14590 49534 14642 49586
rect 14814 49534 14866 49586
rect 15486 49534 15538 49586
rect 15822 49534 15874 49586
rect 18174 49534 18226 49586
rect 20526 49534 20578 49586
rect 21086 49534 21138 49586
rect 30606 49534 30658 49586
rect 39790 49534 39842 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 6302 49198 6354 49250
rect 21870 49198 21922 49250
rect 35982 49198 36034 49250
rect 42142 49198 42194 49250
rect 42926 49198 42978 49250
rect 7870 49086 7922 49138
rect 11342 49086 11394 49138
rect 16718 49086 16770 49138
rect 19966 49086 20018 49138
rect 22766 49086 22818 49138
rect 23774 49086 23826 49138
rect 24334 49086 24386 49138
rect 26014 49086 26066 49138
rect 26798 49086 26850 49138
rect 29598 49086 29650 49138
rect 31166 49086 31218 49138
rect 39566 49086 39618 49138
rect 47742 49086 47794 49138
rect 48302 49086 48354 49138
rect 50990 49086 51042 49138
rect 6078 48974 6130 49026
rect 7198 48974 7250 49026
rect 12686 48974 12738 49026
rect 13470 48974 13522 49026
rect 16606 48974 16658 49026
rect 17166 48974 17218 49026
rect 21310 48974 21362 49026
rect 21534 48974 21586 49026
rect 23102 48974 23154 49026
rect 23214 48974 23266 49026
rect 23886 48974 23938 49026
rect 27358 48974 27410 49026
rect 27582 48974 27634 49026
rect 28478 48974 28530 49026
rect 29038 48974 29090 49026
rect 29486 48974 29538 49026
rect 34078 48974 34130 49026
rect 36094 48974 36146 49026
rect 39342 48974 39394 49026
rect 40798 48974 40850 49026
rect 41470 48974 41522 49026
rect 43262 48974 43314 49026
rect 43710 48974 43762 49026
rect 44942 48974 44994 49026
rect 49310 48974 49362 49026
rect 50654 48974 50706 49026
rect 12798 48862 12850 48914
rect 14142 48862 14194 48914
rect 15150 48862 15202 48914
rect 17838 48862 17890 48914
rect 20302 48862 20354 48914
rect 20638 48862 20690 48914
rect 22766 48862 22818 48914
rect 26686 48862 26738 48914
rect 27246 48862 27298 48914
rect 30046 48862 30098 48914
rect 30830 48862 30882 48914
rect 33294 48862 33346 48914
rect 35982 48862 36034 48914
rect 40126 48862 40178 48914
rect 40686 48862 40738 48914
rect 41134 48862 41186 48914
rect 41806 48862 41858 48914
rect 44046 48862 44098 48914
rect 45614 48862 45666 48914
rect 50318 48862 50370 48914
rect 50878 48862 50930 48914
rect 6638 48750 6690 48802
rect 6974 48750 7026 48802
rect 13022 48750 13074 48802
rect 22542 48750 22594 48802
rect 23662 48750 23714 48802
rect 25566 48750 25618 48802
rect 26462 48750 26514 48802
rect 26910 48750 26962 48802
rect 29710 48750 29762 48802
rect 30382 48750 30434 48802
rect 30718 48750 30770 48802
rect 34526 48750 34578 48802
rect 39006 48750 39058 48802
rect 42030 48750 42082 48802
rect 49086 48750 49138 48802
rect 49646 48750 49698 48802
rect 49982 48750 50034 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 2830 48414 2882 48466
rect 17614 48414 17666 48466
rect 19518 48414 19570 48466
rect 19966 48414 20018 48466
rect 20190 48414 20242 48466
rect 20974 48414 21026 48466
rect 22990 48414 23042 48466
rect 23214 48414 23266 48466
rect 26350 48414 26402 48466
rect 27470 48414 27522 48466
rect 27582 48414 27634 48466
rect 28702 48414 28754 48466
rect 28814 48414 28866 48466
rect 39230 48414 39282 48466
rect 39678 48414 39730 48466
rect 40014 48414 40066 48466
rect 45838 48414 45890 48466
rect 49534 48414 49586 48466
rect 12126 48302 12178 48354
rect 14142 48302 14194 48354
rect 15598 48302 15650 48354
rect 17726 48302 17778 48354
rect 18846 48302 18898 48354
rect 19182 48302 19234 48354
rect 20414 48302 20466 48354
rect 20526 48302 20578 48354
rect 23438 48302 23490 48354
rect 24670 48302 24722 48354
rect 26686 48302 26738 48354
rect 27134 48302 27186 48354
rect 30606 48302 30658 48354
rect 31838 48302 31890 48354
rect 39342 48302 39394 48354
rect 44494 48302 44546 48354
rect 46398 48302 46450 48354
rect 47854 48302 47906 48354
rect 7646 48190 7698 48242
rect 8318 48190 8370 48242
rect 8430 48190 8482 48242
rect 10222 48190 10274 48242
rect 10894 48190 10946 48242
rect 11342 48190 11394 48242
rect 12350 48190 12402 48242
rect 14702 48190 14754 48242
rect 16830 48190 16882 48242
rect 17278 48190 17330 48242
rect 17950 48190 18002 48242
rect 18622 48190 18674 48242
rect 19854 48190 19906 48242
rect 23550 48190 23602 48242
rect 24334 48190 24386 48242
rect 25790 48190 25842 48242
rect 26014 48190 26066 48242
rect 27358 48190 27410 48242
rect 27694 48190 27746 48242
rect 28926 48190 28978 48242
rect 29038 48190 29090 48242
rect 29374 48190 29426 48242
rect 30046 48190 30098 48242
rect 30382 48190 30434 48242
rect 31390 48190 31442 48242
rect 32062 48190 32114 48242
rect 33406 48190 33458 48242
rect 46062 48190 46114 48242
rect 46622 48190 46674 48242
rect 47070 48190 47122 48242
rect 47182 48190 47234 48242
rect 47630 48190 47682 48242
rect 48078 48190 48130 48242
rect 50094 48190 50146 48242
rect 50542 48190 50594 48242
rect 2942 48078 2994 48130
rect 4734 48078 4786 48130
rect 6862 48078 6914 48130
rect 8094 48078 8146 48130
rect 10670 48078 10722 48130
rect 11678 48078 11730 48130
rect 15486 48078 15538 48130
rect 22430 48078 22482 48130
rect 28142 48078 28194 48130
rect 28254 48078 28306 48130
rect 30942 48078 30994 48130
rect 34190 48078 34242 48130
rect 36318 48078 36370 48130
rect 46174 48078 46226 48130
rect 47406 48078 47458 48130
rect 49198 48078 49250 48130
rect 51326 48078 51378 48130
rect 53454 48078 53506 48130
rect 3054 47966 3106 48018
rect 7982 47966 8034 48018
rect 9662 47966 9714 48018
rect 9774 47966 9826 48018
rect 9998 47966 10050 48018
rect 10558 47966 10610 48018
rect 12686 47966 12738 48018
rect 22654 47966 22706 48018
rect 24334 47966 24386 48018
rect 25454 47966 25506 48018
rect 29598 47966 29650 48018
rect 30270 47966 30322 48018
rect 49086 47966 49138 48018
rect 49310 47966 49362 48018
rect 49870 47966 49922 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 19966 47630 20018 47682
rect 29262 47630 29314 47682
rect 50430 47630 50482 47682
rect 50542 47630 50594 47682
rect 50878 47630 50930 47682
rect 1710 47518 1762 47570
rect 3838 47518 3890 47570
rect 8990 47518 9042 47570
rect 11118 47518 11170 47570
rect 12238 47518 12290 47570
rect 18622 47518 18674 47570
rect 23886 47518 23938 47570
rect 32398 47518 32450 47570
rect 33966 47518 34018 47570
rect 34750 47518 34802 47570
rect 34862 47518 34914 47570
rect 44270 47518 44322 47570
rect 44830 47518 44882 47570
rect 45166 47518 45218 47570
rect 47966 47518 48018 47570
rect 48526 47518 48578 47570
rect 48862 47518 48914 47570
rect 49086 47518 49138 47570
rect 4622 47406 4674 47458
rect 6078 47406 6130 47458
rect 7086 47406 7138 47458
rect 8206 47406 8258 47458
rect 11678 47406 11730 47458
rect 12686 47406 12738 47458
rect 13806 47406 13858 47458
rect 15934 47406 15986 47458
rect 18174 47406 18226 47458
rect 20190 47406 20242 47458
rect 6190 47294 6242 47346
rect 7646 47294 7698 47346
rect 13918 47294 13970 47346
rect 16382 47294 16434 47346
rect 20526 47350 20578 47402
rect 22318 47406 22370 47458
rect 22654 47406 22706 47458
rect 24110 47406 24162 47458
rect 27582 47406 27634 47458
rect 27918 47406 27970 47458
rect 28254 47406 28306 47458
rect 33182 47406 33234 47458
rect 33742 47406 33794 47458
rect 35086 47406 35138 47458
rect 41358 47406 41410 47458
rect 45502 47406 45554 47458
rect 45838 47406 45890 47458
rect 46174 47406 46226 47458
rect 46398 47406 46450 47458
rect 47294 47406 47346 47458
rect 47518 47406 47570 47458
rect 50766 47406 50818 47458
rect 22094 47294 22146 47346
rect 29150 47294 29202 47346
rect 29262 47294 29314 47346
rect 34190 47294 34242 47346
rect 34414 47294 34466 47346
rect 42142 47294 42194 47346
rect 46622 47294 46674 47346
rect 48302 47294 48354 47346
rect 5070 47182 5122 47234
rect 6302 47182 6354 47234
rect 11454 47182 11506 47234
rect 12350 47182 12402 47234
rect 12798 47182 12850 47234
rect 13022 47182 13074 47234
rect 15262 47182 15314 47234
rect 19182 47182 19234 47234
rect 19630 47182 19682 47234
rect 20638 47182 20690 47234
rect 20862 47182 20914 47234
rect 22318 47182 22370 47234
rect 24446 47182 24498 47234
rect 24670 47182 24722 47234
rect 24782 47182 24834 47234
rect 25006 47182 25058 47234
rect 25342 47182 25394 47234
rect 25790 47182 25842 47234
rect 26126 47182 26178 47234
rect 26574 47182 26626 47234
rect 27134 47182 27186 47234
rect 27806 47182 27858 47234
rect 35646 47182 35698 47234
rect 45054 47182 45106 47234
rect 45614 47182 45666 47234
rect 46510 47182 46562 47234
rect 49646 47182 49698 47234
rect 49982 47182 50034 47234
rect 51326 47182 51378 47234
rect 51774 47182 51826 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 4286 46846 4338 46898
rect 9886 46846 9938 46898
rect 16382 46846 16434 46898
rect 26798 46846 26850 46898
rect 27582 46846 27634 46898
rect 28254 46846 28306 46898
rect 28702 46846 28754 46898
rect 30830 46846 30882 46898
rect 31390 46846 31442 46898
rect 48078 46846 48130 46898
rect 50206 46846 50258 46898
rect 2158 46734 2210 46786
rect 2270 46734 2322 46786
rect 2606 46734 2658 46786
rect 4510 46734 4562 46786
rect 6302 46734 6354 46786
rect 12910 46734 12962 46786
rect 14366 46734 14418 46786
rect 15710 46734 15762 46786
rect 18734 46734 18786 46786
rect 22542 46734 22594 46786
rect 23886 46734 23938 46786
rect 27022 46734 27074 46786
rect 28814 46734 28866 46786
rect 29486 46734 29538 46786
rect 30046 46734 30098 46786
rect 30718 46734 30770 46786
rect 31726 46734 31778 46786
rect 32062 46734 32114 46786
rect 41134 46734 41186 46786
rect 46734 46734 46786 46786
rect 2718 46622 2770 46674
rect 3054 46622 3106 46674
rect 3950 46622 4002 46674
rect 4174 46622 4226 46674
rect 6638 46622 6690 46674
rect 10222 46622 10274 46674
rect 11678 46622 11730 46674
rect 12014 46622 12066 46674
rect 12686 46622 12738 46674
rect 13470 46622 13522 46674
rect 14030 46622 14082 46674
rect 14478 46622 14530 46674
rect 15038 46622 15090 46674
rect 15822 46622 15874 46674
rect 16270 46622 16322 46674
rect 19406 46622 19458 46674
rect 20078 46622 20130 46674
rect 20750 46622 20802 46674
rect 21198 46622 21250 46674
rect 22318 46622 22370 46674
rect 23214 46622 23266 46674
rect 25678 46622 25730 46674
rect 26462 46622 26514 46674
rect 27358 46622 27410 46674
rect 28478 46622 28530 46674
rect 29262 46622 29314 46674
rect 30606 46622 30658 46674
rect 31166 46622 31218 46674
rect 32174 46622 32226 46674
rect 33070 46622 33122 46674
rect 35870 46622 35922 46674
rect 40350 46622 40402 46674
rect 44942 46622 44994 46674
rect 45614 46622 45666 46674
rect 46622 46622 46674 46674
rect 46846 46622 46898 46674
rect 47294 46622 47346 46674
rect 47966 46622 48018 46674
rect 48078 46622 48130 46674
rect 48862 46622 48914 46674
rect 49086 46622 49138 46674
rect 49758 46622 49810 46674
rect 50094 46622 50146 46674
rect 50542 46622 50594 46674
rect 51774 46622 51826 46674
rect 51886 46622 51938 46674
rect 10446 46510 10498 46562
rect 11230 46510 11282 46562
rect 11902 46510 11954 46562
rect 14254 46510 14306 46562
rect 17390 46510 17442 46562
rect 17614 46510 17666 46562
rect 19518 46510 19570 46562
rect 22542 46510 22594 46562
rect 22990 46510 23042 46562
rect 24446 46510 24498 46562
rect 25342 46510 25394 46562
rect 26238 46510 26290 46562
rect 28142 46510 28194 46562
rect 29822 46510 29874 46562
rect 33518 46510 33570 46562
rect 34078 46510 34130 46562
rect 34526 46510 34578 46562
rect 35646 46510 35698 46562
rect 36654 46510 36706 46562
rect 38782 46510 38834 46562
rect 44382 46510 44434 46562
rect 45278 46510 45330 46562
rect 2158 46398 2210 46450
rect 11566 46398 11618 46450
rect 16382 46398 16434 46450
rect 17950 46398 18002 46450
rect 27134 46398 27186 46450
rect 27694 46398 27746 46450
rect 30158 46398 30210 46450
rect 40910 46398 40962 46450
rect 41246 46398 41298 46450
rect 44606 46398 44658 46450
rect 45390 46398 45442 46450
rect 45726 46398 45778 46450
rect 47742 46398 47794 46450
rect 50318 46398 50370 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 7758 46062 7810 46114
rect 15150 46062 15202 46114
rect 26126 46062 26178 46114
rect 31278 46062 31330 46114
rect 1710 45950 1762 46002
rect 3838 45950 3890 46002
rect 11902 45950 11954 46002
rect 14254 45950 14306 46002
rect 18398 45950 18450 46002
rect 19406 45950 19458 46002
rect 22206 45950 22258 46002
rect 24334 45950 24386 46002
rect 26462 45950 26514 46002
rect 29374 45950 29426 46002
rect 31614 45950 31666 46002
rect 34750 45950 34802 46002
rect 38894 45950 38946 46002
rect 39678 45950 39730 46002
rect 41806 45950 41858 46002
rect 46174 45950 46226 46002
rect 48302 45950 48354 46002
rect 4622 45838 4674 45890
rect 5742 45838 5794 45890
rect 6526 45838 6578 45890
rect 6974 45838 7026 45890
rect 12574 45838 12626 45890
rect 13694 45838 13746 45890
rect 14590 45838 14642 45890
rect 14814 45838 14866 45890
rect 18174 45838 18226 45890
rect 19070 45838 19122 45890
rect 20190 45838 20242 45890
rect 20750 45838 20802 45890
rect 22430 45838 22482 45890
rect 23550 45838 23602 45890
rect 24110 45838 24162 45890
rect 24558 45838 24610 45890
rect 26686 45838 26738 45890
rect 27134 45838 27186 45890
rect 27358 45838 27410 45890
rect 27806 45838 27858 45890
rect 29486 45838 29538 45890
rect 30046 45838 30098 45890
rect 30382 45838 30434 45890
rect 33070 45838 33122 45890
rect 35534 45838 35586 45890
rect 38670 45838 38722 45890
rect 42590 45838 42642 45890
rect 43038 45838 43090 45890
rect 45502 45838 45554 45890
rect 49086 45838 49138 45890
rect 5630 45726 5682 45778
rect 7198 45726 7250 45778
rect 7534 45726 7586 45778
rect 9774 45726 9826 45778
rect 11454 45726 11506 45778
rect 12910 45726 12962 45778
rect 15710 45726 15762 45778
rect 26350 45726 26402 45778
rect 31502 45726 31554 45778
rect 39342 45726 39394 45778
rect 45726 45726 45778 45778
rect 5070 45614 5122 45666
rect 7646 45614 7698 45666
rect 10110 45614 10162 45666
rect 11118 45614 11170 45666
rect 11342 45614 11394 45666
rect 11790 45614 11842 45666
rect 15038 45614 15090 45666
rect 15822 45614 15874 45666
rect 16046 45614 16098 45666
rect 27246 45614 27298 45666
rect 27694 45614 27746 45666
rect 28366 45614 28418 45666
rect 45054 45614 45106 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 5406 45278 5458 45330
rect 9662 45278 9714 45330
rect 12350 45278 12402 45330
rect 13918 45278 13970 45330
rect 14254 45278 14306 45330
rect 14478 45278 14530 45330
rect 14814 45278 14866 45330
rect 28366 45278 28418 45330
rect 38334 45278 38386 45330
rect 44942 45278 44994 45330
rect 49198 45278 49250 45330
rect 2830 45166 2882 45218
rect 4286 45166 4338 45218
rect 14702 45166 14754 45218
rect 16494 45166 16546 45218
rect 17614 45166 17666 45218
rect 18958 45166 19010 45218
rect 19406 45166 19458 45218
rect 21758 45166 21810 45218
rect 22766 45166 22818 45218
rect 24558 45166 24610 45218
rect 25230 45166 25282 45218
rect 26798 45166 26850 45218
rect 29598 45166 29650 45218
rect 30606 45166 30658 45218
rect 31950 45166 32002 45218
rect 33966 45166 34018 45218
rect 35198 45166 35250 45218
rect 37998 45166 38050 45218
rect 40350 45166 40402 45218
rect 50318 45166 50370 45218
rect 1710 45054 1762 45106
rect 3726 45054 3778 45106
rect 5966 45054 6018 45106
rect 10446 45054 10498 45106
rect 10782 45054 10834 45106
rect 12014 45054 12066 45106
rect 14142 45054 14194 45106
rect 16718 45054 16770 45106
rect 17390 45054 17442 45106
rect 19070 45054 19122 45106
rect 19742 45054 19794 45106
rect 20078 45054 20130 45106
rect 20302 45054 20354 45106
rect 20974 45054 21026 45106
rect 21198 45054 21250 45106
rect 24334 45054 24386 45106
rect 25566 45054 25618 45106
rect 26014 45054 26066 45106
rect 27134 45054 27186 45106
rect 27470 45054 27522 45106
rect 27694 45054 27746 45106
rect 27918 45054 27970 45106
rect 28590 45054 28642 45106
rect 29262 45054 29314 45106
rect 31054 45054 31106 45106
rect 31390 45054 31442 45106
rect 32286 45054 32338 45106
rect 33182 45054 33234 45106
rect 33518 45054 33570 45106
rect 33742 45054 33794 45106
rect 34190 45054 34242 45106
rect 34526 45054 34578 45106
rect 39678 45054 39730 45106
rect 41470 45054 41522 45106
rect 49534 45054 49586 45106
rect 6638 44942 6690 44994
rect 8766 44942 8818 44994
rect 10558 44942 10610 44994
rect 11790 44942 11842 44994
rect 15374 44942 15426 44994
rect 15934 44942 15986 44994
rect 18062 44942 18114 44994
rect 26350 44942 26402 44994
rect 27246 44942 27298 44994
rect 28142 44942 28194 44994
rect 28478 44942 28530 44994
rect 29374 44942 29426 44994
rect 31166 44942 31218 44994
rect 32062 44942 32114 44994
rect 37326 44942 37378 44994
rect 40014 44942 40066 44994
rect 41134 44942 41186 44994
rect 42142 44942 42194 44994
rect 44382 44942 44434 44994
rect 52446 44942 52498 44994
rect 10222 44830 10274 44882
rect 15374 44830 15426 44882
rect 15934 44830 15986 44882
rect 18958 44830 19010 44882
rect 20526 44830 20578 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 2046 44494 2098 44546
rect 3278 44494 3330 44546
rect 6190 44494 6242 44546
rect 6526 44494 6578 44546
rect 17278 44494 17330 44546
rect 23102 44494 23154 44546
rect 23326 44494 23378 44546
rect 30046 44494 30098 44546
rect 34414 44494 34466 44546
rect 2494 44382 2546 44434
rect 4622 44382 4674 44434
rect 7646 44382 7698 44434
rect 11006 44382 11058 44434
rect 12686 44382 12738 44434
rect 14030 44382 14082 44434
rect 17390 44382 17442 44434
rect 23550 44382 23602 44434
rect 23886 44382 23938 44434
rect 30942 44382 30994 44434
rect 32622 44382 32674 44434
rect 33630 44382 33682 44434
rect 42366 44382 42418 44434
rect 44830 44382 44882 44434
rect 48190 44382 48242 44434
rect 2382 44270 2434 44322
rect 2606 44270 2658 44322
rect 3054 44270 3106 44322
rect 3614 44270 3666 44322
rect 3838 44270 3890 44322
rect 4174 44270 4226 44322
rect 4398 44270 4450 44322
rect 6302 44270 6354 44322
rect 6750 44270 6802 44322
rect 7086 44270 7138 44322
rect 7422 44270 7474 44322
rect 8206 44270 8258 44322
rect 11902 44270 11954 44322
rect 13582 44270 13634 44322
rect 13806 44270 13858 44322
rect 14254 44270 14306 44322
rect 14478 44270 14530 44322
rect 15038 44270 15090 44322
rect 15262 44270 15314 44322
rect 16382 44270 16434 44322
rect 16606 44270 16658 44322
rect 16830 44270 16882 44322
rect 17502 44270 17554 44322
rect 18062 44270 18114 44322
rect 18734 44270 18786 44322
rect 19294 44270 19346 44322
rect 19518 44270 19570 44322
rect 19630 44270 19682 44322
rect 20414 44270 20466 44322
rect 21534 44270 21586 44322
rect 22094 44270 22146 44322
rect 22542 44270 22594 44322
rect 23998 44270 24050 44322
rect 24446 44270 24498 44322
rect 25006 44270 25058 44322
rect 25790 44270 25842 44322
rect 26574 44270 26626 44322
rect 26910 44270 26962 44322
rect 29374 44270 29426 44322
rect 29710 44270 29762 44322
rect 29934 44270 29986 44322
rect 30606 44270 30658 44322
rect 30830 44270 30882 44322
rect 31166 44270 31218 44322
rect 31838 44270 31890 44322
rect 33406 44270 33458 44322
rect 38558 44270 38610 44322
rect 39454 44270 39506 44322
rect 39902 44270 39954 44322
rect 40126 44270 40178 44322
rect 40462 44270 40514 44322
rect 40798 44270 40850 44322
rect 41358 44270 41410 44322
rect 41694 44270 41746 44322
rect 42142 44270 42194 44322
rect 42478 44270 42530 44322
rect 42702 44270 42754 44322
rect 47630 44270 47682 44322
rect 1934 44158 1986 44210
rect 4734 44158 4786 44210
rect 5742 44158 5794 44210
rect 5854 44158 5906 44210
rect 8878 44158 8930 44210
rect 12350 44158 12402 44210
rect 12574 44158 12626 44210
rect 15598 44158 15650 44210
rect 16158 44158 16210 44210
rect 17726 44158 17778 44210
rect 25454 44158 25506 44210
rect 27358 44158 27410 44210
rect 31614 44158 31666 44210
rect 32286 44158 32338 44210
rect 33182 44158 33234 44210
rect 33630 44158 33682 44210
rect 34638 44158 34690 44210
rect 38334 44158 38386 44210
rect 41806 44158 41858 44210
rect 46958 44158 47010 44210
rect 11566 44046 11618 44098
rect 13694 44046 13746 44098
rect 14702 44046 14754 44098
rect 14926 44046 14978 44098
rect 15486 44046 15538 44098
rect 20750 44046 20802 44098
rect 22766 44046 22818 44098
rect 23774 44046 23826 44098
rect 24782 44046 24834 44098
rect 24894 44046 24946 44098
rect 27134 44046 27186 44098
rect 27806 44046 27858 44098
rect 28590 44046 28642 44098
rect 29038 44046 29090 44098
rect 29150 44046 29202 44098
rect 30382 44046 30434 44098
rect 31390 44046 31442 44098
rect 32510 44046 32562 44098
rect 33742 44046 33794 44098
rect 34526 44046 34578 44098
rect 37550 44046 37602 44098
rect 40910 44046 40962 44098
rect 41022 44046 41074 44098
rect 41918 44046 41970 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 12126 43710 12178 43762
rect 15710 43710 15762 43762
rect 21758 43710 21810 43762
rect 24334 43710 24386 43762
rect 27582 43710 27634 43762
rect 29262 43710 29314 43762
rect 34190 43710 34242 43762
rect 48190 43710 48242 43762
rect 3838 43598 3890 43650
rect 5070 43598 5122 43650
rect 5182 43598 5234 43650
rect 5630 43598 5682 43650
rect 10110 43598 10162 43650
rect 11118 43598 11170 43650
rect 11678 43598 11730 43650
rect 12350 43598 12402 43650
rect 14814 43598 14866 43650
rect 17614 43598 17666 43650
rect 17726 43598 17778 43650
rect 20862 43598 20914 43650
rect 23102 43598 23154 43650
rect 24222 43598 24274 43650
rect 25342 43598 25394 43650
rect 26350 43598 26402 43650
rect 28030 43598 28082 43650
rect 28254 43598 28306 43650
rect 29598 43598 29650 43650
rect 33406 43598 33458 43650
rect 33966 43598 34018 43650
rect 35646 43598 35698 43650
rect 39006 43598 39058 43650
rect 39230 43598 39282 43650
rect 39678 43598 39730 43650
rect 40238 43598 40290 43650
rect 46510 43598 46562 43650
rect 47070 43598 47122 43650
rect 52110 43598 52162 43650
rect 4622 43486 4674 43538
rect 5966 43486 6018 43538
rect 6862 43486 6914 43538
rect 10446 43486 10498 43538
rect 10670 43486 10722 43538
rect 11230 43486 11282 43538
rect 12798 43486 12850 43538
rect 13022 43486 13074 43538
rect 13806 43486 13858 43538
rect 14030 43486 14082 43538
rect 14254 43486 14306 43538
rect 15150 43486 15202 43538
rect 16158 43486 16210 43538
rect 16606 43486 16658 43538
rect 17950 43486 18002 43538
rect 18286 43486 18338 43538
rect 19070 43486 19122 43538
rect 19854 43486 19906 43538
rect 21646 43486 21698 43538
rect 23438 43486 23490 43538
rect 23774 43486 23826 43538
rect 24446 43486 24498 43538
rect 25678 43486 25730 43538
rect 26126 43486 26178 43538
rect 27022 43486 27074 43538
rect 27806 43486 27858 43538
rect 28478 43486 28530 43538
rect 29822 43486 29874 43538
rect 30606 43486 30658 43538
rect 31278 43486 31330 43538
rect 31726 43486 31778 43538
rect 33070 43486 33122 43538
rect 33854 43486 33906 43538
rect 34862 43486 34914 43538
rect 38894 43486 38946 43538
rect 39454 43486 39506 43538
rect 40350 43486 40402 43538
rect 40798 43486 40850 43538
rect 41582 43486 41634 43538
rect 44942 43486 44994 43538
rect 45614 43486 45666 43538
rect 45950 43486 46002 43538
rect 48862 43486 48914 43538
rect 51998 43486 52050 43538
rect 1710 43374 1762 43426
rect 4958 43374 5010 43426
rect 8206 43374 8258 43426
rect 9886 43374 9938 43426
rect 12238 43374 12290 43426
rect 12910 43374 12962 43426
rect 13246 43374 13298 43426
rect 16830 43374 16882 43426
rect 19518 43374 19570 43426
rect 23326 43374 23378 43426
rect 34526 43374 34578 43426
rect 37774 43374 37826 43426
rect 41806 43374 41858 43426
rect 44718 43374 44770 43426
rect 47518 43374 47570 43426
rect 49534 43374 49586 43426
rect 51662 43374 51714 43426
rect 10222 43262 10274 43314
rect 11118 43262 11170 43314
rect 13470 43262 13522 43314
rect 14366 43262 14418 43314
rect 16382 43262 16434 43314
rect 28366 43262 28418 43314
rect 30942 43262 30994 43314
rect 39790 43262 39842 43314
rect 40238 43262 40290 43314
rect 41918 43262 41970 43314
rect 46174 43262 46226 43314
rect 46398 43262 46450 43314
rect 52110 43262 52162 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 3614 42926 3666 42978
rect 11790 42926 11842 42978
rect 14366 42926 14418 42978
rect 15038 42926 15090 42978
rect 16382 42926 16434 42978
rect 18174 42926 18226 42978
rect 18510 42926 18562 42978
rect 19182 42926 19234 42978
rect 27806 42926 27858 42978
rect 34302 42926 34354 42978
rect 52782 42926 52834 42978
rect 4174 42814 4226 42866
rect 5742 42814 5794 42866
rect 8878 42814 8930 42866
rect 11006 42814 11058 42866
rect 11566 42814 11618 42866
rect 13694 42814 13746 42866
rect 15038 42814 15090 42866
rect 15710 42814 15762 42866
rect 18622 42814 18674 42866
rect 22990 42814 23042 42866
rect 27358 42814 27410 42866
rect 29598 42814 29650 42866
rect 35422 42814 35474 42866
rect 50542 42814 50594 42866
rect 3950 42702 4002 42754
rect 8206 42702 8258 42754
rect 12798 42702 12850 42754
rect 13582 42702 13634 42754
rect 14254 42702 14306 42754
rect 21310 42702 21362 42754
rect 21870 42702 21922 42754
rect 22878 42702 22930 42754
rect 23102 42702 23154 42754
rect 23886 42702 23938 42754
rect 24334 42702 24386 42754
rect 25566 42702 25618 42754
rect 27918 42702 27970 42754
rect 29150 42702 29202 42754
rect 29710 42702 29762 42754
rect 30382 42702 30434 42754
rect 30718 42702 30770 42754
rect 34526 42702 34578 42754
rect 35870 42702 35922 42754
rect 40238 42702 40290 42754
rect 40574 42702 40626 42754
rect 40798 42702 40850 42754
rect 41918 42702 41970 42754
rect 42254 42702 42306 42754
rect 43038 42702 43090 42754
rect 48862 42702 48914 42754
rect 49086 42702 49138 42754
rect 49870 42702 49922 42754
rect 50766 42702 50818 42754
rect 52670 42702 52722 42754
rect 12462 42590 12514 42642
rect 16494 42590 16546 42642
rect 16942 42590 16994 42642
rect 17838 42590 17890 42642
rect 18062 42590 18114 42642
rect 19294 42590 19346 42642
rect 24446 42590 24498 42642
rect 25230 42590 25282 42642
rect 25342 42590 25394 42642
rect 25790 42590 25842 42642
rect 27806 42590 27858 42642
rect 30494 42590 30546 42642
rect 34862 42590 34914 42642
rect 36990 42590 37042 42642
rect 40350 42590 40402 42642
rect 40910 42590 40962 42642
rect 42814 42590 42866 42642
rect 46062 42590 46114 42642
rect 49310 42590 49362 42642
rect 51102 42590 51154 42642
rect 51438 42590 51490 42642
rect 51662 42590 51714 42642
rect 51998 42590 52050 42642
rect 4958 42478 5010 42530
rect 12126 42478 12178 42530
rect 12574 42478 12626 42530
rect 13806 42478 13858 42530
rect 14702 42478 14754 42530
rect 16270 42478 16322 42530
rect 16718 42478 16770 42530
rect 17502 42478 17554 42530
rect 18734 42478 18786 42530
rect 22654 42478 22706 42530
rect 25902 42478 25954 42530
rect 29486 42478 29538 42530
rect 32622 42478 32674 42530
rect 33966 42478 34018 42530
rect 34750 42478 34802 42530
rect 34974 42478 35026 42530
rect 36430 42478 36482 42530
rect 37102 42478 37154 42530
rect 37214 42478 37266 42530
rect 41134 42478 41186 42530
rect 42366 42478 42418 42530
rect 42478 42478 42530 42530
rect 43374 42478 43426 42530
rect 45614 42478 45666 42530
rect 47406 42478 47458 42530
rect 47742 42478 47794 42530
rect 50206 42478 50258 42530
rect 51774 42478 51826 42530
rect 52782 42478 52834 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 11566 42142 11618 42194
rect 12910 42142 12962 42194
rect 14590 42142 14642 42194
rect 16270 42142 16322 42194
rect 16718 42142 16770 42194
rect 17614 42142 17666 42194
rect 20750 42142 20802 42194
rect 22206 42142 22258 42194
rect 22990 42142 23042 42194
rect 23998 42142 24050 42194
rect 24110 42142 24162 42194
rect 26910 42142 26962 42194
rect 27134 42142 27186 42194
rect 27918 42142 27970 42194
rect 28142 42142 28194 42194
rect 31166 42142 31218 42194
rect 31950 42142 32002 42194
rect 32174 42142 32226 42194
rect 35422 42142 35474 42194
rect 41806 42142 41858 42194
rect 53118 42142 53170 42194
rect 12798 42030 12850 42082
rect 16830 42030 16882 42082
rect 18398 42030 18450 42082
rect 19742 42030 19794 42082
rect 20638 42030 20690 42082
rect 25118 42030 25170 42082
rect 25342 42030 25394 42082
rect 25454 42030 25506 42082
rect 25902 42030 25954 42082
rect 26350 42030 26402 42082
rect 26798 42030 26850 42082
rect 28926 42030 28978 42082
rect 29822 42030 29874 42082
rect 33294 42030 33346 42082
rect 39790 42030 39842 42082
rect 40126 42030 40178 42082
rect 40238 42030 40290 42082
rect 53006 42030 53058 42082
rect 53790 42030 53842 42082
rect 1822 41918 1874 41970
rect 8430 41918 8482 41970
rect 8878 41918 8930 41970
rect 9662 41918 9714 41970
rect 11006 41918 11058 41970
rect 11230 41918 11282 41970
rect 12462 41918 12514 41970
rect 13246 41918 13298 41970
rect 13470 41918 13522 41970
rect 14142 41918 14194 41970
rect 15486 41918 15538 41970
rect 15934 41918 15986 41970
rect 16158 41918 16210 41970
rect 16494 41918 16546 41970
rect 17390 41918 17442 41970
rect 17502 41918 17554 41970
rect 17950 41918 18002 41970
rect 18846 41918 18898 41970
rect 19966 41918 20018 41970
rect 20302 41918 20354 41970
rect 21646 41918 21698 41970
rect 22430 41918 22482 41970
rect 22766 41918 22818 41970
rect 23886 41918 23938 41970
rect 24558 41918 24610 41970
rect 25790 41918 25842 41970
rect 26462 41918 26514 41970
rect 27694 41918 27746 41970
rect 28366 41918 28418 41970
rect 29262 41918 29314 41970
rect 30830 41918 30882 41970
rect 31502 41918 31554 41970
rect 31726 41918 31778 41970
rect 32062 41918 32114 41970
rect 34190 41918 34242 41970
rect 34750 41918 34802 41970
rect 35198 41918 35250 41970
rect 35758 41918 35810 41970
rect 36542 41918 36594 41970
rect 39006 41918 39058 41970
rect 39230 41918 39282 41970
rect 39678 41918 39730 41970
rect 40462 41918 40514 41970
rect 41694 41918 41746 41970
rect 42254 41918 42306 41970
rect 43374 41918 43426 41970
rect 44158 41918 44210 41970
rect 45054 41918 45106 41970
rect 45502 41918 45554 41970
rect 49422 41918 49474 41970
rect 49758 41918 49810 41970
rect 51774 41918 51826 41970
rect 52334 41918 52386 41970
rect 52782 41918 52834 41970
rect 53678 41918 53730 41970
rect 2494 41806 2546 41858
rect 4622 41806 4674 41858
rect 4958 41806 5010 41858
rect 5518 41806 5570 41858
rect 6078 41806 6130 41858
rect 12238 41806 12290 41858
rect 14702 41806 14754 41858
rect 18958 41806 19010 41858
rect 19406 41806 19458 41858
rect 20078 41806 20130 41858
rect 29934 41806 29986 41858
rect 33182 41806 33234 41858
rect 34526 41806 34578 41858
rect 35310 41806 35362 41858
rect 38670 41806 38722 41858
rect 46734 41806 46786 41858
rect 47182 41806 47234 41858
rect 48750 41806 48802 41858
rect 50766 41806 50818 41858
rect 5294 41694 5346 41746
rect 13022 41694 13074 41746
rect 14254 41694 14306 41746
rect 15374 41694 15426 41746
rect 20862 41694 20914 41746
rect 21870 41694 21922 41746
rect 23102 41694 23154 41746
rect 26350 41694 26402 41746
rect 27806 41694 27858 41746
rect 29598 41694 29650 41746
rect 33070 41694 33122 41746
rect 34190 41694 34242 41746
rect 34638 41694 34690 41746
rect 39454 41694 39506 41746
rect 41806 41694 41858 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 2942 41358 2994 41410
rect 6862 41358 6914 41410
rect 17950 41358 18002 41410
rect 18286 41358 18338 41410
rect 18622 41358 18674 41410
rect 19294 41358 19346 41410
rect 19966 41358 20018 41410
rect 22094 41358 22146 41410
rect 23326 41358 23378 41410
rect 26798 41358 26850 41410
rect 39566 41358 39618 41410
rect 39902 41358 39954 41410
rect 49870 41358 49922 41410
rect 51998 41358 52050 41410
rect 52782 41358 52834 41410
rect 4958 41246 5010 41298
rect 8990 41246 9042 41298
rect 11118 41246 11170 41298
rect 23774 41246 23826 41298
rect 24558 41246 24610 41298
rect 25902 41246 25954 41298
rect 29934 41246 29986 41298
rect 32734 41246 32786 41298
rect 34862 41246 34914 41298
rect 39230 41246 39282 41298
rect 45166 41246 45218 41298
rect 48638 41246 48690 41298
rect 3278 41134 3330 41186
rect 3726 41134 3778 41186
rect 3838 41134 3890 41186
rect 4286 41134 4338 41186
rect 5966 41134 6018 41186
rect 6190 41134 6242 41186
rect 6414 41134 6466 41186
rect 6974 41134 7026 41186
rect 8318 41134 8370 41186
rect 14142 41134 14194 41186
rect 14478 41134 14530 41186
rect 15038 41134 15090 41186
rect 16046 41134 16098 41186
rect 16270 41134 16322 41186
rect 16494 41134 16546 41186
rect 16942 41134 16994 41186
rect 17390 41134 17442 41186
rect 18286 41134 18338 41186
rect 19966 41134 20018 41186
rect 20414 41134 20466 41186
rect 22766 41134 22818 41186
rect 22878 41134 22930 41186
rect 23998 41134 24050 41186
rect 24110 41134 24162 41186
rect 24670 41134 24722 41186
rect 25454 41134 25506 41186
rect 25678 41134 25730 41186
rect 26574 41134 26626 41186
rect 26910 41134 26962 41186
rect 27918 41134 27970 41186
rect 28590 41134 28642 41186
rect 29150 41134 29202 41186
rect 29822 41134 29874 41186
rect 30270 41134 30322 41186
rect 31950 41134 32002 41186
rect 35198 41134 35250 41186
rect 35534 41134 35586 41186
rect 36990 41134 37042 41186
rect 42926 41134 42978 41186
rect 43262 41134 43314 41186
rect 48078 41134 48130 41186
rect 48974 41134 49026 41186
rect 50318 41134 50370 41186
rect 50542 41134 50594 41186
rect 51214 41134 51266 41186
rect 51438 41134 51490 41186
rect 51550 41134 51602 41186
rect 3054 41022 3106 41074
rect 4846 41022 4898 41074
rect 5070 41022 5122 41074
rect 6526 41022 6578 41074
rect 7086 41022 7138 41074
rect 15150 41022 15202 41074
rect 17278 41022 17330 41074
rect 17502 41022 17554 41074
rect 18958 41022 19010 41074
rect 19630 41022 19682 41074
rect 20638 41022 20690 41074
rect 22094 41022 22146 41074
rect 22206 41022 22258 41074
rect 22654 41022 22706 41074
rect 23662 41022 23714 41074
rect 28478 41022 28530 41074
rect 29486 41022 29538 41074
rect 30606 41022 30658 41074
rect 35758 41022 35810 41074
rect 36430 41022 36482 41074
rect 37102 41022 37154 41074
rect 38446 41022 38498 41074
rect 39790 41022 39842 41074
rect 41582 41022 41634 41074
rect 42590 41022 42642 41074
rect 44270 41022 44322 41074
rect 47294 41022 47346 41074
rect 49870 41022 49922 41074
rect 49982 41022 50034 41074
rect 52894 41022 52946 41074
rect 3614 40910 3666 40962
rect 7870 40910 7922 40962
rect 14030 40910 14082 40962
rect 14590 40910 14642 40962
rect 14814 40910 14866 40962
rect 15374 40910 15426 40962
rect 16382 40910 16434 40962
rect 19182 40910 19234 40962
rect 28366 40910 28418 40962
rect 29374 40910 29426 40962
rect 35646 40910 35698 40962
rect 36206 40910 36258 40962
rect 36318 40910 36370 40962
rect 37214 40910 37266 40962
rect 37438 40910 37490 40962
rect 38110 40910 38162 40962
rect 38782 40910 38834 40962
rect 41470 40910 41522 40962
rect 41694 40910 41746 40962
rect 41918 40910 41970 40962
rect 43486 40910 43538 40962
rect 43710 40910 43762 40962
rect 44158 40910 44210 40962
rect 49534 40910 49586 40962
rect 50878 40910 50930 40962
rect 52782 40910 52834 40962
rect 53342 40910 53394 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 4510 40574 4562 40626
rect 11342 40574 11394 40626
rect 11678 40574 11730 40626
rect 15486 40574 15538 40626
rect 17614 40574 17666 40626
rect 21198 40574 21250 40626
rect 22318 40574 22370 40626
rect 22654 40574 22706 40626
rect 24110 40574 24162 40626
rect 25790 40574 25842 40626
rect 28366 40574 28418 40626
rect 28926 40574 28978 40626
rect 29150 40574 29202 40626
rect 29822 40574 29874 40626
rect 31838 40574 31890 40626
rect 34526 40574 34578 40626
rect 45278 40574 45330 40626
rect 46510 40574 46562 40626
rect 46846 40574 46898 40626
rect 47630 40574 47682 40626
rect 49198 40574 49250 40626
rect 51438 40574 51490 40626
rect 53790 40574 53842 40626
rect 7646 40462 7698 40514
rect 12014 40462 12066 40514
rect 12686 40462 12738 40514
rect 13246 40462 13298 40514
rect 13470 40462 13522 40514
rect 16158 40462 16210 40514
rect 18510 40462 18562 40514
rect 22094 40462 22146 40514
rect 25566 40462 25618 40514
rect 26014 40462 26066 40514
rect 27358 40462 27410 40514
rect 27582 40462 27634 40514
rect 27918 40462 27970 40514
rect 30158 40462 30210 40514
rect 30942 40462 30994 40514
rect 32510 40462 32562 40514
rect 35646 40462 35698 40514
rect 40014 40462 40066 40514
rect 42142 40462 42194 40514
rect 44942 40462 44994 40514
rect 46174 40462 46226 40514
rect 47182 40462 47234 40514
rect 51886 40462 51938 40514
rect 52446 40462 52498 40514
rect 4846 40350 4898 40402
rect 8318 40350 8370 40402
rect 12350 40350 12402 40402
rect 13582 40350 13634 40402
rect 13806 40350 13858 40402
rect 14030 40350 14082 40402
rect 14590 40350 14642 40402
rect 14926 40350 14978 40402
rect 15934 40350 15986 40402
rect 17950 40350 18002 40402
rect 19294 40350 19346 40402
rect 19966 40350 20018 40402
rect 21422 40350 21474 40402
rect 21534 40350 21586 40402
rect 21646 40350 21698 40402
rect 21982 40350 22034 40402
rect 22542 40350 22594 40402
rect 24334 40350 24386 40402
rect 25454 40350 25506 40402
rect 26350 40350 26402 40402
rect 28142 40350 28194 40402
rect 28702 40350 28754 40402
rect 31390 40350 31442 40402
rect 31950 40350 32002 40402
rect 34862 40350 34914 40402
rect 40350 40350 40402 40402
rect 41470 40350 41522 40402
rect 41918 40350 41970 40402
rect 42702 40350 42754 40402
rect 44270 40350 44322 40402
rect 44718 40350 44770 40402
rect 45838 40350 45890 40402
rect 48078 40350 48130 40402
rect 48974 40350 49026 40402
rect 49198 40350 49250 40402
rect 49534 40350 49586 40402
rect 50766 40350 50818 40402
rect 50878 40350 50930 40402
rect 51326 40350 51378 40402
rect 51550 40350 51602 40402
rect 52110 40350 52162 40402
rect 53454 40350 53506 40402
rect 5518 40238 5570 40290
rect 8878 40238 8930 40290
rect 19406 40238 19458 40290
rect 26238 40238 26290 40290
rect 27470 40238 27522 40290
rect 28814 40238 28866 40290
rect 37774 40238 37826 40290
rect 43150 40238 43202 40290
rect 44494 40238 44546 40290
rect 49982 40238 50034 40290
rect 52334 40238 52386 40290
rect 52894 40238 52946 40290
rect 4510 40126 4562 40178
rect 4622 40126 4674 40178
rect 15150 40126 15202 40178
rect 19630 40126 19682 40178
rect 19854 40126 19906 40178
rect 23998 40126 24050 40178
rect 28478 40126 28530 40178
rect 43934 40126 43986 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 5742 39790 5794 39842
rect 27022 39790 27074 39842
rect 2494 39678 2546 39730
rect 4622 39678 4674 39730
rect 6526 39678 6578 39730
rect 9438 39678 9490 39730
rect 11566 39678 11618 39730
rect 14366 39678 14418 39730
rect 17390 39678 17442 39730
rect 19070 39678 19122 39730
rect 21758 39678 21810 39730
rect 26350 39678 26402 39730
rect 34302 39678 34354 39730
rect 34750 39678 34802 39730
rect 36430 39678 36482 39730
rect 37774 39678 37826 39730
rect 39902 39678 39954 39730
rect 41694 39678 41746 39730
rect 42814 39678 42866 39730
rect 45614 39678 45666 39730
rect 48190 39678 48242 39730
rect 48974 39678 49026 39730
rect 50206 39678 50258 39730
rect 50542 39678 50594 39730
rect 52670 39678 52722 39730
rect 54798 39678 54850 39730
rect 1822 39566 1874 39618
rect 5518 39566 5570 39618
rect 8654 39566 8706 39618
rect 14254 39566 14306 39618
rect 14926 39566 14978 39618
rect 16942 39566 16994 39618
rect 19406 39566 19458 39618
rect 25230 39566 25282 39618
rect 26910 39566 26962 39618
rect 27582 39566 27634 39618
rect 27918 39566 27970 39618
rect 28254 39566 28306 39618
rect 31502 39566 31554 39618
rect 37102 39566 37154 39618
rect 41358 39566 41410 39618
rect 42590 39566 42642 39618
rect 45390 39566 45442 39618
rect 46062 39566 46114 39618
rect 46286 39566 46338 39618
rect 46734 39566 46786 39618
rect 46846 39566 46898 39618
rect 48526 39566 48578 39618
rect 49870 39566 49922 39618
rect 50878 39566 50930 39618
rect 55470 39566 55522 39618
rect 6638 39454 6690 39506
rect 6862 39454 6914 39506
rect 7198 39454 7250 39506
rect 7534 39454 7586 39506
rect 15150 39454 15202 39506
rect 15486 39454 15538 39506
rect 16606 39454 16658 39506
rect 19966 39454 20018 39506
rect 21534 39454 21586 39506
rect 22542 39454 22594 39506
rect 25454 39454 25506 39506
rect 26798 39454 26850 39506
rect 27694 39454 27746 39506
rect 28478 39454 28530 39506
rect 32174 39454 32226 39506
rect 42030 39454 42082 39506
rect 43486 39454 43538 39506
rect 51102 39454 51154 39506
rect 51886 39454 51938 39506
rect 5070 39342 5122 39394
rect 5854 39342 5906 39394
rect 6078 39342 6130 39394
rect 8318 39342 8370 39394
rect 14478 39342 14530 39394
rect 16158 39342 16210 39394
rect 16718 39342 16770 39394
rect 17278 39342 17330 39394
rect 18062 39342 18114 39394
rect 19518 39342 19570 39394
rect 20078 39342 20130 39394
rect 20750 39342 20802 39394
rect 22206 39342 22258 39394
rect 23438 39342 23490 39394
rect 25902 39342 25954 39394
rect 44270 39342 44322 39394
rect 46622 39342 46674 39394
rect 47518 39342 47570 39394
rect 51438 39342 51490 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 4398 39006 4450 39058
rect 5966 39006 6018 39058
rect 6302 39006 6354 39058
rect 7646 39006 7698 39058
rect 7758 39006 7810 39058
rect 11678 39006 11730 39058
rect 15150 39006 15202 39058
rect 15710 39006 15762 39058
rect 21758 39006 21810 39058
rect 23998 39006 24050 39058
rect 25566 39006 25618 39058
rect 26126 39006 26178 39058
rect 26910 39006 26962 39058
rect 28366 39006 28418 39058
rect 28702 39006 28754 39058
rect 29150 39006 29202 39058
rect 31614 39006 31666 39058
rect 32286 39006 32338 39058
rect 33182 39006 33234 39058
rect 42142 39006 42194 39058
rect 43038 39006 43090 39058
rect 43822 39006 43874 39058
rect 44046 39006 44098 39058
rect 45614 39006 45666 39058
rect 45726 39006 45778 39058
rect 46286 39006 46338 39058
rect 48302 39006 48354 39058
rect 49870 39006 49922 39058
rect 49982 39006 50034 39058
rect 50094 39006 50146 39058
rect 3054 38894 3106 38946
rect 3726 38894 3778 38946
rect 3950 38894 4002 38946
rect 4510 38894 4562 38946
rect 5406 38894 5458 38946
rect 5518 38894 5570 38946
rect 14814 38894 14866 38946
rect 15934 38894 15986 38946
rect 17390 38894 17442 38946
rect 17726 38894 17778 38946
rect 17950 38894 18002 38946
rect 18846 38894 18898 38946
rect 19854 38894 19906 38946
rect 26014 38894 26066 38946
rect 33294 38894 33346 38946
rect 37102 38894 37154 38946
rect 37886 38894 37938 38946
rect 38446 38894 38498 38946
rect 43710 38894 43762 38946
rect 44270 38894 44322 38946
rect 46510 38894 46562 38946
rect 48078 38894 48130 38946
rect 49198 38894 49250 38946
rect 2830 38782 2882 38834
rect 3390 38782 3442 38834
rect 3502 38782 3554 38834
rect 4286 38782 4338 38834
rect 4846 38782 4898 38834
rect 5182 38782 5234 38834
rect 6638 38782 6690 38834
rect 6862 38782 6914 38834
rect 7086 38782 7138 38834
rect 7534 38782 7586 38834
rect 12350 38782 12402 38834
rect 12574 38782 12626 38834
rect 13358 38782 13410 38834
rect 15038 38782 15090 38834
rect 16606 38782 16658 38834
rect 16830 38782 16882 38834
rect 19518 38782 19570 38834
rect 21422 38782 21474 38834
rect 22094 38782 22146 38834
rect 22430 38782 22482 38834
rect 22990 38782 23042 38834
rect 23662 38782 23714 38834
rect 24446 38782 24498 38834
rect 25230 38782 25282 38834
rect 27246 38782 27298 38834
rect 27694 38782 27746 38834
rect 30830 38782 30882 38834
rect 32062 38782 32114 38834
rect 32174 38782 32226 38834
rect 32622 38782 32674 38834
rect 32958 38782 33010 38834
rect 37774 38782 37826 38834
rect 38334 38782 38386 38834
rect 38670 38782 38722 38834
rect 42478 38782 42530 38834
rect 42702 38782 42754 38834
rect 45166 38782 45218 38834
rect 45838 38782 45890 38834
rect 46846 38782 46898 38834
rect 47406 38782 47458 38834
rect 47966 38782 48018 38834
rect 49310 38782 49362 38834
rect 49534 38782 49586 38834
rect 50430 38782 50482 38834
rect 54014 38782 54066 38834
rect 13022 38670 13074 38722
rect 15598 38670 15650 38722
rect 17502 38670 17554 38722
rect 30494 38670 30546 38722
rect 37214 38670 37266 38722
rect 37326 38670 37378 38722
rect 44606 38670 44658 38722
rect 47070 38670 47122 38722
rect 47630 38670 47682 38722
rect 51102 38670 51154 38722
rect 53230 38670 53282 38722
rect 15150 38558 15202 38610
rect 16270 38558 16322 38610
rect 20526 38558 20578 38610
rect 26126 38558 26178 38610
rect 37886 38558 37938 38610
rect 46622 38558 46674 38610
rect 48750 38558 48802 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 31614 38222 31666 38274
rect 50878 38222 50930 38274
rect 2494 38110 2546 38162
rect 4622 38110 4674 38162
rect 5070 38110 5122 38162
rect 6078 38110 6130 38162
rect 8206 38110 8258 38162
rect 10782 38110 10834 38162
rect 12910 38110 12962 38162
rect 13694 38110 13746 38162
rect 17166 38110 17218 38162
rect 18734 38110 18786 38162
rect 21310 38110 21362 38162
rect 23886 38110 23938 38162
rect 25342 38110 25394 38162
rect 27470 38110 27522 38162
rect 36206 38110 36258 38162
rect 38894 38110 38946 38162
rect 40126 38110 40178 38162
rect 44270 38110 44322 38162
rect 45054 38110 45106 38162
rect 1822 37998 1874 38050
rect 8878 37998 8930 38050
rect 10110 37998 10162 38050
rect 14366 37998 14418 38050
rect 14814 37998 14866 38050
rect 15038 37998 15090 38050
rect 15262 37998 15314 38050
rect 15822 37998 15874 38050
rect 19854 37998 19906 38050
rect 22654 37998 22706 38050
rect 23214 37998 23266 38050
rect 23662 37998 23714 38050
rect 28142 37998 28194 38050
rect 29486 37998 29538 38050
rect 31054 37998 31106 38050
rect 31278 37998 31330 38050
rect 34078 37998 34130 38050
rect 34526 37998 34578 38050
rect 38334 37998 38386 38050
rect 39230 37998 39282 38050
rect 42926 37998 42978 38050
rect 43374 37998 43426 38050
rect 44158 37998 44210 38050
rect 44830 37998 44882 38050
rect 45278 37998 45330 38050
rect 45390 37998 45442 38050
rect 45838 37998 45890 38050
rect 46622 37998 46674 38050
rect 47630 37998 47682 38050
rect 48862 37998 48914 38050
rect 49534 37998 49586 38050
rect 50206 37998 50258 38050
rect 51326 37998 51378 38050
rect 51774 37998 51826 38050
rect 52670 37998 52722 38050
rect 53118 37998 53170 38050
rect 13582 37886 13634 37938
rect 14030 37886 14082 37938
rect 14590 37886 14642 37938
rect 18622 37886 18674 37938
rect 19182 37886 19234 37938
rect 24222 37886 24274 37938
rect 24334 37886 24386 37938
rect 24446 37886 24498 37938
rect 29822 37886 29874 37938
rect 30382 37886 30434 37938
rect 30718 37886 30770 37938
rect 33742 37886 33794 37938
rect 37662 37886 37714 37938
rect 42254 37886 42306 37938
rect 43710 37886 43762 37938
rect 44942 37886 44994 37938
rect 9438 37774 9490 37826
rect 14142 37774 14194 37826
rect 14926 37774 14978 37826
rect 19294 37774 19346 37826
rect 19518 37774 19570 37826
rect 19742 37774 19794 37826
rect 20302 37774 20354 37826
rect 21870 37774 21922 37826
rect 25118 37774 25170 37826
rect 33966 37774 34018 37826
rect 34190 37774 34242 37826
rect 34638 37774 34690 37826
rect 34750 37774 34802 37826
rect 46174 37774 46226 37826
rect 47070 37774 47122 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 4398 37438 4450 37490
rect 15822 37438 15874 37490
rect 16158 37438 16210 37490
rect 16382 37438 16434 37490
rect 21422 37438 21474 37490
rect 24446 37438 24498 37490
rect 25342 37438 25394 37490
rect 25790 37438 25842 37490
rect 27022 37438 27074 37490
rect 30830 37438 30882 37490
rect 31502 37438 31554 37490
rect 36430 37438 36482 37490
rect 37662 37438 37714 37490
rect 39678 37438 39730 37490
rect 41022 37438 41074 37490
rect 44606 37438 44658 37490
rect 47630 37438 47682 37490
rect 53790 37438 53842 37490
rect 4622 37326 4674 37378
rect 4846 37326 4898 37378
rect 14702 37326 14754 37378
rect 15038 37326 15090 37378
rect 15598 37326 15650 37378
rect 20078 37326 20130 37378
rect 23774 37326 23826 37378
rect 26798 37326 26850 37378
rect 32174 37326 32226 37378
rect 33854 37326 33906 37378
rect 37102 37326 37154 37378
rect 37214 37326 37266 37378
rect 40238 37326 40290 37378
rect 40350 37326 40402 37378
rect 43262 37326 43314 37378
rect 44830 37326 44882 37378
rect 45726 37326 45778 37378
rect 55694 37326 55746 37378
rect 4174 37214 4226 37266
rect 9662 37214 9714 37266
rect 15262 37214 15314 37266
rect 16494 37214 16546 37266
rect 18062 37214 18114 37266
rect 18286 37214 18338 37266
rect 19070 37214 19122 37266
rect 20862 37214 20914 37266
rect 23326 37214 23378 37266
rect 24110 37214 24162 37266
rect 25566 37214 25618 37266
rect 27582 37214 27634 37266
rect 31166 37214 31218 37266
rect 31950 37214 32002 37266
rect 33070 37214 33122 37266
rect 36206 37214 36258 37266
rect 36542 37214 36594 37266
rect 36878 37214 36930 37266
rect 38446 37214 38498 37266
rect 38894 37214 38946 37266
rect 40014 37214 40066 37266
rect 43150 37214 43202 37266
rect 44270 37214 44322 37266
rect 45166 37214 45218 37266
rect 45390 37214 45442 37266
rect 48190 37214 48242 37266
rect 50094 37214 50146 37266
rect 51214 37214 51266 37266
rect 51774 37214 51826 37266
rect 52222 37214 52274 37266
rect 54686 37214 54738 37266
rect 54910 37214 54962 37266
rect 55358 37214 55410 37266
rect 55806 37214 55858 37266
rect 10334 37102 10386 37154
rect 12462 37102 12514 37154
rect 12910 37102 12962 37154
rect 13358 37102 13410 37154
rect 14478 37102 14530 37154
rect 14814 37102 14866 37154
rect 17614 37102 17666 37154
rect 22094 37102 22146 37154
rect 22878 37102 22930 37154
rect 25678 37102 25730 37154
rect 26462 37102 26514 37154
rect 27134 37102 27186 37154
rect 28254 37102 28306 37154
rect 30382 37102 30434 37154
rect 35982 37102 36034 37154
rect 39006 37102 39058 37154
rect 39454 37102 39506 37154
rect 42814 37102 42866 37154
rect 45614 37102 45666 37154
rect 47070 37102 47122 37154
rect 49982 37102 50034 37154
rect 53454 37102 53506 37154
rect 54238 37102 54290 37154
rect 55134 37102 55186 37154
rect 15934 36990 15986 37042
rect 17838 36990 17890 37042
rect 18734 36990 18786 37042
rect 21982 36990 22034 37042
rect 30606 36990 30658 37042
rect 30942 36990 30994 37042
rect 39790 36990 39842 37042
rect 47070 36990 47122 37042
rect 47518 36990 47570 37042
rect 47854 36990 47906 37042
rect 48190 36990 48242 37042
rect 55694 36990 55746 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 18958 36654 19010 36706
rect 19854 36654 19906 36706
rect 20750 36654 20802 36706
rect 31502 36654 31554 36706
rect 37550 36654 37602 36706
rect 38894 36654 38946 36706
rect 45502 36654 45554 36706
rect 47742 36654 47794 36706
rect 53006 36654 53058 36706
rect 56366 36654 56418 36706
rect 19070 36542 19122 36594
rect 19630 36542 19682 36594
rect 23662 36542 23714 36594
rect 24110 36542 24162 36594
rect 26238 36542 26290 36594
rect 27582 36542 27634 36594
rect 28590 36542 28642 36594
rect 33406 36542 33458 36594
rect 37998 36542 38050 36594
rect 40462 36542 40514 36594
rect 42590 36542 42642 36594
rect 47630 36542 47682 36594
rect 50878 36542 50930 36594
rect 54686 36542 54738 36594
rect 17502 36430 17554 36482
rect 18622 36430 18674 36482
rect 19294 36430 19346 36482
rect 20078 36430 20130 36482
rect 20302 36430 20354 36482
rect 21534 36430 21586 36482
rect 22206 36430 22258 36482
rect 23326 36430 23378 36482
rect 27022 36430 27074 36482
rect 30718 36430 30770 36482
rect 32062 36430 32114 36482
rect 33742 36430 33794 36482
rect 36094 36430 36146 36482
rect 36990 36430 37042 36482
rect 37214 36430 37266 36482
rect 37886 36430 37938 36482
rect 38110 36430 38162 36482
rect 38558 36430 38610 36482
rect 39678 36430 39730 36482
rect 45838 36430 45890 36482
rect 46174 36430 46226 36482
rect 47294 36430 47346 36482
rect 48078 36430 48130 36482
rect 48526 36430 48578 36482
rect 49646 36430 49698 36482
rect 50318 36430 50370 36482
rect 50542 36430 50594 36482
rect 50654 36430 50706 36482
rect 51326 36430 51378 36482
rect 53230 36430 53282 36482
rect 53454 36430 53506 36482
rect 55022 36430 55074 36482
rect 56366 36430 56418 36482
rect 57038 36430 57090 36482
rect 14590 36318 14642 36370
rect 16046 36318 16098 36370
rect 21310 36318 21362 36370
rect 22654 36318 22706 36370
rect 30158 36318 30210 36370
rect 31166 36318 31218 36370
rect 35870 36318 35922 36370
rect 39006 36318 39058 36370
rect 44830 36318 44882 36370
rect 46510 36318 46562 36370
rect 49086 36318 49138 36370
rect 50990 36318 51042 36370
rect 51662 36318 51714 36370
rect 51998 36318 52050 36370
rect 55470 36318 55522 36370
rect 55806 36318 55858 36370
rect 56030 36318 56082 36370
rect 14926 36206 14978 36258
rect 18286 36206 18338 36258
rect 22766 36206 22818 36258
rect 22878 36206 22930 36258
rect 30494 36206 30546 36258
rect 31390 36206 31442 36258
rect 31838 36206 31890 36258
rect 38894 36206 38946 36258
rect 43038 36206 43090 36258
rect 44270 36206 44322 36258
rect 45166 36206 45218 36258
rect 45614 36206 45666 36258
rect 48638 36206 48690 36258
rect 48750 36206 48802 36258
rect 49198 36206 49250 36258
rect 49310 36206 49362 36258
rect 52558 36206 52610 36258
rect 53902 36206 53954 36258
rect 56254 36206 56306 36258
rect 57486 36206 57538 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 16830 35870 16882 35922
rect 17390 35870 17442 35922
rect 18286 35870 18338 35922
rect 21422 35870 21474 35922
rect 21870 35870 21922 35922
rect 24782 35870 24834 35922
rect 25454 35870 25506 35922
rect 30494 35870 30546 35922
rect 31166 35870 31218 35922
rect 31614 35870 31666 35922
rect 40126 35870 40178 35922
rect 45166 35870 45218 35922
rect 48078 35870 48130 35922
rect 57374 35870 57426 35922
rect 16158 35758 16210 35810
rect 20526 35758 20578 35810
rect 22878 35758 22930 35810
rect 25790 35758 25842 35810
rect 26126 35758 26178 35810
rect 26462 35758 26514 35810
rect 34414 35758 34466 35810
rect 37550 35758 37602 35810
rect 44718 35758 44770 35810
rect 47854 35758 47906 35810
rect 48190 35758 48242 35810
rect 54014 35758 54066 35810
rect 56590 35758 56642 35810
rect 12014 35646 12066 35698
rect 15486 35646 15538 35698
rect 15710 35646 15762 35698
rect 15934 35646 15986 35698
rect 16494 35646 16546 35698
rect 17726 35646 17778 35698
rect 17950 35646 18002 35698
rect 18622 35646 18674 35698
rect 20078 35646 20130 35698
rect 22430 35646 22482 35698
rect 23438 35646 23490 35698
rect 23886 35646 23938 35698
rect 27246 35646 27298 35698
rect 29934 35646 29986 35698
rect 30270 35646 30322 35698
rect 31390 35646 31442 35698
rect 34638 35646 34690 35698
rect 36990 35646 37042 35698
rect 38558 35646 38610 35698
rect 39006 35646 39058 35698
rect 39342 35646 39394 35698
rect 39678 35646 39730 35698
rect 44942 35646 44994 35698
rect 46734 35646 46786 35698
rect 47070 35646 47122 35698
rect 47742 35646 47794 35698
rect 48750 35646 48802 35698
rect 49534 35646 49586 35698
rect 50654 35646 50706 35698
rect 52110 35646 52162 35698
rect 53230 35646 53282 35698
rect 54350 35646 54402 35698
rect 55134 35646 55186 35698
rect 56926 35646 56978 35698
rect 12686 35534 12738 35586
rect 14814 35534 14866 35586
rect 15598 35534 15650 35586
rect 19742 35534 19794 35586
rect 23550 35534 23602 35586
rect 30382 35534 30434 35586
rect 31502 35534 31554 35586
rect 36766 35534 36818 35586
rect 38110 35534 38162 35586
rect 43150 35534 43202 35586
rect 44270 35534 44322 35586
rect 45054 35534 45106 35586
rect 45614 35534 45666 35586
rect 51438 35534 51490 35586
rect 55806 35534 55858 35586
rect 56702 35534 56754 35586
rect 57822 35534 57874 35586
rect 34862 35422 34914 35474
rect 35086 35422 35138 35474
rect 35534 35422 35586 35474
rect 39678 35422 39730 35474
rect 57374 35422 57426 35474
rect 58046 35422 58098 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 13470 35086 13522 35138
rect 13806 35086 13858 35138
rect 15038 35086 15090 35138
rect 30382 35086 30434 35138
rect 31390 35086 31442 35138
rect 44046 35086 44098 35138
rect 44158 35086 44210 35138
rect 46174 35086 46226 35138
rect 53118 35086 53170 35138
rect 54574 35086 54626 35138
rect 14590 34974 14642 35026
rect 14814 34974 14866 35026
rect 18622 34974 18674 35026
rect 19070 34974 19122 35026
rect 21534 34974 21586 35026
rect 22430 34974 22482 35026
rect 25902 34974 25954 35026
rect 26238 34974 26290 35026
rect 27134 34974 27186 35026
rect 29710 34974 29762 35026
rect 30046 34974 30098 35026
rect 37550 34974 37602 35026
rect 40014 34974 40066 35026
rect 42142 34974 42194 35026
rect 45278 34974 45330 35026
rect 49422 34974 49474 35026
rect 49758 34974 49810 35026
rect 52894 34974 52946 35026
rect 54462 34974 54514 35026
rect 55246 34974 55298 35026
rect 57374 34974 57426 35026
rect 15822 34862 15874 34914
rect 19518 34862 19570 34914
rect 19966 34862 20018 34914
rect 20750 34862 20802 34914
rect 21982 34862 22034 34914
rect 22654 34862 22706 34914
rect 26798 34862 26850 34914
rect 27582 34862 27634 34914
rect 28142 34862 28194 34914
rect 31054 34862 31106 34914
rect 33518 34862 33570 34914
rect 34078 34862 34130 34914
rect 34414 34862 34466 34914
rect 34862 34862 34914 34914
rect 34974 34862 35026 34914
rect 35310 34862 35362 34914
rect 37214 34862 37266 34914
rect 39342 34862 39394 34914
rect 43822 34862 43874 34914
rect 45054 34862 45106 34914
rect 45502 34862 45554 34914
rect 45726 34862 45778 34914
rect 46062 34862 46114 34914
rect 47854 34862 47906 34914
rect 48414 34862 48466 34914
rect 50206 34862 50258 34914
rect 50654 34862 50706 34914
rect 52110 34862 52162 34914
rect 53342 34862 53394 34914
rect 53790 34862 53842 34914
rect 54798 34862 54850 34914
rect 58046 34862 58098 34914
rect 16494 34750 16546 34802
rect 20190 34750 20242 34802
rect 33854 34750 33906 34802
rect 43710 34750 43762 34802
rect 44830 34750 44882 34802
rect 46622 34750 46674 34802
rect 51102 34750 51154 34802
rect 13582 34638 13634 34690
rect 15374 34638 15426 34690
rect 18958 34638 19010 34690
rect 19854 34638 19906 34690
rect 23214 34638 23266 34690
rect 23550 34638 23602 34690
rect 23998 34638 24050 34690
rect 26350 34638 26402 34690
rect 28590 34638 28642 34690
rect 29150 34638 29202 34690
rect 30158 34638 30210 34690
rect 31278 34638 31330 34690
rect 33966 34638 34018 34690
rect 34750 34638 34802 34690
rect 38446 34638 38498 34690
rect 42590 34638 42642 34690
rect 42926 34638 42978 34690
rect 43374 34638 43426 34690
rect 45614 34638 45666 34690
rect 50990 34638 51042 34690
rect 51998 34638 52050 34690
rect 54462 34638 54514 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 15598 34302 15650 34354
rect 15934 34302 15986 34354
rect 17502 34302 17554 34354
rect 22654 34302 22706 34354
rect 25454 34302 25506 34354
rect 27582 34302 27634 34354
rect 36654 34302 36706 34354
rect 46958 34302 47010 34354
rect 47966 34302 48018 34354
rect 54014 34302 54066 34354
rect 56030 34302 56082 34354
rect 57374 34302 57426 34354
rect 58046 34302 58098 34354
rect 14030 34190 14082 34242
rect 14702 34190 14754 34242
rect 17390 34190 17442 34242
rect 17726 34190 17778 34242
rect 18846 34190 18898 34242
rect 21422 34190 21474 34242
rect 23214 34190 23266 34242
rect 29374 34190 29426 34242
rect 33854 34190 33906 34242
rect 43374 34190 43426 34242
rect 47854 34190 47906 34242
rect 48078 34190 48130 34242
rect 54238 34190 54290 34242
rect 54798 34190 54850 34242
rect 55022 34190 55074 34242
rect 55918 34190 55970 34242
rect 56590 34190 56642 34242
rect 57262 34190 57314 34242
rect 57486 34190 57538 34242
rect 16382 34078 16434 34130
rect 17950 34078 18002 34130
rect 22094 34078 22146 34130
rect 23550 34078 23602 34130
rect 24446 34078 24498 34130
rect 28702 34078 28754 34130
rect 33070 34078 33122 34130
rect 36766 34078 36818 34130
rect 37102 34078 37154 34130
rect 38222 34078 38274 34130
rect 39342 34078 39394 34130
rect 42702 34078 42754 34130
rect 46734 34078 46786 34130
rect 47182 34078 47234 34130
rect 47518 34078 47570 34130
rect 50318 34078 50370 34130
rect 50990 34078 51042 34130
rect 53230 34078 53282 34130
rect 53454 34078 53506 34130
rect 55246 34078 55298 34130
rect 55470 34078 55522 34130
rect 56814 34078 56866 34130
rect 14142 33966 14194 34018
rect 16942 33966 16994 34018
rect 18510 33966 18562 34018
rect 19294 33966 19346 34018
rect 23438 33966 23490 34018
rect 31502 33966 31554 34018
rect 32062 33966 32114 34018
rect 35982 33966 36034 34018
rect 45502 33966 45554 34018
rect 45950 33966 46002 34018
rect 47070 33966 47122 34018
rect 49870 33966 49922 34018
rect 53902 33966 53954 34018
rect 54910 33966 54962 34018
rect 14254 33854 14306 33906
rect 24110 33854 24162 33906
rect 24446 33854 24498 33906
rect 36654 33854 36706 33906
rect 38558 33854 38610 33906
rect 50206 33854 50258 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 17278 33518 17330 33570
rect 43822 33518 43874 33570
rect 48974 33518 49026 33570
rect 49310 33518 49362 33570
rect 50206 33518 50258 33570
rect 54798 33518 54850 33570
rect 14254 33406 14306 33458
rect 16382 33406 16434 33458
rect 16942 33406 16994 33458
rect 20750 33406 20802 33458
rect 24558 33406 24610 33458
rect 26686 33406 26738 33458
rect 31726 33406 31778 33458
rect 33854 33406 33906 33458
rect 40350 33406 40402 33458
rect 43598 33406 43650 33458
rect 49982 33406 50034 33458
rect 55246 33406 55298 33458
rect 57374 33406 57426 33458
rect 13582 33294 13634 33346
rect 18398 33294 18450 33346
rect 18958 33294 19010 33346
rect 19630 33294 19682 33346
rect 21310 33294 21362 33346
rect 21646 33294 21698 33346
rect 21982 33294 22034 33346
rect 22766 33294 22818 33346
rect 23774 33294 23826 33346
rect 27470 33294 27522 33346
rect 27582 33294 27634 33346
rect 31054 33294 31106 33346
rect 35534 33294 35586 33346
rect 37438 33294 37490 33346
rect 40910 33294 40962 33346
rect 42030 33294 42082 33346
rect 43486 33294 43538 33346
rect 46846 33294 46898 33346
rect 50318 33294 50370 33346
rect 53342 33294 53394 33346
rect 54350 33294 54402 33346
rect 58158 33294 58210 33346
rect 17054 33182 17106 33234
rect 27022 33182 27074 33234
rect 27246 33182 27298 33234
rect 35086 33182 35138 33234
rect 35646 33182 35698 33234
rect 38222 33182 38274 33234
rect 41022 33182 41074 33234
rect 42590 33182 42642 33234
rect 45838 33182 45890 33234
rect 46062 33182 46114 33234
rect 46510 33182 46562 33234
rect 49086 33182 49138 33234
rect 52782 33182 52834 33234
rect 54238 33182 54290 33234
rect 54686 33182 54738 33234
rect 17726 33070 17778 33122
rect 17838 33070 17890 33122
rect 17950 33070 18002 33122
rect 20190 33070 20242 33122
rect 21758 33070 21810 33122
rect 23102 33070 23154 33122
rect 23438 33070 23490 33122
rect 27806 33070 27858 33122
rect 34302 33070 34354 33122
rect 36206 33070 36258 33122
rect 37102 33070 37154 33122
rect 41918 33070 41970 33122
rect 43262 33070 43314 33122
rect 45950 33070 46002 33122
rect 46622 33070 46674 33122
rect 51102 33070 51154 33122
rect 52110 33070 52162 33122
rect 53230 33070 53282 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 15598 32734 15650 32786
rect 18510 32734 18562 32786
rect 19294 32734 19346 32786
rect 30046 32734 30098 32786
rect 32174 32734 32226 32786
rect 32510 32734 32562 32786
rect 34190 32734 34242 32786
rect 35086 32734 35138 32786
rect 36990 32734 37042 32786
rect 37662 32734 37714 32786
rect 38110 32734 38162 32786
rect 38558 32734 38610 32786
rect 41246 32734 41298 32786
rect 45054 32734 45106 32786
rect 45390 32734 45442 32786
rect 45726 32734 45778 32786
rect 49086 32734 49138 32786
rect 49870 32734 49922 32786
rect 52222 32734 52274 32786
rect 56702 32734 56754 32786
rect 18846 32622 18898 32674
rect 19630 32622 19682 32674
rect 25566 32622 25618 32674
rect 26014 32622 26066 32674
rect 28814 32622 28866 32674
rect 30830 32622 30882 32674
rect 37438 32622 37490 32674
rect 43262 32622 43314 32674
rect 43486 32622 43538 32674
rect 45278 32622 45330 32674
rect 47406 32622 47458 32674
rect 49534 32622 49586 32674
rect 50318 32622 50370 32674
rect 53342 32622 53394 32674
rect 54798 32622 54850 32674
rect 12350 32510 12402 32562
rect 16270 32510 16322 32562
rect 16382 32510 16434 32562
rect 16606 32510 16658 32562
rect 16830 32510 16882 32562
rect 17502 32510 17554 32562
rect 17614 32510 17666 32562
rect 17726 32510 17778 32562
rect 17838 32510 17890 32562
rect 18062 32510 18114 32562
rect 18398 32510 18450 32562
rect 18622 32510 18674 32562
rect 20078 32510 20130 32562
rect 23326 32510 23378 32562
rect 23550 32510 23602 32562
rect 23774 32510 23826 32562
rect 23998 32510 24050 32562
rect 24334 32510 24386 32562
rect 26126 32510 26178 32562
rect 26350 32510 26402 32562
rect 29598 32510 29650 32562
rect 30606 32510 30658 32562
rect 33518 32510 33570 32562
rect 35310 32510 35362 32562
rect 37326 32510 37378 32562
rect 37886 32510 37938 32562
rect 38334 32510 38386 32562
rect 41582 32510 41634 32562
rect 43038 32510 43090 32562
rect 44830 32510 44882 32562
rect 45614 32510 45666 32562
rect 47070 32510 47122 32562
rect 47630 32510 47682 32562
rect 48862 32510 48914 32562
rect 49758 32510 49810 32562
rect 49982 32510 50034 32562
rect 50542 32510 50594 32562
rect 50878 32510 50930 32562
rect 51662 32510 51714 32562
rect 51774 32510 51826 32562
rect 52110 32510 52162 32562
rect 55918 32510 55970 32562
rect 13022 32398 13074 32450
rect 15150 32398 15202 32450
rect 16494 32398 16546 32450
rect 20750 32398 20802 32450
rect 22878 32398 22930 32450
rect 23662 32398 23714 32450
rect 24446 32398 24498 32450
rect 25678 32398 25730 32450
rect 26686 32398 26738 32450
rect 33182 32398 33234 32450
rect 34750 32398 34802 32450
rect 38222 32398 38274 32450
rect 41806 32398 41858 32450
rect 41918 32398 41970 32450
rect 42702 32398 42754 32450
rect 43150 32398 43202 32450
rect 47518 32398 47570 32450
rect 48190 32398 48242 32450
rect 50766 32398 50818 32450
rect 51438 32398 51490 32450
rect 57150 32398 57202 32450
rect 45838 32286 45890 32338
rect 46062 32286 46114 32338
rect 46286 32286 46338 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 18734 31950 18786 32002
rect 23550 31950 23602 32002
rect 27470 31950 27522 32002
rect 37550 31950 37602 32002
rect 48974 31950 49026 32002
rect 51550 31950 51602 32002
rect 13694 31838 13746 31890
rect 15598 31838 15650 31890
rect 21870 31838 21922 31890
rect 24558 31838 24610 31890
rect 28366 31838 28418 31890
rect 33518 31838 33570 31890
rect 38782 31838 38834 31890
rect 40686 31838 40738 31890
rect 41918 31838 41970 31890
rect 44046 31838 44098 31890
rect 46958 31838 47010 31890
rect 53230 31838 53282 31890
rect 53902 31838 53954 31890
rect 13806 31726 13858 31778
rect 16158 31726 16210 31778
rect 16606 31726 16658 31778
rect 17390 31726 17442 31778
rect 18846 31726 18898 31778
rect 19518 31726 19570 31778
rect 22206 31726 22258 31778
rect 23102 31726 23154 31778
rect 23662 31726 23714 31778
rect 27022 31726 27074 31778
rect 27246 31726 27298 31778
rect 27806 31726 27858 31778
rect 30270 31726 30322 31778
rect 31502 31726 31554 31778
rect 32062 31726 32114 31778
rect 34190 31726 34242 31778
rect 34302 31726 34354 31778
rect 34526 31726 34578 31778
rect 37438 31726 37490 31778
rect 37662 31726 37714 31778
rect 41246 31726 41298 31778
rect 46286 31726 46338 31778
rect 48078 31726 48130 31778
rect 49422 31726 49474 31778
rect 49646 31726 49698 31778
rect 50654 31726 50706 31778
rect 50878 31726 50930 31778
rect 51550 31726 51602 31778
rect 51886 31726 51938 31778
rect 52110 31726 52162 31778
rect 52670 31726 52722 31778
rect 56702 31726 56754 31778
rect 13470 31614 13522 31666
rect 15710 31614 15762 31666
rect 17054 31614 17106 31666
rect 20078 31614 20130 31666
rect 21870 31614 21922 31666
rect 22430 31614 22482 31666
rect 24894 31614 24946 31666
rect 26350 31614 26402 31666
rect 29934 31614 29986 31666
rect 33854 31614 33906 31666
rect 34750 31614 34802 31666
rect 37102 31614 37154 31666
rect 38894 31614 38946 31666
rect 40350 31614 40402 31666
rect 40574 31614 40626 31666
rect 45838 31614 45890 31666
rect 47182 31614 47234 31666
rect 48302 31614 48354 31666
rect 48862 31614 48914 31666
rect 49982 31614 50034 31666
rect 51998 31614 52050 31666
rect 56030 31614 56082 31666
rect 14254 31502 14306 31554
rect 15486 31502 15538 31554
rect 21982 31502 22034 31554
rect 25678 31502 25730 31554
rect 26686 31502 26738 31554
rect 27806 31502 27858 31554
rect 34302 31502 34354 31554
rect 35198 31502 35250 31554
rect 35982 31502 36034 31554
rect 36430 31502 36482 31554
rect 37550 31502 37602 31554
rect 38334 31502 38386 31554
rect 44942 31502 44994 31554
rect 46958 31502 47010 31554
rect 48974 31502 49026 31554
rect 49758 31502 49810 31554
rect 50318 31502 50370 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 13470 31166 13522 31218
rect 14030 31166 14082 31218
rect 17390 31166 17442 31218
rect 19182 31166 19234 31218
rect 22990 31166 23042 31218
rect 24222 31166 24274 31218
rect 47070 31166 47122 31218
rect 47518 31166 47570 31218
rect 53678 31166 53730 31218
rect 13246 31054 13298 31106
rect 16830 31054 16882 31106
rect 17502 31054 17554 31106
rect 18286 31054 18338 31106
rect 23102 31054 23154 31106
rect 23886 31054 23938 31106
rect 24446 31054 24498 31106
rect 34414 31054 34466 31106
rect 37662 31054 37714 31106
rect 41918 31054 41970 31106
rect 43486 31054 43538 31106
rect 43598 31054 43650 31106
rect 43934 31054 43986 31106
rect 44718 31054 44770 31106
rect 45838 31054 45890 31106
rect 48750 31054 48802 31106
rect 54462 31054 54514 31106
rect 9550 30942 9602 30994
rect 16158 30942 16210 30994
rect 18174 30942 18226 30994
rect 19070 30942 19122 30994
rect 19630 30942 19682 30994
rect 23998 30942 24050 30994
rect 24558 30942 24610 30994
rect 32062 30942 32114 30994
rect 32510 30942 32562 30994
rect 33742 30942 33794 30994
rect 36878 30942 36930 30994
rect 41470 30942 41522 30994
rect 42142 30942 42194 30994
rect 43262 30942 43314 30994
rect 44158 30942 44210 30994
rect 44270 30942 44322 30994
rect 44830 30942 44882 30994
rect 45502 30942 45554 30994
rect 46398 30942 46450 30994
rect 48078 30942 48130 30994
rect 48862 30942 48914 30994
rect 49086 30942 49138 30994
rect 49198 30942 49250 30994
rect 51102 30942 51154 30994
rect 51438 30942 51490 30994
rect 52446 30942 52498 30994
rect 52782 30942 52834 30994
rect 53006 30942 53058 30994
rect 53902 30942 53954 30994
rect 10334 30830 10386 30882
rect 12462 30830 12514 30882
rect 12910 30830 12962 30882
rect 16382 30830 16434 30882
rect 20414 30830 20466 30882
rect 22542 30830 22594 30882
rect 29150 30830 29202 30882
rect 31278 30830 31330 30882
rect 36542 30830 36594 30882
rect 39790 30830 39842 30882
rect 41022 30830 41074 30882
rect 49870 30830 49922 30882
rect 51998 30830 52050 30882
rect 13582 30718 13634 30770
rect 13918 30718 13970 30770
rect 14254 30718 14306 30770
rect 42478 30718 42530 30770
rect 44718 30718 44770 30770
rect 45390 30718 45442 30770
rect 45726 30718 45778 30770
rect 46286 30718 46338 30770
rect 46622 30718 46674 30770
rect 53342 30718 53394 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 20414 30382 20466 30434
rect 20750 30382 20802 30434
rect 21310 30382 21362 30434
rect 21646 30382 21698 30434
rect 29822 30382 29874 30434
rect 36094 30382 36146 30434
rect 39566 30382 39618 30434
rect 14254 30270 14306 30322
rect 16382 30270 16434 30322
rect 19294 30270 19346 30322
rect 25230 30270 25282 30322
rect 35758 30270 35810 30322
rect 13470 30158 13522 30210
rect 16830 30158 16882 30210
rect 17502 30158 17554 30210
rect 18622 30158 18674 30210
rect 19742 30158 19794 30210
rect 21310 30158 21362 30210
rect 22990 30158 23042 30210
rect 24334 30158 24386 30210
rect 25454 30158 25506 30210
rect 26574 30158 26626 30210
rect 27022 30158 27074 30210
rect 28254 30158 28306 30210
rect 29822 30158 29874 30210
rect 30270 30158 30322 30210
rect 33630 30158 33682 30210
rect 36990 30158 37042 30210
rect 37326 30158 37378 30210
rect 38110 30158 38162 30210
rect 38782 30158 38834 30210
rect 39454 30158 39506 30210
rect 40126 30158 40178 30210
rect 40798 30158 40850 30210
rect 41134 30158 41186 30210
rect 41806 30158 41858 30210
rect 42478 30158 42530 30210
rect 43150 30158 43202 30210
rect 45054 30158 45106 30210
rect 45614 30158 45666 30210
rect 46286 30158 46338 30210
rect 46846 30158 46898 30210
rect 47630 30158 47682 30210
rect 48974 30158 49026 30210
rect 50206 30158 50258 30210
rect 50542 30158 50594 30210
rect 53118 30158 53170 30210
rect 53790 30158 53842 30210
rect 9550 30046 9602 30098
rect 9886 30046 9938 30098
rect 17950 30046 18002 30098
rect 20526 30046 20578 30098
rect 25790 30046 25842 30098
rect 26462 30046 26514 30098
rect 28590 30046 28642 30098
rect 29486 30046 29538 30098
rect 39230 30046 39282 30098
rect 40462 30046 40514 30098
rect 41470 30046 41522 30098
rect 45166 30046 45218 30098
rect 46958 30046 47010 30098
rect 47966 30046 48018 30098
rect 51550 30046 51602 30098
rect 53566 30046 53618 30098
rect 18398 29934 18450 29986
rect 22094 29934 22146 29986
rect 28478 29934 28530 29986
rect 35982 29934 36034 29986
rect 39790 29934 39842 29986
rect 42142 29934 42194 29986
rect 42814 29934 42866 29986
rect 43486 29934 43538 29986
rect 45278 29934 45330 29986
rect 45726 29934 45778 29986
rect 50878 29934 50930 29986
rect 52894 29934 52946 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 10334 29598 10386 29650
rect 16270 29598 16322 29650
rect 18174 29598 18226 29650
rect 19518 29598 19570 29650
rect 29038 29598 29090 29650
rect 31278 29598 31330 29650
rect 32398 29598 32450 29650
rect 33182 29598 33234 29650
rect 34862 29598 34914 29650
rect 47518 29598 47570 29650
rect 48862 29598 48914 29650
rect 51662 29598 51714 29650
rect 11230 29486 11282 29538
rect 13694 29486 13746 29538
rect 25342 29486 25394 29538
rect 28814 29486 28866 29538
rect 29486 29486 29538 29538
rect 30158 29486 30210 29538
rect 30270 29486 30322 29538
rect 30830 29486 30882 29538
rect 35422 29486 35474 29538
rect 41246 29486 41298 29538
rect 45838 29486 45890 29538
rect 46510 29486 46562 29538
rect 48078 29486 48130 29538
rect 49646 29486 49698 29538
rect 52110 29486 52162 29538
rect 52222 29486 52274 29538
rect 53342 29486 53394 29538
rect 5294 29374 5346 29426
rect 8542 29374 8594 29426
rect 11454 29374 11506 29426
rect 12910 29374 12962 29426
rect 21310 29374 21362 29426
rect 25454 29374 25506 29426
rect 25678 29374 25730 29426
rect 26462 29374 26514 29426
rect 28702 29374 28754 29426
rect 29374 29374 29426 29426
rect 29934 29374 29986 29426
rect 31950 29374 32002 29426
rect 32174 29374 32226 29426
rect 32622 29374 32674 29426
rect 34190 29374 34242 29426
rect 41022 29374 41074 29426
rect 44158 29374 44210 29426
rect 45166 29374 45218 29426
rect 46062 29374 46114 29426
rect 46622 29374 46674 29426
rect 49758 29374 49810 29426
rect 50430 29374 50482 29426
rect 50542 29374 50594 29426
rect 52446 29374 52498 29426
rect 53118 29374 53170 29426
rect 53454 29374 53506 29426
rect 53678 29374 53730 29426
rect 54574 29374 54626 29426
rect 5966 29262 6018 29314
rect 8094 29262 8146 29314
rect 15822 29262 15874 29314
rect 18286 29262 18338 29314
rect 18958 29262 19010 29314
rect 21982 29262 22034 29314
rect 24110 29262 24162 29314
rect 24670 29262 24722 29314
rect 29710 29262 29762 29314
rect 33518 29262 33570 29314
rect 34414 29262 34466 29314
rect 35198 29262 35250 29314
rect 43710 29262 43762 29314
rect 46958 29262 47010 29314
rect 47854 29262 47906 29314
rect 49982 29262 50034 29314
rect 54014 29262 54066 29314
rect 55022 29262 55074 29314
rect 10670 29150 10722 29202
rect 30270 29150 30322 29202
rect 30718 29150 30770 29202
rect 52670 29150 52722 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 21982 28814 22034 28866
rect 27582 28814 27634 28866
rect 28254 28814 28306 28866
rect 33406 28814 33458 28866
rect 35198 28814 35250 28866
rect 46174 28814 46226 28866
rect 46846 28814 46898 28866
rect 12014 28702 12066 28754
rect 16718 28702 16770 28754
rect 19518 28702 19570 28754
rect 23214 28702 23266 28754
rect 23550 28702 23602 28754
rect 27918 28702 27970 28754
rect 28590 28702 28642 28754
rect 29150 28702 29202 28754
rect 31278 28702 31330 28754
rect 37102 28702 37154 28754
rect 37998 28702 38050 28754
rect 39678 28702 39730 28754
rect 45502 28702 45554 28754
rect 45614 28702 45666 28754
rect 48638 28702 48690 28754
rect 55246 28702 55298 28754
rect 57374 28702 57426 28754
rect 6526 28590 6578 28642
rect 7198 28590 7250 28642
rect 7534 28590 7586 28642
rect 9214 28590 9266 28642
rect 12462 28590 12514 28642
rect 15934 28590 15986 28642
rect 23662 28590 23714 28642
rect 26686 28590 26738 28642
rect 26798 28590 26850 28642
rect 27134 28590 27186 28642
rect 32062 28590 32114 28642
rect 32622 28590 32674 28642
rect 32958 28590 33010 28642
rect 33182 28590 33234 28642
rect 33630 28590 33682 28642
rect 33966 28590 34018 28642
rect 34526 28590 34578 28642
rect 34862 28590 34914 28642
rect 36206 28590 36258 28642
rect 37550 28590 37602 28642
rect 38334 28590 38386 28642
rect 40014 28590 40066 28642
rect 40686 28590 40738 28642
rect 42590 28590 42642 28642
rect 43374 28590 43426 28642
rect 43934 28590 43986 28642
rect 45166 28590 45218 28642
rect 45950 28590 46002 28642
rect 49310 28590 49362 28642
rect 50318 28590 50370 28642
rect 50990 28590 51042 28642
rect 52110 28590 52162 28642
rect 52670 28590 52722 28642
rect 53230 28590 53282 28642
rect 53902 28590 53954 28642
rect 54574 28590 54626 28642
rect 6302 28478 6354 28530
rect 7758 28478 7810 28530
rect 8094 28478 8146 28530
rect 9886 28478 9938 28530
rect 21310 28478 21362 28530
rect 22094 28478 22146 28530
rect 22318 28478 22370 28530
rect 26350 28478 26402 28530
rect 27806 28478 27858 28530
rect 28478 28478 28530 28530
rect 32510 28478 32562 28530
rect 35310 28478 35362 28530
rect 38670 28478 38722 28530
rect 41022 28478 41074 28530
rect 46958 28478 47010 28530
rect 51998 28478 52050 28530
rect 52894 28478 52946 28530
rect 18958 28366 19010 28418
rect 21646 28366 21698 28418
rect 27134 28366 27186 28418
rect 32846 28366 32898 28418
rect 34638 28366 34690 28418
rect 35198 28366 35250 28418
rect 35758 28366 35810 28418
rect 40350 28366 40402 28418
rect 40910 28366 40962 28418
rect 42926 28366 42978 28418
rect 46510 28366 46562 28418
rect 51102 28366 51154 28418
rect 52782 28366 52834 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 9774 28030 9826 28082
rect 19742 28030 19794 28082
rect 19854 28030 19906 28082
rect 25454 28030 25506 28082
rect 39342 28030 39394 28082
rect 41694 28030 41746 28082
rect 46286 28030 46338 28082
rect 47630 28030 47682 28082
rect 47854 28030 47906 28082
rect 52110 28030 52162 28082
rect 55134 28030 55186 28082
rect 55582 28030 55634 28082
rect 55694 28030 55746 28082
rect 56590 28030 56642 28082
rect 7870 27918 7922 27970
rect 8430 27918 8482 27970
rect 11454 27918 11506 27970
rect 19294 27918 19346 27970
rect 20526 27918 20578 27970
rect 22318 27918 22370 27970
rect 22654 27918 22706 27970
rect 25342 27918 25394 27970
rect 25566 27918 25618 27970
rect 28142 27918 28194 27970
rect 30158 27918 30210 27970
rect 34526 27918 34578 27970
rect 35982 27918 36034 27970
rect 36206 27918 36258 27970
rect 36654 27918 36706 27970
rect 39230 27918 39282 27970
rect 46734 27918 46786 27970
rect 52670 27918 52722 27970
rect 53006 27918 53058 27970
rect 3502 27806 3554 27858
rect 7758 27806 7810 27858
rect 10110 27806 10162 27858
rect 10558 27806 10610 27858
rect 11342 27806 11394 27858
rect 19070 27806 19122 27858
rect 20750 27806 20802 27858
rect 21086 27806 21138 27858
rect 21646 27806 21698 27858
rect 22878 27806 22930 27858
rect 23998 27806 24050 27858
rect 24446 27806 24498 27858
rect 24558 27806 24610 27858
rect 28814 27806 28866 27858
rect 29374 27806 29426 27858
rect 33406 27806 33458 27858
rect 34078 27806 34130 27858
rect 34302 27806 34354 27858
rect 34750 27806 34802 27858
rect 34862 27806 34914 27858
rect 35534 27806 35586 27858
rect 36542 27806 36594 27858
rect 38670 27806 38722 27858
rect 41806 27806 41858 27858
rect 41918 27806 41970 27858
rect 43038 27806 43090 27858
rect 46846 27806 46898 27858
rect 46958 27806 47010 27858
rect 47406 27806 47458 27858
rect 49198 27806 49250 27858
rect 51662 27806 51714 27858
rect 51886 27806 51938 27858
rect 52782 27806 52834 27858
rect 54350 27806 54402 27858
rect 54686 27806 54738 27858
rect 54910 27806 54962 27858
rect 56702 27806 56754 27858
rect 4174 27694 4226 27746
rect 6302 27694 6354 27746
rect 7086 27694 7138 27746
rect 18734 27694 18786 27746
rect 21422 27694 21474 27746
rect 24222 27694 24274 27746
rect 26014 27694 26066 27746
rect 32398 27694 32450 27746
rect 33294 27694 33346 27746
rect 36094 27694 36146 27746
rect 42142 27694 42194 27746
rect 43710 27694 43762 27746
rect 45838 27694 45890 27746
rect 47518 27694 47570 27746
rect 50430 27694 50482 27746
rect 51774 27694 51826 27746
rect 53790 27694 53842 27746
rect 55470 27694 55522 27746
rect 6750 27582 6802 27634
rect 8318 27582 8370 27634
rect 10894 27582 10946 27634
rect 19966 27582 20018 27634
rect 20414 27582 20466 27634
rect 35758 27582 35810 27634
rect 42366 27582 42418 27634
rect 54798 27582 54850 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 34526 27246 34578 27298
rect 37438 27246 37490 27298
rect 7086 27134 7138 27186
rect 16270 27134 16322 27186
rect 18398 27134 18450 27186
rect 18734 27134 18786 27186
rect 19406 27134 19458 27186
rect 20302 27134 20354 27186
rect 26574 27160 26626 27212
rect 33518 27134 33570 27186
rect 38782 27134 38834 27186
rect 40910 27134 40962 27186
rect 42366 27134 42418 27186
rect 46734 27134 46786 27186
rect 49422 27134 49474 27186
rect 49646 27134 49698 27186
rect 50206 27134 50258 27186
rect 50542 27134 50594 27186
rect 51998 27134 52050 27186
rect 53006 27134 53058 27186
rect 57038 27134 57090 27186
rect 4958 27022 5010 27074
rect 15486 27022 15538 27074
rect 20078 27022 20130 27074
rect 21310 27022 21362 27074
rect 21870 27022 21922 27074
rect 22542 27022 22594 27074
rect 23774 27022 23826 27074
rect 27022 27022 27074 27074
rect 29262 27022 29314 27074
rect 33406 27022 33458 27074
rect 34414 27022 34466 27074
rect 34638 27022 34690 27074
rect 36094 27022 36146 27074
rect 37214 27022 37266 27074
rect 37550 27022 37602 27074
rect 37998 27022 38050 27074
rect 41694 27022 41746 27074
rect 42254 27022 42306 27074
rect 42926 27022 42978 27074
rect 43710 27022 43762 27074
rect 44158 27022 44210 27074
rect 44830 27022 44882 27074
rect 48526 27022 48578 27074
rect 48862 27022 48914 27074
rect 49870 27022 49922 27074
rect 50654 27022 50706 27074
rect 51550 27022 51602 27074
rect 52782 27022 52834 27074
rect 53230 27022 53282 27074
rect 54126 27022 54178 27074
rect 4622 26910 4674 26962
rect 5630 26910 5682 26962
rect 5966 26910 6018 26962
rect 13470 26910 13522 26962
rect 13806 26910 13858 26962
rect 18846 26910 18898 26962
rect 19070 26910 19122 26962
rect 21198 26910 21250 26962
rect 21534 26910 21586 26962
rect 24446 26910 24498 26962
rect 29710 26910 29762 26962
rect 33854 26910 33906 26962
rect 34190 26910 34242 26962
rect 35870 26910 35922 26962
rect 36990 26910 37042 26962
rect 42478 26910 42530 26962
rect 43150 26910 43202 26962
rect 43262 26910 43314 26962
rect 43486 26910 43538 26962
rect 44046 26910 44098 26962
rect 45950 26910 46002 26962
rect 48638 26910 48690 26962
rect 49198 26910 49250 26962
rect 53342 26910 53394 26962
rect 53454 26910 53506 26962
rect 54910 26910 54962 26962
rect 6526 26798 6578 26850
rect 6974 26798 7026 26850
rect 15150 26798 15202 26850
rect 23438 26798 23490 26850
rect 35086 26798 35138 26850
rect 35534 26798 35586 26850
rect 37102 26798 37154 26850
rect 38334 26798 38386 26850
rect 49982 26798 50034 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 15374 26462 15426 26514
rect 16606 26462 16658 26514
rect 24222 26462 24274 26514
rect 25566 26462 25618 26514
rect 32510 26462 32562 26514
rect 34862 26462 34914 26514
rect 41918 26462 41970 26514
rect 44718 26462 44770 26514
rect 46398 26462 46450 26514
rect 47182 26462 47234 26514
rect 55582 26462 55634 26514
rect 4846 26350 4898 26402
rect 7982 26350 8034 26402
rect 10110 26350 10162 26402
rect 11678 26350 11730 26402
rect 12910 26350 12962 26402
rect 19518 26350 19570 26402
rect 21982 26350 22034 26402
rect 24446 26350 24498 26402
rect 25230 26350 25282 26402
rect 26462 26350 26514 26402
rect 34750 26350 34802 26402
rect 35086 26350 35138 26402
rect 35198 26350 35250 26402
rect 36430 26350 36482 26402
rect 40126 26350 40178 26402
rect 45390 26350 45442 26402
rect 46622 26350 46674 26402
rect 46846 26350 46898 26402
rect 47742 26350 47794 26402
rect 48302 26350 48354 26402
rect 48750 26350 48802 26402
rect 4174 26238 4226 26290
rect 8318 26238 8370 26290
rect 9886 26238 9938 26290
rect 10558 26238 10610 26290
rect 10894 26238 10946 26290
rect 11454 26238 11506 26290
rect 12238 26238 12290 26290
rect 15710 26238 15762 26290
rect 18286 26238 18338 26290
rect 18622 26238 18674 26290
rect 19966 26238 20018 26290
rect 20414 26238 20466 26290
rect 21534 26238 21586 26290
rect 22206 26238 22258 26290
rect 22430 26238 22482 26290
rect 22878 26238 22930 26290
rect 23662 26238 23714 26290
rect 23998 26238 24050 26290
rect 24110 26238 24162 26290
rect 26238 26238 26290 26290
rect 29598 26238 29650 26290
rect 33070 26238 33122 26290
rect 33294 26238 33346 26290
rect 33518 26238 33570 26290
rect 33742 26238 33794 26290
rect 33966 26238 34018 26290
rect 34190 26238 34242 26290
rect 34526 26238 34578 26290
rect 35758 26238 35810 26290
rect 38894 26238 38946 26290
rect 39790 26238 39842 26290
rect 40350 26238 40402 26290
rect 40910 26238 40962 26290
rect 42814 26238 42866 26290
rect 44046 26238 44098 26290
rect 44382 26238 44434 26290
rect 46286 26238 46338 26290
rect 49086 26238 49138 26290
rect 49422 26238 49474 26290
rect 49758 26238 49810 26290
rect 50766 26238 50818 26290
rect 51438 26238 51490 26290
rect 52334 26238 52386 26290
rect 6974 26126 7026 26178
rect 7422 26126 7474 26178
rect 15038 26126 15090 26178
rect 16158 26126 16210 26178
rect 17838 26126 17890 26178
rect 19182 26126 19234 26178
rect 21086 26126 21138 26178
rect 23326 26126 23378 26178
rect 29150 26126 29202 26178
rect 33182 26126 33234 26178
rect 38558 26126 38610 26178
rect 39902 26126 39954 26178
rect 41358 26126 41410 26178
rect 49646 26126 49698 26178
rect 50094 26126 50146 26178
rect 50878 26126 50930 26178
rect 51550 26126 51602 26178
rect 53006 26126 53058 26178
rect 55134 26126 55186 26178
rect 7198 26014 7250 26066
rect 7758 26014 7810 26066
rect 21870 26014 21922 26066
rect 38894 26014 38946 26066
rect 39230 26014 39282 26066
rect 47518 26014 47570 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 13582 25678 13634 25730
rect 13918 25678 13970 25730
rect 23438 25678 23490 25730
rect 49758 25678 49810 25730
rect 50094 25678 50146 25730
rect 6974 25566 7026 25618
rect 9102 25566 9154 25618
rect 10222 25566 10274 25618
rect 12350 25566 12402 25618
rect 16046 25566 16098 25618
rect 18174 25566 18226 25618
rect 24446 25566 24498 25618
rect 30718 25566 30770 25618
rect 32846 25566 32898 25618
rect 33630 25566 33682 25618
rect 38446 25566 38498 25618
rect 40574 25566 40626 25618
rect 42478 25566 42530 25618
rect 43262 25566 43314 25618
rect 45838 25566 45890 25618
rect 46734 25566 46786 25618
rect 47742 25566 47794 25618
rect 52894 25566 52946 25618
rect 54686 25566 54738 25618
rect 6302 25454 6354 25506
rect 9550 25454 9602 25506
rect 15262 25454 15314 25506
rect 18734 25454 18786 25506
rect 18846 25454 18898 25506
rect 20750 25454 20802 25506
rect 21422 25454 21474 25506
rect 22094 25454 22146 25506
rect 22766 25454 22818 25506
rect 23102 25454 23154 25506
rect 23774 25454 23826 25506
rect 23998 25454 24050 25506
rect 27918 25454 27970 25506
rect 28254 25454 28306 25506
rect 29934 25454 29986 25506
rect 34190 25454 34242 25506
rect 36430 25454 36482 25506
rect 36990 25454 37042 25506
rect 37662 25454 37714 25506
rect 41918 25454 41970 25506
rect 42366 25454 42418 25506
rect 43150 25454 43202 25506
rect 44830 25454 44882 25506
rect 45278 25454 45330 25506
rect 45502 25454 45554 25506
rect 47518 25454 47570 25506
rect 47966 25454 48018 25506
rect 48078 25454 48130 25506
rect 48862 25454 48914 25506
rect 49982 25454 50034 25506
rect 50430 25454 50482 25506
rect 50878 25454 50930 25506
rect 51102 25454 51154 25506
rect 52110 25454 52162 25506
rect 52670 25454 52722 25506
rect 53566 25454 53618 25506
rect 14142 25342 14194 25394
rect 14478 25342 14530 25394
rect 18510 25342 18562 25394
rect 19742 25342 19794 25394
rect 20190 25342 20242 25394
rect 22542 25342 22594 25394
rect 22990 25342 23042 25394
rect 33966 25342 34018 25394
rect 34862 25342 34914 25394
rect 37326 25342 37378 25394
rect 41022 25342 41074 25394
rect 41694 25342 41746 25394
rect 46398 25342 46450 25394
rect 51438 25342 51490 25394
rect 51998 25342 52050 25394
rect 12798 25230 12850 25282
rect 21534 25230 21586 25282
rect 24894 25230 24946 25282
rect 27582 25230 27634 25282
rect 28590 25230 28642 25282
rect 29598 25230 29650 25282
rect 37214 25230 37266 25282
rect 41918 25230 41970 25282
rect 45390 25230 45442 25282
rect 47294 25230 47346 25282
rect 48638 25230 48690 25282
rect 48974 25230 49026 25282
rect 49086 25230 49138 25282
rect 50094 25230 50146 25282
rect 50766 25230 50818 25282
rect 54238 25230 54290 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 6078 24894 6130 24946
rect 7758 24894 7810 24946
rect 9662 24894 9714 24946
rect 11678 24894 11730 24946
rect 18398 24894 18450 24946
rect 26238 24894 26290 24946
rect 41022 24894 41074 24946
rect 41134 24894 41186 24946
rect 44718 24894 44770 24946
rect 53678 24894 53730 24946
rect 54126 24894 54178 24946
rect 2718 24782 2770 24834
rect 3390 24782 3442 24834
rect 7198 24782 7250 24834
rect 8878 24782 8930 24834
rect 14030 24782 14082 24834
rect 18846 24782 18898 24834
rect 22206 24782 22258 24834
rect 24558 24782 24610 24834
rect 28702 24782 28754 24834
rect 30158 24782 30210 24834
rect 37886 24782 37938 24834
rect 39118 24782 39170 24834
rect 45726 24782 45778 24834
rect 46622 24782 46674 24834
rect 2942 24670 2994 24722
rect 3726 24670 3778 24722
rect 6414 24670 6466 24722
rect 6862 24670 6914 24722
rect 8094 24670 8146 24722
rect 8654 24670 8706 24722
rect 12014 24670 12066 24722
rect 13806 24670 13858 24722
rect 17950 24670 18002 24722
rect 19854 24670 19906 24722
rect 22766 24670 22818 24722
rect 23438 24670 23490 24722
rect 24446 24670 24498 24722
rect 24782 24670 24834 24722
rect 25678 24670 25730 24722
rect 29374 24670 29426 24722
rect 29934 24670 29986 24722
rect 36318 24670 36370 24722
rect 37214 24670 37266 24722
rect 38558 24670 38610 24722
rect 40910 24670 40962 24722
rect 41470 24670 41522 24722
rect 42254 24670 42306 24722
rect 42814 24670 42866 24722
rect 44942 24670 44994 24722
rect 46846 24670 46898 24722
rect 47294 24670 47346 24722
rect 47518 24670 47570 24722
rect 47742 24670 47794 24722
rect 48750 24670 48802 24722
rect 49086 24670 49138 24722
rect 50654 24670 50706 24722
rect 52110 24670 52162 24722
rect 12462 24558 12514 24610
rect 13134 24558 13186 24610
rect 14926 24558 14978 24610
rect 17502 24558 17554 24610
rect 20078 24558 20130 24610
rect 22430 24558 22482 24610
rect 25230 24558 25282 24610
rect 26574 24558 26626 24610
rect 33966 24558 34018 24610
rect 35758 24558 35810 24610
rect 40014 24558 40066 24610
rect 41918 24558 41970 24610
rect 47070 24558 47122 24610
rect 48862 24558 48914 24610
rect 52222 24558 52274 24610
rect 48078 24446 48130 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 12350 24110 12402 24162
rect 25566 24110 25618 24162
rect 41806 24110 41858 24162
rect 43262 24110 43314 24162
rect 45390 24110 45442 24162
rect 50318 24110 50370 24162
rect 2942 23998 2994 24050
rect 5070 23998 5122 24050
rect 5742 23998 5794 24050
rect 7310 23998 7362 24050
rect 9550 23998 9602 24050
rect 12910 23998 12962 24050
rect 14254 23998 14306 24050
rect 16382 23998 16434 24050
rect 18734 23998 18786 24050
rect 24334 23998 24386 24050
rect 33182 23998 33234 24050
rect 36094 23998 36146 24050
rect 42590 23998 42642 24050
rect 46286 23998 46338 24050
rect 47182 23998 47234 24050
rect 47630 23998 47682 24050
rect 48750 23998 48802 24050
rect 54350 23998 54402 24050
rect 2270 23886 2322 23938
rect 7646 23886 7698 23938
rect 7982 23886 8034 23938
rect 12686 23886 12738 23938
rect 13470 23886 13522 23938
rect 18398 23886 18450 23938
rect 20750 23886 20802 23938
rect 22990 23886 23042 23938
rect 23214 23886 23266 23938
rect 24894 23886 24946 23938
rect 25342 23886 25394 23938
rect 26126 23886 26178 23938
rect 29262 23886 29314 23938
rect 34302 23886 34354 23938
rect 34638 23886 34690 23938
rect 35198 23886 35250 23938
rect 35646 23886 35698 23938
rect 36990 23886 37042 23938
rect 40798 23886 40850 23938
rect 41358 23886 41410 23938
rect 41806 23886 41858 23938
rect 42254 23886 42306 23938
rect 43822 23886 43874 23938
rect 43934 23886 43986 23938
rect 44942 23886 44994 23938
rect 45166 23886 45218 23938
rect 45950 23886 46002 23938
rect 46510 23886 46562 23938
rect 47518 23886 47570 23938
rect 48302 23886 48354 23938
rect 49086 23886 49138 23938
rect 49534 23886 49586 23938
rect 51102 23886 51154 23938
rect 51662 23886 51714 23938
rect 53342 23886 53394 23938
rect 53902 23886 53954 23938
rect 18062 23774 18114 23826
rect 19070 23774 19122 23826
rect 22766 23774 22818 23826
rect 23998 23774 24050 23826
rect 36206 23774 36258 23826
rect 37102 23774 37154 23826
rect 40686 23774 40738 23826
rect 43710 23774 43762 23826
rect 45614 23774 45666 23826
rect 49198 23774 49250 23826
rect 49758 23774 49810 23826
rect 49870 23774 49922 23826
rect 51774 23774 51826 23826
rect 52670 23774 52722 23826
rect 52894 23774 52946 23826
rect 53566 23774 53618 23826
rect 7422 23662 7474 23714
rect 7870 23662 7922 23714
rect 8542 23662 8594 23714
rect 9662 23662 9714 23714
rect 26350 23662 26402 23714
rect 27918 23662 27970 23714
rect 28366 23662 28418 23714
rect 29486 23662 29538 23714
rect 37214 23662 37266 23714
rect 45502 23662 45554 23714
rect 53006 23662 53058 23714
rect 53678 23662 53730 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 5406 23326 5458 23378
rect 13582 23326 13634 23378
rect 21870 23326 21922 23378
rect 23438 23326 23490 23378
rect 33630 23326 33682 23378
rect 34974 23326 35026 23378
rect 38446 23326 38498 23378
rect 39006 23326 39058 23378
rect 41358 23326 41410 23378
rect 42590 23326 42642 23378
rect 47406 23326 47458 23378
rect 48190 23326 48242 23378
rect 2606 23214 2658 23266
rect 6414 23214 6466 23266
rect 7534 23214 7586 23266
rect 7646 23214 7698 23266
rect 8206 23214 8258 23266
rect 15262 23214 15314 23266
rect 16382 23214 16434 23266
rect 16718 23214 16770 23266
rect 17502 23214 17554 23266
rect 19854 23214 19906 23266
rect 20974 23214 21026 23266
rect 23886 23214 23938 23266
rect 27358 23214 27410 23266
rect 30718 23214 30770 23266
rect 33854 23214 33906 23266
rect 38558 23214 38610 23266
rect 42030 23214 42082 23266
rect 42926 23214 42978 23266
rect 44718 23214 44770 23266
rect 45726 23214 45778 23266
rect 50430 23214 50482 23266
rect 1934 23102 1986 23154
rect 6526 23102 6578 23154
rect 7310 23102 7362 23154
rect 9662 23102 9714 23154
rect 13694 23102 13746 23154
rect 14478 23102 14530 23154
rect 15150 23102 15202 23154
rect 18062 23102 18114 23154
rect 20526 23102 20578 23154
rect 23326 23102 23378 23154
rect 23662 23102 23714 23154
rect 28142 23102 28194 23154
rect 31390 23102 31442 23154
rect 34078 23102 34130 23154
rect 34526 23102 34578 23154
rect 37438 23102 37490 23154
rect 39790 23102 39842 23154
rect 39902 23102 39954 23154
rect 41694 23102 41746 23154
rect 41806 23102 41858 23154
rect 42366 23102 42418 23154
rect 43710 23102 43762 23154
rect 45166 23102 45218 23154
rect 45950 23102 46002 23154
rect 46398 23102 46450 23154
rect 47182 23102 47234 23154
rect 47742 23102 47794 23154
rect 49310 23102 49362 23154
rect 49646 23102 49698 23154
rect 50094 23102 50146 23154
rect 50878 23102 50930 23154
rect 4734 22990 4786 23042
rect 8766 22990 8818 23042
rect 10334 22990 10386 23042
rect 12462 22990 12514 23042
rect 13134 22990 13186 23042
rect 15822 22990 15874 23042
rect 19630 22990 19682 23042
rect 22206 22990 22258 23042
rect 24110 22990 24162 23042
rect 25230 22990 25282 23042
rect 28590 22990 28642 23042
rect 34302 22990 34354 23042
rect 35086 22990 35138 23042
rect 36318 22990 36370 23042
rect 39566 22990 39618 23042
rect 46174 22990 46226 23042
rect 46734 22990 46786 23042
rect 47294 22990 47346 23042
rect 48750 22990 48802 23042
rect 51550 22990 51602 23042
rect 53678 22990 53730 23042
rect 5742 22878 5794 22930
rect 7982 22878 8034 22930
rect 8318 22878 8370 22930
rect 13582 22878 13634 22930
rect 14142 22878 14194 22930
rect 18286 22878 18338 22930
rect 19742 22878 19794 22930
rect 24446 22878 24498 22930
rect 34750 22878 34802 22930
rect 38334 22878 38386 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 6078 22542 6130 22594
rect 7310 22542 7362 22594
rect 11790 22542 11842 22594
rect 14030 22542 14082 22594
rect 14366 22542 14418 22594
rect 20302 22542 20354 22594
rect 20638 22542 20690 22594
rect 21758 22542 21810 22594
rect 22542 22542 22594 22594
rect 26574 22542 26626 22594
rect 26910 22542 26962 22594
rect 29262 22542 29314 22594
rect 46622 22542 46674 22594
rect 46958 22542 47010 22594
rect 47518 22542 47570 22594
rect 51438 22542 51490 22594
rect 52670 22542 52722 22594
rect 5070 22430 5122 22482
rect 13694 22430 13746 22482
rect 18510 22430 18562 22482
rect 21534 22430 21586 22482
rect 25678 22430 25730 22482
rect 28478 22430 28530 22482
rect 29598 22430 29650 22482
rect 34078 22430 34130 22482
rect 36206 22430 36258 22482
rect 37102 22430 37154 22482
rect 40350 22430 40402 22482
rect 42590 22430 42642 22482
rect 44270 22430 44322 22482
rect 44830 22430 44882 22482
rect 45726 22430 45778 22482
rect 47182 22430 47234 22482
rect 47854 22430 47906 22482
rect 48414 22430 48466 22482
rect 49646 22430 49698 22482
rect 50430 22430 50482 22482
rect 50878 22430 50930 22482
rect 5742 22318 5794 22370
rect 6526 22318 6578 22370
rect 10670 22318 10722 22370
rect 11454 22318 11506 22370
rect 12574 22318 12626 22370
rect 17950 22318 18002 22370
rect 18846 22318 18898 22370
rect 19182 22318 19234 22370
rect 20526 22318 20578 22370
rect 22430 22318 22482 22370
rect 22878 22318 22930 22370
rect 23102 22318 23154 22370
rect 23774 22318 23826 22370
rect 24222 22318 24274 22370
rect 27694 22318 27746 22370
rect 31166 22318 31218 22370
rect 34638 22318 34690 22370
rect 35534 22318 35586 22370
rect 35758 22318 35810 22370
rect 35982 22318 36034 22370
rect 37326 22318 37378 22370
rect 37998 22318 38050 22370
rect 38222 22318 38274 22370
rect 40574 22318 40626 22370
rect 40798 22318 40850 22370
rect 43486 22318 43538 22370
rect 43710 22318 43762 22370
rect 45278 22318 45330 22370
rect 46062 22318 46114 22370
rect 48862 22318 48914 22370
rect 51214 22318 51266 22370
rect 51774 22318 51826 22370
rect 52782 22318 52834 22370
rect 3614 22206 3666 22258
rect 6862 22206 6914 22258
rect 10334 22206 10386 22258
rect 12462 22206 12514 22258
rect 14590 22206 14642 22258
rect 14926 22206 14978 22258
rect 16718 22206 16770 22258
rect 17166 22206 17218 22258
rect 18062 22206 18114 22258
rect 18398 22206 18450 22258
rect 19070 22206 19122 22258
rect 19742 22206 19794 22258
rect 23326 22206 23378 22258
rect 24894 22206 24946 22258
rect 25230 22206 25282 22258
rect 27470 22206 27522 22258
rect 29822 22206 29874 22258
rect 30382 22206 30434 22258
rect 31950 22206 32002 22258
rect 36430 22206 36482 22258
rect 40350 22206 40402 22258
rect 41582 22206 41634 22258
rect 43374 22206 43426 22258
rect 45838 22206 45890 22258
rect 47630 22206 47682 22258
rect 48302 22206 48354 22258
rect 48526 22206 48578 22258
rect 49198 22206 49250 22258
rect 51998 22206 52050 22258
rect 3278 22094 3330 22146
rect 7422 22094 7474 22146
rect 7534 22094 7586 22146
rect 15710 22094 15762 22146
rect 16046 22094 16098 22146
rect 16382 22094 16434 22146
rect 17502 22094 17554 22146
rect 22094 22094 22146 22146
rect 22990 22094 23042 22146
rect 23886 22094 23938 22146
rect 25006 22094 25058 22146
rect 25790 22094 25842 22146
rect 28590 22094 28642 22146
rect 34414 22094 34466 22146
rect 35198 22094 35250 22146
rect 36542 22094 36594 22146
rect 42926 22094 42978 22146
rect 51662 22094 51714 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 7758 21758 7810 21810
rect 8878 21758 8930 21810
rect 14590 21758 14642 21810
rect 20302 21758 20354 21810
rect 20750 21758 20802 21810
rect 21422 21758 21474 21810
rect 22654 21758 22706 21810
rect 27022 21758 27074 21810
rect 27694 21758 27746 21810
rect 28478 21758 28530 21810
rect 30270 21758 30322 21810
rect 32062 21758 32114 21810
rect 34974 21758 35026 21810
rect 35198 21758 35250 21810
rect 35534 21758 35586 21810
rect 35758 21758 35810 21810
rect 39230 21758 39282 21810
rect 45166 21758 45218 21810
rect 46846 21758 46898 21810
rect 47406 21758 47458 21810
rect 47854 21758 47906 21810
rect 3054 21646 3106 21698
rect 6974 21646 7026 21698
rect 8094 21646 8146 21698
rect 10558 21646 10610 21698
rect 10894 21646 10946 21698
rect 11118 21646 11170 21698
rect 11678 21646 11730 21698
rect 12126 21646 12178 21698
rect 13806 21646 13858 21698
rect 15934 21646 15986 21698
rect 19070 21646 19122 21698
rect 20190 21646 20242 21698
rect 20862 21646 20914 21698
rect 21646 21646 21698 21698
rect 22318 21646 22370 21698
rect 22990 21646 23042 21698
rect 24558 21646 24610 21698
rect 25566 21646 25618 21698
rect 26238 21646 26290 21698
rect 28030 21646 28082 21698
rect 29822 21646 29874 21698
rect 33742 21646 33794 21698
rect 34078 21646 34130 21698
rect 35310 21646 35362 21698
rect 35870 21646 35922 21698
rect 36990 21646 37042 21698
rect 40350 21646 40402 21698
rect 40910 21646 40962 21698
rect 44382 21646 44434 21698
rect 47966 21646 48018 21698
rect 2270 21534 2322 21586
rect 7198 21534 7250 21586
rect 7422 21534 7474 21586
rect 7758 21534 7810 21586
rect 8318 21534 8370 21586
rect 8542 21534 8594 21586
rect 8654 21534 8706 21586
rect 12350 21534 12402 21586
rect 14030 21534 14082 21586
rect 14254 21534 14306 21586
rect 14366 21534 14418 21586
rect 16158 21534 16210 21586
rect 16718 21534 16770 21586
rect 19182 21534 19234 21586
rect 20526 21534 20578 21586
rect 24334 21534 24386 21586
rect 25230 21534 25282 21586
rect 26574 21534 26626 21586
rect 29598 21534 29650 21586
rect 32398 21534 32450 21586
rect 33182 21534 33234 21586
rect 36318 21534 36370 21586
rect 39790 21534 39842 21586
rect 42142 21534 42194 21586
rect 42478 21534 42530 21586
rect 42926 21534 42978 21586
rect 43150 21534 43202 21586
rect 43710 21534 43762 21586
rect 43934 21534 43986 21586
rect 44494 21534 44546 21586
rect 47182 21534 47234 21586
rect 47630 21534 47682 21586
rect 5182 21422 5234 21474
rect 5630 21422 5682 21474
rect 13246 21422 13298 21474
rect 21534 21422 21586 21474
rect 25902 21422 25954 21474
rect 30830 21422 30882 21474
rect 40238 21422 40290 21474
rect 43038 21422 43090 21474
rect 43374 21422 43426 21474
rect 44158 21422 44210 21474
rect 45278 21422 45330 21474
rect 50878 21422 50930 21474
rect 5406 21310 5458 21362
rect 5742 21310 5794 21362
rect 10782 21310 10834 21362
rect 12686 21310 12738 21362
rect 18174 21310 18226 21362
rect 18510 21310 18562 21362
rect 23102 21310 23154 21362
rect 23998 21310 24050 21362
rect 33518 21310 33570 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 5742 20974 5794 21026
rect 9102 20974 9154 21026
rect 10110 20974 10162 21026
rect 13918 20974 13970 21026
rect 38222 20974 38274 21026
rect 38446 20974 38498 21026
rect 38558 20974 38610 21026
rect 43598 20974 43650 21026
rect 4622 20862 4674 20914
rect 8094 20862 8146 20914
rect 11342 20862 11394 20914
rect 19742 20862 19794 20914
rect 22654 20862 22706 20914
rect 23438 20862 23490 20914
rect 25790 20862 25842 20914
rect 27918 20862 27970 20914
rect 37326 20862 37378 20914
rect 37662 20862 37714 20914
rect 39678 20862 39730 20914
rect 41806 20862 41858 20914
rect 42254 20862 42306 20914
rect 42814 20862 42866 20914
rect 43598 20862 43650 20914
rect 45614 20862 45666 20914
rect 47742 20862 47794 20914
rect 48190 20862 48242 20914
rect 1822 20750 1874 20802
rect 6078 20750 6130 20802
rect 7646 20750 7698 20802
rect 8206 20750 8258 20802
rect 9102 20750 9154 20802
rect 9662 20750 9714 20802
rect 10222 20750 10274 20802
rect 11006 20750 11058 20802
rect 13470 20750 13522 20802
rect 13694 20750 13746 20802
rect 14030 20750 14082 20802
rect 15150 20750 15202 20802
rect 15374 20750 15426 20802
rect 15598 20750 15650 20802
rect 16942 20750 16994 20802
rect 20638 20750 20690 20802
rect 22990 20750 23042 20802
rect 24110 20750 24162 20802
rect 25118 20750 25170 20802
rect 29374 20750 29426 20802
rect 32846 20750 32898 20802
rect 34526 20750 34578 20802
rect 35198 20750 35250 20802
rect 35534 20750 35586 20802
rect 38110 20750 38162 20802
rect 39006 20750 39058 20802
rect 42142 20750 42194 20802
rect 42366 20750 42418 20802
rect 42814 20750 42866 20802
rect 44942 20750 44994 20802
rect 2494 20638 2546 20690
rect 6302 20638 6354 20690
rect 6750 20638 6802 20690
rect 7870 20638 7922 20690
rect 8766 20638 8818 20690
rect 9886 20638 9938 20690
rect 10558 20638 10610 20690
rect 10894 20638 10946 20690
rect 11230 20638 11282 20690
rect 17614 20638 17666 20690
rect 20302 20638 20354 20690
rect 23662 20638 23714 20690
rect 33070 20638 33122 20690
rect 33630 20638 33682 20690
rect 35758 20638 35810 20690
rect 36094 20638 36146 20690
rect 5070 20526 5122 20578
rect 8094 20526 8146 20578
rect 10110 20526 10162 20578
rect 13582 20526 13634 20578
rect 16382 20526 16434 20578
rect 20526 20526 20578 20578
rect 21422 20526 21474 20578
rect 24558 20526 24610 20578
rect 28366 20526 28418 20578
rect 29150 20526 29202 20578
rect 32510 20526 32562 20578
rect 34750 20526 34802 20578
rect 43262 20526 43314 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 2494 20190 2546 20242
rect 11006 20190 11058 20242
rect 15934 20190 15986 20242
rect 17502 20190 17554 20242
rect 22206 20190 22258 20242
rect 22766 20190 22818 20242
rect 26798 20190 26850 20242
rect 39118 20190 39170 20242
rect 41246 20190 41298 20242
rect 48190 20190 48242 20242
rect 5966 20078 6018 20130
rect 7086 20078 7138 20130
rect 7310 20078 7362 20130
rect 7982 20078 8034 20130
rect 13806 20078 13858 20130
rect 17838 20078 17890 20130
rect 19294 20078 19346 20130
rect 21422 20078 21474 20130
rect 21534 20078 21586 20130
rect 21646 20078 21698 20130
rect 22094 20078 22146 20130
rect 22430 20078 22482 20130
rect 24110 20078 24162 20130
rect 24558 20078 24610 20130
rect 25566 20078 25618 20130
rect 27694 20078 27746 20130
rect 29150 20078 29202 20130
rect 32062 20078 32114 20130
rect 32398 20078 32450 20130
rect 35310 20078 35362 20130
rect 40350 20078 40402 20130
rect 41134 20078 41186 20130
rect 45614 20078 45666 20130
rect 2830 19966 2882 20018
rect 5070 19966 5122 20018
rect 5406 19966 5458 20018
rect 6190 19966 6242 20018
rect 10558 19966 10610 20018
rect 10782 19966 10834 20018
rect 11006 19966 11058 20018
rect 11118 19966 11170 20018
rect 14142 19966 14194 20018
rect 14702 19966 14754 20018
rect 14926 19966 14978 20018
rect 15822 19966 15874 20018
rect 16046 19966 16098 20018
rect 19182 19966 19234 20018
rect 23102 19966 23154 20018
rect 24222 19966 24274 20018
rect 24670 19966 24722 20018
rect 25230 19966 25282 20018
rect 27134 19966 27186 20018
rect 27918 19966 27970 20018
rect 28366 19966 28418 20018
rect 34638 19966 34690 20018
rect 39790 19966 39842 20018
rect 44942 19966 44994 20018
rect 7422 19854 7474 19906
rect 14814 19854 14866 19906
rect 15598 19854 15650 19906
rect 18174 19854 18226 19906
rect 18734 19854 18786 19906
rect 20862 19854 20914 19906
rect 23550 19854 23602 19906
rect 25902 19854 25954 19906
rect 31278 19854 31330 19906
rect 34302 19854 34354 19906
rect 37438 19854 37490 19906
rect 37886 19854 37938 19906
rect 38558 19854 38610 19906
rect 39454 19854 39506 19906
rect 47742 19854 47794 19906
rect 7646 19742 7698 19794
rect 8094 19742 8146 19794
rect 13358 19742 13410 19794
rect 13470 19742 13522 19794
rect 13694 19742 13746 19794
rect 14366 19742 14418 19794
rect 18510 19742 18562 19794
rect 19966 19742 20018 19794
rect 20302 19742 20354 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 11118 19406 11170 19458
rect 12574 19406 12626 19458
rect 14926 19406 14978 19458
rect 15262 19406 15314 19458
rect 23550 19406 23602 19458
rect 27022 19406 27074 19458
rect 29262 19406 29314 19458
rect 29598 19406 29650 19458
rect 7198 19294 7250 19346
rect 23326 19294 23378 19346
rect 24334 19294 24386 19346
rect 26686 19294 26738 19346
rect 31950 19294 32002 19346
rect 34078 19294 34130 19346
rect 37214 19294 37266 19346
rect 8430 19182 8482 19234
rect 9774 19182 9826 19234
rect 11006 19182 11058 19234
rect 11342 19182 11394 19234
rect 12686 19182 12738 19234
rect 14254 19182 14306 19234
rect 14702 19182 14754 19234
rect 15150 19182 15202 19234
rect 16158 19182 16210 19234
rect 16494 19182 16546 19234
rect 19182 19182 19234 19234
rect 19854 19182 19906 19234
rect 21982 19182 22034 19234
rect 22318 19182 22370 19234
rect 31166 19182 31218 19234
rect 35534 19182 35586 19234
rect 4062 19070 4114 19122
rect 6862 19070 6914 19122
rect 7086 19070 7138 19122
rect 7646 19070 7698 19122
rect 7758 19070 7810 19122
rect 8094 19070 8146 19122
rect 8766 19070 8818 19122
rect 9102 19070 9154 19122
rect 9998 19070 10050 19122
rect 10670 19070 10722 19122
rect 12126 19070 12178 19122
rect 12350 19070 12402 19122
rect 14030 19070 14082 19122
rect 22654 19070 22706 19122
rect 26798 19070 26850 19122
rect 29822 19070 29874 19122
rect 30382 19070 30434 19122
rect 35758 19070 35810 19122
rect 36094 19070 36146 19122
rect 3726 18958 3778 19010
rect 5742 18958 5794 19010
rect 7422 18958 7474 19010
rect 8206 18958 8258 19010
rect 10894 18958 10946 19010
rect 12910 18958 12962 19010
rect 15822 18958 15874 19010
rect 16606 18958 16658 19010
rect 19406 18958 19458 19010
rect 21646 18958 21698 19010
rect 23886 18958 23938 19010
rect 24894 18958 24946 19010
rect 28030 18958 28082 19010
rect 35198 18958 35250 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 8318 18622 8370 18674
rect 9998 18622 10050 18674
rect 11566 18622 11618 18674
rect 13022 18622 13074 18674
rect 14366 18622 14418 18674
rect 23214 18622 23266 18674
rect 25230 18622 25282 18674
rect 30830 18622 30882 18674
rect 2270 18510 2322 18562
rect 3390 18510 3442 18562
rect 6862 18510 6914 18562
rect 7534 18510 7586 18562
rect 8990 18510 9042 18562
rect 9550 18510 9602 18562
rect 14478 18510 14530 18562
rect 15374 18510 15426 18562
rect 19518 18510 19570 18562
rect 23550 18510 23602 18562
rect 24222 18510 24274 18562
rect 26014 18510 26066 18562
rect 29710 18510 29762 18562
rect 29934 18510 29986 18562
rect 34078 18510 34130 18562
rect 35198 18510 35250 18562
rect 2046 18398 2098 18450
rect 2718 18398 2770 18450
rect 5966 18398 6018 18450
rect 6302 18398 6354 18450
rect 7086 18398 7138 18450
rect 7758 18398 7810 18450
rect 7982 18398 8034 18450
rect 8318 18398 8370 18450
rect 8766 18398 8818 18450
rect 9774 18398 9826 18450
rect 10110 18398 10162 18450
rect 11118 18398 11170 18450
rect 11342 18398 11394 18450
rect 11566 18398 11618 18450
rect 11678 18398 11730 18450
rect 12238 18398 12290 18450
rect 12462 18398 12514 18450
rect 12686 18398 12738 18450
rect 12798 18398 12850 18450
rect 13694 18398 13746 18450
rect 14142 18398 14194 18450
rect 14814 18398 14866 18450
rect 15038 18398 15090 18450
rect 18734 18398 18786 18450
rect 22094 18398 22146 18450
rect 23998 18398 24050 18450
rect 25230 18398 25282 18450
rect 25566 18398 25618 18450
rect 25678 18398 25730 18450
rect 28366 18398 28418 18450
rect 33742 18398 33794 18450
rect 34974 18398 35026 18450
rect 37662 18398 37714 18450
rect 38446 18398 38498 18450
rect 5518 18286 5570 18338
rect 21646 18286 21698 18338
rect 35534 18286 35586 18338
rect 38894 18286 38946 18338
rect 10110 18174 10162 18226
rect 13918 18174 13970 18226
rect 15262 18174 15314 18226
rect 28030 18174 28082 18226
rect 28366 18174 28418 18226
rect 29598 18174 29650 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 5742 17838 5794 17890
rect 6078 17838 6130 17890
rect 12462 17838 12514 17890
rect 14030 17838 14082 17890
rect 14254 17838 14306 17890
rect 24446 17838 24498 17890
rect 25342 17838 25394 17890
rect 26350 17838 26402 17890
rect 29598 17838 29650 17890
rect 2494 17726 2546 17778
rect 4622 17726 4674 17778
rect 9886 17726 9938 17778
rect 17166 17726 17218 17778
rect 27694 17726 27746 17778
rect 33406 17726 33458 17778
rect 35534 17726 35586 17778
rect 1822 17614 1874 17666
rect 6862 17614 6914 17666
rect 8766 17614 8818 17666
rect 9438 17614 9490 17666
rect 12350 17614 12402 17666
rect 12574 17614 12626 17666
rect 13806 17614 13858 17666
rect 16606 17614 16658 17666
rect 21534 17614 21586 17666
rect 22542 17614 22594 17666
rect 24110 17614 24162 17666
rect 26126 17614 26178 17666
rect 26462 17614 26514 17666
rect 29150 17614 29202 17666
rect 29374 17614 29426 17666
rect 29710 17614 29762 17666
rect 32174 17614 32226 17666
rect 36206 17614 36258 17666
rect 37102 17614 37154 17666
rect 6750 17502 6802 17554
rect 8430 17502 8482 17554
rect 9102 17502 9154 17554
rect 11342 17502 11394 17554
rect 12014 17502 12066 17554
rect 15598 17502 15650 17554
rect 15934 17502 15986 17554
rect 16382 17502 16434 17554
rect 22990 17502 23042 17554
rect 23326 17502 23378 17554
rect 24670 17502 24722 17554
rect 24894 17502 24946 17554
rect 25454 17502 25506 17554
rect 26798 17502 26850 17554
rect 30382 17502 30434 17554
rect 31838 17502 31890 17554
rect 32398 17502 32450 17554
rect 32734 17502 32786 17554
rect 5070 17390 5122 17442
rect 11678 17390 11730 17442
rect 12798 17390 12850 17442
rect 13918 17390 13970 17442
rect 21198 17390 21250 17442
rect 21422 17390 21474 17442
rect 21982 17390 22034 17442
rect 22318 17390 22370 17442
rect 24110 17390 24162 17442
rect 25342 17390 25394 17442
rect 26686 17390 26738 17442
rect 27134 17390 27186 17442
rect 29262 17390 29314 17442
rect 30718 17390 30770 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 6302 17054 6354 17106
rect 7086 17054 7138 17106
rect 8094 17054 8146 17106
rect 8542 17054 8594 17106
rect 10334 17054 10386 17106
rect 11006 17054 11058 17106
rect 13358 17054 13410 17106
rect 13694 17054 13746 17106
rect 14814 17054 14866 17106
rect 15374 17054 15426 17106
rect 16494 17054 16546 17106
rect 20750 17054 20802 17106
rect 22878 17054 22930 17106
rect 23214 17054 23266 17106
rect 23774 17054 23826 17106
rect 24782 17054 24834 17106
rect 33630 17054 33682 17106
rect 7758 16942 7810 16994
rect 15038 16942 15090 16994
rect 16158 16942 16210 16994
rect 16830 16942 16882 16994
rect 23998 16942 24050 16994
rect 24558 16942 24610 16994
rect 26014 16942 26066 16994
rect 28142 16942 28194 16994
rect 28366 16942 28418 16994
rect 31726 16942 31778 16994
rect 34190 16942 34242 16994
rect 34526 16942 34578 16994
rect 6974 16830 7026 16882
rect 15934 16830 15986 16882
rect 17502 16830 17554 16882
rect 23550 16830 23602 16882
rect 24446 16830 24498 16882
rect 27806 16830 27858 16882
rect 28590 16830 28642 16882
rect 28702 16830 28754 16882
rect 32510 16830 32562 16882
rect 33182 16830 33234 16882
rect 6190 16718 6242 16770
rect 10222 16718 10274 16770
rect 11118 16718 11170 16770
rect 18174 16718 18226 16770
rect 20302 16718 20354 16770
rect 23662 16718 23714 16770
rect 28254 16718 28306 16770
rect 29598 16718 29650 16770
rect 33966 16606 34018 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 14926 16270 14978 16322
rect 16158 16270 16210 16322
rect 19518 16270 19570 16322
rect 26350 16270 26402 16322
rect 26686 16270 26738 16322
rect 29486 16270 29538 16322
rect 30382 16270 30434 16322
rect 30718 16270 30770 16322
rect 11342 16158 11394 16210
rect 11790 16158 11842 16210
rect 17502 16158 17554 16210
rect 23998 16158 24050 16210
rect 24894 16158 24946 16210
rect 25790 16158 25842 16210
rect 6078 16046 6130 16098
rect 6862 16046 6914 16098
rect 7198 16046 7250 16098
rect 7534 16046 7586 16098
rect 7870 16046 7922 16098
rect 8542 16046 8594 16098
rect 12798 16046 12850 16098
rect 14142 16046 14194 16098
rect 15150 16046 15202 16098
rect 15822 16046 15874 16098
rect 17054 16046 17106 16098
rect 20302 16046 20354 16098
rect 22878 16046 22930 16098
rect 25230 16046 25282 16098
rect 25678 16046 25730 16098
rect 27358 16046 27410 16098
rect 29150 16046 29202 16098
rect 35534 16046 35586 16098
rect 4062 15934 4114 15986
rect 6750 15934 6802 15986
rect 7422 15934 7474 15986
rect 9214 15934 9266 15986
rect 13806 15934 13858 15986
rect 16270 15934 16322 15986
rect 16718 15934 16770 15986
rect 18286 15934 18338 15986
rect 18622 15934 18674 15986
rect 19182 15934 19234 15986
rect 20078 15934 20130 15986
rect 23662 15934 23714 15986
rect 24558 15934 24610 15986
rect 27470 15934 27522 15986
rect 29710 15934 29762 15986
rect 29934 15934 29986 15986
rect 30942 15934 30994 15986
rect 31278 15934 31330 15986
rect 35758 15934 35810 15986
rect 36318 15934 36370 15986
rect 3726 15822 3778 15874
rect 5742 15822 5794 15874
rect 7982 15822 8034 15874
rect 8206 15822 8258 15874
rect 12238 15822 12290 15874
rect 12462 15822 12514 15874
rect 12686 15822 12738 15874
rect 13582 15822 13634 15874
rect 14590 15822 14642 15874
rect 15486 15822 15538 15874
rect 22654 15822 22706 15874
rect 23214 15822 23266 15874
rect 23886 15822 23938 15874
rect 24110 15822 24162 15874
rect 24782 15822 24834 15874
rect 25006 15822 25058 15874
rect 25902 15822 25954 15874
rect 28030 15822 28082 15874
rect 29150 15822 29202 15874
rect 35198 15822 35250 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 6078 15486 6130 15538
rect 7870 15486 7922 15538
rect 8990 15486 9042 15538
rect 13582 15486 13634 15538
rect 14478 15486 14530 15538
rect 15486 15486 15538 15538
rect 16158 15486 16210 15538
rect 16494 15486 16546 15538
rect 17390 15486 17442 15538
rect 23774 15486 23826 15538
rect 27246 15486 27298 15538
rect 2382 15374 2434 15426
rect 3502 15374 3554 15426
rect 7198 15374 7250 15426
rect 8430 15374 8482 15426
rect 13694 15374 13746 15426
rect 14926 15374 14978 15426
rect 16830 15374 16882 15426
rect 17726 15374 17778 15426
rect 26238 15374 26290 15426
rect 28590 15374 28642 15426
rect 29038 15374 29090 15426
rect 31390 15374 31442 15426
rect 31726 15374 31778 15426
rect 35422 15374 35474 15426
rect 37886 15374 37938 15426
rect 2158 15262 2210 15314
rect 2830 15262 2882 15314
rect 6414 15262 6466 15314
rect 6862 15262 6914 15314
rect 8766 15262 8818 15314
rect 9998 15262 10050 15314
rect 20190 15262 20242 15314
rect 24222 15262 24274 15314
rect 25678 15262 25730 15314
rect 26574 15262 26626 15314
rect 27022 15262 27074 15314
rect 27358 15262 27410 15314
rect 27918 15262 27970 15314
rect 28254 15262 28306 15314
rect 35086 15262 35138 15314
rect 38670 15262 38722 15314
rect 39118 15262 39170 15314
rect 5630 15150 5682 15202
rect 11790 15150 11842 15202
rect 12574 15150 12626 15202
rect 20862 15150 20914 15202
rect 22990 15150 23042 15202
rect 24558 15150 24610 15202
rect 25790 15150 25842 15202
rect 35758 15150 35810 15202
rect 13582 15038 13634 15090
rect 26798 15038 26850 15090
rect 30830 15038 30882 15090
rect 31166 15038 31218 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 11118 14702 11170 14754
rect 11454 14702 11506 14754
rect 28030 14702 28082 14754
rect 35198 14702 35250 14754
rect 2494 14590 2546 14642
rect 4622 14590 4674 14642
rect 5070 14590 5122 14642
rect 5854 14590 5906 14642
rect 9774 14590 9826 14642
rect 19854 14590 19906 14642
rect 22878 14590 22930 14642
rect 24446 14590 24498 14642
rect 31166 14590 31218 14642
rect 1822 14478 1874 14530
rect 6974 14478 7026 14530
rect 12238 14478 12290 14530
rect 14030 14478 14082 14530
rect 14478 14478 14530 14530
rect 16606 14478 16658 14530
rect 16942 14478 16994 14530
rect 20414 14478 20466 14530
rect 22206 14478 22258 14530
rect 22542 14478 22594 14530
rect 22766 14478 22818 14530
rect 23550 14478 23602 14530
rect 26238 14478 26290 14530
rect 26574 14478 26626 14530
rect 26798 14478 26850 14530
rect 27694 14478 27746 14530
rect 28254 14478 28306 14530
rect 28478 14478 28530 14530
rect 30606 14478 30658 14530
rect 33966 14478 34018 14530
rect 34526 14478 34578 14530
rect 35534 14478 35586 14530
rect 7646 14366 7698 14418
rect 10446 14366 10498 14418
rect 12014 14366 12066 14418
rect 13470 14366 13522 14418
rect 16046 14366 16098 14418
rect 17726 14366 17778 14418
rect 20638 14366 20690 14418
rect 22990 14366 23042 14418
rect 27022 14366 27074 14418
rect 30830 14366 30882 14418
rect 33294 14366 33346 14418
rect 35758 14366 35810 14418
rect 36094 14366 36146 14418
rect 10110 14254 10162 14306
rect 12910 14254 12962 14306
rect 14702 14254 14754 14306
rect 26238 14254 26290 14306
rect 27694 14254 27746 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 7982 13918 8034 13970
rect 9102 13918 9154 13970
rect 11454 13918 11506 13970
rect 16718 13918 16770 13970
rect 21422 13918 21474 13970
rect 22654 13918 22706 13970
rect 23998 13918 24050 13970
rect 25566 13918 25618 13970
rect 26686 13918 26738 13970
rect 27022 13918 27074 13970
rect 28814 13918 28866 13970
rect 29150 13918 29202 13970
rect 29486 13918 29538 13970
rect 33182 13918 33234 13970
rect 2606 13806 2658 13858
rect 6078 13806 6130 13858
rect 10782 13806 10834 13858
rect 12462 13806 12514 13858
rect 15150 13806 15202 13858
rect 19518 13806 19570 13858
rect 20302 13806 20354 13858
rect 26126 13806 26178 13858
rect 33742 13806 33794 13858
rect 34190 13806 34242 13858
rect 36318 13806 36370 13858
rect 36542 13806 36594 13858
rect 2942 13694 2994 13746
rect 6190 13694 6242 13746
rect 8318 13694 8370 13746
rect 9774 13694 9826 13746
rect 10110 13694 10162 13746
rect 10894 13694 10946 13746
rect 12574 13694 12626 13746
rect 15822 13694 15874 13746
rect 19742 13694 19794 13746
rect 20526 13694 20578 13746
rect 21086 13694 21138 13746
rect 21870 13694 21922 13746
rect 22206 13694 22258 13746
rect 22654 13694 22706 13746
rect 23550 13694 23602 13746
rect 23886 13694 23938 13746
rect 24110 13694 24162 13746
rect 25902 13694 25954 13746
rect 26462 13694 26514 13746
rect 27246 13694 27298 13746
rect 27470 13694 27522 13746
rect 27806 13694 27858 13746
rect 33518 13694 33570 13746
rect 35646 13694 35698 13746
rect 35982 13694 36034 13746
rect 13022 13582 13074 13634
rect 5070 13470 5122 13522
rect 5406 13470 5458 13522
rect 11790 13470 11842 13522
rect 18622 13470 18674 13522
rect 18958 13470 19010 13522
rect 22318 13470 22370 13522
rect 23998 13470 24050 13522
rect 26462 13470 26514 13522
rect 27358 13470 27410 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 5742 13134 5794 13186
rect 8654 13134 8706 13186
rect 8990 13134 9042 13186
rect 14366 13134 14418 13186
rect 14702 13134 14754 13186
rect 19070 13134 19122 13186
rect 20302 13134 20354 13186
rect 22206 13134 22258 13186
rect 24334 13134 24386 13186
rect 27022 13134 27074 13186
rect 2494 13022 2546 13074
rect 4622 13022 4674 13074
rect 6078 13022 6130 13074
rect 12574 13022 12626 13074
rect 21310 13022 21362 13074
rect 22318 13022 22370 13074
rect 25454 13022 25506 13074
rect 26238 13022 26290 13074
rect 29150 13022 29202 13074
rect 1822 12910 1874 12962
rect 7534 12910 7586 12962
rect 9550 12910 9602 12962
rect 10782 12910 10834 12962
rect 18286 12910 18338 12962
rect 19742 12910 19794 12962
rect 21646 12910 21698 12962
rect 22542 12910 22594 12962
rect 23438 12910 23490 12962
rect 23662 12910 23714 12962
rect 23774 12910 23826 12962
rect 25230 12910 25282 12962
rect 26686 12910 26738 12962
rect 27358 12910 27410 12962
rect 28366 12910 28418 12962
rect 32062 12910 32114 12962
rect 32510 12910 32562 12962
rect 36318 12910 36370 12962
rect 6302 12798 6354 12850
rect 6750 12798 6802 12850
rect 9774 12798 9826 12850
rect 13806 12798 13858 12850
rect 14030 12798 14082 12850
rect 17950 12798 18002 12850
rect 18958 12798 19010 12850
rect 19518 12798 19570 12850
rect 21870 12798 21922 12850
rect 22766 12798 22818 12850
rect 22990 12798 23042 12850
rect 23214 12798 23266 12850
rect 25790 12798 25842 12850
rect 27134 12798 27186 12850
rect 28590 12798 28642 12850
rect 31278 12798 31330 12850
rect 35534 12798 35586 12850
rect 5070 12686 5122 12738
rect 7310 12686 7362 12738
rect 20638 12686 20690 12738
rect 23998 12686 24050 12738
rect 24446 12686 24498 12738
rect 24558 12686 24610 12738
rect 35870 12686 35922 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 13134 12350 13186 12402
rect 15038 12350 15090 12402
rect 19966 12350 20018 12402
rect 23550 12350 23602 12402
rect 25790 12350 25842 12402
rect 28254 12350 28306 12402
rect 29598 12350 29650 12402
rect 39678 12350 39730 12402
rect 6862 12238 6914 12290
rect 10334 12238 10386 12290
rect 14030 12238 14082 12290
rect 14478 12238 14530 12290
rect 28814 12238 28866 12290
rect 30270 12238 30322 12290
rect 30494 12238 30546 12290
rect 32510 12238 32562 12290
rect 33854 12238 33906 12290
rect 38446 12238 38498 12290
rect 2382 12126 2434 12178
rect 5630 12126 5682 12178
rect 6190 12126 6242 12178
rect 9550 12126 9602 12178
rect 23102 12126 23154 12178
rect 26126 12126 26178 12178
rect 26350 12126 26402 12178
rect 28254 12126 28306 12178
rect 29038 12126 29090 12178
rect 29934 12126 29986 12178
rect 32286 12126 32338 12178
rect 33070 12126 33122 12178
rect 39118 12126 39170 12178
rect 3054 12014 3106 12066
rect 5182 12014 5234 12066
rect 8990 12014 9042 12066
rect 12462 12014 12514 12066
rect 13470 12014 13522 12066
rect 15598 12014 15650 12066
rect 20190 12014 20242 12066
rect 22318 12014 22370 12066
rect 26910 12014 26962 12066
rect 35982 12014 36034 12066
rect 36318 12014 36370 12066
rect 14702 11902 14754 11954
rect 28478 11902 28530 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 7310 11566 7362 11618
rect 7646 11566 7698 11618
rect 11230 11566 11282 11618
rect 11566 11566 11618 11618
rect 23886 11566 23938 11618
rect 31950 11566 32002 11618
rect 33182 11566 33234 11618
rect 33518 11566 33570 11618
rect 35198 11566 35250 11618
rect 9214 11454 9266 11506
rect 18510 11454 18562 11506
rect 19966 11454 20018 11506
rect 20750 11454 20802 11506
rect 21422 11454 21474 11506
rect 25678 11454 25730 11506
rect 26126 11454 26178 11506
rect 29262 11454 29314 11506
rect 29710 11454 29762 11506
rect 3726 11342 3778 11394
rect 8094 11342 8146 11394
rect 12014 11342 12066 11394
rect 13694 11342 13746 11394
rect 15262 11342 15314 11394
rect 15598 11342 15650 11394
rect 20078 11342 20130 11394
rect 22206 11342 22258 11394
rect 24222 11342 24274 11394
rect 24894 11342 24946 11394
rect 26238 11342 26290 11394
rect 34302 11342 34354 11394
rect 35534 11342 35586 11394
rect 3390 11230 3442 11282
rect 8206 11230 8258 11282
rect 12126 11230 12178 11282
rect 16382 11230 16434 11282
rect 19182 11230 19234 11282
rect 19518 11230 19570 11282
rect 22542 11230 22594 11282
rect 22878 11230 22930 11282
rect 25006 11230 25058 11282
rect 26798 11230 26850 11282
rect 32062 11230 32114 11282
rect 32286 11230 32338 11282
rect 34190 11230 34242 11282
rect 35758 11230 35810 11282
rect 36318 11230 36370 11282
rect 13470 11118 13522 11170
rect 18846 11118 18898 11170
rect 22990 11118 23042 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 11566 10782 11618 10834
rect 12126 10782 12178 10834
rect 16382 10782 16434 10834
rect 19182 10782 19234 10834
rect 24222 10782 24274 10834
rect 27134 10782 27186 10834
rect 29486 10782 29538 10834
rect 7982 10670 8034 10722
rect 11790 10670 11842 10722
rect 13246 10670 13298 10722
rect 15710 10670 15762 10722
rect 18398 10670 18450 10722
rect 19742 10670 19794 10722
rect 20302 10670 20354 10722
rect 22766 10670 22818 10722
rect 25342 10670 25394 10722
rect 26798 10670 26850 10722
rect 28590 10670 28642 10722
rect 28926 10670 28978 10722
rect 29822 10670 29874 10722
rect 30494 10670 30546 10722
rect 31502 10670 31554 10722
rect 32062 10670 32114 10722
rect 8094 10558 8146 10610
rect 12462 10558 12514 10610
rect 16046 10558 16098 10610
rect 16718 10558 16770 10610
rect 17502 10558 17554 10610
rect 18622 10558 18674 10610
rect 22990 10558 23042 10610
rect 25566 10558 25618 10610
rect 26014 10558 26066 10610
rect 26462 10558 26514 10610
rect 30270 10558 30322 10610
rect 31278 10558 31330 10610
rect 11006 10446 11058 10498
rect 15374 10446 15426 10498
rect 19518 10446 19570 10498
rect 20862 10446 20914 10498
rect 24670 10446 24722 10498
rect 27246 10446 27298 10498
rect 30942 10446 30994 10498
rect 7086 10334 7138 10386
rect 7422 10334 7474 10386
rect 17838 10334 17890 10386
rect 27918 10334 27970 10386
rect 28254 10334 28306 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 11678 9998 11730 10050
rect 13694 9998 13746 10050
rect 29934 9998 29986 10050
rect 11230 9886 11282 9938
rect 12014 9886 12066 9938
rect 16382 9886 16434 9938
rect 18398 9886 18450 9938
rect 20526 9886 20578 9938
rect 22206 9886 22258 9938
rect 24334 9886 24386 9938
rect 27582 9886 27634 9938
rect 29822 9886 29874 9938
rect 31054 9886 31106 9938
rect 33182 9886 33234 9938
rect 6862 9774 6914 9826
rect 8430 9774 8482 9826
rect 12798 9774 12850 9826
rect 14030 9774 14082 9826
rect 17726 9774 17778 9826
rect 21534 9774 21586 9826
rect 24782 9774 24834 9826
rect 28030 9774 28082 9826
rect 29486 9774 29538 9826
rect 30270 9774 30322 9826
rect 9102 9662 9154 9714
rect 12574 9662 12626 9714
rect 14254 9662 14306 9714
rect 14702 9662 14754 9714
rect 25454 9662 25506 9714
rect 6526 9550 6578 9602
rect 28366 9550 28418 9602
rect 29150 9550 29202 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 9550 9214 9602 9266
rect 12238 9214 12290 9266
rect 19294 9214 19346 9266
rect 22206 9214 22258 9266
rect 25342 9214 25394 9266
rect 6414 9102 6466 9154
rect 11342 9102 11394 9154
rect 12798 9102 12850 9154
rect 13358 9102 13410 9154
rect 21534 9102 21586 9154
rect 23214 9102 23266 9154
rect 26910 9102 26962 9154
rect 28478 9102 28530 9154
rect 5742 8990 5794 9042
rect 8990 8990 9042 9042
rect 9886 8990 9938 9042
rect 10446 8990 10498 9042
rect 10782 8990 10834 9042
rect 11566 8990 11618 9042
rect 18622 8990 18674 9042
rect 21646 8990 21698 9042
rect 23326 8990 23378 9042
rect 23774 8990 23826 9042
rect 24110 8990 24162 9042
rect 26798 8990 26850 9042
rect 27806 8990 27858 9042
rect 8542 8878 8594 8930
rect 18062 8878 18114 8930
rect 18398 8878 18450 8930
rect 19742 8878 19794 8930
rect 23998 8878 24050 8930
rect 30606 8878 30658 8930
rect 12574 8766 12626 8818
rect 19070 8766 19122 8818
rect 19406 8766 19458 8818
rect 19742 8766 19794 8818
rect 20526 8766 20578 8818
rect 20862 8766 20914 8818
rect 22542 8766 22594 8818
rect 25790 8766 25842 8818
rect 26126 8766 26178 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 22206 8430 22258 8482
rect 11454 8318 11506 8370
rect 15262 8318 15314 8370
rect 18510 8318 18562 8370
rect 19518 8318 19570 8370
rect 20750 8318 20802 8370
rect 21646 8318 21698 8370
rect 22766 8318 22818 8370
rect 23102 8318 23154 8370
rect 24446 8318 24498 8370
rect 15598 8206 15650 8258
rect 19406 8206 19458 8258
rect 21982 8206 22034 8258
rect 23886 8206 23938 8258
rect 25790 8206 25842 8258
rect 29934 8206 29986 8258
rect 16382 8094 16434 8146
rect 18846 8094 18898 8146
rect 20078 8094 20130 8146
rect 23662 8094 23714 8146
rect 25454 8094 25506 8146
rect 27358 7982 27410 8034
rect 27806 7982 27858 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 14702 7646 14754 7698
rect 16382 7646 16434 7698
rect 22878 7646 22930 7698
rect 23326 7646 23378 7698
rect 26350 7646 26402 7698
rect 29150 7646 29202 7698
rect 10222 7534 10274 7586
rect 12238 7534 12290 7586
rect 14142 7534 14194 7586
rect 15822 7534 15874 7586
rect 18062 7534 18114 7586
rect 18510 7534 18562 7586
rect 25342 7534 25394 7586
rect 28254 7534 28306 7586
rect 28702 7534 28754 7586
rect 10558 7422 10610 7474
rect 11118 7422 11170 7474
rect 11454 7422 11506 7474
rect 12126 7422 12178 7474
rect 13358 7422 13410 7474
rect 14030 7422 14082 7474
rect 15710 7422 15762 7474
rect 16718 7422 16770 7474
rect 17502 7422 17554 7474
rect 17838 7422 17890 7474
rect 19518 7422 19570 7474
rect 25678 7422 25730 7474
rect 27918 7422 27970 7474
rect 20190 7310 20242 7362
rect 22318 7310 22370 7362
rect 26462 7310 26514 7362
rect 29262 7310 29314 7362
rect 13022 7198 13074 7250
rect 15038 7198 15090 7250
rect 27582 7198 27634 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 17166 6862 17218 6914
rect 10110 6750 10162 6802
rect 12238 6750 12290 6802
rect 19854 6750 19906 6802
rect 25342 6750 25394 6802
rect 27470 6750 27522 6802
rect 28590 6750 28642 6802
rect 9326 6638 9378 6690
rect 12686 6638 12738 6690
rect 13694 6638 13746 6690
rect 17950 6638 18002 6690
rect 20638 6638 20690 6690
rect 22542 6638 22594 6690
rect 24670 6638 24722 6690
rect 27806 6638 27858 6690
rect 17726 6526 17778 6578
rect 20414 6526 20466 6578
rect 13470 6414 13522 6466
rect 16270 6414 16322 6466
rect 16830 6414 16882 6466
rect 28142 6414 28194 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 11790 6078 11842 6130
rect 25678 6078 25730 6130
rect 12910 5966 12962 6018
rect 16382 5966 16434 6018
rect 16718 5966 16770 6018
rect 21982 5966 22034 6018
rect 23326 5966 23378 6018
rect 23886 5966 23938 6018
rect 26574 5966 26626 6018
rect 28030 5966 28082 6018
rect 12126 5854 12178 5906
rect 21422 5854 21474 5906
rect 22206 5854 22258 5906
rect 23102 5854 23154 5906
rect 26014 5854 26066 5906
rect 26686 5854 26738 5906
rect 27246 5854 27298 5906
rect 15038 5742 15090 5794
rect 30158 5742 30210 5794
rect 21086 5630 21138 5682
rect 22766 5630 22818 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 15374 5182 15426 5234
rect 16382 5182 16434 5234
rect 18510 5182 18562 5234
rect 24894 5182 24946 5234
rect 25342 5182 25394 5234
rect 26910 5182 26962 5234
rect 15598 5070 15650 5122
rect 20414 5070 20466 5122
rect 21310 5070 21362 5122
rect 22094 5070 22146 5122
rect 22766 5070 22818 5122
rect 21646 4958 21698 5010
rect 20750 4846 20802 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 23774 4510 23826 4562
rect 21198 4398 21250 4450
rect 20526 4286 20578 4338
rect 23326 4174 23378 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 4032 59200 4144 60000
rect 4480 59200 4592 60000
rect 4928 59200 5040 60000
rect 5376 59200 5488 60000
rect 5824 59200 5936 60000
rect 6272 59200 6384 60000
rect 6720 59200 6832 60000
rect 7168 59200 7280 60000
rect 7616 59200 7728 60000
rect 8064 59200 8176 60000
rect 8512 59200 8624 60000
rect 8960 59200 9072 60000
rect 9408 59200 9520 60000
rect 9856 59200 9968 60000
rect 10304 59200 10416 60000
rect 10752 59200 10864 60000
rect 11200 59200 11312 60000
rect 11648 59200 11760 60000
rect 12096 59200 12208 60000
rect 12544 59200 12656 60000
rect 12992 59200 13104 60000
rect 13440 59200 13552 60000
rect 13888 59200 14000 60000
rect 14336 59200 14448 60000
rect 14784 59200 14896 60000
rect 15232 59200 15344 60000
rect 15680 59200 15792 60000
rect 16128 59200 16240 60000
rect 16576 59200 16688 60000
rect 17024 59200 17136 60000
rect 17472 59200 17584 60000
rect 17920 59200 18032 60000
rect 18368 59200 18480 60000
rect 18816 59200 18928 60000
rect 19264 59200 19376 60000
rect 19712 59200 19824 60000
rect 20160 59200 20272 60000
rect 20608 59200 20720 60000
rect 21056 59200 21168 60000
rect 21504 59200 21616 60000
rect 21952 59200 22064 60000
rect 22400 59200 22512 60000
rect 22848 59200 22960 60000
rect 23296 59200 23408 60000
rect 23744 59200 23856 60000
rect 24192 59200 24304 60000
rect 24640 59200 24752 60000
rect 25088 59200 25200 60000
rect 25536 59200 25648 60000
rect 25984 59200 26096 60000
rect 26432 59200 26544 60000
rect 26880 59200 26992 60000
rect 27328 59200 27440 60000
rect 27776 59200 27888 60000
rect 28224 59200 28336 60000
rect 28672 59200 28784 60000
rect 29120 59200 29232 60000
rect 29568 59200 29680 60000
rect 30016 59200 30128 60000
rect 30464 59200 30576 60000
rect 30912 59200 31024 60000
rect 31360 59200 31472 60000
rect 31808 59200 31920 60000
rect 32256 59200 32368 60000
rect 32704 59200 32816 60000
rect 33152 59200 33264 60000
rect 33600 59200 33712 60000
rect 34048 59200 34160 60000
rect 34496 59200 34608 60000
rect 34944 59200 35056 60000
rect 35392 59200 35504 60000
rect 35840 59200 35952 60000
rect 36288 59200 36400 60000
rect 36736 59200 36848 60000
rect 37184 59200 37296 60000
rect 37632 59200 37744 60000
rect 38080 59200 38192 60000
rect 38528 59200 38640 60000
rect 38976 59200 39088 60000
rect 39424 59200 39536 60000
rect 39872 59200 39984 60000
rect 40320 59200 40432 60000
rect 40768 59200 40880 60000
rect 41216 59200 41328 60000
rect 41664 59200 41776 60000
rect 42112 59200 42224 60000
rect 42560 59200 42672 60000
rect 43008 59200 43120 60000
rect 43456 59200 43568 60000
rect 43904 59200 44016 60000
rect 44352 59200 44464 60000
rect 44800 59200 44912 60000
rect 45248 59200 45360 60000
rect 45696 59200 45808 60000
rect 46144 59200 46256 60000
rect 46592 59200 46704 60000
rect 47040 59200 47152 60000
rect 47488 59200 47600 60000
rect 47936 59200 48048 60000
rect 48384 59200 48496 60000
rect 48832 59200 48944 60000
rect 49280 59200 49392 60000
rect 49728 59200 49840 60000
rect 50176 59200 50288 60000
rect 50624 59200 50736 60000
rect 51072 59200 51184 60000
rect 51520 59200 51632 60000
rect 51968 59200 52080 60000
rect 52416 59200 52528 60000
rect 52864 59200 52976 60000
rect 53312 59200 53424 60000
rect 53760 59200 53872 60000
rect 54208 59200 54320 60000
rect 54656 59200 54768 60000
rect 55104 59200 55216 60000
rect 55552 59200 55664 60000
rect 1820 55298 1876 55310
rect 1820 55246 1822 55298
rect 1874 55246 1876 55298
rect 1820 53730 1876 55246
rect 2492 55186 2548 55198
rect 2492 55134 2494 55186
rect 2546 55134 2548 55186
rect 2492 54738 2548 55134
rect 4060 54852 4116 59200
rect 4508 56308 4564 59200
rect 5404 56868 5460 59200
rect 5852 57764 5908 59200
rect 5852 57708 6244 57764
rect 4956 56812 5460 56868
rect 4620 56308 4676 56318
rect 4508 56252 4620 56308
rect 4620 56214 4676 56252
rect 4956 55970 5012 56812
rect 5516 56308 5572 56318
rect 5516 56194 5572 56252
rect 6188 56306 6244 57708
rect 6188 56254 6190 56306
rect 6242 56254 6244 56306
rect 6188 56242 6244 56254
rect 5516 56142 5518 56194
rect 5570 56142 5572 56194
rect 5516 56130 5572 56142
rect 5852 56196 5908 56206
rect 5852 56102 5908 56140
rect 4956 55918 4958 55970
rect 5010 55918 5012 55970
rect 4956 55906 5012 55918
rect 6748 55972 6804 59200
rect 7196 56308 7252 59200
rect 7420 56308 7476 56318
rect 7196 56306 7476 56308
rect 7196 56254 7422 56306
rect 7474 56254 7476 56306
rect 7196 56252 7476 56254
rect 7420 56242 7476 56252
rect 6972 55972 7028 55982
rect 6748 55970 7028 55972
rect 6748 55918 6974 55970
rect 7026 55918 7028 55970
rect 6748 55916 7028 55918
rect 8092 55972 8148 59200
rect 8540 56308 8596 59200
rect 8652 56308 8708 56318
rect 8540 56306 8708 56308
rect 8540 56254 8654 56306
rect 8706 56254 8708 56306
rect 8540 56252 8708 56254
rect 8652 56242 8708 56252
rect 8428 56196 8484 56206
rect 8204 55972 8260 55982
rect 8092 55970 8260 55972
rect 8092 55918 8206 55970
rect 8258 55918 8260 55970
rect 8092 55916 8260 55918
rect 6972 55906 7028 55916
rect 8204 55906 8260 55916
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4060 54786 4116 54796
rect 4620 55410 4676 55422
rect 4620 55358 4622 55410
rect 4674 55358 4676 55410
rect 4620 54740 4676 55358
rect 5964 55410 6020 55422
rect 5964 55358 5966 55410
rect 6018 55358 6020 55410
rect 2492 54686 2494 54738
rect 2546 54686 2548 54738
rect 2492 54674 2548 54686
rect 4172 54684 4676 54740
rect 5068 55074 5124 55086
rect 5068 55022 5070 55074
rect 5122 55022 5124 55074
rect 1820 53678 1822 53730
rect 1874 53678 1876 53730
rect 1820 52162 1876 53678
rect 2380 54628 2436 54638
rect 2380 53172 2436 54572
rect 2604 54516 2660 54526
rect 2940 54516 2996 54526
rect 2604 54514 2996 54516
rect 2604 54462 2606 54514
rect 2658 54462 2942 54514
rect 2994 54462 2996 54514
rect 2604 54460 2996 54462
rect 2604 54450 2660 54460
rect 2940 54450 2996 54460
rect 3724 54516 3780 54526
rect 4172 54516 4228 54684
rect 4396 54516 4452 54526
rect 3724 54514 4228 54516
rect 3724 54462 3726 54514
rect 3778 54462 4228 54514
rect 3724 54460 4228 54462
rect 4284 54514 4452 54516
rect 4284 54462 4398 54514
rect 4450 54462 4452 54514
rect 4284 54460 4452 54462
rect 3612 54402 3668 54414
rect 3612 54350 3614 54402
rect 3666 54350 3668 54402
rect 3612 53732 3668 54350
rect 3500 53676 3612 53732
rect 2492 53620 2548 53630
rect 2492 53618 2884 53620
rect 2492 53566 2494 53618
rect 2546 53566 2884 53618
rect 2492 53564 2884 53566
rect 2492 53554 2548 53564
rect 2380 53116 2772 53172
rect 2716 53058 2772 53116
rect 2828 53170 2884 53564
rect 2828 53118 2830 53170
rect 2882 53118 2884 53170
rect 2828 53106 2884 53118
rect 3388 53060 3444 53070
rect 3500 53060 3556 53676
rect 3612 53666 3668 53676
rect 2716 53006 2718 53058
rect 2770 53006 2772 53058
rect 2716 52994 2772 53006
rect 3052 53058 3556 53060
rect 3052 53006 3390 53058
rect 3442 53006 3556 53058
rect 3052 53004 3556 53006
rect 3612 53170 3668 53182
rect 3612 53118 3614 53170
rect 3666 53118 3668 53170
rect 3052 52946 3108 53004
rect 3388 52966 3444 53004
rect 3052 52894 3054 52946
rect 3106 52894 3108 52946
rect 3052 52882 3108 52894
rect 1820 52110 1822 52162
rect 1874 52110 1876 52162
rect 1820 49810 1876 52110
rect 2492 52052 2548 52062
rect 2492 51958 2548 51996
rect 3612 51716 3668 53118
rect 3724 52946 3780 54460
rect 4284 53956 4340 54460
rect 4396 54450 4452 54460
rect 4956 54402 5012 54414
rect 4956 54350 4958 54402
rect 5010 54350 5012 54402
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4284 53900 4676 53956
rect 4508 53058 4564 53900
rect 4620 53842 4676 53900
rect 4620 53790 4622 53842
rect 4674 53790 4676 53842
rect 4620 53778 4676 53790
rect 4508 53006 4510 53058
rect 4562 53006 4564 53058
rect 4508 52994 4564 53006
rect 4956 53732 5012 54350
rect 5068 53844 5124 55022
rect 5964 54516 6020 55358
rect 8092 55188 8148 55198
rect 7756 55186 8148 55188
rect 7756 55134 8094 55186
rect 8146 55134 8148 55186
rect 7756 55132 8148 55134
rect 6972 54628 7028 54638
rect 6636 54516 6692 54526
rect 5964 54514 6692 54516
rect 5964 54462 6638 54514
rect 6690 54462 6692 54514
rect 5964 54460 6692 54462
rect 5068 53842 5236 53844
rect 5068 53790 5070 53842
rect 5122 53790 5236 53842
rect 5068 53788 5236 53790
rect 5068 53778 5124 53788
rect 3724 52894 3726 52946
rect 3778 52894 3780 52946
rect 3724 52724 3780 52894
rect 3836 52948 3892 52958
rect 3836 52854 3892 52892
rect 4396 52946 4452 52958
rect 4396 52894 4398 52946
rect 4450 52894 4452 52946
rect 4396 52724 4452 52894
rect 4620 52948 4676 52958
rect 4676 52892 4900 52948
rect 4620 52854 4676 52892
rect 3724 52668 4452 52724
rect 3724 51940 3780 52668
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4844 52388 4900 52892
rect 4620 52332 4900 52388
rect 4620 52300 4676 52332
rect 4620 52248 4622 52300
rect 4674 52248 4676 52300
rect 4620 52236 4676 52248
rect 4844 52276 4900 52332
rect 4844 52210 4900 52220
rect 4620 52164 4676 52174
rect 3724 51874 3780 51884
rect 4508 52052 4564 52062
rect 3612 51660 4452 51716
rect 4396 51378 4452 51660
rect 4508 51602 4564 51996
rect 4508 51550 4510 51602
rect 4562 51550 4564 51602
rect 4508 51538 4564 51550
rect 4396 51326 4398 51378
rect 4450 51326 4452 51378
rect 4396 51314 4452 51326
rect 4620 51378 4676 52108
rect 4956 52164 5012 53676
rect 5180 53732 5236 53788
rect 5068 52722 5124 52734
rect 5068 52670 5070 52722
rect 5122 52670 5124 52722
rect 5068 52500 5124 52670
rect 5068 52434 5124 52444
rect 4956 52098 5012 52108
rect 5068 52276 5124 52286
rect 5180 52276 5236 53676
rect 6412 52946 6468 52958
rect 6412 52894 6414 52946
rect 6466 52894 6468 52946
rect 5964 52724 6020 52734
rect 5964 52722 6132 52724
rect 5964 52670 5966 52722
rect 6018 52670 6132 52722
rect 5964 52668 6132 52670
rect 5964 52658 6020 52668
rect 5068 52274 5460 52276
rect 5068 52222 5070 52274
rect 5122 52222 5460 52274
rect 5068 52220 5460 52222
rect 4620 51326 4622 51378
rect 4674 51326 4676 51378
rect 4620 51314 4676 51326
rect 4844 51156 4900 51166
rect 4844 51062 4900 51100
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 2492 50484 2548 50494
rect 2492 49922 2548 50428
rect 2492 49870 2494 49922
rect 2546 49870 2548 49922
rect 2492 49858 2548 49870
rect 1820 49758 1822 49810
rect 1874 49758 1876 49810
rect 1820 48692 1876 49758
rect 4620 49700 4676 49710
rect 4620 49606 4676 49644
rect 5068 49698 5124 52220
rect 5404 51378 5460 52220
rect 5628 52164 5684 52174
rect 5628 52070 5684 52108
rect 5740 52050 5796 52062
rect 5740 51998 5742 52050
rect 5794 51998 5796 52050
rect 5740 51940 5796 51998
rect 5740 51874 5796 51884
rect 5404 51326 5406 51378
rect 5458 51326 5460 51378
rect 5404 51314 5460 51326
rect 5740 51156 5796 51166
rect 5740 50820 5796 51100
rect 5068 49646 5070 49698
rect 5122 49646 5124 49698
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 1820 48626 1876 48636
rect 4732 48804 4788 48814
rect 2828 48580 2884 48590
rect 2828 48466 2884 48524
rect 2828 48414 2830 48466
rect 2882 48414 2884 48466
rect 2828 48402 2884 48414
rect 2940 48132 2996 48142
rect 2940 48038 2996 48076
rect 3836 48132 3892 48142
rect 3052 48018 3108 48030
rect 3052 47966 3054 48018
rect 3106 47966 3108 48018
rect 1708 47570 1764 47582
rect 1708 47518 1710 47570
rect 1762 47518 1764 47570
rect 1596 46676 1652 46686
rect 1596 46116 1652 46620
rect 1708 46228 1764 47518
rect 3052 47236 3108 47966
rect 3836 47570 3892 48076
rect 4732 48130 4788 48748
rect 4732 48078 4734 48130
rect 4786 48078 4788 48130
rect 4732 48066 4788 48078
rect 5068 48692 5124 49646
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 3836 47518 3838 47570
rect 3890 47518 3892 47570
rect 3836 47506 3892 47518
rect 4620 47460 4676 47470
rect 5068 47460 5124 48636
rect 5404 50818 5796 50820
rect 5404 50766 5742 50818
rect 5794 50766 5796 50818
rect 5404 50764 5796 50766
rect 5404 48356 5460 50764
rect 5740 50754 5796 50764
rect 5964 50594 6020 50606
rect 5964 50542 5966 50594
rect 6018 50542 6020 50594
rect 5628 50484 5684 50522
rect 5628 50418 5684 50428
rect 5740 50372 5796 50382
rect 5740 49812 5796 50316
rect 5964 50036 6020 50542
rect 6076 50372 6132 52668
rect 6412 52500 6468 52894
rect 6524 52948 6580 52958
rect 6636 52948 6692 54460
rect 6860 54402 6916 54414
rect 6860 54350 6862 54402
rect 6914 54350 6916 54402
rect 6748 53732 6804 53742
rect 6748 53638 6804 53676
rect 6748 52948 6804 52958
rect 6636 52946 6804 52948
rect 6636 52894 6750 52946
rect 6802 52894 6804 52946
rect 6636 52892 6804 52894
rect 6860 52948 6916 54350
rect 6972 53172 7028 54572
rect 7644 54628 7700 54638
rect 7644 54534 7700 54572
rect 7084 54516 7140 54526
rect 7420 54516 7476 54526
rect 7084 54514 7476 54516
rect 7084 54462 7086 54514
rect 7138 54462 7422 54514
rect 7474 54462 7476 54514
rect 7084 54460 7476 54462
rect 7084 54450 7140 54460
rect 7420 54450 7476 54460
rect 7756 54402 7812 55132
rect 8092 55122 8148 55132
rect 7756 54350 7758 54402
rect 7810 54350 7812 54402
rect 7756 54338 7812 54350
rect 7532 53618 7588 53630
rect 7532 53566 7534 53618
rect 7586 53566 7588 53618
rect 7532 53172 7588 53566
rect 6972 53116 7140 53172
rect 6972 52948 7028 52958
rect 6860 52946 7028 52948
rect 6860 52894 6974 52946
rect 7026 52894 7028 52946
rect 6860 52892 7028 52894
rect 6524 52854 6580 52892
rect 6748 52836 6804 52892
rect 6748 52770 6804 52780
rect 6412 52434 6468 52444
rect 6972 52500 7028 52892
rect 6972 52434 7028 52444
rect 7084 52276 7140 53116
rect 7532 53106 7588 53116
rect 7420 52946 7476 52958
rect 7420 52894 7422 52946
rect 7474 52894 7476 52946
rect 6748 52220 7140 52276
rect 7196 52834 7252 52846
rect 7196 52782 7198 52834
rect 7250 52782 7252 52834
rect 6188 51268 6244 51278
rect 6188 51266 6580 51268
rect 6188 51214 6190 51266
rect 6242 51214 6580 51266
rect 6188 51212 6580 51214
rect 6188 51202 6244 51212
rect 6524 50818 6580 51212
rect 6524 50766 6526 50818
rect 6578 50766 6580 50818
rect 6524 50754 6580 50766
rect 6636 51156 6692 51166
rect 6636 50818 6692 51100
rect 6636 50766 6638 50818
rect 6690 50766 6692 50818
rect 6636 50754 6692 50766
rect 6076 50306 6132 50316
rect 6188 50594 6244 50606
rect 6188 50542 6190 50594
rect 6242 50542 6244 50594
rect 6188 50260 6244 50542
rect 6188 50194 6244 50204
rect 6076 50036 6132 50046
rect 5964 50034 6468 50036
rect 5964 49982 6078 50034
rect 6130 49982 6468 50034
rect 5964 49980 6468 49982
rect 6076 49970 6132 49980
rect 5740 49718 5796 49756
rect 5404 48290 5460 48300
rect 5516 49700 5572 49710
rect 4620 47458 5124 47460
rect 4620 47406 4622 47458
rect 4674 47406 5124 47458
rect 4620 47404 5124 47406
rect 5516 47460 5572 49644
rect 6300 49250 6356 49980
rect 6412 49922 6468 49980
rect 6412 49870 6414 49922
rect 6466 49870 6468 49922
rect 6412 49858 6468 49870
rect 6636 49922 6692 49934
rect 6636 49870 6638 49922
rect 6690 49870 6692 49922
rect 6300 49198 6302 49250
rect 6354 49198 6356 49250
rect 6300 49186 6356 49198
rect 6524 49698 6580 49710
rect 6524 49646 6526 49698
rect 6578 49646 6580 49698
rect 6076 49028 6132 49038
rect 6076 48804 6132 48972
rect 6076 48738 6132 48748
rect 6188 48916 6244 48926
rect 6076 47460 6132 47470
rect 5516 47458 6132 47460
rect 5516 47406 6078 47458
rect 6130 47406 6132 47458
rect 5516 47404 6132 47406
rect 4620 47394 4676 47404
rect 2604 47180 3108 47236
rect 5068 47234 5124 47404
rect 6076 47394 6132 47404
rect 6188 47346 6244 48860
rect 6300 48356 6356 48366
rect 6356 48300 6468 48356
rect 6300 48290 6356 48300
rect 6188 47294 6190 47346
rect 6242 47294 6244 47346
rect 6188 47282 6244 47294
rect 6412 48132 6468 48300
rect 6524 48244 6580 49646
rect 6636 49028 6692 49870
rect 6636 48962 6692 48972
rect 6636 48802 6692 48814
rect 6636 48750 6638 48802
rect 6690 48750 6692 48802
rect 6636 48356 6692 48750
rect 6748 48804 6804 52220
rect 6972 51938 7028 51950
rect 6972 51886 6974 51938
rect 7026 51886 7028 51938
rect 6860 50594 6916 50606
rect 6860 50542 6862 50594
rect 6914 50542 6916 50594
rect 6860 50372 6916 50542
rect 6860 50306 6916 50316
rect 6972 49252 7028 51886
rect 7084 50596 7140 50606
rect 7196 50596 7252 52782
rect 7420 52836 7476 52894
rect 7420 52770 7476 52780
rect 7532 52948 7588 52958
rect 7532 51492 7588 52892
rect 8316 52836 8372 52846
rect 7756 52276 7812 52286
rect 7756 52162 7812 52220
rect 7756 52110 7758 52162
rect 7810 52110 7812 52162
rect 7756 52098 7812 52110
rect 8316 52050 8372 52780
rect 8316 51998 8318 52050
rect 8370 51998 8372 52050
rect 8316 51986 8372 51998
rect 7532 51436 8372 51492
rect 7532 50706 7588 51436
rect 7532 50654 7534 50706
rect 7586 50654 7588 50706
rect 7532 50642 7588 50654
rect 8092 51268 8148 51278
rect 7084 50594 7252 50596
rect 7084 50542 7086 50594
rect 7138 50542 7252 50594
rect 7084 50540 7252 50542
rect 8092 50594 8148 51212
rect 8316 51266 8372 51436
rect 8316 51214 8318 51266
rect 8370 51214 8372 51266
rect 8316 51202 8372 51214
rect 8092 50542 8094 50594
rect 8146 50542 8148 50594
rect 7084 50530 7140 50540
rect 7420 50370 7476 50382
rect 7420 50318 7422 50370
rect 7474 50318 7476 50370
rect 7196 50260 7252 50270
rect 7196 50034 7252 50204
rect 7196 49982 7198 50034
rect 7250 49982 7252 50034
rect 7196 49970 7252 49982
rect 7308 49922 7364 49934
rect 7308 49870 7310 49922
rect 7362 49870 7364 49922
rect 7084 49812 7140 49822
rect 7084 49718 7140 49756
rect 7308 49700 7364 49870
rect 7308 49634 7364 49644
rect 6972 49196 7364 49252
rect 7196 49026 7252 49038
rect 7196 48974 7198 49026
rect 7250 48974 7252 49026
rect 6972 48804 7028 48814
rect 6748 48802 7028 48804
rect 6748 48750 6974 48802
rect 7026 48750 7028 48802
rect 6748 48748 7028 48750
rect 6972 48580 7028 48748
rect 6972 48514 7028 48524
rect 7084 48804 7140 48814
rect 6636 48290 6692 48300
rect 6524 48178 6580 48188
rect 5068 47182 5070 47234
rect 5122 47182 5124 47234
rect 2156 46786 2212 46798
rect 2156 46734 2158 46786
rect 2210 46734 2212 46786
rect 2156 46676 2212 46734
rect 2268 46788 2324 46798
rect 2268 46694 2324 46732
rect 2604 46786 2660 47180
rect 4284 46900 4340 46910
rect 3836 46898 4340 46900
rect 3836 46846 4286 46898
rect 4338 46846 4340 46898
rect 3836 46844 4340 46846
rect 2604 46734 2606 46786
rect 2658 46734 2660 46786
rect 2604 46722 2660 46734
rect 3276 46788 3332 46798
rect 2156 46610 2212 46620
rect 2716 46674 2772 46686
rect 2716 46622 2718 46674
rect 2770 46622 2772 46674
rect 2156 46450 2212 46462
rect 2156 46398 2158 46450
rect 2210 46398 2212 46450
rect 2156 46340 2212 46398
rect 2716 46340 2772 46622
rect 2156 46284 2772 46340
rect 3052 46674 3108 46686
rect 3052 46622 3054 46674
rect 3106 46622 3108 46674
rect 3052 46228 3108 46622
rect 1708 46172 3108 46228
rect 1596 46060 1764 46116
rect 1708 46002 1764 46060
rect 1708 45950 1710 46002
rect 1762 45950 1764 46002
rect 1708 45556 1764 45950
rect 1708 45106 1764 45500
rect 2604 45556 2660 45566
rect 2492 45444 2548 45454
rect 1708 45054 1710 45106
rect 1762 45054 1764 45106
rect 1708 45042 1764 45054
rect 2044 45108 2100 45118
rect 2044 44546 2100 45052
rect 2044 44494 2046 44546
rect 2098 44494 2100 44546
rect 2044 44482 2100 44494
rect 2380 44548 2436 44558
rect 2380 44322 2436 44492
rect 2492 44434 2548 45388
rect 2492 44382 2494 44434
rect 2546 44382 2548 44434
rect 2492 44370 2548 44382
rect 2380 44270 2382 44322
rect 2434 44270 2436 44322
rect 2380 44258 2436 44270
rect 2604 44322 2660 45500
rect 2828 45220 2884 45230
rect 3052 45220 3108 46172
rect 2828 45218 3108 45220
rect 2828 45166 2830 45218
rect 2882 45166 3108 45218
rect 2828 45164 3108 45166
rect 2828 45154 2884 45164
rect 3276 44548 3332 46732
rect 3836 46002 3892 46844
rect 4284 46834 4340 46844
rect 4508 46788 4564 46798
rect 4508 46694 4564 46732
rect 3836 45950 3838 46002
rect 3890 45950 3892 46002
rect 3836 45938 3892 45950
rect 3948 46674 4004 46686
rect 3948 46622 3950 46674
rect 4002 46622 4004 46674
rect 3948 45444 4004 46622
rect 4172 46676 4228 46686
rect 4172 46582 4228 46620
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4620 45892 4676 45902
rect 5068 45892 5124 47182
rect 6300 47234 6356 47246
rect 6300 47182 6302 47234
rect 6354 47182 6356 47234
rect 6300 47012 6356 47182
rect 5740 46956 6356 47012
rect 4620 45890 5124 45892
rect 4620 45838 4622 45890
rect 4674 45838 5124 45890
rect 4620 45836 5124 45838
rect 4620 45826 4676 45836
rect 3948 45378 4004 45388
rect 5068 45666 5124 45836
rect 5068 45614 5070 45666
rect 5122 45614 5124 45666
rect 5068 45332 5124 45614
rect 5068 45266 5124 45276
rect 5404 45892 5460 45902
rect 5404 45330 5460 45836
rect 5740 45890 5796 46956
rect 6300 46788 6356 46798
rect 6412 46788 6468 48076
rect 6860 48130 6916 48142
rect 6860 48078 6862 48130
rect 6914 48078 6916 48130
rect 6860 48020 6916 48078
rect 6972 48020 7028 48030
rect 6860 47964 6972 48020
rect 6972 47954 7028 47964
rect 6636 47908 6692 47918
rect 6300 46786 6468 46788
rect 6300 46734 6302 46786
rect 6354 46734 6468 46786
rect 6300 46732 6468 46734
rect 6524 47852 6636 47908
rect 6300 46722 6356 46732
rect 5740 45838 5742 45890
rect 5794 45838 5796 45890
rect 5740 45826 5796 45838
rect 6524 45890 6580 47852
rect 6636 47842 6692 47852
rect 7084 47458 7140 48748
rect 7084 47406 7086 47458
rect 7138 47406 7140 47458
rect 7084 47394 7140 47406
rect 7196 47124 7252 48974
rect 7308 47908 7364 49196
rect 7420 48916 7476 50318
rect 7868 49140 7924 49150
rect 8092 49140 8148 50542
rect 8428 50428 8484 56140
rect 9436 55972 9492 59200
rect 9884 56308 9940 59200
rect 10108 56308 10164 56318
rect 9884 56306 10164 56308
rect 9884 56254 10110 56306
rect 10162 56254 10164 56306
rect 9884 56252 10164 56254
rect 10108 56242 10164 56252
rect 9660 55972 9716 55982
rect 9436 55970 9716 55972
rect 9436 55918 9662 55970
rect 9714 55918 9716 55970
rect 9436 55916 9716 55918
rect 10780 55972 10836 59200
rect 11228 56308 11284 59200
rect 11452 56308 11508 56318
rect 11228 56306 11508 56308
rect 11228 56254 11454 56306
rect 11506 56254 11508 56306
rect 11228 56252 11508 56254
rect 11452 56242 11508 56252
rect 11004 55972 11060 55982
rect 10780 55970 11060 55972
rect 10780 55918 11006 55970
rect 11058 55918 11060 55970
rect 10780 55916 11060 55918
rect 12124 55972 12180 59200
rect 12572 57090 12628 59200
rect 12572 57038 12574 57090
rect 12626 57038 12628 57090
rect 12572 57026 12628 57038
rect 13132 57090 13188 57102
rect 13132 57038 13134 57090
rect 13186 57038 13188 57090
rect 13132 56306 13188 57038
rect 13132 56254 13134 56306
rect 13186 56254 13188 56306
rect 13132 56242 13188 56254
rect 12348 55972 12404 55982
rect 12124 55970 12404 55972
rect 12124 55918 12350 55970
rect 12402 55918 12404 55970
rect 12124 55916 12404 55918
rect 13468 55972 13524 59200
rect 13916 56308 13972 59200
rect 14028 56308 14084 56318
rect 13916 56306 14084 56308
rect 13916 56254 14030 56306
rect 14082 56254 14084 56306
rect 13916 56252 14084 56254
rect 14028 56242 14084 56252
rect 13580 55972 13636 55982
rect 13468 55970 13636 55972
rect 13468 55918 13582 55970
rect 13634 55918 13636 55970
rect 13468 55916 13636 55918
rect 9660 55906 9716 55916
rect 11004 55906 11060 55916
rect 12348 55906 12404 55916
rect 13580 55906 13636 55916
rect 14588 55972 14644 55982
rect 14812 55972 14868 59200
rect 15036 56308 15092 56318
rect 15260 56308 15316 59200
rect 15708 56644 15764 59200
rect 15036 56306 15316 56308
rect 15036 56254 15038 56306
rect 15090 56254 15316 56306
rect 15036 56252 15316 56254
rect 15484 56588 15764 56644
rect 16044 56754 16100 56766
rect 16044 56702 16046 56754
rect 16098 56702 16100 56754
rect 15036 56242 15092 56252
rect 14588 55970 14868 55972
rect 14588 55918 14590 55970
rect 14642 55918 14868 55970
rect 14588 55916 14868 55918
rect 15484 56082 15540 56588
rect 15708 56196 15764 56206
rect 16044 56196 16100 56702
rect 15708 56102 15764 56140
rect 15932 56194 16100 56196
rect 15932 56142 16046 56194
rect 16098 56142 16100 56194
rect 15932 56140 16100 56142
rect 15484 56030 15486 56082
rect 15538 56030 15540 56082
rect 14588 55906 14644 55916
rect 8876 55298 8932 55310
rect 8876 55246 8878 55298
rect 8930 55246 8932 55298
rect 8876 55076 8932 55246
rect 15484 55188 15540 56030
rect 15932 55972 15988 56140
rect 16044 56130 16100 56140
rect 15596 55916 15988 55972
rect 15596 55410 15652 55916
rect 15932 55524 15988 55534
rect 16156 55524 16212 59200
rect 16380 56196 16436 56206
rect 15932 55522 16212 55524
rect 15932 55470 15934 55522
rect 15986 55470 16212 55522
rect 15932 55468 16212 55470
rect 16268 56194 16436 56196
rect 16268 56142 16382 56194
rect 16434 56142 16436 56194
rect 16268 56140 16436 56142
rect 15932 55458 15988 55468
rect 15596 55358 15598 55410
rect 15650 55358 15652 55410
rect 15596 55346 15652 55358
rect 16268 55188 16324 56140
rect 16380 56130 16436 56140
rect 16604 55860 16660 59200
rect 17052 56754 17108 59200
rect 17052 56702 17054 56754
rect 17106 56702 17108 56754
rect 17052 56690 17108 56702
rect 17164 56642 17220 56654
rect 17164 56590 17166 56642
rect 17218 56590 17220 56642
rect 17164 56306 17220 56590
rect 17164 56254 17166 56306
rect 17218 56254 17220 56306
rect 17164 56242 17220 56254
rect 15484 55132 15988 55188
rect 9324 55076 9380 55086
rect 8876 55074 9380 55076
rect 8876 55022 9326 55074
rect 9378 55022 9380 55074
rect 8876 55020 9380 55022
rect 9100 54852 9156 54862
rect 8764 51268 8820 51278
rect 8764 51174 8820 51212
rect 8876 50484 8932 50522
rect 8428 50372 8596 50428
rect 8876 50418 8932 50428
rect 7420 48850 7476 48860
rect 7644 49138 8092 49140
rect 7644 49086 7870 49138
rect 7922 49086 8092 49138
rect 7644 49084 8092 49086
rect 8148 49084 8260 49140
rect 7644 48242 7700 49084
rect 7868 49074 7924 49084
rect 8092 49074 8148 49084
rect 7644 48190 7646 48242
rect 7698 48190 7700 48242
rect 7644 48178 7700 48190
rect 7756 48356 7812 48366
rect 7308 47842 7364 47852
rect 7644 47348 7700 47358
rect 6524 45838 6526 45890
rect 6578 45838 6580 45890
rect 6524 45826 6580 45838
rect 6636 47068 7252 47124
rect 7532 47346 7700 47348
rect 7532 47294 7646 47346
rect 7698 47294 7700 47346
rect 7532 47292 7700 47294
rect 6636 46674 6692 47068
rect 6636 46622 6638 46674
rect 6690 46622 6692 46674
rect 5628 45780 5684 45790
rect 5404 45278 5406 45330
rect 5458 45278 5460 45330
rect 5404 45266 5460 45278
rect 5516 45778 5684 45780
rect 5516 45726 5630 45778
rect 5682 45726 5684 45778
rect 5516 45724 5684 45726
rect 4284 45218 4340 45230
rect 4284 45166 4286 45218
rect 4338 45166 4340 45218
rect 3724 45108 3780 45118
rect 3724 45014 3780 45052
rect 3276 44454 3332 44492
rect 4172 44548 4228 44558
rect 2604 44270 2606 44322
rect 2658 44270 2660 44322
rect 2604 44258 2660 44270
rect 3052 44322 3108 44334
rect 3052 44270 3054 44322
rect 3106 44270 3108 44322
rect 1932 44210 1988 44222
rect 1932 44158 1934 44210
rect 1986 44158 1988 44210
rect 1932 43876 1988 44158
rect 3052 44212 3108 44270
rect 3052 44146 3108 44156
rect 3612 44322 3668 44334
rect 3836 44324 3892 44334
rect 3612 44270 3614 44322
rect 3666 44270 3668 44322
rect 1932 43708 1988 43820
rect 1708 43652 1988 43708
rect 1708 43426 1764 43652
rect 1708 43374 1710 43426
rect 1762 43374 1764 43426
rect 1708 43362 1764 43374
rect 3612 43428 3668 44270
rect 3724 44268 3836 44324
rect 3724 43876 3780 44268
rect 3836 44230 3892 44268
rect 4172 44322 4228 44492
rect 4172 44270 4174 44322
rect 4226 44270 4228 44322
rect 4172 44258 4228 44270
rect 4060 43988 4116 43998
rect 3724 43810 3780 43820
rect 3836 43932 4060 43988
rect 3836 43650 3892 43932
rect 4060 43922 4116 43932
rect 3836 43598 3838 43650
rect 3890 43598 3892 43650
rect 3836 43586 3892 43598
rect 3612 42980 3668 43372
rect 3388 42978 3668 42980
rect 3388 42926 3614 42978
rect 3666 42926 3668 42978
rect 3388 42924 3668 42926
rect 1820 42532 1876 42542
rect 1820 41970 1876 42476
rect 3388 42420 3444 42924
rect 3612 42914 3668 42924
rect 4172 42868 4228 42878
rect 4284 42868 4340 45166
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4620 44436 4676 44446
rect 4620 44342 4676 44380
rect 4396 44322 4452 44334
rect 4396 44270 4398 44322
rect 4450 44270 4452 44322
rect 4396 43652 4452 44270
rect 4956 44324 5012 44334
rect 4732 44210 4788 44222
rect 4732 44158 4734 44210
rect 4786 44158 4788 44210
rect 4732 43988 4788 44158
rect 4732 43922 4788 43932
rect 4956 43876 5012 44268
rect 4956 43820 5236 43876
rect 4396 43586 4452 43596
rect 5068 43652 5124 43662
rect 5068 43558 5124 43596
rect 5180 43650 5236 43820
rect 5180 43598 5182 43650
rect 5234 43598 5236 43650
rect 5180 43586 5236 43598
rect 4620 43540 4676 43550
rect 4620 43446 4676 43484
rect 4956 43428 5012 43438
rect 4956 43334 5012 43372
rect 4844 43316 4900 43326
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4172 42866 4676 42868
rect 4172 42814 4174 42866
rect 4226 42814 4676 42866
rect 4172 42812 4676 42814
rect 4172 42802 4228 42812
rect 1820 41918 1822 41970
rect 1874 41918 1876 41970
rect 1820 39618 1876 41918
rect 3164 42364 3444 42420
rect 3948 42754 4004 42766
rect 3948 42702 3950 42754
rect 4002 42702 4004 42754
rect 2492 41860 2548 41870
rect 2492 41858 2996 41860
rect 2492 41806 2494 41858
rect 2546 41806 2996 41858
rect 2492 41804 2996 41806
rect 2492 41794 2548 41804
rect 2940 41410 2996 41804
rect 2940 41358 2942 41410
rect 2994 41358 2996 41410
rect 2940 41346 2996 41358
rect 3052 41076 3108 41086
rect 3164 41076 3220 42364
rect 3948 41860 4004 42702
rect 3948 41794 4004 41804
rect 4172 41860 4228 41870
rect 3836 41748 3892 41758
rect 3276 41188 3332 41198
rect 3724 41188 3780 41198
rect 3276 41186 3780 41188
rect 3276 41134 3278 41186
rect 3330 41134 3726 41186
rect 3778 41134 3780 41186
rect 3276 41132 3780 41134
rect 3276 41122 3332 41132
rect 3724 41122 3780 41132
rect 3836 41186 3892 41692
rect 3836 41134 3838 41186
rect 3890 41134 3892 41186
rect 3836 41122 3892 41134
rect 3052 41074 3220 41076
rect 3052 41022 3054 41074
rect 3106 41022 3220 41074
rect 3052 41020 3220 41022
rect 3052 41010 3108 41020
rect 3612 40964 3668 40974
rect 3612 40870 3668 40908
rect 4172 40964 4228 41804
rect 4620 41858 4676 42812
rect 4620 41806 4622 41858
rect 4674 41806 4676 41858
rect 4620 41748 4676 41806
rect 4620 41682 4676 41692
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4844 41524 4900 43260
rect 5516 43316 5572 45724
rect 5628 45714 5684 45724
rect 6636 45556 6692 46622
rect 6972 45892 7028 45930
rect 6972 45826 7028 45836
rect 7196 45780 7252 45790
rect 7196 45686 7252 45724
rect 7532 45778 7588 47292
rect 7644 47282 7700 47292
rect 7532 45726 7534 45778
rect 7586 45726 7588 45778
rect 6860 45668 6916 45678
rect 5852 45500 6692 45556
rect 6748 45612 6860 45668
rect 5516 43250 5572 43260
rect 5628 44324 5684 44334
rect 5628 43650 5684 44268
rect 5740 44212 5796 44222
rect 5740 44118 5796 44156
rect 5852 44210 5908 45500
rect 5964 45332 6020 45342
rect 5964 45108 6020 45276
rect 5964 45106 6132 45108
rect 5964 45054 5966 45106
rect 6018 45054 6132 45106
rect 5964 45052 6132 45054
rect 5964 45042 6020 45052
rect 5852 44158 5854 44210
rect 5906 44158 5908 44210
rect 5628 43598 5630 43650
rect 5682 43598 5684 43650
rect 5628 42644 5684 43598
rect 5852 43540 5908 44158
rect 5964 43540 6020 43550
rect 5852 43538 6020 43540
rect 5852 43486 5966 43538
rect 6018 43486 6020 43538
rect 5852 43484 6020 43486
rect 5964 43428 6020 43484
rect 5964 43362 6020 43372
rect 6076 43540 6132 45052
rect 6636 44996 6692 45006
rect 6188 44994 6692 44996
rect 6188 44942 6638 44994
rect 6690 44942 6692 44994
rect 6188 44940 6692 44942
rect 6188 44546 6244 44940
rect 6636 44930 6692 44940
rect 6748 44772 6804 45612
rect 6860 45602 6916 45612
rect 6188 44494 6190 44546
rect 6242 44494 6244 44546
rect 6188 44482 6244 44494
rect 6524 44716 6804 44772
rect 7532 44996 7588 45726
rect 7756 46114 7812 48300
rect 8092 48132 8148 48142
rect 8092 48038 8148 48076
rect 7980 48020 8036 48030
rect 7980 47926 8036 47964
rect 7756 46062 7758 46114
rect 7810 46062 7812 46114
rect 7644 45668 7700 45678
rect 7644 45574 7700 45612
rect 6524 44546 6580 44716
rect 6524 44494 6526 44546
rect 6578 44494 6580 44546
rect 6524 44482 6580 44494
rect 7532 44436 7588 44940
rect 7644 44436 7700 44446
rect 7532 44434 7700 44436
rect 7532 44382 7646 44434
rect 7698 44382 7700 44434
rect 7532 44380 7700 44382
rect 7644 44370 7700 44380
rect 6300 44324 6356 44334
rect 6300 44230 6356 44268
rect 6748 44324 6804 44334
rect 7084 44324 7140 44334
rect 6748 44322 7140 44324
rect 6748 44270 6750 44322
rect 6802 44270 7086 44322
rect 7138 44270 7140 44322
rect 6748 44268 7140 44270
rect 6076 43204 6132 43484
rect 5740 43148 6132 43204
rect 5740 42866 5796 43148
rect 5740 42814 5742 42866
rect 5794 42814 5796 42866
rect 5740 42802 5796 42814
rect 5628 42588 5908 42644
rect 4956 42532 5012 42542
rect 4956 42084 5012 42476
rect 4956 42018 5012 42028
rect 4956 41860 5012 41870
rect 4956 41766 5012 41804
rect 5516 41858 5572 41870
rect 5516 41806 5518 41858
rect 5570 41806 5572 41858
rect 5292 41746 5348 41758
rect 5292 41694 5294 41746
rect 5346 41694 5348 41746
rect 4844 41468 5012 41524
rect 4844 41300 4900 41310
rect 4284 41188 4340 41198
rect 4284 41094 4340 41132
rect 4732 41188 4788 41198
rect 4172 40898 4228 40908
rect 2492 40628 2548 40638
rect 2492 39730 2548 40572
rect 4508 40628 4564 40638
rect 4508 40534 4564 40572
rect 4508 40180 4564 40190
rect 2492 39678 2494 39730
rect 2546 39678 2548 39730
rect 2492 39666 2548 39678
rect 4284 40178 4564 40180
rect 4284 40126 4510 40178
rect 4562 40126 4564 40178
rect 4284 40124 4564 40126
rect 3948 39620 4004 39630
rect 1820 39566 1822 39618
rect 1874 39566 1876 39618
rect 1820 38724 1876 39566
rect 3836 39564 3948 39620
rect 2828 39060 2884 39070
rect 1820 38050 1876 38668
rect 2492 38836 2548 38846
rect 2492 38162 2548 38780
rect 2828 38834 2884 39004
rect 3052 38948 3108 38958
rect 3052 38854 3108 38892
rect 3724 38948 3780 38958
rect 3724 38854 3780 38892
rect 2828 38782 2830 38834
rect 2882 38782 2884 38834
rect 2828 38770 2884 38782
rect 3388 38834 3444 38846
rect 3388 38782 3390 38834
rect 3442 38782 3444 38834
rect 3388 38668 3444 38782
rect 3500 38836 3556 38846
rect 3500 38742 3556 38780
rect 3836 38668 3892 39564
rect 3948 39554 4004 39564
rect 4284 39396 4340 40124
rect 4508 40114 4564 40124
rect 4620 40180 4676 40218
rect 4732 40180 4788 41132
rect 4844 41074 4900 41244
rect 4956 41298 5012 41468
rect 5292 41412 5348 41694
rect 5292 41346 5348 41356
rect 4956 41246 4958 41298
rect 5010 41246 5012 41298
rect 4956 41234 5012 41246
rect 5516 41300 5572 41806
rect 4844 41022 4846 41074
rect 4898 41022 4900 41074
rect 4844 41010 4900 41022
rect 5068 41076 5124 41086
rect 5068 41074 5460 41076
rect 5068 41022 5070 41074
rect 5122 41022 5460 41074
rect 5068 41020 5460 41022
rect 5068 41010 5124 41020
rect 4844 40404 4900 40414
rect 4844 40310 4900 40348
rect 4732 40124 4900 40180
rect 4620 40114 4676 40124
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4620 39732 4676 39742
rect 4620 39638 4676 39676
rect 4284 39340 4676 39396
rect 3948 39116 4340 39172
rect 3948 38946 4004 39116
rect 4284 39060 4340 39116
rect 4396 39060 4452 39070
rect 4284 39058 4452 39060
rect 4284 39006 4398 39058
rect 4450 39006 4452 39058
rect 4284 39004 4452 39006
rect 4396 38994 4452 39004
rect 3948 38894 3950 38946
rect 4002 38894 4004 38946
rect 3948 38882 4004 38894
rect 4508 38948 4564 38958
rect 4508 38854 4564 38892
rect 4284 38836 4340 38846
rect 4172 38834 4340 38836
rect 4172 38782 4286 38834
rect 4338 38782 4340 38834
rect 4172 38780 4340 38782
rect 4172 38668 4228 38780
rect 4284 38770 4340 38780
rect 4620 38668 4676 39340
rect 4844 39172 4900 40124
rect 5404 40068 5460 41020
rect 5516 40290 5572 41244
rect 5852 40404 5908 42588
rect 6076 42084 6132 42094
rect 5964 41860 6020 41870
rect 5964 41186 6020 41804
rect 6076 41858 6132 42028
rect 6076 41806 6078 41858
rect 6130 41806 6132 41858
rect 6076 41794 6132 41806
rect 5964 41134 5966 41186
rect 6018 41134 6020 41186
rect 5964 41122 6020 41134
rect 6076 41412 6132 41422
rect 5852 40338 5908 40348
rect 5516 40238 5518 40290
rect 5570 40238 5572 40290
rect 5516 40226 5572 40238
rect 6076 40180 6132 41356
rect 6188 41188 6244 41198
rect 6188 41094 6244 41132
rect 6412 41186 6468 41198
rect 6412 41134 6414 41186
rect 6466 41134 6468 41186
rect 6412 40404 6468 41134
rect 6524 41074 6580 41086
rect 6524 41022 6526 41074
rect 6578 41022 6580 41074
rect 6524 40516 6580 41022
rect 6524 40450 6580 40460
rect 6412 40338 6468 40348
rect 5964 40124 6076 40180
rect 5404 40012 5796 40068
rect 5740 39842 5796 40012
rect 5740 39790 5742 39842
rect 5794 39790 5796 39842
rect 5740 39778 5796 39790
rect 4844 38834 4900 39116
rect 4844 38782 4846 38834
rect 4898 38782 4900 38834
rect 4844 38770 4900 38782
rect 4956 39732 5012 39742
rect 4956 38668 5012 39676
rect 5516 39732 5572 39742
rect 5516 39620 5572 39676
rect 5404 39618 5572 39620
rect 5404 39566 5518 39618
rect 5570 39566 5572 39618
rect 5404 39564 5572 39566
rect 3388 38612 4228 38668
rect 2492 38110 2494 38162
rect 2546 38110 2548 38162
rect 2492 38098 2548 38110
rect 1820 37998 1822 38050
rect 1874 37998 1876 38050
rect 1820 37986 1876 37998
rect 4172 37266 4228 38612
rect 4284 38612 4676 38668
rect 4844 38612 5012 38668
rect 5068 39396 5124 39406
rect 5068 38724 5124 39340
rect 4284 37492 4340 38612
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4620 38276 4676 38286
rect 4620 38162 4676 38220
rect 4620 38110 4622 38162
rect 4674 38110 4676 38162
rect 4620 38098 4676 38110
rect 4396 37492 4452 37502
rect 4284 37490 4452 37492
rect 4284 37438 4398 37490
rect 4450 37438 4452 37490
rect 4284 37436 4452 37438
rect 4396 37426 4452 37436
rect 4620 37380 4676 37390
rect 4620 37286 4676 37324
rect 4844 37378 4900 38612
rect 5068 38162 5124 38668
rect 5068 38110 5070 38162
rect 5122 38110 5124 38162
rect 5068 38098 5124 38110
rect 5180 38948 5236 38958
rect 5180 38834 5236 38892
rect 5404 38946 5460 39564
rect 5516 39554 5572 39564
rect 5852 39394 5908 39406
rect 5852 39342 5854 39394
rect 5906 39342 5908 39394
rect 5852 39060 5908 39342
rect 5404 38894 5406 38946
rect 5458 38894 5460 38946
rect 5404 38882 5460 38894
rect 5516 38948 5572 38958
rect 5516 38854 5572 38892
rect 5180 38782 5182 38834
rect 5234 38782 5236 38834
rect 4844 37326 4846 37378
rect 4898 37326 4900 37378
rect 4844 37314 4900 37326
rect 5180 37380 5236 38782
rect 5852 38836 5908 39004
rect 5964 39058 6020 40124
rect 6076 40114 6132 40124
rect 6524 39730 6580 39742
rect 6524 39678 6526 39730
rect 6578 39678 6580 39730
rect 6300 39508 6356 39518
rect 5964 39006 5966 39058
rect 6018 39006 6020 39058
rect 5964 38994 6020 39006
rect 6076 39394 6132 39406
rect 6076 39342 6078 39394
rect 6130 39342 6132 39394
rect 5852 38770 5908 38780
rect 6076 38836 6132 39342
rect 6300 39058 6356 39452
rect 6300 39006 6302 39058
rect 6354 39006 6356 39058
rect 6300 38948 6356 39006
rect 6300 38882 6356 38892
rect 6076 38162 6132 38780
rect 6076 38110 6078 38162
rect 6130 38110 6132 38162
rect 6076 38098 6132 38110
rect 6524 38164 6580 39678
rect 6636 39620 6692 39630
rect 6636 39506 6692 39564
rect 6636 39454 6638 39506
rect 6690 39454 6692 39506
rect 6636 39442 6692 39454
rect 6748 39060 6804 44268
rect 7084 44258 7140 44268
rect 7420 44322 7476 44334
rect 7420 44270 7422 44322
rect 7474 44270 7476 44322
rect 7420 44212 7476 44270
rect 7756 44212 7812 46062
rect 7420 44156 7812 44212
rect 8204 47458 8260 49084
rect 8428 48356 8484 48366
rect 8316 48244 8372 48254
rect 8316 48150 8372 48188
rect 8428 48242 8484 48300
rect 8428 48190 8430 48242
rect 8482 48190 8484 48242
rect 8428 48178 8484 48190
rect 8204 47406 8206 47458
rect 8258 47406 8260 47458
rect 8204 45332 8260 47406
rect 8204 44322 8260 45276
rect 8204 44270 8206 44322
rect 8258 44270 8260 44322
rect 6860 43538 6916 43550
rect 6860 43486 6862 43538
rect 6914 43486 6916 43538
rect 6860 41972 6916 43486
rect 8204 43426 8260 44270
rect 8204 43374 8206 43426
rect 8258 43374 8260 43426
rect 8204 42754 8260 43374
rect 8204 42702 8206 42754
rect 8258 42702 8260 42754
rect 8204 42690 8260 42702
rect 6860 41906 6916 41916
rect 8428 41972 8484 41982
rect 8428 41878 8484 41916
rect 6860 41412 6916 41422
rect 6860 41318 6916 41356
rect 7084 41300 7140 41310
rect 6972 41188 7028 41198
rect 6972 41094 7028 41132
rect 7084 41074 7140 41244
rect 7084 41022 7086 41074
rect 7138 41022 7140 41074
rect 7084 41010 7140 41022
rect 8316 41186 8372 41198
rect 8316 41134 8318 41186
rect 8370 41134 8372 41186
rect 7868 40964 7924 40974
rect 8316 40964 8372 41134
rect 7868 40962 8372 40964
rect 7868 40910 7870 40962
rect 7922 40910 8372 40962
rect 7868 40908 8372 40910
rect 7868 40898 7924 40908
rect 7644 40516 7700 40526
rect 7644 40422 7700 40460
rect 8316 40402 8372 40908
rect 8540 40628 8596 50372
rect 9100 48132 9156 54796
rect 9324 54404 9380 55020
rect 15932 54738 15988 55132
rect 16268 55122 16324 55132
rect 16380 55804 16660 55860
rect 17052 56196 17108 56206
rect 16380 55186 16436 55804
rect 16828 55524 16884 55534
rect 16828 55412 16884 55468
rect 16380 55134 16382 55186
rect 16434 55134 16436 55186
rect 16380 55122 16436 55134
rect 16716 55356 16884 55412
rect 16940 55412 16996 55422
rect 16604 55076 16660 55086
rect 15932 54686 15934 54738
rect 15986 54686 15988 54738
rect 15932 54674 15988 54686
rect 16492 55074 16660 55076
rect 16492 55022 16606 55074
rect 16658 55022 16660 55074
rect 16492 55020 16660 55022
rect 16380 54628 16436 54638
rect 16492 54628 16548 55020
rect 16604 55010 16660 55020
rect 16716 54964 16772 55356
rect 16940 55298 16996 55356
rect 16940 55246 16942 55298
rect 16994 55246 16996 55298
rect 16940 55234 16996 55246
rect 16828 55188 16884 55198
rect 16828 55094 16884 55132
rect 16716 54908 16884 54964
rect 16604 54740 16660 54750
rect 16604 54646 16660 54684
rect 16828 54738 16884 54908
rect 16828 54686 16830 54738
rect 16882 54686 16884 54738
rect 16828 54674 16884 54686
rect 16380 54626 16548 54628
rect 16380 54574 16382 54626
rect 16434 54574 16548 54626
rect 16380 54572 16548 54574
rect 16380 54562 16436 54572
rect 11900 54516 11956 54526
rect 12236 54516 12292 54526
rect 11900 54514 12292 54516
rect 11900 54462 11902 54514
rect 11954 54462 12238 54514
rect 12290 54462 12292 54514
rect 11900 54460 12292 54462
rect 11900 54450 11956 54460
rect 9884 54404 9940 54414
rect 9324 54402 9940 54404
rect 9324 54350 9886 54402
rect 9938 54350 9940 54402
rect 9324 54348 9940 54350
rect 9660 53844 9716 53854
rect 9660 53750 9716 53788
rect 9884 53732 9940 54348
rect 11452 53844 11508 53854
rect 9996 53732 10052 53742
rect 9884 53730 10052 53732
rect 9884 53678 9998 53730
rect 10050 53678 10052 53730
rect 9884 53676 10052 53678
rect 9660 52836 9716 52846
rect 9884 52836 9940 53676
rect 9996 53666 10052 53676
rect 10780 53620 10836 53630
rect 10780 53526 10836 53564
rect 9996 53172 10052 53182
rect 9996 53058 10052 53116
rect 9996 53006 9998 53058
rect 10050 53006 10052 53058
rect 9996 52994 10052 53006
rect 10332 53116 11396 53172
rect 10332 52946 10388 53116
rect 10332 52894 10334 52946
rect 10386 52894 10388 52946
rect 10332 52882 10388 52894
rect 9660 52834 9940 52836
rect 9660 52782 9662 52834
rect 9714 52782 9940 52834
rect 9660 52780 9940 52782
rect 9660 51268 9716 52780
rect 10108 52722 10164 52734
rect 10108 52670 10110 52722
rect 10162 52670 10164 52722
rect 10108 51828 10164 52670
rect 10444 52722 10500 52734
rect 10444 52670 10446 52722
rect 10498 52670 10500 52722
rect 10444 52500 10500 52670
rect 10444 52434 10500 52444
rect 10892 52500 10948 52510
rect 10892 52386 10948 52444
rect 10892 52334 10894 52386
rect 10946 52334 10948 52386
rect 10892 52322 10948 52334
rect 11340 52274 11396 53116
rect 11340 52222 11342 52274
rect 11394 52222 11396 52274
rect 11340 52210 11396 52222
rect 10332 52164 10388 52174
rect 10332 52070 10388 52108
rect 10556 52162 10612 52174
rect 10556 52110 10558 52162
rect 10610 52110 10612 52162
rect 9996 51772 10164 51828
rect 9996 51380 10052 51772
rect 10556 51716 10612 52110
rect 11452 52164 11508 53788
rect 11564 53060 11620 53070
rect 11564 52966 11620 53004
rect 11676 52724 11732 52734
rect 11676 52630 11732 52668
rect 11564 52164 11620 52174
rect 11452 52108 11564 52164
rect 11620 52108 11844 52164
rect 11564 52070 11620 52108
rect 11228 52050 11284 52062
rect 11228 51998 11230 52050
rect 11282 51998 11284 52050
rect 11228 51716 11284 51998
rect 11788 51940 11844 52108
rect 11788 51874 11844 51884
rect 10332 51660 11284 51716
rect 12012 51716 12068 54460
rect 12236 54450 12292 54460
rect 13020 54404 13076 54414
rect 13020 54402 13300 54404
rect 13020 54350 13022 54402
rect 13074 54350 13300 54402
rect 13020 54348 13300 54350
rect 13020 54338 13076 54348
rect 12908 53842 12964 53854
rect 12908 53790 12910 53842
rect 12962 53790 12964 53842
rect 12908 53732 12964 53790
rect 12796 53676 12908 53732
rect 12796 53060 12852 53676
rect 12908 53666 12964 53676
rect 12460 52946 12516 52958
rect 12460 52894 12462 52946
rect 12514 52894 12516 52946
rect 12460 52724 12516 52894
rect 12460 52276 12516 52668
rect 12460 52210 12516 52220
rect 12572 52164 12628 52174
rect 12572 52070 12628 52108
rect 12796 52162 12852 53004
rect 12908 52946 12964 52958
rect 12908 52894 12910 52946
rect 12962 52894 12964 52946
rect 12908 52500 12964 52894
rect 13020 52836 13076 52846
rect 13020 52742 13076 52780
rect 12908 52434 12964 52444
rect 12796 52110 12798 52162
rect 12850 52110 12852 52162
rect 12796 52098 12852 52110
rect 12908 52162 12964 52174
rect 12908 52110 12910 52162
rect 12962 52110 12964 52162
rect 12460 51940 12516 51950
rect 12012 51660 12404 51716
rect 10108 51604 10164 51614
rect 10332 51604 10388 51660
rect 10108 51602 10388 51604
rect 10108 51550 10110 51602
rect 10162 51550 10388 51602
rect 10108 51548 10388 51550
rect 10108 51538 10164 51548
rect 11004 51492 11060 51502
rect 10444 51490 11060 51492
rect 10444 51438 11006 51490
rect 11058 51438 11060 51490
rect 10444 51436 11060 51438
rect 9996 51324 10164 51380
rect 9660 51202 9716 51212
rect 10108 48356 10164 51324
rect 10444 51378 10500 51436
rect 11004 51426 11060 51436
rect 10444 51326 10446 51378
rect 10498 51326 10500 51378
rect 10444 50428 10500 51326
rect 10668 51268 10724 51278
rect 10668 51266 10948 51268
rect 10668 51214 10670 51266
rect 10722 51214 10948 51266
rect 10668 51212 10948 51214
rect 10668 51202 10724 51212
rect 8876 48076 9156 48132
rect 9772 48300 10164 48356
rect 10220 50372 10500 50428
rect 10892 50428 10948 51212
rect 11004 50706 11060 50718
rect 11004 50654 11006 50706
rect 11058 50654 11060 50706
rect 11004 50428 11060 50654
rect 11228 50596 11284 51660
rect 11340 51380 11396 51390
rect 11788 51380 11844 51390
rect 11340 51378 11844 51380
rect 11340 51326 11342 51378
rect 11394 51326 11790 51378
rect 11842 51326 11844 51378
rect 11340 51324 11844 51326
rect 11340 51314 11396 51324
rect 11340 51156 11396 51166
rect 11340 51154 11620 51156
rect 11340 51102 11342 51154
rect 11394 51102 11620 51154
rect 11340 51100 11620 51102
rect 11340 51090 11396 51100
rect 11564 50818 11620 51100
rect 11564 50766 11566 50818
rect 11618 50766 11620 50818
rect 11564 50754 11620 50766
rect 11340 50596 11396 50606
rect 11228 50594 11396 50596
rect 11228 50542 11342 50594
rect 11394 50542 11396 50594
rect 11228 50540 11396 50542
rect 11340 50530 11396 50540
rect 11676 50428 11732 51324
rect 11788 51314 11844 51324
rect 11788 50820 11844 50830
rect 12124 50820 12180 50830
rect 11788 50818 12180 50820
rect 11788 50766 11790 50818
rect 11842 50766 12126 50818
rect 12178 50766 12180 50818
rect 11788 50764 12180 50766
rect 11788 50754 11844 50764
rect 12124 50754 12180 50764
rect 12348 50706 12404 51660
rect 12348 50654 12350 50706
rect 12402 50654 12404 50706
rect 12124 50596 12180 50606
rect 10892 50372 11060 50428
rect 8876 47348 8932 48076
rect 9660 48020 9716 48030
rect 8988 48018 9716 48020
rect 8988 47966 9662 48018
rect 9714 47966 9716 48018
rect 8988 47964 9716 47966
rect 8988 47570 9044 47964
rect 9660 47954 9716 47964
rect 9772 48018 9828 48300
rect 10220 48244 10276 50372
rect 10892 49810 10948 50372
rect 11004 50306 11060 50316
rect 11564 50372 11732 50428
rect 11900 50484 11956 50522
rect 11900 50418 11956 50428
rect 11788 50372 11844 50382
rect 10892 49758 10894 49810
rect 10946 49758 10948 49810
rect 10892 49746 10948 49758
rect 11340 49698 11396 49710
rect 11340 49646 11342 49698
rect 11394 49646 11396 49698
rect 11340 49364 11396 49646
rect 11564 49364 11620 50372
rect 11788 49924 11844 50316
rect 11900 49924 11956 49934
rect 11788 49922 11956 49924
rect 11788 49870 11902 49922
rect 11954 49870 11956 49922
rect 11788 49868 11956 49870
rect 11900 49858 11956 49868
rect 12124 49810 12180 50540
rect 12124 49758 12126 49810
rect 12178 49758 12180 49810
rect 12124 49746 12180 49758
rect 11340 49308 11620 49364
rect 11340 49140 11396 49150
rect 11340 49046 11396 49084
rect 11340 48468 11396 48478
rect 9772 47966 9774 48018
rect 9826 47966 9828 48018
rect 8988 47518 8990 47570
rect 9042 47518 9044 47570
rect 8988 47506 9044 47518
rect 8876 47292 9156 47348
rect 8764 44996 8820 45006
rect 8764 44902 8820 44940
rect 8876 44210 8932 44222
rect 8876 44158 8878 44210
rect 8930 44158 8932 44210
rect 8876 43652 8932 44158
rect 8876 43586 8932 43596
rect 8876 43316 8932 43326
rect 8876 42866 8932 43260
rect 8876 42814 8878 42866
rect 8930 42814 8932 42866
rect 8876 42802 8932 42814
rect 8988 42196 9044 42206
rect 8876 41972 8932 41982
rect 8876 41878 8932 41916
rect 8988 41298 9044 42140
rect 8988 41246 8990 41298
rect 9042 41246 9044 41298
rect 8988 41234 9044 41246
rect 8540 40562 8596 40572
rect 8316 40350 8318 40402
rect 8370 40350 8372 40402
rect 7196 39620 7252 39630
rect 6860 39508 6916 39518
rect 6860 39506 7140 39508
rect 6860 39454 6862 39506
rect 6914 39454 7140 39506
rect 6860 39452 7140 39454
rect 6860 39442 6916 39452
rect 6860 39172 6916 39182
rect 7084 39172 7140 39452
rect 7196 39506 7252 39564
rect 7196 39454 7198 39506
rect 7250 39454 7252 39506
rect 7196 39442 7252 39454
rect 7532 39508 7588 39518
rect 7532 39414 7588 39452
rect 8316 39396 8372 40350
rect 8876 40290 8932 40302
rect 8876 40238 8878 40290
rect 8930 40238 8932 40290
rect 8652 39620 8708 39630
rect 8876 39620 8932 40238
rect 8652 39618 8932 39620
rect 8652 39566 8654 39618
rect 8706 39566 8932 39618
rect 8652 39564 8932 39566
rect 8652 39396 8708 39564
rect 8372 39340 8708 39396
rect 6916 39116 7028 39172
rect 7084 39116 7700 39172
rect 6860 39106 6916 39116
rect 6636 38836 6692 38846
rect 6748 38836 6804 39004
rect 6636 38834 6804 38836
rect 6636 38782 6638 38834
rect 6690 38782 6804 38834
rect 6636 38780 6804 38782
rect 6860 38836 6916 38846
rect 6972 38836 7028 39116
rect 7644 39058 7700 39116
rect 7644 39006 7646 39058
rect 7698 39006 7700 39058
rect 7644 38994 7700 39006
rect 7756 39060 7812 39070
rect 7756 38966 7812 39004
rect 7084 38836 7140 38846
rect 6972 38834 7140 38836
rect 6972 38782 7086 38834
rect 7138 38782 7140 38834
rect 6972 38780 7140 38782
rect 6636 38770 6692 38780
rect 6860 38742 6916 38780
rect 7084 38770 7140 38780
rect 7532 38836 7588 38846
rect 7532 38742 7588 38780
rect 8316 38668 8372 39340
rect 9100 38668 9156 47292
rect 9772 46676 9828 47966
rect 9884 48242 10276 48244
rect 9884 48190 10222 48242
rect 10274 48190 10276 48242
rect 9884 48188 10276 48190
rect 9884 46898 9940 48188
rect 10220 48178 10276 48188
rect 10892 48242 10948 48254
rect 11340 48244 11396 48412
rect 10892 48190 10894 48242
rect 10946 48190 10948 48242
rect 10668 48130 10724 48142
rect 10668 48078 10670 48130
rect 10722 48078 10724 48130
rect 9996 48020 10052 48030
rect 10556 48020 10612 48030
rect 9996 47926 10052 47964
rect 10220 48018 10612 48020
rect 10220 47966 10558 48018
rect 10610 47966 10612 48018
rect 10220 47964 10612 47966
rect 9884 46846 9886 46898
rect 9938 46846 9940 46898
rect 9884 46834 9940 46846
rect 9772 46620 10164 46676
rect 10108 46452 10164 46620
rect 10108 46386 10164 46396
rect 10220 46674 10276 47964
rect 10556 47954 10612 47964
rect 10668 48020 10724 48078
rect 10668 47954 10724 47964
rect 10892 47236 10948 48190
rect 11116 48242 11396 48244
rect 11116 48190 11342 48242
rect 11394 48190 11396 48242
rect 11116 48188 11396 48190
rect 11116 47570 11172 48188
rect 11340 48178 11396 48188
rect 11116 47518 11118 47570
rect 11170 47518 11172 47570
rect 11116 47506 11172 47518
rect 11452 47236 11508 47246
rect 10892 47234 11508 47236
rect 10892 47182 11454 47234
rect 11506 47182 11508 47234
rect 10892 47180 11508 47182
rect 10220 46622 10222 46674
rect 10274 46622 10276 46674
rect 9772 45780 9828 45790
rect 9772 45686 9828 45724
rect 10108 45666 10164 45678
rect 10108 45614 10110 45666
rect 10162 45614 10164 45666
rect 9660 45332 9716 45342
rect 9660 45238 9716 45276
rect 10108 43876 10164 45614
rect 10220 44884 10276 46622
rect 10444 46562 10500 46574
rect 10444 46510 10446 46562
rect 10498 46510 10500 46562
rect 10444 46340 10500 46510
rect 11228 46564 11284 46602
rect 11228 46498 11284 46508
rect 10444 46274 10500 46284
rect 11228 46340 11284 46350
rect 11452 46340 11508 47180
rect 11564 46788 11620 49308
rect 12348 49140 12404 50654
rect 12460 50708 12516 51884
rect 12908 51156 12964 52110
rect 13244 51490 13300 54348
rect 15148 54402 15204 54414
rect 15148 54350 15150 54402
rect 15202 54350 15204 54402
rect 13468 53732 13524 53742
rect 13468 53638 13524 53676
rect 14364 53620 14420 53630
rect 13804 53506 13860 53518
rect 13804 53454 13806 53506
rect 13858 53454 13860 53506
rect 13356 52946 13412 52958
rect 13356 52894 13358 52946
rect 13410 52894 13412 52946
rect 13356 52500 13412 52894
rect 13692 52948 13748 52958
rect 13804 52948 13860 53454
rect 14364 53170 14420 53564
rect 14364 53118 14366 53170
rect 14418 53118 14420 53170
rect 14364 53106 14420 53118
rect 14476 53058 14532 53070
rect 14476 53006 14478 53058
rect 14530 53006 14532 53058
rect 13692 52946 13860 52948
rect 13692 52894 13694 52946
rect 13746 52894 13860 52946
rect 13692 52892 13860 52894
rect 13916 52946 13972 52958
rect 13916 52894 13918 52946
rect 13970 52894 13972 52946
rect 13356 52434 13412 52444
rect 13468 52834 13524 52846
rect 13468 52782 13470 52834
rect 13522 52782 13524 52834
rect 13244 51438 13246 51490
rect 13298 51438 13300 51490
rect 13244 51426 13300 51438
rect 13468 51380 13524 52782
rect 13580 52162 13636 52174
rect 13580 52110 13582 52162
rect 13634 52110 13636 52162
rect 13580 51940 13636 52110
rect 13580 51874 13636 51884
rect 13692 52162 13748 52892
rect 13692 52110 13694 52162
rect 13746 52110 13748 52162
rect 13580 51380 13636 51390
rect 13468 51378 13636 51380
rect 13468 51326 13582 51378
rect 13634 51326 13636 51378
rect 13468 51324 13636 51326
rect 13580 51314 13636 51324
rect 12908 51090 12964 51100
rect 13356 51154 13412 51166
rect 13356 51102 13358 51154
rect 13410 51102 13412 51154
rect 12572 50820 12628 50830
rect 13356 50820 13412 51102
rect 12572 50818 13412 50820
rect 12572 50766 12574 50818
rect 12626 50766 13412 50818
rect 12572 50764 13412 50766
rect 12572 50754 12628 50764
rect 12460 50428 12516 50652
rect 12796 50596 12852 50606
rect 12796 50502 12852 50540
rect 12908 50482 12964 50494
rect 12908 50430 12910 50482
rect 12962 50430 12964 50482
rect 12908 50428 12964 50430
rect 12460 50372 12964 50428
rect 13356 50036 13412 50764
rect 13580 51156 13636 51166
rect 13468 50596 13524 50634
rect 13468 50530 13524 50540
rect 13580 50428 13636 51100
rect 13244 49980 13412 50036
rect 13468 50372 13636 50428
rect 13692 50428 13748 52110
rect 13804 52500 13860 52510
rect 13804 52162 13860 52444
rect 13804 52110 13806 52162
rect 13858 52110 13860 52162
rect 13804 52098 13860 52110
rect 13916 51940 13972 52894
rect 14252 52836 14308 52846
rect 14252 52742 14308 52780
rect 13916 51874 13972 51884
rect 14252 51938 14308 51950
rect 14252 51886 14254 51938
rect 14306 51886 14308 51938
rect 13804 51378 13860 51390
rect 13804 51326 13806 51378
rect 13858 51326 13860 51378
rect 13804 51268 13860 51326
rect 13804 51202 13860 51212
rect 14252 51268 14308 51886
rect 14252 51202 14308 51212
rect 14476 51156 14532 53006
rect 15148 52276 15204 54350
rect 16940 54292 16996 54302
rect 16940 54198 16996 54236
rect 17052 53732 17108 56140
rect 17500 56084 17556 59200
rect 17948 56642 18004 59200
rect 17948 56590 17950 56642
rect 18002 56590 18004 56642
rect 17948 56578 18004 56590
rect 18396 56644 18452 59200
rect 18508 56644 18564 56654
rect 18396 56642 18564 56644
rect 18396 56590 18510 56642
rect 18562 56590 18564 56642
rect 18396 56588 18564 56590
rect 18508 56578 18564 56588
rect 17612 56196 17668 56206
rect 17612 56102 17668 56140
rect 17948 56196 18004 56206
rect 17500 56018 17556 56028
rect 17724 55970 17780 55982
rect 17724 55918 17726 55970
rect 17778 55918 17780 55970
rect 17500 55524 17556 55534
rect 17500 55298 17556 55468
rect 17500 55246 17502 55298
rect 17554 55246 17556 55298
rect 17500 55234 17556 55246
rect 17724 55524 17780 55918
rect 17836 55860 17892 55870
rect 17948 55860 18004 56140
rect 18620 56196 18676 56206
rect 18620 56102 18676 56140
rect 17836 55858 18004 55860
rect 17836 55806 17838 55858
rect 17890 55806 18004 55858
rect 17836 55804 18004 55806
rect 17836 55794 17892 55804
rect 17836 55524 17892 55534
rect 17724 55522 17892 55524
rect 17724 55470 17838 55522
rect 17890 55470 17892 55522
rect 17724 55468 17892 55470
rect 17276 55186 17332 55198
rect 17276 55134 17278 55186
rect 17330 55134 17332 55186
rect 17276 54292 17332 55134
rect 17276 54226 17332 54236
rect 17612 55186 17668 55198
rect 17612 55134 17614 55186
rect 17666 55134 17668 55186
rect 17500 53956 17556 53966
rect 17500 53862 17556 53900
rect 17276 53732 17332 53742
rect 17052 53676 17276 53732
rect 17276 53638 17332 53676
rect 16604 52834 16660 52846
rect 16604 52782 16606 52834
rect 16658 52782 16660 52834
rect 16492 52724 16548 52734
rect 15820 52722 16548 52724
rect 15820 52670 16494 52722
rect 16546 52670 16548 52722
rect 15820 52668 16548 52670
rect 15036 52220 15204 52276
rect 14588 52164 14644 52174
rect 15036 52164 15092 52220
rect 14644 52108 15092 52164
rect 14588 52070 14644 52108
rect 14812 51940 14868 51950
rect 14924 51940 14980 51950
rect 14868 51938 14980 51940
rect 14868 51886 14926 51938
rect 14978 51886 14980 51938
rect 14868 51884 14980 51886
rect 14588 51156 14644 51166
rect 14476 51100 14588 51156
rect 14588 51090 14644 51100
rect 14476 50708 14532 50718
rect 13692 50372 13972 50428
rect 12460 49812 12516 49822
rect 12460 49698 12516 49756
rect 12460 49646 12462 49698
rect 12514 49646 12516 49698
rect 12460 49634 12516 49646
rect 12348 49074 12404 49084
rect 12460 49476 12516 49486
rect 12124 48916 12180 48926
rect 11564 46722 11620 46732
rect 11676 48356 11732 48366
rect 11676 48130 11732 48300
rect 11676 48078 11678 48130
rect 11730 48078 11732 48130
rect 11676 47458 11732 48078
rect 11676 47406 11678 47458
rect 11730 47406 11732 47458
rect 11676 46674 11732 47406
rect 12124 48354 12180 48860
rect 12124 48302 12126 48354
rect 12178 48302 12180 48354
rect 11676 46622 11678 46674
rect 11730 46622 11732 46674
rect 11676 46610 11732 46622
rect 12012 46676 12068 46686
rect 12012 46582 12068 46620
rect 11900 46564 11956 46574
rect 11788 46508 11900 46564
rect 11284 46284 11508 46340
rect 11564 46450 11620 46462
rect 11564 46398 11566 46450
rect 11618 46398 11620 46450
rect 11004 45892 11060 45902
rect 10556 45780 10612 45790
rect 10444 45108 10500 45118
rect 10444 45014 10500 45052
rect 10556 44994 10612 45724
rect 10780 45668 10836 45678
rect 10780 45106 10836 45612
rect 10780 45054 10782 45106
rect 10834 45054 10836 45106
rect 10780 45042 10836 45054
rect 10892 45332 10948 45342
rect 10556 44942 10558 44994
rect 10610 44942 10612 44994
rect 10556 44930 10612 44942
rect 10220 44882 10500 44884
rect 10220 44830 10222 44882
rect 10274 44830 10500 44882
rect 10220 44828 10500 44830
rect 10220 44818 10276 44828
rect 10108 43820 10276 43876
rect 10108 43652 10164 43662
rect 10108 43558 10164 43596
rect 10220 43540 10276 43820
rect 10220 43474 10276 43484
rect 10444 43538 10500 44828
rect 10444 43486 10446 43538
rect 10498 43486 10500 43538
rect 10444 43474 10500 43486
rect 10668 44100 10724 44110
rect 10668 43538 10724 44044
rect 10668 43486 10670 43538
rect 10722 43486 10724 43538
rect 10668 43474 10724 43486
rect 9884 43426 9940 43438
rect 9884 43374 9886 43426
rect 9938 43374 9940 43426
rect 9884 43316 9940 43374
rect 10220 43316 10276 43326
rect 9884 43314 10276 43316
rect 9884 43262 10222 43314
rect 10274 43262 10276 43314
rect 9884 43260 10276 43262
rect 10220 42308 10276 43260
rect 10220 42242 10276 42252
rect 9660 41972 9716 41982
rect 10892 41972 10948 45276
rect 11004 44434 11060 45836
rect 11116 45666 11172 45678
rect 11116 45614 11118 45666
rect 11170 45614 11172 45666
rect 11116 45220 11172 45614
rect 11228 45556 11284 46284
rect 11452 45778 11508 45790
rect 11452 45726 11454 45778
rect 11506 45726 11508 45778
rect 11228 45490 11284 45500
rect 11340 45666 11396 45678
rect 11340 45614 11342 45666
rect 11394 45614 11396 45666
rect 11340 45220 11396 45614
rect 11452 45444 11508 45726
rect 11564 45668 11620 46398
rect 11788 45892 11844 46508
rect 11900 46470 11956 46508
rect 11900 46004 11956 46014
rect 12124 46004 12180 48302
rect 12236 48244 12292 48254
rect 12236 47570 12292 48188
rect 12348 48244 12404 48254
rect 12460 48244 12516 49420
rect 12796 49252 12852 49262
rect 12684 49028 12740 49038
rect 12684 48934 12740 48972
rect 12796 48914 12852 49196
rect 12796 48862 12798 48914
rect 12850 48862 12852 48914
rect 12796 48850 12852 48862
rect 12908 49140 12964 49150
rect 12348 48242 12628 48244
rect 12348 48190 12350 48242
rect 12402 48190 12628 48242
rect 12348 48188 12628 48190
rect 12348 48178 12404 48188
rect 12236 47518 12238 47570
rect 12290 47518 12292 47570
rect 12236 47506 12292 47518
rect 12572 47460 12628 48188
rect 12684 48018 12740 48030
rect 12684 47966 12686 48018
rect 12738 47966 12740 48018
rect 12684 47908 12740 47966
rect 12684 47842 12740 47852
rect 12684 47460 12740 47470
rect 12572 47458 12740 47460
rect 12572 47406 12686 47458
rect 12738 47406 12740 47458
rect 12572 47404 12740 47406
rect 12348 47234 12404 47246
rect 12348 47182 12350 47234
rect 12402 47182 12404 47234
rect 12348 46900 12404 47182
rect 12684 47012 12740 47404
rect 12348 46834 12404 46844
rect 12460 46956 12684 47012
rect 11900 46002 12180 46004
rect 11900 45950 11902 46002
rect 11954 45950 12180 46002
rect 11900 45948 12180 45950
rect 11900 45938 11956 45948
rect 11564 45602 11620 45612
rect 11676 45836 11844 45892
rect 12124 45892 12180 45948
rect 11452 45378 11508 45388
rect 11116 45164 11284 45220
rect 11228 45108 11284 45164
rect 11340 45154 11396 45164
rect 11228 45042 11284 45052
rect 11004 44382 11006 44434
rect 11058 44382 11060 44434
rect 11004 44370 11060 44382
rect 11564 44098 11620 44110
rect 11564 44046 11566 44098
rect 11618 44046 11620 44098
rect 11004 43764 11060 43774
rect 11564 43708 11620 44046
rect 11004 43092 11060 43708
rect 11116 43652 11620 43708
rect 11116 43650 11172 43652
rect 11116 43598 11118 43650
rect 11170 43598 11172 43650
rect 11116 43586 11172 43598
rect 11228 43540 11284 43550
rect 11228 43446 11284 43484
rect 11116 43428 11172 43438
rect 11116 43314 11172 43372
rect 11116 43262 11118 43314
rect 11170 43262 11172 43314
rect 11116 43250 11172 43262
rect 11004 43036 11172 43092
rect 11004 42868 11060 42878
rect 11004 42774 11060 42812
rect 11004 41972 11060 41982
rect 10892 41970 11060 41972
rect 10892 41918 11006 41970
rect 11058 41918 11060 41970
rect 10892 41916 11060 41918
rect 9660 41878 9716 41916
rect 11004 41906 11060 41916
rect 11116 41972 11172 43036
rect 11340 42756 11396 43652
rect 11676 43650 11732 45836
rect 12124 45826 12180 45836
rect 11788 45668 11844 45678
rect 11788 45574 11844 45612
rect 12012 45444 12068 45454
rect 11900 45332 11956 45342
rect 11788 45220 11844 45230
rect 11788 44994 11844 45164
rect 11788 44942 11790 44994
rect 11842 44942 11844 44994
rect 11788 43764 11844 44942
rect 11900 44322 11956 45276
rect 12012 45106 12068 45388
rect 12348 45332 12404 45342
rect 12460 45332 12516 46956
rect 12684 46946 12740 46956
rect 12796 47234 12852 47246
rect 12796 47182 12798 47234
rect 12850 47182 12852 47234
rect 12684 46674 12740 46686
rect 12684 46622 12686 46674
rect 12738 46622 12740 46674
rect 12572 45892 12628 45902
rect 12572 45798 12628 45836
rect 12684 45444 12740 46622
rect 12796 45892 12852 47182
rect 12908 46786 12964 49084
rect 13020 48804 13076 48814
rect 13020 48802 13188 48804
rect 13020 48750 13022 48802
rect 13074 48750 13188 48802
rect 13020 48748 13188 48750
rect 13020 48738 13076 48748
rect 13132 47348 13188 48748
rect 13132 47282 13188 47292
rect 13020 47236 13076 47246
rect 13020 47142 13076 47180
rect 12908 46734 12910 46786
rect 12962 46734 12964 46786
rect 12908 46722 12964 46734
rect 12796 45780 12852 45836
rect 12908 45780 12964 45790
rect 12796 45778 12964 45780
rect 12796 45726 12910 45778
rect 12962 45726 12964 45778
rect 12796 45724 12964 45726
rect 12908 45714 12964 45724
rect 12684 45378 12740 45388
rect 13020 45444 13076 45454
rect 12348 45330 12516 45332
rect 12348 45278 12350 45330
rect 12402 45278 12516 45330
rect 12348 45276 12516 45278
rect 12348 45266 12404 45276
rect 12684 45108 12740 45118
rect 12012 45054 12014 45106
rect 12066 45054 12068 45106
rect 12012 45042 12068 45054
rect 12572 45052 12684 45108
rect 11900 44270 11902 44322
rect 11954 44270 11956 44322
rect 11900 44258 11956 44270
rect 12460 44324 12516 44334
rect 12348 44212 12404 44222
rect 11788 43698 11844 43708
rect 12012 44210 12404 44212
rect 12012 44158 12350 44210
rect 12402 44158 12404 44210
rect 12012 44156 12404 44158
rect 11676 43598 11678 43650
rect 11730 43598 11732 43650
rect 11340 42690 11396 42700
rect 11564 42868 11620 42878
rect 11676 42868 11732 43598
rect 11788 43540 11844 43550
rect 11788 42978 11844 43484
rect 11788 42926 11790 42978
rect 11842 42926 11844 42978
rect 11788 42914 11844 42926
rect 12012 43540 12068 44156
rect 12348 44146 12404 44156
rect 12124 43764 12180 43774
rect 12124 43670 12180 43708
rect 12348 43652 12404 43662
rect 12460 43652 12516 44268
rect 12572 44210 12628 45052
rect 12684 45042 12740 45052
rect 12684 44436 12740 44446
rect 12684 44342 12740 44380
rect 12572 44158 12574 44210
rect 12626 44158 12628 44210
rect 12572 44146 12628 44158
rect 12348 43650 12516 43652
rect 12348 43598 12350 43650
rect 12402 43598 12516 43650
rect 12348 43596 12516 43598
rect 12348 43586 12404 43596
rect 11564 42866 11732 42868
rect 11564 42814 11566 42866
rect 11618 42814 11732 42866
rect 11564 42812 11732 42814
rect 12012 42868 12068 43484
rect 12796 43538 12852 43550
rect 12796 43486 12798 43538
rect 12850 43486 12852 43538
rect 12236 43426 12292 43438
rect 12236 43374 12238 43426
rect 12290 43374 12292 43426
rect 12236 42868 12292 43374
rect 12012 42812 12180 42868
rect 12236 42812 12740 42868
rect 11564 42194 11620 42812
rect 12124 42756 12180 42812
rect 12124 42700 12516 42756
rect 12460 42642 12516 42700
rect 12460 42590 12462 42642
rect 12514 42590 12516 42642
rect 12460 42578 12516 42590
rect 12124 42532 12180 42542
rect 12124 42530 12404 42532
rect 12124 42478 12126 42530
rect 12178 42478 12404 42530
rect 12124 42476 12404 42478
rect 12124 42466 12180 42476
rect 11564 42142 11566 42194
rect 11618 42142 11620 42194
rect 11228 41972 11284 41982
rect 11116 41970 11284 41972
rect 11116 41918 11230 41970
rect 11282 41918 11284 41970
rect 11116 41916 11284 41918
rect 11116 41298 11172 41916
rect 11228 41906 11284 41916
rect 11564 41860 11620 42142
rect 12348 41972 12404 42476
rect 12572 42530 12628 42542
rect 12572 42478 12574 42530
rect 12626 42478 12628 42530
rect 12460 41972 12516 41982
rect 12348 41970 12516 41972
rect 12348 41918 12462 41970
rect 12514 41918 12516 41970
rect 12348 41916 12516 41918
rect 12460 41906 12516 41916
rect 11564 41794 11620 41804
rect 12236 41860 12292 41870
rect 12236 41766 12292 41804
rect 12572 41860 12628 42478
rect 12684 41860 12740 42812
rect 12796 42754 12852 43486
rect 13020 43538 13076 45388
rect 13244 43708 13300 49980
rect 13356 49810 13412 49822
rect 13356 49758 13358 49810
rect 13410 49758 13412 49810
rect 13356 49476 13412 49758
rect 13356 49410 13412 49420
rect 13468 49026 13524 50372
rect 13468 48974 13470 49026
rect 13522 48974 13524 49026
rect 13468 48962 13524 48974
rect 13692 49810 13748 49822
rect 13692 49758 13694 49810
rect 13746 49758 13748 49810
rect 13692 48804 13748 49758
rect 13804 49812 13860 49822
rect 13804 49698 13860 49756
rect 13804 49646 13806 49698
rect 13858 49646 13860 49698
rect 13804 49634 13860 49646
rect 13916 49028 13972 50372
rect 13916 48962 13972 48972
rect 14140 49810 14196 49822
rect 14140 49758 14142 49810
rect 14194 49758 14196 49810
rect 14140 48914 14196 49758
rect 14364 49812 14420 49822
rect 14364 49718 14420 49756
rect 14140 48862 14142 48914
rect 14194 48862 14196 48914
rect 14140 48850 14196 48862
rect 13692 48738 13748 48748
rect 14140 48354 14196 48366
rect 14140 48302 14142 48354
rect 14194 48302 14196 48354
rect 14140 47908 14196 48302
rect 14140 47842 14196 47852
rect 13804 47458 13860 47470
rect 13804 47406 13806 47458
rect 13858 47406 13860 47458
rect 13692 47012 13748 47022
rect 13804 47012 13860 47406
rect 13916 47348 13972 47358
rect 13916 47254 13972 47292
rect 13804 46956 14196 47012
rect 13468 46900 13524 46910
rect 13468 46674 13524 46844
rect 13468 46622 13470 46674
rect 13522 46622 13524 46674
rect 13468 46610 13524 46622
rect 13468 46452 13524 46462
rect 13468 45332 13524 46396
rect 13468 45266 13524 45276
rect 13580 45892 13636 45902
rect 13580 44322 13636 45836
rect 13692 45890 13748 46956
rect 13692 45838 13694 45890
rect 13746 45838 13748 45890
rect 13692 45826 13748 45838
rect 13916 46788 13972 46798
rect 14140 46788 14196 46956
rect 14364 46788 14420 46798
rect 14140 46786 14420 46788
rect 14140 46734 14366 46786
rect 14418 46734 14420 46786
rect 14140 46732 14420 46734
rect 13916 46452 13972 46732
rect 14364 46722 14420 46732
rect 14028 46676 14084 46686
rect 14028 46582 14084 46620
rect 14476 46674 14532 50652
rect 14700 50706 14756 50718
rect 14700 50654 14702 50706
rect 14754 50654 14756 50706
rect 14588 49586 14644 49598
rect 14588 49534 14590 49586
rect 14642 49534 14644 49586
rect 14588 47908 14644 49534
rect 14700 48244 14756 50654
rect 14812 49812 14868 51884
rect 14924 51874 14980 51884
rect 15148 51156 15204 52220
rect 15372 52276 15428 52286
rect 15372 51940 15428 52220
rect 15484 52164 15540 52174
rect 15484 52070 15540 52108
rect 15372 51884 15540 51940
rect 15372 51492 15428 51502
rect 15372 51398 15428 51436
rect 15260 51380 15316 51390
rect 15260 51286 15316 51324
rect 15484 51156 15540 51884
rect 15820 51490 15876 52668
rect 16492 52658 16548 52668
rect 16156 52052 16212 52062
rect 16156 52050 16324 52052
rect 16156 51998 16158 52050
rect 16210 51998 16324 52050
rect 16156 51996 16324 51998
rect 16156 51986 16212 51996
rect 16268 51602 16324 51996
rect 16268 51550 16270 51602
rect 16322 51550 16324 51602
rect 16268 51538 16324 51550
rect 15820 51438 15822 51490
rect 15874 51438 15876 51490
rect 15820 51426 15876 51438
rect 15596 51380 15652 51390
rect 15596 51286 15652 51324
rect 16492 51380 16548 51390
rect 16044 51268 16100 51278
rect 15148 51100 15428 51156
rect 15484 51100 15988 51156
rect 15036 50932 15092 50942
rect 14924 50484 14980 50522
rect 14924 50418 14980 50428
rect 14812 49756 14980 49812
rect 14812 49588 14868 49598
rect 14812 49494 14868 49532
rect 14812 49252 14868 49262
rect 14924 49252 14980 49756
rect 15036 49810 15092 50876
rect 15372 50596 15428 51100
rect 15372 50594 15876 50596
rect 15372 50542 15374 50594
rect 15426 50542 15876 50594
rect 15372 50540 15876 50542
rect 15372 50530 15428 50540
rect 15820 50148 15876 50540
rect 15932 50482 15988 51100
rect 16044 51044 16100 51212
rect 16044 50978 16100 50988
rect 16268 51156 16324 51166
rect 15932 50430 15934 50482
rect 15986 50430 15988 50482
rect 15932 50418 15988 50430
rect 15820 50092 16212 50148
rect 16156 50034 16212 50092
rect 16156 49982 16158 50034
rect 16210 49982 16212 50034
rect 16156 49970 16212 49982
rect 15036 49758 15038 49810
rect 15090 49758 15092 49810
rect 15036 49746 15092 49758
rect 15932 49922 15988 49934
rect 15932 49870 15934 49922
rect 15986 49870 15988 49922
rect 15484 49588 15540 49598
rect 14868 49196 14980 49252
rect 15372 49586 15540 49588
rect 15372 49534 15486 49586
rect 15538 49534 15540 49586
rect 15372 49532 15540 49534
rect 14812 49186 14868 49196
rect 15148 48914 15204 48926
rect 15148 48862 15150 48914
rect 15202 48862 15204 48914
rect 15148 48468 15204 48862
rect 15148 48402 15204 48412
rect 14700 48150 14756 48188
rect 14588 47842 14644 47852
rect 15036 47684 15092 47694
rect 14476 46622 14478 46674
rect 14530 46622 14532 46674
rect 14476 46610 14532 46622
rect 14588 47348 14644 47358
rect 14252 46564 14308 46574
rect 14252 46470 14308 46508
rect 13916 45330 13972 46396
rect 13916 45278 13918 45330
rect 13970 45278 13972 45330
rect 13916 45266 13972 45278
rect 14252 46004 14308 46014
rect 14588 46004 14644 47292
rect 15036 46900 15092 47628
rect 15260 47234 15316 47246
rect 15260 47182 15262 47234
rect 15314 47182 15316 47234
rect 15036 46844 15204 46900
rect 14252 46002 14644 46004
rect 14252 45950 14254 46002
rect 14306 45950 14644 46002
rect 14252 45948 14644 45950
rect 14252 45330 14308 45948
rect 14588 45890 14644 45948
rect 15036 46674 15092 46686
rect 15036 46622 15038 46674
rect 15090 46622 15092 46674
rect 14588 45838 14590 45890
rect 14642 45838 14644 45890
rect 14252 45278 14254 45330
rect 14306 45278 14308 45330
rect 14252 45266 14308 45278
rect 14476 45780 14532 45790
rect 14476 45330 14532 45724
rect 14476 45278 14478 45330
rect 14530 45278 14532 45330
rect 14476 45266 14532 45278
rect 14140 45108 14196 45118
rect 14140 45014 14196 45052
rect 14588 44548 14644 45838
rect 14812 45892 14868 45902
rect 15036 45892 15092 46622
rect 15148 46114 15204 46844
rect 15148 46062 15150 46114
rect 15202 46062 15204 46114
rect 15148 46050 15204 46062
rect 14868 45836 15092 45892
rect 14812 45798 14868 45836
rect 15036 45666 15092 45678
rect 15036 45614 15038 45666
rect 15090 45614 15092 45666
rect 14700 45556 14756 45566
rect 14700 45218 14756 45500
rect 15036 45556 15092 45614
rect 15036 45490 15092 45500
rect 15260 45556 15316 47182
rect 15372 46116 15428 49532
rect 15484 49522 15540 49532
rect 15820 49588 15876 49598
rect 15820 49494 15876 49532
rect 15596 48356 15652 48366
rect 15932 48356 15988 49870
rect 16156 48804 16212 48814
rect 15652 48300 15988 48356
rect 16044 48748 16156 48804
rect 15596 48262 15652 48300
rect 15372 45668 15428 46060
rect 15372 45602 15428 45612
rect 15484 48130 15540 48142
rect 15484 48078 15486 48130
rect 15538 48078 15540 48130
rect 15260 45490 15316 45500
rect 14812 45444 14868 45454
rect 14812 45330 14868 45388
rect 14812 45278 14814 45330
rect 14866 45278 14868 45330
rect 14812 45266 14868 45278
rect 15260 45332 15316 45342
rect 14700 45166 14702 45218
rect 14754 45166 14756 45218
rect 14700 45154 14756 45166
rect 14028 44492 14420 44548
rect 14588 44492 14980 44548
rect 13580 44270 13582 44322
rect 13634 44270 13636 44322
rect 13580 44258 13636 44270
rect 13804 44436 13860 44446
rect 13804 44324 13860 44380
rect 14028 44434 14084 44492
rect 14028 44382 14030 44434
rect 14082 44382 14084 44434
rect 14028 44370 14084 44382
rect 13804 44322 13972 44324
rect 13804 44270 13806 44322
rect 13858 44270 13972 44322
rect 13804 44268 13972 44270
rect 13804 44258 13860 44268
rect 13692 44100 13748 44110
rect 13692 44006 13748 44044
rect 13244 43652 13748 43708
rect 13020 43486 13022 43538
rect 13074 43486 13076 43538
rect 12908 43428 12964 43438
rect 12908 43334 12964 43372
rect 13020 42868 13076 43486
rect 13244 43426 13300 43438
rect 13244 43374 13246 43426
rect 13298 43374 13300 43426
rect 13244 42980 13300 43374
rect 13468 43314 13524 43326
rect 13468 43262 13470 43314
rect 13522 43262 13524 43314
rect 13468 43204 13524 43262
rect 13580 43204 13636 43214
rect 13468 43148 13580 43204
rect 13580 43138 13636 43148
rect 13580 42980 13636 42990
rect 13244 42924 13580 42980
rect 13020 42802 13076 42812
rect 12796 42702 12798 42754
rect 12850 42702 12852 42754
rect 12796 42082 12852 42702
rect 13580 42754 13636 42924
rect 13692 42866 13748 43652
rect 13804 43538 13860 43550
rect 13804 43486 13806 43538
rect 13858 43486 13860 43538
rect 13804 43428 13860 43486
rect 13916 43540 13972 44268
rect 14252 44322 14308 44334
rect 14252 44270 14254 44322
rect 14306 44270 14308 44322
rect 14252 44212 14308 44270
rect 14028 44156 14308 44212
rect 14028 43764 14084 44156
rect 14364 44100 14420 44492
rect 14476 44324 14532 44334
rect 14924 44324 14980 44492
rect 15036 44324 15092 44334
rect 14924 44322 15092 44324
rect 14924 44270 15038 44322
rect 15090 44270 15092 44322
rect 14924 44268 15092 44270
rect 14476 44230 14532 44268
rect 15036 44258 15092 44268
rect 15260 44322 15316 45276
rect 15372 44994 15428 45006
rect 15372 44942 15374 44994
rect 15426 44942 15428 44994
rect 15372 44882 15428 44942
rect 15372 44830 15374 44882
rect 15426 44830 15428 44882
rect 15372 44818 15428 44830
rect 15484 44324 15540 48078
rect 15708 47796 15764 47806
rect 15708 46786 15764 47740
rect 15932 47460 15988 47470
rect 16044 47460 16100 48748
rect 16156 48738 16212 48748
rect 15932 47458 16100 47460
rect 15932 47406 15934 47458
rect 15986 47406 16100 47458
rect 15932 47404 16100 47406
rect 15932 47394 15988 47404
rect 16268 47012 16324 51100
rect 16492 51156 16548 51324
rect 16492 51090 16548 51100
rect 16604 50932 16660 52782
rect 17612 52724 17668 55134
rect 17724 54740 17780 55468
rect 17836 55458 17892 55468
rect 17724 54674 17780 54684
rect 17948 54516 18004 55804
rect 18284 55860 18340 55870
rect 18284 55766 18340 55804
rect 18844 55860 18900 59200
rect 18956 56642 19012 56654
rect 18956 56590 18958 56642
rect 19010 56590 19012 56642
rect 18956 56196 19012 56590
rect 19292 56308 19348 59200
rect 19740 57092 19796 59200
rect 20188 57428 20244 59200
rect 20188 57372 20468 57428
rect 19740 57036 20244 57092
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19404 56308 19460 56318
rect 19292 56306 19460 56308
rect 19292 56254 19406 56306
rect 19458 56254 19460 56306
rect 19292 56252 19460 56254
rect 19404 56242 19460 56252
rect 18956 56194 19236 56196
rect 18956 56142 18958 56194
rect 19010 56142 19236 56194
rect 18956 56140 19236 56142
rect 18956 56130 19012 56140
rect 18844 55794 18900 55804
rect 18396 55524 18452 55534
rect 18508 55524 18564 55534
rect 18452 55522 18564 55524
rect 18452 55470 18510 55522
rect 18562 55470 18564 55522
rect 18452 55468 18564 55470
rect 17948 54450 18004 54460
rect 18060 55298 18116 55310
rect 18060 55246 18062 55298
rect 18114 55246 18116 55298
rect 18060 54180 18116 55246
rect 17836 54124 18116 54180
rect 18284 54516 18340 54526
rect 17836 53954 17892 54124
rect 17836 53902 17838 53954
rect 17890 53902 17892 53954
rect 17836 53890 17892 53902
rect 18172 53956 18228 53966
rect 18284 53956 18340 54460
rect 18396 54402 18452 55468
rect 18508 55458 18564 55468
rect 18844 55412 18900 55422
rect 18844 55318 18900 55356
rect 19180 55300 19236 56140
rect 19852 56194 19908 56206
rect 19852 56142 19854 56194
rect 19906 56142 19908 56194
rect 19404 56084 19460 56094
rect 19404 55522 19460 56028
rect 19404 55470 19406 55522
rect 19458 55470 19460 55522
rect 19404 55458 19460 55470
rect 19852 55412 19908 56142
rect 20188 56196 20244 57036
rect 20188 56102 20244 56140
rect 20412 55522 20468 57372
rect 20636 56308 20692 59200
rect 21532 57204 21588 59200
rect 21532 57148 21812 57204
rect 20748 56308 20804 56318
rect 20636 56306 20804 56308
rect 20636 56254 20750 56306
rect 20802 56254 20804 56306
rect 20636 56252 20804 56254
rect 20748 56242 20804 56252
rect 21308 56196 21364 56206
rect 21308 56102 21364 56140
rect 20412 55470 20414 55522
rect 20466 55470 20468 55522
rect 20412 55458 20468 55470
rect 19852 55346 19908 55356
rect 19180 55234 19236 55244
rect 19068 55188 19124 55198
rect 18956 55132 19068 55188
rect 18508 54516 18564 54526
rect 18508 54514 18788 54516
rect 18508 54462 18510 54514
rect 18562 54462 18788 54514
rect 18508 54460 18788 54462
rect 18508 54450 18564 54460
rect 18396 54350 18398 54402
rect 18450 54350 18452 54402
rect 18396 54338 18452 54350
rect 18228 53900 18340 53956
rect 18172 53890 18228 53900
rect 18396 53844 18452 53854
rect 18396 53750 18452 53788
rect 18620 53732 18676 53742
rect 18732 53732 18788 54460
rect 18676 53676 18788 53732
rect 18844 54290 18900 54302
rect 18844 54238 18846 54290
rect 18898 54238 18900 54290
rect 18620 53638 18676 53676
rect 17052 52668 17668 52724
rect 16828 51380 16884 51390
rect 16828 51286 16884 51324
rect 16604 50866 16660 50876
rect 16828 50372 16884 50382
rect 16380 49810 16436 49822
rect 16380 49758 16382 49810
rect 16434 49758 16436 49810
rect 16380 49028 16436 49758
rect 16716 49138 16772 49150
rect 16716 49086 16718 49138
rect 16770 49086 16772 49138
rect 16380 48962 16436 48972
rect 16604 49028 16660 49038
rect 16604 48934 16660 48972
rect 16716 47460 16772 49086
rect 16828 48804 16884 50316
rect 16828 48242 16884 48748
rect 16828 48190 16830 48242
rect 16882 48190 16884 48242
rect 16828 48178 16884 48190
rect 16716 47394 16772 47404
rect 16380 47348 16436 47358
rect 16380 47254 16436 47292
rect 16604 47348 16660 47358
rect 15708 46734 15710 46786
rect 15762 46734 15764 46786
rect 15708 46452 15764 46734
rect 15932 46956 16324 47012
rect 15708 46386 15764 46396
rect 15820 46676 15876 46686
rect 15820 46228 15876 46620
rect 15596 46172 15876 46228
rect 15596 45444 15652 46172
rect 15708 45780 15764 45790
rect 15708 45686 15764 45724
rect 15820 45668 15876 45678
rect 15820 45574 15876 45612
rect 15932 45444 15988 46956
rect 16380 46900 16436 46910
rect 16156 46898 16436 46900
rect 16156 46846 16382 46898
rect 16434 46846 16436 46898
rect 16156 46844 16436 46846
rect 16156 46676 16212 46844
rect 16380 46834 16436 46844
rect 16156 46610 16212 46620
rect 16268 46676 16324 46686
rect 16604 46676 16660 47292
rect 16268 46674 16660 46676
rect 16268 46622 16270 46674
rect 16322 46622 16660 46674
rect 16268 46620 16660 46622
rect 16268 46610 16324 46620
rect 16380 46452 16436 46462
rect 16380 46358 16436 46396
rect 16044 45668 16100 45678
rect 16044 45574 16100 45612
rect 15932 45388 16100 45444
rect 15596 45378 15652 45388
rect 15932 44994 15988 45006
rect 15932 44942 15934 44994
rect 15986 44942 15988 44994
rect 15932 44882 15988 44942
rect 15932 44830 15934 44882
rect 15986 44830 15988 44882
rect 15932 44548 15988 44830
rect 15260 44270 15262 44322
rect 15314 44270 15316 44322
rect 15260 44258 15316 44270
rect 15372 44268 15540 44324
rect 15820 44324 15876 44334
rect 14028 43698 14084 43708
rect 14140 44044 14420 44100
rect 14700 44098 14756 44110
rect 14700 44046 14702 44098
rect 14754 44046 14756 44098
rect 14028 43540 14084 43550
rect 13916 43538 14084 43540
rect 13916 43486 14030 43538
rect 14082 43486 14084 43538
rect 13916 43484 14084 43486
rect 14028 43474 14084 43484
rect 13804 43362 13860 43372
rect 14028 43204 14084 43214
rect 14140 43204 14196 44044
rect 14700 43988 14756 44046
rect 14924 44100 14980 44110
rect 14924 44006 14980 44044
rect 15372 43988 15428 44268
rect 15596 44212 15652 44222
rect 15596 44210 15764 44212
rect 15596 44158 15598 44210
rect 15650 44158 15764 44210
rect 15596 44156 15764 44158
rect 15596 44146 15652 44156
rect 14252 43932 14756 43988
rect 15260 43932 15428 43988
rect 15484 44100 15540 44110
rect 14252 43538 14308 43932
rect 15260 43876 15316 43932
rect 14252 43486 14254 43538
rect 14306 43486 14308 43538
rect 14252 43474 14308 43486
rect 14476 43820 15316 43876
rect 14364 43316 14420 43326
rect 14364 43222 14420 43260
rect 14084 43148 14196 43204
rect 14028 43138 14084 43148
rect 14364 42980 14420 42990
rect 13692 42814 13694 42866
rect 13746 42814 13748 42866
rect 13692 42802 13748 42814
rect 14252 42978 14420 42980
rect 14252 42926 14366 42978
rect 14418 42926 14420 42978
rect 14252 42924 14420 42926
rect 13580 42702 13582 42754
rect 13634 42702 13636 42754
rect 13580 42690 13636 42702
rect 14252 42754 14308 42924
rect 14364 42914 14420 42924
rect 14476 42756 14532 43820
rect 15484 43764 15540 44044
rect 15260 43708 15540 43764
rect 15708 43762 15764 44156
rect 15708 43710 15710 43762
rect 15762 43710 15764 43762
rect 14812 43650 14868 43662
rect 14812 43598 14814 43650
rect 14866 43598 14868 43650
rect 14812 43092 14868 43598
rect 15036 43652 15316 43708
rect 15708 43698 15764 43710
rect 14924 43092 14980 43102
rect 14812 43036 14924 43092
rect 14924 43026 14980 43036
rect 15036 42978 15092 43652
rect 15148 43538 15204 43550
rect 15148 43486 15150 43538
rect 15202 43486 15204 43538
rect 15148 43428 15204 43486
rect 15148 43362 15204 43372
rect 15036 42926 15038 42978
rect 15090 42926 15092 42978
rect 15036 42866 15092 42926
rect 15036 42814 15038 42866
rect 15090 42814 15092 42866
rect 15036 42802 15092 42814
rect 15372 43092 15428 43102
rect 14252 42702 14254 42754
rect 14306 42702 14308 42754
rect 14252 42690 14308 42702
rect 14364 42700 14980 42756
rect 13804 42532 13860 42542
rect 13804 42438 13860 42476
rect 13468 42308 13524 42318
rect 14364 42308 14420 42700
rect 14476 42532 14532 42542
rect 14700 42532 14756 42542
rect 14532 42476 14644 42532
rect 14476 42466 14532 42476
rect 12908 42196 12964 42206
rect 13468 42196 13524 42252
rect 12908 42102 12964 42140
rect 13356 42140 13524 42196
rect 14140 42252 14420 42308
rect 12796 42030 12798 42082
rect 12850 42030 12852 42082
rect 12796 42018 12852 42030
rect 13244 41972 13300 41982
rect 12908 41970 13300 41972
rect 12908 41918 13246 41970
rect 13298 41918 13300 41970
rect 12908 41916 13300 41918
rect 12908 41860 12964 41916
rect 13244 41906 13300 41916
rect 12684 41804 12964 41860
rect 12572 41794 12628 41804
rect 13020 41748 13076 41758
rect 13020 41654 13076 41692
rect 13356 41412 13412 42140
rect 13468 41970 13524 41982
rect 13468 41918 13470 41970
rect 13522 41918 13524 41970
rect 13468 41860 13524 41918
rect 14140 41970 14196 42252
rect 14140 41918 14142 41970
rect 14194 41918 14196 41970
rect 14140 41906 14196 41918
rect 14476 42196 14532 42206
rect 13804 41860 13860 41870
rect 13468 41804 13804 41860
rect 13804 41794 13860 41804
rect 14252 41746 14308 41758
rect 14252 41694 14254 41746
rect 14306 41694 14308 41746
rect 13356 41356 13524 41412
rect 11116 41246 11118 41298
rect 11170 41246 11172 41298
rect 11116 41234 11172 41246
rect 13244 40964 13300 40974
rect 11340 40628 11396 40638
rect 11676 40628 11732 40638
rect 11396 40626 11732 40628
rect 11396 40574 11678 40626
rect 11730 40574 11732 40626
rect 11396 40572 11732 40574
rect 11340 40534 11396 40572
rect 9436 40404 9492 40414
rect 9436 39730 9492 40348
rect 9436 39678 9438 39730
rect 9490 39678 9492 39730
rect 9436 39666 9492 39678
rect 11564 39732 11620 39742
rect 11564 39638 11620 39676
rect 11676 39060 11732 40572
rect 12012 40516 12068 40526
rect 12012 40422 12068 40460
rect 12684 40514 12740 40526
rect 12684 40462 12686 40514
rect 12738 40462 12740 40514
rect 12348 40402 12404 40414
rect 12348 40350 12350 40402
rect 12402 40350 12404 40402
rect 12348 39732 12404 40350
rect 12684 40180 12740 40462
rect 13244 40514 13300 40908
rect 13244 40462 13246 40514
rect 13298 40462 13300 40514
rect 13244 40450 13300 40462
rect 13468 40740 13524 41356
rect 14252 41300 14308 41694
rect 14252 41234 14308 41244
rect 14140 41188 14196 41198
rect 14476 41188 14532 42140
rect 14588 42194 14644 42476
rect 14700 42530 14868 42532
rect 14700 42478 14702 42530
rect 14754 42478 14868 42530
rect 14700 42476 14868 42478
rect 14700 42466 14756 42476
rect 14588 42142 14590 42194
rect 14642 42142 14644 42194
rect 14588 42130 14644 42142
rect 14700 41860 14756 41870
rect 14140 41094 14196 41132
rect 14364 41186 14532 41188
rect 14364 41134 14478 41186
rect 14530 41134 14532 41186
rect 14364 41132 14532 41134
rect 14028 41076 14084 41086
rect 14028 40964 14084 41020
rect 13468 40514 13524 40684
rect 13468 40462 13470 40514
rect 13522 40462 13524 40514
rect 13468 40450 13524 40462
rect 13804 40962 14084 40964
rect 13804 40910 14030 40962
rect 14082 40910 14084 40962
rect 13804 40908 14084 40910
rect 13580 40404 13636 40414
rect 13580 40310 13636 40348
rect 13804 40402 13860 40908
rect 14028 40898 14084 40908
rect 13804 40350 13806 40402
rect 13858 40350 13860 40402
rect 13804 40338 13860 40350
rect 13916 40740 13972 40750
rect 14364 40740 14420 41132
rect 14476 41122 14532 41132
rect 14588 41188 14644 41198
rect 14588 40964 14644 41132
rect 13916 40404 13972 40684
rect 13916 40338 13972 40348
rect 14028 40684 14420 40740
rect 14476 40962 14644 40964
rect 14476 40910 14590 40962
rect 14642 40910 14644 40962
rect 14476 40908 14644 40910
rect 14028 40402 14084 40684
rect 14028 40350 14030 40402
rect 14082 40350 14084 40402
rect 14028 40338 14084 40350
rect 14476 40180 14532 40908
rect 14588 40898 14644 40908
rect 14588 40404 14644 40414
rect 14588 40310 14644 40348
rect 14588 40180 14644 40190
rect 14476 40124 14588 40180
rect 12684 40114 12740 40124
rect 14588 40114 14644 40124
rect 11676 39058 12292 39060
rect 11676 39006 11678 39058
rect 11730 39006 12292 39058
rect 11676 39004 12292 39006
rect 11676 38994 11732 39004
rect 10780 38724 10836 38734
rect 8316 38612 8932 38668
rect 9100 38612 9828 38668
rect 6524 38098 6580 38108
rect 8204 38164 8260 38174
rect 8204 38070 8260 38108
rect 5180 37314 5236 37324
rect 8876 38050 8932 38612
rect 8876 37998 8878 38050
rect 8930 37998 8932 38050
rect 8876 37828 8932 37998
rect 9436 37828 9492 37838
rect 8876 37826 9492 37828
rect 8876 37774 9438 37826
rect 9490 37774 9492 37826
rect 8876 37772 9492 37774
rect 4172 37214 4174 37266
rect 4226 37214 4228 37266
rect 4172 37202 4228 37214
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5292 29428 5348 29438
rect 5292 29334 5348 29372
rect 8540 29428 8596 29438
rect 8876 29428 8932 37772
rect 9436 37762 9492 37772
rect 9660 37266 9716 37278
rect 9660 37214 9662 37266
rect 9714 37214 9716 37266
rect 9660 37156 9716 37214
rect 9660 37090 9716 37100
rect 9548 30996 9604 31006
rect 8596 29372 8932 29428
rect 9212 30994 9604 30996
rect 9212 30942 9550 30994
rect 9602 30942 9604 30994
rect 9212 30940 9604 30942
rect 5964 29316 6020 29326
rect 8092 29316 8148 29326
rect 5964 29314 6356 29316
rect 5964 29262 5966 29314
rect 6018 29262 6356 29314
rect 5964 29260 6356 29262
rect 5964 29250 6020 29260
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 6300 28530 6356 29260
rect 8092 29314 8260 29316
rect 8092 29262 8094 29314
rect 8146 29262 8260 29314
rect 8092 29260 8260 29262
rect 8092 29250 8148 29260
rect 6524 28644 6580 28654
rect 6524 28550 6580 28588
rect 7196 28644 7252 28654
rect 7196 28550 7252 28588
rect 7532 28642 7588 28654
rect 7532 28590 7534 28642
rect 7586 28590 7588 28642
rect 6300 28478 6302 28530
rect 6354 28478 6356 28530
rect 6300 28466 6356 28478
rect 7532 27972 7588 28590
rect 7532 27906 7588 27916
rect 7756 28530 7812 28542
rect 7756 28478 7758 28530
rect 7810 28478 7812 28530
rect 3500 27858 3556 27870
rect 3500 27806 3502 27858
rect 3554 27806 3556 27858
rect 2268 26516 2324 26526
rect 2268 23940 2324 26460
rect 3500 26516 3556 27806
rect 6636 27860 6692 27870
rect 4172 27748 4228 27758
rect 6300 27748 6356 27758
rect 4172 27746 4340 27748
rect 4172 27694 4174 27746
rect 4226 27694 4340 27746
rect 4172 27692 4340 27694
rect 4172 27682 4228 27692
rect 4284 27300 4340 27692
rect 6300 27654 6356 27692
rect 4956 27636 5012 27646
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 27244 4676 27300
rect 4620 26962 4676 27244
rect 4956 27074 5012 27580
rect 4956 27022 4958 27074
rect 5010 27022 5012 27074
rect 4956 27010 5012 27022
rect 4620 26910 4622 26962
rect 4674 26910 4676 26962
rect 4620 26898 4676 26910
rect 4844 26964 4900 26974
rect 3500 26180 3556 26460
rect 4844 26402 4900 26908
rect 5628 26964 5684 27002
rect 5628 26898 5684 26908
rect 5964 26962 6020 26974
rect 5964 26910 5966 26962
rect 6018 26910 6020 26962
rect 4844 26350 4846 26402
rect 4898 26350 4900 26402
rect 4844 26338 4900 26350
rect 3500 26114 3556 26124
rect 4172 26290 4228 26302
rect 4172 26238 4174 26290
rect 4226 26238 4228 26290
rect 4172 26180 4228 26238
rect 4172 26114 4228 26124
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 5964 24948 6020 26910
rect 6524 26850 6580 26862
rect 6524 26798 6526 26850
rect 6578 26798 6580 26850
rect 6524 26180 6580 26798
rect 6300 26124 6524 26180
rect 6300 25508 6356 26124
rect 6524 26114 6580 26124
rect 6188 25506 6356 25508
rect 6188 25454 6302 25506
rect 6354 25454 6356 25506
rect 6188 25452 6356 25454
rect 6076 24948 6132 24958
rect 5964 24946 6132 24948
rect 5964 24894 6078 24946
rect 6130 24894 6132 24946
rect 5964 24892 6132 24894
rect 6076 24882 6132 24892
rect 1932 23938 2324 23940
rect 1932 23886 2270 23938
rect 2322 23886 2324 23938
rect 1932 23884 2324 23886
rect 1932 23154 1988 23884
rect 2268 23874 2324 23884
rect 2716 24834 2772 24846
rect 3388 24836 3444 24846
rect 2716 24782 2718 24834
rect 2770 24782 2772 24834
rect 2604 23268 2660 23278
rect 2716 23268 2772 24782
rect 3164 24834 3444 24836
rect 3164 24782 3390 24834
rect 3442 24782 3444 24834
rect 3164 24780 3444 24782
rect 2940 24724 2996 24734
rect 2604 23266 2772 23268
rect 2604 23214 2606 23266
rect 2658 23214 2772 23266
rect 2604 23212 2772 23214
rect 2828 24722 2996 24724
rect 2828 24670 2942 24722
rect 2994 24670 2996 24722
rect 2828 24668 2996 24670
rect 2604 23202 2660 23212
rect 1932 23102 1934 23154
rect 1986 23102 1988 23154
rect 1932 23090 1988 23102
rect 2828 22372 2884 24668
rect 2940 24658 2996 24668
rect 3164 24276 3220 24780
rect 3388 24770 3444 24780
rect 2940 24220 3220 24276
rect 3724 24722 3780 24734
rect 6188 24724 6244 25452
rect 6300 25442 6356 25452
rect 3724 24670 3726 24722
rect 3778 24670 3780 24722
rect 2940 24050 2996 24220
rect 2940 23998 2942 24050
rect 2994 23998 2996 24050
rect 2940 23986 2996 23998
rect 3724 23380 3780 24670
rect 5740 24668 6244 24724
rect 6412 24724 6468 24734
rect 6636 24724 6692 27804
rect 7756 27858 7812 28478
rect 8092 28530 8148 28542
rect 8092 28478 8094 28530
rect 8146 28478 8148 28530
rect 7756 27806 7758 27858
rect 7810 27806 7812 27858
rect 7084 27748 7140 27758
rect 7756 27748 7812 27806
rect 6748 27636 6804 27646
rect 6748 27542 6804 27580
rect 7084 27186 7140 27692
rect 7084 27134 7086 27186
rect 7138 27134 7140 27186
rect 7084 27122 7140 27134
rect 7532 27692 7812 27748
rect 7868 27970 7924 27982
rect 7868 27918 7870 27970
rect 7922 27918 7924 27970
rect 7868 27748 7924 27918
rect 6972 26852 7028 26862
rect 6860 26850 7028 26852
rect 6860 26798 6974 26850
rect 7026 26798 7028 26850
rect 6860 26796 7028 26798
rect 6860 25396 6916 26796
rect 6972 26786 7028 26796
rect 7084 26236 7364 26292
rect 6972 26180 7028 26190
rect 7084 26180 7140 26236
rect 6972 26178 7140 26180
rect 6972 26126 6974 26178
rect 7026 26126 7140 26178
rect 6972 26124 7140 26126
rect 6972 26114 7028 26124
rect 7196 26066 7252 26078
rect 7196 26014 7198 26066
rect 7250 26014 7252 26066
rect 6972 25620 7028 25630
rect 7196 25620 7252 26014
rect 6972 25618 7252 25620
rect 6972 25566 6974 25618
rect 7026 25566 7252 25618
rect 6972 25564 7252 25566
rect 6972 25554 7028 25564
rect 6860 25340 7028 25396
rect 6412 24722 6692 24724
rect 6412 24670 6414 24722
rect 6466 24670 6692 24722
rect 6412 24668 6692 24670
rect 6860 25172 6916 25182
rect 6860 24722 6916 25116
rect 6860 24670 6862 24722
rect 6914 24670 6916 24722
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 3724 23314 3780 23324
rect 5068 24050 5124 24062
rect 5740 24052 5796 24668
rect 6412 24658 6468 24668
rect 6860 24658 6916 24670
rect 5068 23998 5070 24050
rect 5122 23998 5124 24050
rect 4732 23042 4788 23054
rect 4732 22990 4734 23042
rect 4786 22990 4788 23042
rect 4732 22932 4788 22990
rect 5068 23044 5124 23998
rect 5068 22978 5124 22988
rect 5180 24050 5796 24052
rect 5180 23998 5742 24050
rect 5794 23998 5796 24050
rect 5180 23996 5796 23998
rect 4732 22866 4788 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 5068 22484 5124 22494
rect 5180 22484 5236 23996
rect 5740 23986 5796 23996
rect 5404 23380 5460 23390
rect 5404 23286 5460 23324
rect 6412 23266 6468 23278
rect 6412 23214 6414 23266
rect 6466 23214 6468 23266
rect 5740 23044 5796 23054
rect 5740 22930 5796 22988
rect 5740 22878 5742 22930
rect 5794 22878 5796 22930
rect 5740 22596 5796 22878
rect 5740 22530 5796 22540
rect 6076 22932 6132 22942
rect 6076 22594 6132 22876
rect 6076 22542 6078 22594
rect 6130 22542 6132 22594
rect 6076 22530 6132 22542
rect 6412 22708 6468 23214
rect 5068 22482 5236 22484
rect 5068 22430 5070 22482
rect 5122 22430 5236 22482
rect 5068 22428 5236 22430
rect 5068 22418 5124 22428
rect 2828 22306 2884 22316
rect 5740 22372 5796 22382
rect 5740 22278 5796 22316
rect 3612 22258 3668 22270
rect 3612 22206 3614 22258
rect 3666 22206 3668 22258
rect 3276 22148 3332 22158
rect 3052 22146 3332 22148
rect 3052 22094 3278 22146
rect 3330 22094 3332 22146
rect 3052 22092 3332 22094
rect 3052 21698 3108 22092
rect 3276 22082 3332 22092
rect 3052 21646 3054 21698
rect 3106 21646 3108 21698
rect 3052 21634 3108 21646
rect 2268 21586 2324 21598
rect 2268 21534 2270 21586
rect 2322 21534 2324 21586
rect 1820 20802 1876 20814
rect 1820 20750 1822 20802
rect 1874 20750 1876 20802
rect 1820 20188 1876 20750
rect 2268 20188 2324 21534
rect 3612 21028 3668 22206
rect 6412 22148 6468 22652
rect 6524 23156 6580 23166
rect 6524 22370 6580 23100
rect 6524 22318 6526 22370
rect 6578 22318 6580 22370
rect 6524 22306 6580 22318
rect 6860 22258 6916 22270
rect 6860 22206 6862 22258
rect 6914 22206 6916 22258
rect 6860 22148 6916 22206
rect 6412 22092 6804 22148
rect 5180 21474 5236 21486
rect 5180 21422 5182 21474
rect 5234 21422 5236 21474
rect 5180 21364 5236 21422
rect 5628 21474 5684 21486
rect 5628 21422 5630 21474
rect 5682 21422 5684 21474
rect 5404 21364 5460 21374
rect 5180 21362 5460 21364
rect 5180 21310 5406 21362
rect 5458 21310 5460 21362
rect 5180 21308 5460 21310
rect 5404 21298 5460 21308
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 3612 20962 3668 20972
rect 4620 20914 4676 20926
rect 4620 20862 4622 20914
rect 4674 20862 4676 20914
rect 2492 20690 2548 20702
rect 2492 20638 2494 20690
rect 2546 20638 2548 20690
rect 2492 20242 2548 20638
rect 4620 20356 4676 20862
rect 5068 20580 5124 20590
rect 5628 20580 5684 21422
rect 5740 21364 5796 21374
rect 5740 21362 5908 21364
rect 5740 21310 5742 21362
rect 5794 21310 5908 21362
rect 5740 21308 5908 21310
rect 5740 21298 5796 21308
rect 5740 21028 5796 21038
rect 5740 20934 5796 20972
rect 5852 20804 5908 21308
rect 6076 20804 6132 20814
rect 5852 20802 6132 20804
rect 5852 20750 6078 20802
rect 6130 20750 6132 20802
rect 5852 20748 6132 20750
rect 5068 20578 5684 20580
rect 5068 20526 5070 20578
rect 5122 20526 5684 20578
rect 5068 20524 5684 20526
rect 5068 20514 5124 20524
rect 4620 20290 4676 20300
rect 2492 20190 2494 20242
rect 2546 20190 2548 20242
rect 1820 20132 2436 20188
rect 2492 20178 2548 20190
rect 2268 18562 2324 18574
rect 2268 18510 2270 18562
rect 2322 18510 2324 18562
rect 2044 18450 2100 18462
rect 2044 18398 2046 18450
rect 2098 18398 2100 18450
rect 2044 17892 2100 18398
rect 2044 17826 2100 17836
rect 2268 17780 2324 18510
rect 2380 18452 2436 20132
rect 2828 20020 2884 20030
rect 2828 19926 2884 19964
rect 5068 20020 5124 20030
rect 5068 19926 5124 19964
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4060 19122 4116 19134
rect 4060 19070 4062 19122
rect 4114 19070 4116 19122
rect 3724 19012 3780 19022
rect 3388 19010 3780 19012
rect 3388 18958 3726 19010
rect 3778 18958 3780 19010
rect 3388 18956 3780 18958
rect 3388 18562 3444 18956
rect 3724 18946 3780 18956
rect 3388 18510 3390 18562
rect 3442 18510 3444 18562
rect 3388 18498 3444 18510
rect 2716 18452 2772 18462
rect 2380 18450 2772 18452
rect 2380 18398 2718 18450
rect 2770 18398 2772 18450
rect 2380 18396 2772 18398
rect 2492 17780 2548 17790
rect 2268 17778 2548 17780
rect 2268 17726 2494 17778
rect 2546 17726 2548 17778
rect 2268 17724 2548 17726
rect 2492 17714 2548 17724
rect 1820 17666 1876 17678
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1820 15092 1876 17614
rect 2156 15876 2212 15886
rect 2156 15314 2212 15820
rect 2156 15262 2158 15314
rect 2210 15262 2212 15314
rect 2156 15250 2212 15262
rect 2380 15426 2436 15438
rect 2380 15374 2382 15426
rect 2434 15374 2436 15426
rect 1820 14530 1876 15036
rect 2380 14644 2436 15374
rect 2716 15316 2772 18396
rect 4060 18452 4116 19070
rect 5180 19012 5236 20524
rect 5404 20356 5460 20366
rect 5404 20018 5460 20300
rect 5404 19966 5406 20018
rect 5458 19966 5460 20018
rect 5404 19954 5460 19966
rect 5964 20130 6020 20142
rect 5964 20078 5966 20130
rect 6018 20078 6020 20130
rect 5964 20020 6020 20078
rect 6076 20132 6132 20748
rect 6300 20692 6356 20702
rect 6076 20066 6132 20076
rect 6188 20690 6356 20692
rect 6188 20638 6302 20690
rect 6354 20638 6356 20690
rect 6188 20636 6356 20638
rect 5964 19954 6020 19964
rect 6188 20018 6244 20636
rect 6300 20626 6356 20636
rect 6748 20690 6804 22092
rect 6748 20638 6750 20690
rect 6802 20638 6804 20690
rect 6748 20626 6804 20638
rect 6188 19966 6190 20018
rect 6242 19966 6244 20018
rect 6188 19908 6244 19966
rect 6860 20020 6916 22092
rect 6972 21698 7028 25340
rect 7196 24836 7252 24846
rect 7308 24836 7364 26236
rect 7420 26180 7476 26190
rect 7420 26086 7476 26124
rect 7196 24834 7364 24836
rect 7196 24782 7198 24834
rect 7250 24782 7364 24834
rect 7196 24780 7364 24782
rect 7196 24770 7252 24780
rect 7308 24050 7364 24780
rect 7308 23998 7310 24050
rect 7362 23998 7364 24050
rect 7308 23986 7364 23998
rect 7532 23940 7588 27692
rect 7868 27682 7924 27692
rect 8092 26964 8148 28478
rect 8204 27972 8260 29260
rect 8428 27972 8484 27982
rect 8204 27916 8428 27972
rect 8428 27878 8484 27916
rect 8316 27636 8372 27646
rect 8316 27542 8372 27580
rect 8540 27188 8596 29372
rect 8092 26898 8148 26908
rect 8204 27132 8596 27188
rect 9212 28642 9268 30940
rect 9548 30930 9604 30940
rect 9548 30100 9604 30110
rect 9548 30006 9604 30044
rect 9772 29988 9828 38612
rect 10780 38162 10836 38668
rect 12236 38668 12292 39004
rect 12348 38834 12404 39676
rect 14364 39732 14420 39742
rect 14700 39732 14756 41804
rect 14812 41748 14868 42476
rect 14812 41300 14868 41692
rect 14812 41234 14868 41244
rect 14924 41188 14980 42700
rect 15372 41972 15428 43036
rect 15708 42868 15764 42878
rect 15708 42774 15764 42812
rect 15820 42196 15876 44268
rect 15932 44100 15988 44492
rect 15932 44034 15988 44044
rect 16044 43988 16100 45388
rect 16492 45218 16548 45230
rect 16492 45166 16494 45218
rect 16546 45166 16548 45218
rect 16492 45108 16548 45166
rect 16156 45052 16548 45108
rect 16716 45106 16772 45118
rect 16716 45054 16718 45106
rect 16770 45054 16772 45106
rect 16156 44212 16212 45052
rect 16380 44884 16436 44894
rect 16156 44118 16212 44156
rect 16268 44828 16380 44884
rect 16268 44100 16324 44828
rect 16380 44818 16436 44828
rect 16716 44884 16772 45054
rect 16716 44818 16772 44828
rect 16380 44324 16436 44334
rect 16380 44230 16436 44268
rect 16604 44324 16660 44334
rect 16604 44322 16772 44324
rect 16604 44270 16606 44322
rect 16658 44270 16772 44322
rect 16604 44268 16772 44270
rect 16604 44258 16660 44268
rect 16716 44100 16772 44268
rect 16268 44044 16660 44100
rect 16044 43932 16436 43988
rect 16380 43764 16436 43932
rect 16268 43708 16436 43764
rect 16156 43652 16212 43662
rect 16156 43538 16212 43596
rect 16156 43486 16158 43538
rect 16210 43486 16212 43538
rect 16156 43474 16212 43486
rect 15596 42140 15876 42196
rect 15932 42868 15988 42878
rect 15484 41972 15540 41982
rect 15148 41970 15540 41972
rect 15148 41918 15486 41970
rect 15538 41918 15540 41970
rect 15148 41916 15540 41918
rect 15036 41188 15092 41198
rect 14924 41186 15092 41188
rect 14924 41134 15038 41186
rect 15090 41134 15092 41186
rect 14924 41132 15092 41134
rect 15036 41122 15092 41132
rect 15148 41074 15204 41916
rect 15484 41906 15540 41916
rect 15372 41748 15428 41758
rect 15372 41654 15428 41692
rect 15148 41022 15150 41074
rect 15202 41022 15204 41074
rect 15148 41010 15204 41022
rect 14364 39730 14756 39732
rect 14364 39678 14366 39730
rect 14418 39678 14756 39730
rect 14364 39676 14756 39678
rect 14812 40962 14868 40974
rect 14812 40910 14814 40962
rect 14866 40910 14868 40962
rect 14364 39666 14420 39676
rect 14252 39620 14308 39630
rect 14252 39526 14308 39564
rect 12908 39508 12964 39518
rect 12348 38782 12350 38834
rect 12402 38782 12404 38834
rect 12348 38770 12404 38782
rect 12572 38834 12628 38846
rect 12572 38782 12574 38834
rect 12626 38782 12628 38834
rect 12572 38668 12628 38782
rect 12236 38612 12628 38668
rect 10780 38110 10782 38162
rect 10834 38110 10836 38162
rect 10780 38098 10836 38110
rect 12908 38162 12964 39452
rect 14476 39396 14532 39406
rect 14812 39396 14868 40910
rect 15372 40962 15428 40974
rect 15372 40910 15374 40962
rect 15426 40910 15428 40962
rect 14924 40404 14980 40414
rect 14924 40310 14980 40348
rect 15148 40404 15204 40414
rect 15204 40348 15316 40404
rect 15148 40338 15204 40348
rect 15036 40292 15092 40302
rect 15036 40180 15092 40236
rect 15148 40180 15204 40190
rect 15036 40178 15204 40180
rect 15036 40126 15150 40178
rect 15202 40126 15204 40178
rect 15036 40124 15204 40126
rect 15148 40114 15204 40124
rect 14924 39620 14980 39630
rect 14924 39526 14980 39564
rect 15148 39508 15204 39518
rect 15260 39508 15316 40348
rect 15148 39506 15316 39508
rect 15148 39454 15150 39506
rect 15202 39454 15316 39506
rect 15148 39452 15316 39454
rect 15148 39442 15204 39452
rect 14476 39394 14756 39396
rect 14476 39342 14478 39394
rect 14530 39342 14756 39394
rect 14476 39340 14756 39342
rect 14812 39340 15092 39396
rect 12908 38110 12910 38162
rect 12962 38110 12964 38162
rect 12908 38098 12964 38110
rect 13020 39284 13076 39294
rect 13020 38722 13076 39228
rect 13356 38836 13412 38846
rect 13356 38742 13412 38780
rect 13020 38670 13022 38722
rect 13074 38670 13076 38722
rect 10108 38050 10164 38062
rect 10108 37998 10110 38050
rect 10162 37998 10164 38050
rect 10108 37156 10164 37998
rect 13020 37940 13076 38670
rect 14364 38276 14420 38286
rect 13692 38164 13748 38174
rect 13692 38162 14308 38164
rect 13692 38110 13694 38162
rect 13746 38110 14308 38162
rect 13692 38108 14308 38110
rect 13692 38098 13748 38108
rect 12796 37884 13076 37940
rect 13580 37940 13636 37950
rect 14028 37940 14084 37950
rect 13580 37938 14084 37940
rect 13580 37886 13582 37938
rect 13634 37886 14030 37938
rect 14082 37886 14084 37938
rect 13580 37884 14084 37886
rect 10108 37090 10164 37100
rect 10332 37154 10388 37166
rect 10332 37102 10334 37154
rect 10386 37102 10388 37154
rect 10332 37044 10388 37102
rect 12460 37156 12516 37166
rect 12796 37156 12852 37884
rect 13580 37874 13636 37884
rect 14028 37828 14084 37884
rect 14028 37762 14084 37772
rect 14140 37826 14196 37838
rect 14140 37774 14142 37826
rect 14194 37774 14196 37826
rect 14140 37604 14196 37774
rect 14252 37828 14308 38108
rect 14364 38050 14420 38220
rect 14476 38164 14532 39340
rect 14700 39172 14756 39340
rect 15036 39284 15092 39340
rect 15036 39228 15316 39284
rect 14700 39116 15204 39172
rect 15148 39058 15204 39116
rect 15148 39006 15150 39058
rect 15202 39006 15204 39058
rect 15148 38994 15204 39006
rect 14812 38948 14868 38958
rect 14812 38854 14868 38892
rect 15036 38834 15092 38846
rect 15036 38782 15038 38834
rect 15090 38782 15092 38834
rect 15036 38276 15092 38782
rect 15148 38612 15204 38622
rect 15148 38518 15204 38556
rect 15260 38388 15316 39228
rect 15036 38210 15092 38220
rect 15148 38332 15316 38388
rect 14476 38108 14868 38164
rect 14364 37998 14366 38050
rect 14418 37998 14420 38050
rect 14364 37986 14420 37998
rect 14812 38050 14868 38108
rect 14812 37998 14814 38050
rect 14866 37998 14868 38050
rect 14588 37938 14644 37950
rect 14588 37886 14590 37938
rect 14642 37886 14644 37938
rect 14588 37828 14644 37886
rect 14252 37772 14644 37828
rect 14812 37716 14868 37998
rect 15036 38052 15092 38062
rect 15036 37958 15092 37996
rect 14140 37538 14196 37548
rect 14588 37660 14812 37716
rect 12460 37154 12852 37156
rect 12460 37102 12462 37154
rect 12514 37102 12852 37154
rect 12460 37100 12852 37102
rect 12908 37156 12964 37166
rect 13356 37156 13412 37166
rect 12964 37154 13412 37156
rect 12964 37102 13358 37154
rect 13410 37102 13412 37154
rect 12964 37100 13412 37102
rect 12460 37090 12516 37100
rect 10332 36978 10388 36988
rect 12012 35698 12068 35710
rect 12012 35646 12014 35698
rect 12066 35646 12068 35698
rect 12012 35364 12068 35646
rect 12012 35298 12068 35308
rect 12684 35586 12740 35598
rect 12684 35534 12686 35586
rect 12738 35534 12740 35586
rect 12684 35140 12740 35534
rect 12908 35364 12964 37100
rect 13356 37090 13412 37100
rect 14476 37156 14532 37166
rect 14476 37062 14532 37100
rect 14588 36370 14644 37660
rect 14812 37650 14868 37660
rect 14924 37826 14980 37838
rect 14924 37774 14926 37826
rect 14978 37774 14980 37826
rect 14700 37380 14756 37390
rect 14924 37380 14980 37774
rect 15148 37716 15204 38332
rect 15260 38050 15316 38062
rect 15260 37998 15262 38050
rect 15314 37998 15316 38050
rect 15260 37940 15316 37998
rect 15260 37874 15316 37884
rect 15372 37828 15428 40910
rect 15484 40628 15540 40638
rect 15596 40628 15652 42140
rect 15484 40626 15652 40628
rect 15484 40574 15486 40626
rect 15538 40574 15652 40626
rect 15484 40572 15652 40574
rect 15484 40562 15540 40572
rect 15484 39508 15540 39518
rect 15484 39414 15540 39452
rect 15596 39284 15652 40572
rect 15708 41972 15764 41982
rect 15708 39620 15764 41916
rect 15932 41970 15988 42812
rect 16268 42756 16324 43708
rect 16604 43538 16660 44044
rect 16716 44034 16772 44044
rect 16828 44322 16884 44334
rect 16828 44270 16830 44322
rect 16882 44270 16884 44322
rect 16828 43652 16884 44270
rect 16828 43586 16884 43596
rect 16604 43486 16606 43538
rect 16658 43486 16660 43538
rect 16604 43474 16660 43486
rect 16828 43428 16884 43438
rect 16380 43316 16436 43326
rect 16380 43222 16436 43260
rect 16380 42980 16436 42990
rect 16380 42886 16436 42924
rect 16828 42756 16884 43372
rect 16268 42700 16436 42756
rect 16268 42530 16324 42542
rect 16268 42478 16270 42530
rect 16322 42478 16324 42530
rect 16268 42420 16324 42478
rect 15932 41918 15934 41970
rect 15986 41918 15988 41970
rect 15932 40628 15988 41918
rect 16044 42364 16324 42420
rect 16044 41748 16100 42364
rect 16268 42196 16324 42206
rect 16380 42196 16436 42700
rect 16604 42700 16884 42756
rect 16492 42644 16548 42654
rect 16492 42550 16548 42588
rect 16268 42194 16436 42196
rect 16268 42142 16270 42194
rect 16322 42142 16436 42194
rect 16268 42140 16436 42142
rect 16268 42130 16324 42140
rect 16156 41972 16212 41982
rect 16492 41972 16548 41982
rect 16156 41970 16548 41972
rect 16156 41918 16158 41970
rect 16210 41918 16494 41970
rect 16546 41918 16548 41970
rect 16156 41916 16548 41918
rect 16156 41906 16212 41916
rect 16492 41906 16548 41916
rect 16492 41748 16548 41758
rect 16100 41692 16212 41748
rect 16044 41654 16100 41692
rect 16044 41188 16100 41198
rect 16044 41094 16100 41132
rect 16156 40740 16212 41692
rect 16268 41636 16324 41646
rect 16268 41186 16324 41580
rect 16268 41134 16270 41186
rect 16322 41134 16324 41186
rect 16268 41122 16324 41134
rect 16492 41188 16548 41692
rect 16492 41094 16548 41132
rect 16380 40964 16436 40974
rect 16380 40870 16436 40908
rect 16156 40684 16324 40740
rect 15932 40562 15988 40572
rect 16156 40514 16212 40526
rect 16156 40462 16158 40514
rect 16210 40462 16212 40514
rect 15932 40402 15988 40414
rect 15932 40350 15934 40402
rect 15986 40350 15988 40402
rect 15932 40292 15988 40350
rect 15932 40226 15988 40236
rect 16156 40180 16212 40462
rect 16268 40404 16324 40684
rect 16268 40338 16324 40348
rect 16604 40292 16660 42700
rect 16940 42642 16996 42654
rect 16940 42590 16942 42642
rect 16994 42590 16996 42642
rect 16716 42530 16772 42542
rect 16716 42478 16718 42530
rect 16770 42478 16772 42530
rect 16716 42194 16772 42478
rect 16716 42142 16718 42194
rect 16770 42142 16772 42194
rect 16716 41972 16772 42142
rect 16828 42196 16884 42206
rect 16940 42196 16996 42590
rect 16884 42140 16996 42196
rect 16828 42082 16884 42140
rect 16828 42030 16830 42082
rect 16882 42030 16884 42082
rect 16828 42018 16884 42030
rect 16716 41906 16772 41916
rect 17052 41860 17108 52668
rect 17724 52276 17780 52286
rect 17724 51602 17780 52220
rect 18284 52276 18340 52286
rect 18284 52182 18340 52220
rect 18732 52164 18788 52174
rect 18508 52108 18732 52164
rect 17724 51550 17726 51602
rect 17778 51550 17780 51602
rect 17724 51538 17780 51550
rect 18172 51940 18228 51950
rect 17612 51492 17668 51502
rect 17388 51436 17612 51492
rect 17388 49922 17444 51436
rect 17612 51398 17668 51436
rect 18172 51490 18228 51884
rect 18172 51438 18174 51490
rect 18226 51438 18228 51490
rect 17948 51378 18004 51390
rect 17948 51326 17950 51378
rect 18002 51326 18004 51378
rect 17388 49870 17390 49922
rect 17442 49870 17444 49922
rect 17388 49858 17444 49870
rect 17612 51044 17668 51054
rect 17612 49810 17668 50988
rect 17948 50932 18004 51326
rect 17948 50866 18004 50876
rect 18172 51380 18228 51438
rect 18172 50594 18228 51324
rect 18396 51492 18452 51502
rect 18396 51378 18452 51436
rect 18396 51326 18398 51378
rect 18450 51326 18452 51378
rect 18396 51314 18452 51326
rect 18508 50820 18564 52108
rect 18732 52070 18788 52108
rect 18732 51268 18788 51278
rect 18732 51174 18788 51212
rect 18732 51044 18788 51054
rect 18508 50764 18676 50820
rect 18172 50542 18174 50594
rect 18226 50542 18228 50594
rect 18172 50530 18228 50542
rect 18396 50596 18452 50606
rect 18396 50482 18452 50540
rect 18396 50430 18398 50482
rect 18450 50430 18452 50482
rect 18396 50418 18452 50430
rect 18508 50372 18564 50382
rect 18508 50278 18564 50316
rect 17948 50036 18004 50046
rect 18284 50036 18340 50046
rect 17948 50034 18340 50036
rect 17948 49982 17950 50034
rect 18002 49982 18286 50034
rect 18338 49982 18340 50034
rect 17948 49980 18340 49982
rect 17948 49970 18004 49980
rect 18284 49970 18340 49980
rect 17612 49758 17614 49810
rect 17666 49758 17668 49810
rect 17612 49746 17668 49758
rect 18508 49810 18564 49822
rect 18508 49758 18510 49810
rect 18562 49758 18564 49810
rect 18172 49588 18228 49598
rect 17948 49586 18228 49588
rect 17948 49534 18174 49586
rect 18226 49534 18228 49586
rect 17948 49532 18228 49534
rect 17052 41794 17108 41804
rect 17164 49028 17220 49038
rect 16940 41524 16996 41534
rect 16380 40236 16660 40292
rect 16828 41468 16940 41524
rect 16380 40180 16436 40236
rect 16156 40124 16436 40180
rect 16156 39620 16212 40124
rect 15708 39564 15876 39620
rect 15484 39228 15652 39284
rect 15484 38612 15540 39228
rect 15708 39060 15764 39070
rect 15708 38966 15764 39004
rect 15596 38724 15652 38762
rect 15596 38658 15652 38668
rect 15820 38724 15876 39564
rect 16044 39564 16156 39620
rect 15932 39396 15988 39406
rect 15932 38946 15988 39340
rect 15932 38894 15934 38946
rect 15986 38894 15988 38946
rect 15932 38882 15988 38894
rect 15484 38546 15540 38556
rect 15820 38050 15876 38668
rect 15820 37998 15822 38050
rect 15874 37998 15876 38050
rect 15820 37986 15876 37998
rect 15596 37828 15652 37838
rect 15372 37772 15596 37828
rect 15148 37660 15316 37716
rect 15036 37604 15092 37614
rect 15092 37548 15204 37604
rect 15036 37538 15092 37548
rect 14700 37378 14980 37380
rect 14700 37326 14702 37378
rect 14754 37326 14980 37378
rect 14700 37324 14980 37326
rect 15036 37380 15092 37390
rect 14700 37314 14756 37324
rect 15036 37286 15092 37324
rect 14812 37154 14868 37166
rect 14812 37102 14814 37154
rect 14866 37102 14868 37154
rect 14812 37044 14868 37102
rect 15148 37044 15204 37548
rect 15260 37492 15316 37660
rect 15260 37426 15316 37436
rect 15596 37378 15652 37772
rect 15820 37716 15876 37726
rect 15820 37490 15876 37660
rect 15820 37438 15822 37490
rect 15874 37438 15876 37490
rect 15820 37426 15876 37438
rect 16044 37492 16100 39564
rect 16156 39554 16212 39564
rect 16268 39956 16324 39966
rect 16156 39396 16212 39406
rect 16268 39396 16324 39900
rect 16604 39508 16660 39518
rect 16156 39394 16324 39396
rect 16156 39342 16158 39394
rect 16210 39342 16324 39394
rect 16156 39340 16324 39342
rect 16492 39506 16660 39508
rect 16492 39454 16606 39506
rect 16658 39454 16660 39506
rect 16492 39452 16660 39454
rect 16156 39060 16212 39340
rect 16156 38994 16212 39004
rect 16492 38668 16548 39452
rect 16604 39442 16660 39452
rect 16716 39396 16772 39406
rect 16716 39302 16772 39340
rect 16828 39172 16884 41468
rect 16940 41458 16996 41468
rect 17052 41412 17108 41422
rect 17052 41300 17108 41356
rect 16940 41244 17108 41300
rect 16940 41186 16996 41244
rect 16940 41134 16942 41186
rect 16994 41134 16996 41186
rect 16940 41122 16996 41134
rect 16940 40852 16996 40862
rect 16940 39618 16996 40796
rect 16940 39566 16942 39618
rect 16994 39566 16996 39618
rect 16940 39554 16996 39566
rect 17052 40068 17108 40078
rect 16604 39116 16884 39172
rect 16604 38948 16660 39116
rect 16604 38834 16660 38892
rect 16604 38782 16606 38834
rect 16658 38782 16660 38834
rect 16604 38770 16660 38782
rect 16828 38836 16884 38846
rect 17052 38836 17108 40012
rect 16828 38834 17108 38836
rect 16828 38782 16830 38834
rect 16882 38782 17108 38834
rect 16828 38780 17108 38782
rect 16828 38770 16884 38780
rect 16268 38610 16324 38622
rect 16268 38558 16270 38610
rect 16322 38558 16324 38610
rect 16044 37426 16100 37436
rect 16156 37604 16212 37614
rect 16156 37490 16212 37548
rect 16156 37438 16158 37490
rect 16210 37438 16212 37490
rect 16156 37426 16212 37438
rect 15596 37326 15598 37378
rect 15650 37326 15652 37378
rect 15596 37314 15652 37326
rect 14812 36978 14868 36988
rect 15036 36988 15204 37044
rect 15260 37266 15316 37278
rect 15260 37214 15262 37266
rect 15314 37214 15316 37266
rect 15260 37156 15316 37214
rect 16268 37268 16324 38558
rect 16492 38612 16660 38668
rect 16492 38546 16548 38556
rect 16380 38052 16436 38062
rect 16380 37490 16436 37996
rect 16380 37438 16382 37490
rect 16434 37438 16436 37490
rect 16380 37426 16436 37438
rect 16268 37202 16324 37212
rect 16492 37266 16548 37278
rect 16492 37214 16494 37266
rect 16546 37214 16548 37266
rect 14588 36318 14590 36370
rect 14642 36318 14644 36370
rect 14588 36306 14644 36318
rect 14924 36258 14980 36270
rect 14924 36206 14926 36258
rect 14978 36206 14980 36258
rect 14924 35812 14980 36206
rect 14812 35700 14868 35710
rect 14812 35586 14868 35644
rect 14812 35534 14814 35586
rect 14866 35534 14868 35586
rect 14812 35522 14868 35534
rect 12908 35298 12964 35308
rect 13804 35476 13860 35486
rect 12684 35074 12740 35084
rect 13468 35140 13524 35150
rect 13468 35046 13524 35084
rect 13804 35138 13860 35420
rect 13804 35086 13806 35138
rect 13858 35086 13860 35138
rect 13804 35074 13860 35086
rect 14588 35252 14644 35262
rect 14588 35026 14644 35196
rect 14588 34974 14590 35026
rect 14642 34974 14644 35026
rect 14588 34962 14644 34974
rect 14812 35028 14868 35038
rect 14924 35028 14980 35756
rect 15036 35138 15092 36988
rect 15036 35086 15038 35138
rect 15090 35086 15092 35138
rect 15036 35074 15092 35086
rect 14812 35026 14980 35028
rect 14812 34974 14814 35026
rect 14866 34974 14980 35026
rect 14812 34972 14980 34974
rect 14812 34962 14868 34972
rect 13580 34690 13636 34702
rect 13580 34638 13582 34690
rect 13634 34638 13636 34690
rect 13580 33684 13636 34638
rect 13468 33628 13580 33684
rect 12348 33348 12404 33358
rect 12348 32562 12404 33292
rect 13468 32676 13524 33628
rect 13580 33618 13636 33628
rect 14028 34244 14084 34254
rect 14700 34244 14756 34254
rect 14028 34242 14756 34244
rect 14028 34190 14030 34242
rect 14082 34190 14702 34242
rect 14754 34190 14756 34242
rect 14028 34188 14756 34190
rect 13580 33348 13636 33358
rect 13580 33254 13636 33292
rect 13468 32620 13636 32676
rect 12348 32510 12350 32562
rect 12402 32510 12404 32562
rect 12348 32498 12404 32510
rect 13020 32450 13076 32462
rect 13020 32398 13022 32450
rect 13074 32398 13076 32450
rect 13020 31892 13076 32398
rect 13020 31826 13076 31836
rect 13468 31668 13524 31678
rect 13244 31612 13468 31668
rect 13244 31106 13300 31612
rect 13468 31574 13524 31612
rect 13468 31220 13524 31230
rect 13580 31220 13636 32620
rect 13692 31892 13748 31902
rect 13692 31798 13748 31836
rect 13804 31778 13860 31790
rect 13804 31726 13806 31778
rect 13858 31726 13860 31778
rect 13804 31556 13860 31726
rect 14028 31556 14084 34188
rect 14700 34178 14756 34188
rect 15260 34132 15316 37100
rect 15708 37156 15764 37166
rect 15484 36708 15540 36718
rect 15484 35700 15540 36652
rect 15484 35606 15540 35644
rect 15708 35698 15764 37100
rect 15708 35646 15710 35698
rect 15762 35646 15764 35698
rect 15708 35634 15764 35646
rect 15932 37042 15988 37054
rect 15932 36990 15934 37042
rect 15986 36990 15988 37042
rect 15932 35698 15988 36990
rect 16492 36932 16548 37214
rect 16604 37044 16660 38612
rect 16604 36978 16660 36988
rect 15932 35646 15934 35698
rect 15986 35646 15988 35698
rect 15932 35634 15988 35646
rect 16044 36370 16100 36382
rect 16044 36318 16046 36370
rect 16098 36318 16100 36370
rect 15596 35588 15652 35598
rect 15596 35494 15652 35532
rect 15820 35252 15876 35262
rect 15820 34914 15876 35196
rect 15820 34862 15822 34914
rect 15874 34862 15876 34914
rect 15820 34850 15876 34862
rect 15372 34690 15428 34702
rect 15372 34638 15374 34690
rect 15426 34638 15428 34690
rect 15372 34356 15428 34638
rect 15596 34356 15652 34366
rect 15932 34356 15988 34366
rect 16044 34356 16100 36318
rect 16156 35924 16212 35934
rect 16156 35810 16212 35868
rect 16156 35758 16158 35810
rect 16210 35758 16212 35810
rect 16156 35746 16212 35758
rect 16492 35698 16548 36876
rect 17052 36260 17108 38780
rect 17052 36194 17108 36204
rect 17164 38162 17220 48972
rect 17836 48916 17892 48926
rect 17612 48914 17892 48916
rect 17612 48862 17838 48914
rect 17890 48862 17892 48914
rect 17612 48860 17892 48862
rect 17500 48468 17556 48478
rect 17388 48412 17500 48468
rect 17276 48242 17332 48254
rect 17276 48190 17278 48242
rect 17330 48190 17332 48242
rect 17276 47124 17332 48190
rect 17276 47058 17332 47068
rect 17388 46900 17444 48412
rect 17500 48402 17556 48412
rect 17612 48466 17668 48860
rect 17836 48850 17892 48860
rect 17948 48692 18004 49532
rect 18172 49522 18228 49532
rect 17612 48414 17614 48466
rect 17666 48414 17668 48466
rect 17612 48402 17668 48414
rect 17724 48636 18004 48692
rect 17724 48354 17780 48636
rect 18508 48468 18564 49758
rect 18620 49028 18676 50764
rect 18732 49922 18788 50988
rect 18732 49870 18734 49922
rect 18786 49870 18788 49922
rect 18732 49858 18788 49870
rect 18620 48962 18676 48972
rect 18844 48804 18900 54238
rect 18956 53954 19012 55132
rect 19068 55094 19124 55132
rect 21756 55186 21812 57148
rect 21980 55970 22036 59200
rect 22428 56084 22484 56094
rect 22428 56082 22820 56084
rect 22428 56030 22430 56082
rect 22482 56030 22820 56082
rect 22428 56028 22820 56030
rect 22428 56018 22484 56028
rect 21980 55918 21982 55970
rect 22034 55918 22036 55970
rect 21980 55906 22036 55918
rect 21756 55134 21758 55186
rect 21810 55134 21812 55186
rect 21756 55122 21812 55134
rect 21868 55300 21924 55310
rect 19964 55076 20020 55114
rect 19628 55020 19964 55076
rect 19628 54516 19684 55020
rect 19964 55010 20020 55020
rect 21420 55076 21476 55086
rect 21420 54982 21476 55020
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19516 54514 19684 54516
rect 19516 54462 19630 54514
rect 19682 54462 19684 54514
rect 19516 54460 19684 54462
rect 18956 53902 18958 53954
rect 19010 53902 19012 53954
rect 18956 53890 19012 53902
rect 19292 54404 19348 54414
rect 19180 53730 19236 53742
rect 19180 53678 19182 53730
rect 19234 53678 19236 53730
rect 19180 53508 19236 53678
rect 19180 53442 19236 53452
rect 19292 53506 19348 54348
rect 19292 53454 19294 53506
rect 19346 53454 19348 53506
rect 19292 53442 19348 53454
rect 19404 52948 19460 52958
rect 19516 52948 19572 54460
rect 19628 54450 19684 54460
rect 20412 54404 20468 54414
rect 20412 54310 20468 54348
rect 19852 54292 19908 54302
rect 19740 53620 19796 53630
rect 19740 53526 19796 53564
rect 19404 52946 19572 52948
rect 19404 52894 19406 52946
rect 19458 52894 19572 52946
rect 19404 52892 19572 52894
rect 19628 53508 19684 53518
rect 19068 52836 19124 52846
rect 19404 52836 19460 52892
rect 19068 52834 19460 52836
rect 19068 52782 19070 52834
rect 19122 52782 19460 52834
rect 19068 52780 19460 52782
rect 19068 52164 19124 52780
rect 19068 52098 19124 52108
rect 19180 52276 19236 52286
rect 19180 52050 19236 52220
rect 19180 51998 19182 52050
rect 19234 51998 19236 52050
rect 19068 51940 19124 51950
rect 19068 51846 19124 51884
rect 19068 51492 19124 51502
rect 19068 51398 19124 51436
rect 19180 51268 19236 51998
rect 19628 52164 19684 53452
rect 19852 53506 19908 54236
rect 20636 53844 20692 53854
rect 20692 53788 20804 53844
rect 20636 53778 20692 53788
rect 20300 53730 20356 53742
rect 20300 53678 20302 53730
rect 20354 53678 20356 53730
rect 19852 53454 19854 53506
rect 19906 53454 19908 53506
rect 19852 53442 19908 53454
rect 20188 53620 20244 53630
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 20188 53058 20244 53564
rect 20188 53006 20190 53058
rect 20242 53006 20244 53058
rect 20188 52994 20244 53006
rect 20300 52386 20356 53678
rect 20300 52334 20302 52386
rect 20354 52334 20356 52386
rect 20300 52322 20356 52334
rect 20636 53508 20692 53518
rect 20524 52276 20580 52286
rect 20412 52220 20524 52276
rect 19852 52164 19908 52174
rect 20412 52164 20468 52220
rect 20524 52210 20580 52220
rect 19628 52162 20244 52164
rect 19628 52110 19854 52162
rect 19906 52110 20244 52162
rect 19628 52108 20244 52110
rect 19068 51212 19236 51268
rect 19292 51378 19348 51390
rect 19292 51326 19294 51378
rect 19346 51326 19348 51378
rect 18956 50706 19012 50718
rect 18956 50654 18958 50706
rect 19010 50654 19012 50706
rect 18956 49588 19012 50654
rect 19068 50482 19124 51212
rect 19292 50596 19348 51326
rect 19628 50932 19684 52108
rect 19852 52098 19908 52108
rect 20188 51828 20244 52108
rect 20300 52108 20468 52164
rect 20300 52050 20356 52108
rect 20636 52052 20692 53452
rect 20300 51998 20302 52050
rect 20354 51998 20356 52050
rect 20300 51986 20356 51998
rect 20412 51996 20692 52052
rect 20412 51994 20468 51996
rect 20412 51942 20414 51994
rect 20466 51942 20468 51994
rect 20412 51828 20468 51942
rect 20748 51940 20804 53788
rect 21868 53730 21924 55244
rect 22316 55298 22372 55310
rect 22316 55246 22318 55298
rect 22370 55246 22372 55298
rect 22316 55076 22372 55246
rect 22316 55010 22372 55020
rect 22540 54404 22596 54414
rect 21868 53678 21870 53730
rect 21922 53678 21924 53730
rect 21868 53666 21924 53678
rect 22428 54402 22596 54404
rect 22428 54350 22542 54402
rect 22594 54350 22596 54402
rect 22428 54348 22596 54350
rect 21420 53508 21476 53518
rect 21420 53414 21476 53452
rect 21868 52948 21924 52958
rect 19836 51772 20100 51782
rect 20188 51772 20468 51828
rect 20636 51884 20804 51940
rect 21532 52276 21588 52286
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19852 51378 19908 51390
rect 19852 51326 19854 51378
rect 19906 51326 19908 51378
rect 19740 51268 19796 51278
rect 19852 51268 19908 51326
rect 20188 51378 20244 51390
rect 20188 51326 20190 51378
rect 20242 51326 20244 51378
rect 19796 51212 19908 51268
rect 20076 51268 20132 51278
rect 19740 51202 19796 51212
rect 20076 51174 20132 51212
rect 19964 51156 20020 51166
rect 19292 50530 19348 50540
rect 19404 50876 19684 50932
rect 19740 50932 19796 50942
rect 19068 50430 19070 50482
rect 19122 50430 19124 50482
rect 19068 50418 19124 50430
rect 19404 50428 19460 50876
rect 19180 50372 19236 50382
rect 19180 49810 19236 50316
rect 19180 49758 19182 49810
rect 19234 49758 19236 49810
rect 19180 49746 19236 49758
rect 19292 50372 19460 50428
rect 19516 50596 19572 50606
rect 18956 49140 19012 49532
rect 18956 49074 19012 49084
rect 18508 48402 18564 48412
rect 18620 48748 18900 48804
rect 17724 48302 17726 48354
rect 17778 48302 17780 48354
rect 17724 48290 17780 48302
rect 17948 48242 18004 48254
rect 17948 48190 17950 48242
rect 18002 48190 18004 48242
rect 17948 47236 18004 48190
rect 18620 48244 18676 48748
rect 18620 48150 18676 48188
rect 18844 48356 18900 48366
rect 19180 48356 19236 48366
rect 18844 48354 19236 48356
rect 18844 48302 18846 48354
rect 18898 48302 19182 48354
rect 19234 48302 19236 48354
rect 18844 48300 19236 48302
rect 18620 47570 18676 47582
rect 18620 47518 18622 47570
rect 18674 47518 18676 47570
rect 17948 47170 18004 47180
rect 18172 47460 18228 47470
rect 17276 46844 17444 46900
rect 17276 44546 17332 46844
rect 17388 46564 17444 46574
rect 17388 45106 17444 46508
rect 17612 46564 17668 46574
rect 17612 46470 17668 46508
rect 17948 46452 18004 46462
rect 17836 46450 18004 46452
rect 17836 46398 17950 46450
rect 18002 46398 18004 46450
rect 17836 46396 18004 46398
rect 17388 45054 17390 45106
rect 17442 45054 17444 45106
rect 17388 45042 17444 45054
rect 17612 45218 17668 45230
rect 17612 45166 17614 45218
rect 17666 45166 17668 45218
rect 17612 44772 17668 45166
rect 17612 44706 17668 44716
rect 17724 45108 17780 45118
rect 17276 44494 17278 44546
rect 17330 44494 17332 44546
rect 17276 44482 17332 44494
rect 17500 44660 17556 44670
rect 17388 44436 17444 44446
rect 17388 44342 17444 44380
rect 17500 44322 17556 44604
rect 17500 44270 17502 44322
rect 17554 44270 17556 44322
rect 17500 44258 17556 44270
rect 17724 44210 17780 45052
rect 17724 44158 17726 44210
rect 17778 44158 17780 44210
rect 17276 43876 17332 43886
rect 17276 42644 17332 43820
rect 17724 43876 17780 44158
rect 17724 43810 17780 43820
rect 17612 43652 17668 43662
rect 17612 43558 17668 43596
rect 17724 43650 17780 43662
rect 17724 43598 17726 43650
rect 17778 43598 17780 43650
rect 17724 43540 17780 43598
rect 17724 43474 17780 43484
rect 17836 42868 17892 46396
rect 17948 46386 18004 46396
rect 18172 45890 18228 47404
rect 18508 46676 18564 46686
rect 18172 45838 18174 45890
rect 18226 45838 18228 45890
rect 18172 45826 18228 45838
rect 18396 46002 18452 46014
rect 18396 45950 18398 46002
rect 18450 45950 18452 46002
rect 18172 45444 18228 45454
rect 18060 45108 18116 45118
rect 18060 44994 18116 45052
rect 18060 44942 18062 44994
rect 18114 44942 18116 44994
rect 18060 44930 18116 44942
rect 18060 44324 18116 44334
rect 17276 42578 17332 42588
rect 17724 42812 17892 42868
rect 17948 44322 18116 44324
rect 17948 44270 18062 44322
rect 18114 44270 18116 44322
rect 17948 44268 18116 44270
rect 17948 43538 18004 44268
rect 18060 44258 18116 44268
rect 18172 44100 18228 45388
rect 17948 43486 17950 43538
rect 18002 43486 18004 43538
rect 17500 42532 17556 42542
rect 17500 42530 17668 42532
rect 17500 42478 17502 42530
rect 17554 42478 17668 42530
rect 17500 42476 17668 42478
rect 17500 42466 17556 42476
rect 17612 42308 17668 42476
rect 17612 42194 17668 42252
rect 17612 42142 17614 42194
rect 17666 42142 17668 42194
rect 17388 41970 17444 41982
rect 17388 41918 17390 41970
rect 17442 41918 17444 41970
rect 17388 41636 17444 41918
rect 17500 41972 17556 41982
rect 17500 41878 17556 41916
rect 17612 41748 17668 42142
rect 17612 41682 17668 41692
rect 17444 41580 17556 41636
rect 17388 41570 17444 41580
rect 17500 41524 17556 41580
rect 17724 41524 17780 42812
rect 17500 41468 17668 41524
rect 17388 41412 17444 41422
rect 17388 41186 17444 41356
rect 17388 41134 17390 41186
rect 17442 41134 17444 41186
rect 17388 41122 17444 41134
rect 17276 41076 17332 41086
rect 17276 40982 17332 41020
rect 17500 41074 17556 41086
rect 17500 41022 17502 41074
rect 17554 41022 17556 41074
rect 17388 40964 17444 40974
rect 17500 40964 17556 41022
rect 17444 40908 17556 40964
rect 17388 39730 17444 40908
rect 17612 40628 17668 41468
rect 17724 41458 17780 41468
rect 17836 42642 17892 42654
rect 17836 42590 17838 42642
rect 17890 42590 17892 42642
rect 17612 40534 17668 40572
rect 17388 39678 17390 39730
rect 17442 39678 17444 39730
rect 17388 39666 17444 39678
rect 17836 39508 17892 42590
rect 17948 42196 18004 43486
rect 18060 44044 18228 44100
rect 18284 44660 18340 44670
rect 18060 42642 18116 44044
rect 18284 43538 18340 44604
rect 18396 44436 18452 45950
rect 18396 44370 18452 44380
rect 18284 43486 18286 43538
rect 18338 43486 18340 43538
rect 18284 43474 18340 43486
rect 18508 43204 18564 46620
rect 18620 45892 18676 47518
rect 18620 45826 18676 45836
rect 18732 46786 18788 46798
rect 18732 46734 18734 46786
rect 18786 46734 18788 46786
rect 18732 44660 18788 46734
rect 18732 44594 18788 44604
rect 18620 44324 18676 44334
rect 18620 44100 18676 44268
rect 18620 44034 18676 44044
rect 18732 44322 18788 44334
rect 18732 44270 18734 44322
rect 18786 44270 18788 44322
rect 18732 43540 18788 44270
rect 18284 43148 18564 43204
rect 18620 43316 18676 43326
rect 18172 42980 18228 42990
rect 18172 42886 18228 42924
rect 18060 42590 18062 42642
rect 18114 42590 18116 42642
rect 18060 42578 18116 42590
rect 17948 42140 18228 42196
rect 17948 41970 18004 41982
rect 17948 41918 17950 41970
rect 18002 41918 18004 41970
rect 17948 41860 18004 41918
rect 17948 41794 18004 41804
rect 18060 41972 18116 41982
rect 17948 41412 18004 41422
rect 18060 41412 18116 41916
rect 17948 41410 18116 41412
rect 17948 41358 17950 41410
rect 18002 41358 18116 41410
rect 17948 41356 18116 41358
rect 17948 41346 18004 41356
rect 17948 40964 18004 40974
rect 17948 40516 18004 40908
rect 17948 40402 18004 40460
rect 17948 40350 17950 40402
rect 18002 40350 18004 40402
rect 17948 40068 18004 40350
rect 17948 40002 18004 40012
rect 17388 39452 17892 39508
rect 17948 39844 18004 39854
rect 17164 38110 17166 38162
rect 17218 38110 17220 38162
rect 17164 36036 17220 38110
rect 17276 39394 17332 39406
rect 17276 39342 17278 39394
rect 17330 39342 17332 39394
rect 17276 37156 17332 39342
rect 17276 37090 17332 37100
rect 17388 38946 17444 39452
rect 17388 38894 17390 38946
rect 17442 38894 17444 38946
rect 16492 35646 16494 35698
rect 16546 35646 16548 35698
rect 16492 35634 16548 35646
rect 16828 35980 17220 36036
rect 16828 35922 16884 35980
rect 16828 35870 16830 35922
rect 16882 35870 16884 35922
rect 16828 35252 16884 35870
rect 17388 35924 17444 38894
rect 17724 39060 17780 39070
rect 17724 38946 17780 39004
rect 17724 38894 17726 38946
rect 17778 38894 17780 38946
rect 17724 38882 17780 38894
rect 17948 38946 18004 39788
rect 17948 38894 17950 38946
rect 18002 38894 18004 38946
rect 17948 38882 18004 38894
rect 18060 39394 18116 39406
rect 18060 39342 18062 39394
rect 18114 39342 18116 39394
rect 17500 38722 17556 38734
rect 17500 38670 17502 38722
rect 17554 38670 17556 38722
rect 17500 38668 17556 38670
rect 18060 38724 18116 39342
rect 17500 38612 17892 38668
rect 17724 38052 17780 38062
rect 17612 37828 17668 37838
rect 17500 37772 17612 37828
rect 17500 36482 17556 37772
rect 17612 37762 17668 37772
rect 17500 36430 17502 36482
rect 17554 36430 17556 36482
rect 17500 36418 17556 36430
rect 17612 37268 17668 37278
rect 17612 37154 17668 37212
rect 17612 37102 17614 37154
rect 17666 37102 17668 37154
rect 17612 36372 17668 37102
rect 17612 36306 17668 36316
rect 17388 35830 17444 35868
rect 17724 35698 17780 37996
rect 17836 37268 17892 38612
rect 18060 37828 18116 38668
rect 18060 37762 18116 37772
rect 18060 37268 18116 37278
rect 17836 37266 18116 37268
rect 17836 37214 18062 37266
rect 18114 37214 18116 37266
rect 17836 37212 18116 37214
rect 18060 37202 18116 37212
rect 17836 37044 17892 37054
rect 17836 36950 17892 36988
rect 18172 36484 18228 42140
rect 18284 41636 18340 43148
rect 18508 42980 18564 42990
rect 18508 42886 18564 42924
rect 18620 42866 18676 43260
rect 18732 42980 18788 43484
rect 18844 42980 18900 48300
rect 19180 48290 19236 48300
rect 19180 47236 19236 47246
rect 19180 47142 19236 47180
rect 19292 47012 19348 50372
rect 19516 49810 19572 50540
rect 19740 50594 19796 50876
rect 19964 50706 20020 51100
rect 19964 50654 19966 50706
rect 20018 50654 20020 50706
rect 19964 50642 20020 50654
rect 19740 50542 19742 50594
rect 19794 50542 19796 50594
rect 19740 50530 19796 50542
rect 20188 50596 20244 51326
rect 20188 50502 20244 50540
rect 20412 51378 20468 51390
rect 20412 51326 20414 51378
rect 20466 51326 20468 51378
rect 20412 50594 20468 51326
rect 20412 50542 20414 50594
rect 20466 50542 20468 50594
rect 19628 50484 19684 50494
rect 20412 50428 20468 50542
rect 19628 50036 19684 50428
rect 20300 50372 20468 50428
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19628 49980 20020 50036
rect 19516 49758 19518 49810
rect 19570 49758 19572 49810
rect 19404 49700 19460 49710
rect 19404 49606 19460 49644
rect 19516 48468 19572 49758
rect 19852 49812 19908 49822
rect 19852 49718 19908 49756
rect 19628 49252 19684 49262
rect 19628 48468 19684 49196
rect 19964 49138 20020 49980
rect 19964 49086 19966 49138
rect 20018 49086 20020 49138
rect 19964 49074 20020 49086
rect 20300 49812 20356 50372
rect 20188 48916 20244 48926
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19964 48468 20020 48478
rect 19628 48466 20020 48468
rect 19628 48414 19966 48466
rect 20018 48414 20020 48466
rect 19628 48412 20020 48414
rect 19516 48374 19572 48412
rect 19964 48402 20020 48412
rect 20188 48466 20244 48860
rect 20300 48914 20356 49756
rect 20524 49588 20580 49598
rect 20524 49494 20580 49532
rect 20636 49140 20692 51884
rect 20748 50484 20804 50494
rect 20748 49922 20804 50428
rect 21532 50428 21588 52220
rect 21868 51602 21924 52892
rect 22316 52836 22372 52846
rect 22204 52834 22372 52836
rect 22204 52782 22318 52834
rect 22370 52782 22372 52834
rect 22204 52780 22372 52782
rect 22204 52388 22260 52780
rect 22316 52770 22372 52780
rect 22428 52612 22484 54348
rect 22540 54338 22596 54348
rect 22540 53508 22596 53518
rect 22540 53414 22596 53452
rect 22204 52322 22260 52332
rect 22316 52556 22484 52612
rect 21868 51550 21870 51602
rect 21922 51550 21924 51602
rect 21868 51538 21924 51550
rect 22092 51380 22148 51390
rect 22092 51286 22148 51324
rect 21756 51268 21812 51278
rect 21756 51174 21812 51212
rect 21980 51044 22036 51054
rect 21532 50372 21812 50428
rect 20748 49870 20750 49922
rect 20802 49870 20804 49922
rect 20748 49858 20804 49870
rect 20860 49810 20916 49822
rect 20860 49758 20862 49810
rect 20914 49758 20916 49810
rect 20636 49084 20804 49140
rect 20300 48862 20302 48914
rect 20354 48862 20356 48914
rect 20300 48850 20356 48862
rect 20636 48914 20692 48926
rect 20636 48862 20638 48914
rect 20690 48862 20692 48914
rect 20636 48804 20692 48862
rect 20636 48738 20692 48748
rect 20188 48414 20190 48466
rect 20242 48414 20244 48466
rect 20188 48402 20244 48414
rect 20412 48468 20468 48478
rect 20636 48468 20692 48478
rect 20412 48354 20468 48412
rect 20412 48302 20414 48354
rect 20466 48302 20468 48354
rect 20412 48290 20468 48302
rect 20524 48412 20636 48468
rect 20524 48354 20580 48412
rect 20636 48402 20692 48412
rect 20524 48302 20526 48354
rect 20578 48302 20580 48354
rect 20524 48290 20580 48302
rect 19852 48242 19908 48254
rect 19852 48190 19854 48242
rect 19906 48190 19908 48242
rect 19180 46956 19348 47012
rect 19516 47236 19572 47246
rect 19068 45892 19124 45902
rect 19068 45332 19124 45836
rect 19068 45266 19124 45276
rect 18956 45220 19012 45230
rect 18956 45126 19012 45164
rect 19068 45106 19124 45118
rect 19068 45054 19070 45106
rect 19122 45054 19124 45106
rect 18956 44996 19012 45006
rect 18956 44882 19012 44940
rect 18956 44830 18958 44882
rect 19010 44830 19012 44882
rect 18956 44818 19012 44830
rect 19068 43540 19124 45054
rect 19180 44100 19236 46956
rect 19404 46674 19460 46686
rect 19404 46622 19406 46674
rect 19458 46622 19460 46674
rect 19404 46004 19460 46622
rect 19516 46562 19572 47180
rect 19628 47236 19684 47246
rect 19852 47236 19908 48190
rect 19964 48244 20020 48254
rect 19964 47684 20020 48188
rect 19964 47682 20580 47684
rect 19964 47630 19966 47682
rect 20018 47630 20580 47682
rect 19964 47628 20580 47630
rect 19964 47618 20020 47628
rect 19628 47234 19908 47236
rect 19628 47182 19630 47234
rect 19682 47182 19908 47234
rect 19628 47180 19908 47182
rect 20188 47458 20244 47470
rect 20188 47406 20190 47458
rect 20242 47406 20244 47458
rect 19628 46788 19684 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20076 46788 20132 46798
rect 19628 46732 20076 46788
rect 20076 46674 20132 46732
rect 20076 46622 20078 46674
rect 20130 46622 20132 46674
rect 20076 46610 20132 46622
rect 19516 46510 19518 46562
rect 19570 46510 19572 46562
rect 19516 46498 19572 46510
rect 19404 45444 19460 45948
rect 20188 45890 20244 47406
rect 20524 47402 20580 47628
rect 20524 47350 20526 47402
rect 20578 47350 20580 47402
rect 20524 47338 20580 47350
rect 20636 47234 20692 47246
rect 20636 47182 20638 47234
rect 20690 47182 20692 47234
rect 20636 47068 20692 47182
rect 20188 45838 20190 45890
rect 20242 45838 20244 45890
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19404 45378 19460 45388
rect 19516 45276 20132 45332
rect 19404 45218 19460 45230
rect 19404 45166 19406 45218
rect 19458 45166 19460 45218
rect 19404 44884 19460 45166
rect 19404 44818 19460 44828
rect 19516 44660 19572 45276
rect 19404 44604 19572 44660
rect 19740 45106 19796 45118
rect 19740 45054 19742 45106
rect 19794 45054 19796 45106
rect 19740 44660 19796 45054
rect 20076 45106 20132 45276
rect 20076 45054 20078 45106
rect 20130 45054 20132 45106
rect 20076 45042 20132 45054
rect 19292 44324 19348 44334
rect 19292 44230 19348 44268
rect 19180 44044 19348 44100
rect 19068 43538 19236 43540
rect 19068 43486 19070 43538
rect 19122 43486 19236 43538
rect 19068 43484 19236 43486
rect 19068 43474 19124 43484
rect 19068 43204 19124 43214
rect 18844 42924 19012 42980
rect 18732 42914 18788 42924
rect 18620 42814 18622 42866
rect 18674 42814 18676 42866
rect 18620 42802 18676 42814
rect 18956 42644 19012 42924
rect 18844 42588 19012 42644
rect 18732 42532 18788 42542
rect 18396 42308 18452 42318
rect 18396 42082 18452 42252
rect 18732 42084 18788 42476
rect 18396 42030 18398 42082
rect 18450 42030 18452 42082
rect 18396 41972 18452 42030
rect 18396 41906 18452 41916
rect 18508 42028 18788 42084
rect 18284 41570 18340 41580
rect 18284 41412 18340 41422
rect 18284 41318 18340 41356
rect 18284 41186 18340 41198
rect 18284 41134 18286 41186
rect 18338 41134 18340 41186
rect 18284 40964 18340 41134
rect 18284 40898 18340 40908
rect 18508 40740 18564 42028
rect 18844 41970 18900 42588
rect 18844 41918 18846 41970
rect 18898 41918 18900 41970
rect 18844 41860 18900 41918
rect 18620 41804 18844 41860
rect 18620 41410 18676 41804
rect 18844 41794 18900 41804
rect 18956 41858 19012 41870
rect 18956 41806 18958 41858
rect 19010 41806 19012 41858
rect 18956 41636 19012 41806
rect 18956 41570 19012 41580
rect 18620 41358 18622 41410
rect 18674 41358 18676 41410
rect 18620 41346 18676 41358
rect 18956 41076 19012 41086
rect 18956 40982 19012 41020
rect 18284 40684 18564 40740
rect 18284 39844 18340 40684
rect 18620 40628 18676 40638
rect 18508 40572 18620 40628
rect 18508 40514 18564 40572
rect 18620 40562 18676 40572
rect 18508 40462 18510 40514
rect 18562 40462 18564 40514
rect 18508 40450 18564 40462
rect 18284 39778 18340 39788
rect 18396 39732 18452 39742
rect 18284 38948 18340 38958
rect 18284 38724 18340 38892
rect 18284 38658 18340 38668
rect 18396 38668 18452 39676
rect 19068 39730 19124 43148
rect 19180 42978 19236 43484
rect 19292 43428 19348 44044
rect 19292 43362 19348 43372
rect 19180 42926 19182 42978
rect 19234 42926 19236 42978
rect 19180 42914 19236 42926
rect 19292 42644 19348 42654
rect 19180 42642 19348 42644
rect 19180 42590 19294 42642
rect 19346 42590 19348 42642
rect 19180 42588 19348 42590
rect 19180 42084 19236 42588
rect 19292 42578 19348 42588
rect 19404 42308 19460 44604
rect 19740 44594 19796 44604
rect 19516 44436 19572 44446
rect 19516 44322 19572 44380
rect 19516 44270 19518 44322
rect 19570 44270 19572 44322
rect 19516 43652 19572 44270
rect 19516 43586 19572 43596
rect 19628 44322 19684 44334
rect 19628 44270 19630 44322
rect 19682 44270 19684 44322
rect 19628 43540 19684 44270
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19852 43540 19908 43550
rect 19628 43538 19908 43540
rect 19628 43486 19854 43538
rect 19906 43486 19908 43538
rect 19628 43484 19908 43486
rect 19516 43428 19572 43438
rect 19516 43334 19572 43372
rect 19852 42532 19908 43484
rect 20188 43204 20244 45838
rect 20300 47012 20692 47068
rect 20300 45892 20356 47012
rect 20748 46900 20804 49084
rect 20860 48468 20916 49758
rect 21084 49586 21140 49598
rect 21084 49534 21086 49586
rect 21138 49534 21140 49586
rect 20860 48402 20916 48412
rect 20972 49028 21028 49038
rect 21084 49028 21140 49534
rect 21644 49140 21700 49150
rect 21308 49028 21364 49038
rect 21532 49028 21588 49038
rect 21084 49026 21364 49028
rect 21084 48974 21310 49026
rect 21362 48974 21364 49026
rect 21084 48972 21364 48974
rect 20972 48466 21028 48972
rect 21308 48916 21364 48972
rect 21308 48850 21364 48860
rect 21420 49026 21588 49028
rect 21420 48974 21534 49026
rect 21586 48974 21588 49026
rect 21420 48972 21588 48974
rect 20972 48414 20974 48466
rect 21026 48414 21028 48466
rect 20972 48402 21028 48414
rect 21420 48804 21476 48972
rect 21532 48962 21588 48972
rect 21308 48132 21364 48142
rect 20300 45106 20356 45836
rect 20300 45054 20302 45106
rect 20354 45054 20356 45106
rect 20300 45042 20356 45054
rect 20636 46844 20804 46900
rect 20860 47234 20916 47246
rect 20860 47182 20862 47234
rect 20914 47182 20916 47234
rect 20636 44996 20692 46844
rect 20748 46674 20804 46686
rect 20748 46622 20750 46674
rect 20802 46622 20804 46674
rect 20748 45892 20804 46622
rect 20748 45798 20804 45836
rect 20636 44930 20692 44940
rect 20748 45668 20804 45678
rect 20524 44882 20580 44894
rect 20524 44830 20526 44882
rect 20578 44830 20580 44882
rect 20412 44772 20468 44782
rect 20412 44322 20468 44716
rect 20412 44270 20414 44322
rect 20466 44270 20468 44322
rect 20412 44258 20468 44270
rect 20524 44660 20580 44830
rect 20748 44884 20804 45612
rect 20860 45444 20916 47182
rect 21196 46676 21252 46686
rect 21196 46582 21252 46620
rect 20860 45378 20916 45388
rect 20972 45108 21028 45118
rect 21196 45108 21252 45118
rect 20972 45106 21252 45108
rect 20972 45054 20974 45106
rect 21026 45054 21198 45106
rect 21250 45054 21252 45106
rect 20972 45052 21252 45054
rect 20972 45042 21028 45052
rect 21196 45042 21252 45052
rect 20748 44828 21252 44884
rect 20524 44100 20580 44604
rect 20748 44100 20804 44110
rect 20524 44098 20804 44100
rect 20524 44046 20750 44098
rect 20802 44046 20804 44098
rect 20524 44044 20804 44046
rect 20300 43876 20356 43886
rect 20356 43820 20468 43876
rect 20300 43810 20356 43820
rect 20188 43138 20244 43148
rect 19852 42466 19908 42476
rect 20188 42980 20244 42990
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19404 42242 19460 42252
rect 20188 42196 20244 42924
rect 20076 42140 20244 42196
rect 19740 42084 19796 42094
rect 19180 42018 19236 42028
rect 19292 42082 19796 42084
rect 19292 42030 19742 42082
rect 19794 42030 19796 42082
rect 19292 42028 19796 42030
rect 19292 41410 19348 42028
rect 19740 42018 19796 42028
rect 19964 41972 20020 41982
rect 19852 41970 20020 41972
rect 19852 41918 19966 41970
rect 20018 41918 20020 41970
rect 19852 41916 20020 41918
rect 19292 41358 19294 41410
rect 19346 41358 19348 41410
rect 19292 41346 19348 41358
rect 19404 41860 19460 41870
rect 19404 41412 19460 41804
rect 19404 41346 19460 41356
rect 19852 41300 19908 41916
rect 19964 41906 20020 41916
rect 20076 41858 20132 42140
rect 20300 41972 20356 41982
rect 20076 41806 20078 41858
rect 20130 41806 20132 41858
rect 20076 41794 20132 41806
rect 20188 41916 20300 41972
rect 19964 41412 20020 41422
rect 20188 41412 20244 41916
rect 20300 41878 20356 41916
rect 20412 41748 20468 43820
rect 20748 43092 20804 44044
rect 20860 43652 20916 43662
rect 21196 43652 21252 44828
rect 20916 43596 21140 43652
rect 20860 43558 20916 43596
rect 20748 43036 21028 43092
rect 20748 42196 20804 42206
rect 20748 42102 20804 42140
rect 19964 41410 20244 41412
rect 19964 41358 19966 41410
rect 20018 41358 20244 41410
rect 19964 41356 20244 41358
rect 20300 41692 20468 41748
rect 20636 42084 20692 42094
rect 19964 41346 20020 41356
rect 19516 41244 19908 41300
rect 19180 40964 19236 40974
rect 19180 40870 19236 40908
rect 19068 39678 19070 39730
rect 19122 39678 19124 39730
rect 19068 39620 19124 39678
rect 19292 40402 19348 40414
rect 19292 40350 19294 40402
rect 19346 40350 19348 40402
rect 19292 39732 19348 40350
rect 19404 40292 19460 40302
rect 19404 40198 19460 40236
rect 19292 39666 19348 39676
rect 19068 39554 19124 39564
rect 19404 39618 19460 39630
rect 19404 39566 19406 39618
rect 19458 39566 19460 39618
rect 19404 39508 19460 39566
rect 18844 38948 18900 38958
rect 18844 38854 18900 38892
rect 18396 38612 18564 38668
rect 18508 38388 18564 38612
rect 18284 38332 18564 38388
rect 18732 38612 18788 38622
rect 18284 37266 18340 38332
rect 18732 38162 18788 38556
rect 18732 38110 18734 38162
rect 18786 38110 18788 38162
rect 18732 38098 18788 38110
rect 18620 37940 18676 37950
rect 18620 37846 18676 37884
rect 19180 37938 19236 37950
rect 19180 37886 19182 37938
rect 19234 37886 19236 37938
rect 19068 37268 19124 37278
rect 18284 37214 18286 37266
rect 18338 37214 18340 37266
rect 18284 37202 18340 37214
rect 18620 37266 19124 37268
rect 18620 37214 19070 37266
rect 19122 37214 19124 37266
rect 18620 37212 19124 37214
rect 18620 36484 18676 37212
rect 19068 37202 19124 37212
rect 18732 37044 18788 37054
rect 19180 37044 19236 37886
rect 19292 37826 19348 37838
rect 19292 37774 19294 37826
rect 19346 37774 19348 37826
rect 19292 37268 19348 37774
rect 19404 37380 19460 39452
rect 19516 39394 19572 41244
rect 19964 41188 20020 41198
rect 19964 41186 20244 41188
rect 19964 41134 19966 41186
rect 20018 41134 20244 41186
rect 19964 41132 20244 41134
rect 19964 41122 20020 41132
rect 19628 41074 19684 41086
rect 19628 41022 19630 41074
rect 19682 41022 19684 41074
rect 19628 40852 19684 41022
rect 20188 41076 20244 41132
rect 19628 40786 19684 40796
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19964 40404 20020 40414
rect 19964 40310 20020 40348
rect 19628 40180 19684 40190
rect 19628 40086 19684 40124
rect 19852 40178 19908 40190
rect 19852 40126 19854 40178
rect 19906 40126 19908 40178
rect 19852 40068 19908 40126
rect 20188 40068 20244 41020
rect 19852 40012 20244 40068
rect 19516 39342 19518 39394
rect 19570 39342 19572 39394
rect 19516 38834 19572 39342
rect 19516 38782 19518 38834
rect 19570 38782 19572 38834
rect 19516 38770 19572 38782
rect 19628 39620 19684 39630
rect 19516 37826 19572 37838
rect 19516 37774 19518 37826
rect 19570 37774 19572 37826
rect 19516 37604 19572 37774
rect 19516 37538 19572 37548
rect 19628 37492 19684 39564
rect 19964 39508 20020 39518
rect 19964 39414 20020 39452
rect 20076 39396 20132 39434
rect 20076 39330 20132 39340
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19852 38948 19908 38958
rect 19852 38854 19908 38892
rect 20188 38724 20244 40012
rect 20300 39060 20356 41692
rect 20412 41186 20468 41198
rect 20412 41134 20414 41186
rect 20466 41134 20468 41186
rect 20412 41076 20468 41134
rect 20412 41010 20468 41020
rect 20636 41074 20692 42028
rect 20860 41746 20916 41758
rect 20860 41694 20862 41746
rect 20914 41694 20916 41746
rect 20636 41022 20638 41074
rect 20690 41022 20692 41074
rect 20636 41010 20692 41022
rect 20748 41412 20804 41422
rect 20748 40740 20804 41356
rect 20748 40674 20804 40684
rect 20860 40628 20916 41694
rect 20860 40562 20916 40572
rect 20972 40404 21028 43036
rect 20972 40338 21028 40348
rect 20860 40068 20916 40078
rect 20748 39620 20804 39630
rect 20636 39564 20748 39620
rect 20636 39172 20692 39564
rect 20748 39554 20804 39564
rect 20748 39396 20804 39406
rect 20860 39396 20916 40012
rect 20748 39394 20916 39396
rect 20748 39342 20750 39394
rect 20802 39342 20916 39394
rect 20748 39340 20916 39342
rect 20748 39330 20804 39340
rect 20860 39172 20916 39340
rect 20636 39116 20804 39172
rect 20300 39004 20692 39060
rect 20412 38724 20468 38734
rect 20188 38668 20412 38724
rect 20412 38658 20468 38668
rect 20524 38610 20580 38622
rect 20524 38558 20526 38610
rect 20578 38558 20580 38610
rect 19852 38052 19908 38062
rect 19852 37958 19908 37996
rect 19740 37828 19796 37838
rect 20300 37828 20356 37838
rect 19740 37826 20244 37828
rect 19740 37774 19742 37826
rect 19794 37774 20244 37826
rect 19740 37772 20244 37774
rect 19740 37762 19796 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37436 19908 37492
rect 19404 37324 19684 37380
rect 19292 37202 19348 37212
rect 18732 37042 18900 37044
rect 18732 36990 18734 37042
rect 18786 36990 18900 37042
rect 18732 36988 18900 36990
rect 18732 36978 18788 36988
rect 18172 36428 18452 36484
rect 18284 36260 18340 36270
rect 18284 36166 18340 36204
rect 18284 35924 18340 35934
rect 17724 35646 17726 35698
rect 17778 35646 17780 35698
rect 17724 35634 17780 35646
rect 17948 35868 18284 35924
rect 17948 35698 18004 35868
rect 18284 35830 18340 35868
rect 17948 35646 17950 35698
rect 18002 35646 18004 35698
rect 17948 35634 18004 35646
rect 16828 35186 16884 35196
rect 16492 34804 16548 34814
rect 16492 34710 16548 34748
rect 17500 34804 17556 34814
rect 15372 34300 15596 34356
rect 15596 34262 15652 34300
rect 15708 34354 16100 34356
rect 15708 34302 15934 34354
rect 15986 34302 16100 34354
rect 15708 34300 16100 34302
rect 17388 34356 17444 34366
rect 15260 34066 15316 34076
rect 14140 34018 14196 34030
rect 14140 33966 14142 34018
rect 14194 33966 14196 34018
rect 14140 33460 14196 33966
rect 14252 33908 14308 33918
rect 14252 33906 14420 33908
rect 14252 33854 14254 33906
rect 14306 33854 14420 33906
rect 14252 33852 14420 33854
rect 14252 33842 14308 33852
rect 14364 33572 14420 33852
rect 14364 33506 14420 33516
rect 14252 33460 14308 33470
rect 14140 33458 14308 33460
rect 14140 33406 14254 33458
rect 14306 33406 14308 33458
rect 14140 33404 14308 33406
rect 14252 33394 14308 33404
rect 15708 33348 15764 34300
rect 15932 34290 15988 34300
rect 17388 34242 17444 34300
rect 17500 34354 17556 34748
rect 17500 34302 17502 34354
rect 17554 34302 17556 34354
rect 17500 34290 17556 34302
rect 17724 34692 17780 34702
rect 17388 34190 17390 34242
rect 17442 34190 17444 34242
rect 17388 34178 17444 34190
rect 17724 34242 17780 34636
rect 17724 34190 17726 34242
rect 17778 34190 17780 34242
rect 17724 34178 17780 34190
rect 16380 34132 16436 34142
rect 16380 34038 16436 34076
rect 17948 34132 18004 34142
rect 17948 34038 18004 34076
rect 16940 34018 16996 34030
rect 16940 33966 16942 34018
rect 16994 33966 16996 34018
rect 16940 33796 16996 33966
rect 17164 34020 17220 34030
rect 18396 34020 18452 36428
rect 18508 36482 18676 36484
rect 18508 36430 18622 36482
rect 18674 36430 18676 36482
rect 18508 36428 18676 36430
rect 18508 35028 18564 36428
rect 18620 36418 18676 36428
rect 18620 35700 18676 35710
rect 18620 35698 18788 35700
rect 18620 35646 18622 35698
rect 18674 35646 18788 35698
rect 18620 35644 18788 35646
rect 18620 35634 18676 35644
rect 18732 35588 18788 35644
rect 18620 35028 18676 35038
rect 18508 35026 18676 35028
rect 18508 34974 18622 35026
rect 18674 34974 18676 35026
rect 18508 34972 18676 34974
rect 18620 34962 18676 34972
rect 18508 34020 18564 34030
rect 18396 33964 18508 34020
rect 16996 33740 17108 33796
rect 16940 33730 16996 33740
rect 15596 32788 15652 32798
rect 15708 32788 15764 33292
rect 16380 33458 16436 33470
rect 16380 33406 16382 33458
rect 16434 33406 16436 33458
rect 16380 32788 16436 33406
rect 16940 33460 16996 33470
rect 16940 33366 16996 33404
rect 15596 32786 15764 32788
rect 15596 32734 15598 32786
rect 15650 32734 15764 32786
rect 15596 32732 15764 32734
rect 16044 32732 16436 32788
rect 16716 33348 16772 33358
rect 15596 32722 15652 32732
rect 15148 32450 15204 32462
rect 15148 32398 15150 32450
rect 15202 32398 15204 32450
rect 15148 31892 15204 32398
rect 16044 32452 16100 32732
rect 15148 31826 15204 31836
rect 15596 32004 15652 32014
rect 15596 31890 15652 31948
rect 15596 31838 15598 31890
rect 15650 31838 15652 31890
rect 15596 31826 15652 31838
rect 15708 31666 15764 31678
rect 15708 31614 15710 31666
rect 15762 31614 15764 31666
rect 14252 31556 14308 31566
rect 13804 31554 14420 31556
rect 13804 31502 14254 31554
rect 14306 31502 14420 31554
rect 13804 31500 14420 31502
rect 14252 31490 14308 31500
rect 14028 31220 14084 31230
rect 13468 31218 14084 31220
rect 13468 31166 13470 31218
rect 13522 31166 14030 31218
rect 14082 31166 14084 31218
rect 13468 31164 14084 31166
rect 13468 31154 13524 31164
rect 14028 31154 14084 31164
rect 13244 31054 13246 31106
rect 13298 31054 13300 31106
rect 13244 31042 13300 31054
rect 10332 30884 10388 30894
rect 9884 30882 10388 30884
rect 9884 30830 10334 30882
rect 10386 30830 10388 30882
rect 9884 30828 10388 30830
rect 9884 30098 9940 30828
rect 10332 30818 10388 30828
rect 12460 30882 12516 30894
rect 12460 30830 12462 30882
rect 12514 30830 12516 30882
rect 9884 30046 9886 30098
rect 9938 30046 9940 30098
rect 9884 30034 9940 30046
rect 10332 30100 10388 30110
rect 9772 29922 9828 29932
rect 10332 29650 10388 30044
rect 10332 29598 10334 29650
rect 10386 29598 10388 29650
rect 10332 29586 10388 29598
rect 11228 29540 11284 29550
rect 9212 28590 9214 28642
rect 9266 28590 9268 28642
rect 7644 26852 7700 26862
rect 7644 24724 7700 26796
rect 7980 26404 8036 26414
rect 7756 26402 8036 26404
rect 7756 26350 7982 26402
rect 8034 26350 8036 26402
rect 7756 26348 8036 26350
rect 7756 26066 7812 26348
rect 7980 26338 8036 26348
rect 8204 26180 8260 27132
rect 9212 26908 9268 28590
rect 10668 29202 10724 29214
rect 10668 29150 10670 29202
rect 10722 29150 10724 29202
rect 9884 28532 9940 28542
rect 9772 28530 9940 28532
rect 9772 28478 9886 28530
rect 9938 28478 9940 28530
rect 9772 28476 9940 28478
rect 9772 28082 9828 28476
rect 9884 28466 9940 28476
rect 9772 28030 9774 28082
rect 9826 28030 9828 28082
rect 9772 28018 9828 28030
rect 10108 27860 10164 27870
rect 10556 27860 10612 27870
rect 10108 27858 10612 27860
rect 10108 27806 10110 27858
rect 10162 27806 10558 27858
rect 10610 27806 10612 27858
rect 10108 27804 10612 27806
rect 10108 27794 10164 27804
rect 10556 27794 10612 27804
rect 10668 27748 10724 29150
rect 11228 29092 11284 29484
rect 12460 29540 12516 30830
rect 12460 29474 12516 29484
rect 12908 30882 12964 30894
rect 12908 30830 12910 30882
rect 12962 30830 12964 30882
rect 11452 29428 11508 29438
rect 10668 27682 10724 27692
rect 11116 29036 11284 29092
rect 11340 29372 11452 29428
rect 10892 27634 10948 27646
rect 10892 27582 10894 27634
rect 10946 27582 10948 27634
rect 10892 26908 10948 27582
rect 11116 26908 11172 29036
rect 11340 27858 11396 29372
rect 11452 29334 11508 29372
rect 12908 29428 12964 30830
rect 13580 30770 13636 30782
rect 13580 30718 13582 30770
rect 13634 30718 13636 30770
rect 13580 30548 13636 30718
rect 13580 30482 13636 30492
rect 13916 30770 13972 30782
rect 13916 30718 13918 30770
rect 13970 30718 13972 30770
rect 13468 30210 13524 30222
rect 13468 30158 13470 30210
rect 13522 30158 13524 30210
rect 13468 29428 13524 30158
rect 13916 29988 13972 30718
rect 14252 30772 14308 30782
rect 14252 30678 14308 30716
rect 14364 30660 14420 31500
rect 15484 31554 15540 31566
rect 15484 31502 15486 31554
rect 15538 31502 15540 31554
rect 15484 31220 15540 31502
rect 15708 31332 15764 31614
rect 15708 31266 15764 31276
rect 15484 31154 15540 31164
rect 16044 30996 16100 32396
rect 16268 32562 16324 32574
rect 16268 32510 16270 32562
rect 16322 32510 16324 32562
rect 16268 32340 16324 32510
rect 16268 32274 16324 32284
rect 16380 32562 16436 32574
rect 16380 32510 16382 32562
rect 16434 32510 16436 32562
rect 16268 32004 16324 32014
rect 16156 31778 16212 31790
rect 16156 31726 16158 31778
rect 16210 31726 16212 31778
rect 16156 31332 16212 31726
rect 16156 31266 16212 31276
rect 16156 30996 16212 31006
rect 16044 30994 16212 30996
rect 16044 30942 16158 30994
rect 16210 30942 16212 30994
rect 16044 30940 16212 30942
rect 16156 30930 16212 30940
rect 16268 30884 16324 31948
rect 16380 31892 16436 32510
rect 16604 32562 16660 32574
rect 16604 32510 16606 32562
rect 16658 32510 16660 32562
rect 16380 31108 16436 31836
rect 16492 32450 16548 32462
rect 16492 32398 16494 32450
rect 16546 32398 16548 32450
rect 16492 31668 16548 32398
rect 16604 32228 16660 32510
rect 16604 32162 16660 32172
rect 16492 31602 16548 31612
rect 16604 31778 16660 31790
rect 16604 31726 16606 31778
rect 16658 31726 16660 31778
rect 16604 31220 16660 31726
rect 16604 31154 16660 31164
rect 16380 31042 16436 31052
rect 16380 30884 16436 30894
rect 16268 30882 16436 30884
rect 16268 30830 16382 30882
rect 16434 30830 16436 30882
rect 16268 30828 16436 30830
rect 16380 30818 16436 30828
rect 14364 30594 14420 30604
rect 14252 30548 14308 30558
rect 14252 30322 14308 30492
rect 16380 30324 16436 30334
rect 14252 30270 14254 30322
rect 14306 30270 14308 30322
rect 14252 30258 14308 30270
rect 16156 30322 16436 30324
rect 16156 30270 16382 30322
rect 16434 30270 16436 30322
rect 16156 30268 16436 30270
rect 13692 29932 13972 29988
rect 13692 29538 13748 29932
rect 13692 29486 13694 29538
rect 13746 29486 13748 29538
rect 13692 29474 13748 29486
rect 12908 29426 13468 29428
rect 12908 29374 12910 29426
rect 12962 29374 13468 29426
rect 12908 29372 13468 29374
rect 12012 28754 12068 28766
rect 12012 28702 12014 28754
rect 12066 28702 12068 28754
rect 11340 27806 11342 27858
rect 11394 27806 11396 27858
rect 11340 27794 11396 27806
rect 11452 27972 11508 27982
rect 12012 27972 12068 28702
rect 11452 27970 12068 27972
rect 11452 27918 11454 27970
rect 11506 27918 12068 27970
rect 11452 27916 12068 27918
rect 12460 28644 12516 28654
rect 12908 28644 12964 29372
rect 13468 29334 13524 29372
rect 15932 29428 15988 29438
rect 12460 28642 12964 28644
rect 12460 28590 12462 28642
rect 12514 28590 12964 28642
rect 12460 28588 12964 28590
rect 15820 29314 15876 29326
rect 15820 29262 15822 29314
rect 15874 29262 15876 29314
rect 11452 26908 11508 27916
rect 12460 26908 12516 28588
rect 13916 27748 13972 27758
rect 13468 26962 13524 26974
rect 13468 26910 13470 26962
rect 13522 26910 13524 26962
rect 13468 26908 13524 26910
rect 13804 26962 13860 26974
rect 13804 26910 13806 26962
rect 13858 26910 13860 26962
rect 13804 26908 13860 26910
rect 9212 26852 9604 26908
rect 8204 26114 8260 26124
rect 8316 26290 8372 26302
rect 8316 26238 8318 26290
rect 8370 26238 8372 26290
rect 7756 26014 7758 26066
rect 7810 26014 7812 26066
rect 7756 26002 7812 26014
rect 8316 25508 8372 26238
rect 9436 26180 9492 26190
rect 7756 25452 8372 25508
rect 9100 25618 9156 25630
rect 9100 25566 9102 25618
rect 9154 25566 9156 25618
rect 7756 24946 7812 25452
rect 8652 25172 8708 25182
rect 7756 24894 7758 24946
rect 7810 24894 7812 24946
rect 7756 24882 7812 24894
rect 8316 25060 8372 25070
rect 8092 24724 8148 24734
rect 7644 24722 8148 24724
rect 7644 24670 8094 24722
rect 8146 24670 8148 24722
rect 7644 24668 8148 24670
rect 8092 24658 8148 24668
rect 7644 23940 7700 23950
rect 7980 23940 8036 23950
rect 7532 23938 7700 23940
rect 7532 23886 7646 23938
rect 7698 23886 7700 23938
rect 7532 23884 7700 23886
rect 7644 23874 7700 23884
rect 7756 23884 7980 23940
rect 6972 21646 6974 21698
rect 7026 21646 7028 21698
rect 6972 21634 7028 21646
rect 7084 23716 7140 23726
rect 7084 20356 7140 23660
rect 7420 23714 7476 23726
rect 7420 23662 7422 23714
rect 7474 23662 7476 23714
rect 7308 23156 7364 23166
rect 7308 23062 7364 23100
rect 7308 22596 7364 22606
rect 7308 22502 7364 22540
rect 7420 22372 7476 23662
rect 7532 23266 7588 23278
rect 7532 23214 7534 23266
rect 7586 23214 7588 23266
rect 7532 23044 7588 23214
rect 7644 23268 7700 23278
rect 7756 23268 7812 23884
rect 7980 23846 8036 23884
rect 7868 23716 7924 23726
rect 7868 23622 7924 23660
rect 8316 23548 8372 25004
rect 8652 24722 8708 25116
rect 8652 24670 8654 24722
rect 8706 24670 8708 24722
rect 8652 24658 8708 24670
rect 8876 24836 8932 24846
rect 9100 24836 9156 25566
rect 9436 24948 9492 26124
rect 9548 25506 9604 26852
rect 10556 26852 10948 26908
rect 10556 26786 10612 26796
rect 10108 26402 10164 26414
rect 10108 26350 10110 26402
rect 10162 26350 10164 26402
rect 9884 26292 9940 26302
rect 9884 26198 9940 26236
rect 10108 25620 10164 26350
rect 10556 26292 10612 26302
rect 10556 26198 10612 26236
rect 10892 26290 10948 26852
rect 10892 26238 10894 26290
rect 10946 26238 10948 26290
rect 10220 25620 10276 25630
rect 10108 25618 10276 25620
rect 10108 25566 10222 25618
rect 10274 25566 10276 25618
rect 10108 25564 10276 25566
rect 10220 25554 10276 25564
rect 9548 25454 9550 25506
rect 9602 25454 9604 25506
rect 9548 25284 9604 25454
rect 9772 25284 9828 25294
rect 9548 25228 9772 25284
rect 9660 24948 9716 24958
rect 9436 24946 9716 24948
rect 9436 24894 9662 24946
rect 9714 24894 9716 24946
rect 9436 24892 9716 24894
rect 9660 24882 9716 24892
rect 8876 24834 9156 24836
rect 8876 24782 8878 24834
rect 8930 24782 9156 24834
rect 8876 24780 9156 24782
rect 8876 24052 8932 24780
rect 9548 24052 9604 24062
rect 8876 24050 9604 24052
rect 8876 23998 9550 24050
rect 9602 23998 9604 24050
rect 8876 23996 9604 23998
rect 9548 23986 9604 23996
rect 8540 23716 8596 23726
rect 8540 23622 8596 23660
rect 9660 23714 9716 23726
rect 9660 23662 9662 23714
rect 9714 23662 9716 23714
rect 7644 23266 7812 23268
rect 7644 23214 7646 23266
rect 7698 23214 7812 23266
rect 7644 23212 7812 23214
rect 8092 23492 8372 23548
rect 7644 23202 7700 23212
rect 7532 22978 7588 22988
rect 7980 22932 8036 22942
rect 7980 22838 8036 22876
rect 7420 22316 7700 22372
rect 7420 22146 7476 22158
rect 7420 22094 7422 22146
rect 7474 22094 7476 22146
rect 7420 22036 7476 22094
rect 7308 21980 7476 22036
rect 7532 22146 7588 22158
rect 7532 22094 7534 22146
rect 7586 22094 7588 22146
rect 7196 21586 7252 21598
rect 7196 21534 7198 21586
rect 7250 21534 7252 21586
rect 7196 20692 7252 21534
rect 7308 21588 7364 21980
rect 7420 21588 7476 21598
rect 7308 21586 7476 21588
rect 7308 21534 7422 21586
rect 7474 21534 7476 21586
rect 7308 21532 7476 21534
rect 7420 21522 7476 21532
rect 7420 20692 7476 20702
rect 7196 20636 7420 20692
rect 7420 20626 7476 20636
rect 6860 19954 6916 19964
rect 6972 20300 7140 20356
rect 6188 19842 6244 19852
rect 6300 19124 6356 19134
rect 6860 19124 6916 19134
rect 5740 19012 5796 19022
rect 5180 19010 5796 19012
rect 5180 18958 5742 19010
rect 5794 18958 5796 19010
rect 5180 18956 5796 18958
rect 4060 18386 4116 18396
rect 5516 18564 5572 18574
rect 5516 18338 5572 18508
rect 5516 18286 5518 18338
rect 5570 18286 5572 18338
rect 5516 18274 5572 18286
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4620 17780 4676 17790
rect 4620 17686 4676 17724
rect 5068 17444 5124 17454
rect 5628 17444 5684 18956
rect 5740 18946 5796 18956
rect 6300 18564 6356 19068
rect 6748 19122 6916 19124
rect 6748 19070 6862 19122
rect 6914 19070 6916 19122
rect 6748 19068 6916 19070
rect 6524 18564 6580 18574
rect 5964 18452 6020 18462
rect 5964 18358 6020 18396
rect 6300 18450 6356 18508
rect 6300 18398 6302 18450
rect 6354 18398 6356 18450
rect 6300 18386 6356 18398
rect 6412 18508 6524 18564
rect 5740 17892 5796 17902
rect 5740 17798 5796 17836
rect 6076 17892 6132 17902
rect 6076 17798 6132 17836
rect 5068 17442 5684 17444
rect 5068 17390 5070 17442
rect 5122 17390 5684 17442
rect 5068 17388 5684 17390
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4844 16100 4900 16110
rect 4060 15986 4116 15998
rect 4060 15934 4062 15986
rect 4114 15934 4116 15986
rect 3724 15876 3780 15886
rect 3500 15874 3780 15876
rect 3500 15822 3726 15874
rect 3778 15822 3780 15874
rect 3500 15820 3780 15822
rect 3500 15426 3556 15820
rect 3724 15810 3780 15820
rect 4060 15540 4116 15934
rect 4060 15474 4116 15484
rect 3500 15374 3502 15426
rect 3554 15374 3556 15426
rect 3500 15362 3556 15374
rect 2828 15316 2884 15326
rect 2716 15314 2884 15316
rect 2716 15262 2830 15314
rect 2882 15262 2884 15314
rect 2716 15260 2884 15262
rect 2828 15092 2884 15260
rect 2828 15026 2884 15036
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 2492 14644 2548 14654
rect 2380 14642 2548 14644
rect 2380 14590 2494 14642
rect 2546 14590 2548 14642
rect 2380 14588 2548 14590
rect 2492 14578 2548 14588
rect 4620 14644 4676 14654
rect 4844 14644 4900 16044
rect 4620 14642 4900 14644
rect 4620 14590 4622 14642
rect 4674 14590 4900 14642
rect 4620 14588 4900 14590
rect 5068 15092 5124 17388
rect 6300 17108 6356 17118
rect 6412 17108 6468 18508
rect 6524 18498 6580 18508
rect 6748 17892 6804 19068
rect 6860 19058 6916 19068
rect 6972 18676 7028 20300
rect 7084 20132 7140 20142
rect 7308 20132 7364 20142
rect 7532 20132 7588 22094
rect 7644 20802 7700 22316
rect 7756 21812 7812 21822
rect 7756 21718 7812 21756
rect 8092 21698 8148 23492
rect 9660 23380 9716 23662
rect 9548 23324 9716 23380
rect 8204 23266 8260 23278
rect 8204 23214 8206 23266
rect 8258 23214 8260 23266
rect 8204 21924 8260 23214
rect 8764 23044 8820 23054
rect 8316 22932 8372 22942
rect 8316 22930 8484 22932
rect 8316 22878 8318 22930
rect 8370 22878 8484 22930
rect 8316 22876 8484 22878
rect 8316 22866 8372 22876
rect 8316 21924 8372 21934
rect 8204 21868 8316 21924
rect 8316 21858 8372 21868
rect 8092 21646 8094 21698
rect 8146 21646 8148 21698
rect 8092 21634 8148 21646
rect 7756 21588 7812 21598
rect 7756 21494 7812 21532
rect 8204 21588 8260 21598
rect 8092 20916 8148 20926
rect 7644 20750 7646 20802
rect 7698 20750 7700 20802
rect 7644 20738 7700 20750
rect 7756 20914 8148 20916
rect 7756 20862 8094 20914
rect 8146 20862 8148 20914
rect 7756 20860 8148 20862
rect 7756 20468 7812 20860
rect 8092 20850 8148 20860
rect 8204 20802 8260 21532
rect 8204 20750 8206 20802
rect 8258 20750 8260 20802
rect 8204 20738 8260 20750
rect 8316 21586 8372 21598
rect 8316 21534 8318 21586
rect 8370 21534 8372 21586
rect 7084 20038 7140 20076
rect 7196 20076 7308 20132
rect 7364 20076 7588 20132
rect 7644 20412 7812 20468
rect 7868 20692 7924 20702
rect 7196 19908 7252 20076
rect 7308 20038 7364 20076
rect 7644 20020 7700 20412
rect 7084 19852 7252 19908
rect 7420 19964 7700 20020
rect 7420 19906 7476 19964
rect 7420 19854 7422 19906
rect 7474 19854 7476 19906
rect 7084 19122 7140 19852
rect 7420 19842 7476 19854
rect 7868 19908 7924 20636
rect 8092 20580 8148 20590
rect 8092 20486 8148 20524
rect 8204 20468 8260 20478
rect 7980 20132 8036 20142
rect 8204 20132 8260 20412
rect 7980 20130 8260 20132
rect 7980 20078 7982 20130
rect 8034 20078 8260 20130
rect 7980 20076 8260 20078
rect 7980 20066 8036 20076
rect 7868 19852 8036 19908
rect 7644 19794 7700 19806
rect 7644 19742 7646 19794
rect 7698 19742 7700 19794
rect 7196 19348 7252 19358
rect 7196 19346 7588 19348
rect 7196 19294 7198 19346
rect 7250 19294 7588 19346
rect 7196 19292 7588 19294
rect 7196 19282 7252 19292
rect 7084 19070 7086 19122
rect 7138 19070 7140 19122
rect 7084 19058 7140 19070
rect 7420 19012 7476 19022
rect 7196 19010 7476 19012
rect 7196 18958 7422 19010
rect 7474 18958 7476 19010
rect 7196 18956 7476 18958
rect 7196 18788 7252 18956
rect 7420 18946 7476 18956
rect 6972 18610 7028 18620
rect 7084 18732 7252 18788
rect 7532 18788 7588 19292
rect 7644 19122 7700 19742
rect 7980 19572 8036 19852
rect 8092 19794 8148 20076
rect 8092 19742 8094 19794
rect 8146 19742 8148 19794
rect 8092 19730 8148 19742
rect 8316 19572 8372 21534
rect 8428 21588 8484 22876
rect 8540 21588 8596 21598
rect 8428 21586 8596 21588
rect 8428 21534 8542 21586
rect 8594 21534 8596 21586
rect 8428 21532 8596 21534
rect 8540 21522 8596 21532
rect 8652 21588 8708 21598
rect 8652 21494 8708 21532
rect 8764 21252 8820 22988
rect 9212 21924 9268 21934
rect 8652 21196 8820 21252
rect 8876 21810 8932 21822
rect 8876 21758 8878 21810
rect 8930 21758 8932 21810
rect 8876 21252 8932 21758
rect 8652 20468 8708 21196
rect 8876 21186 8932 21196
rect 9100 21028 9156 21038
rect 9100 20934 9156 20972
rect 9100 20804 9156 20814
rect 9212 20804 9268 21868
rect 9100 20802 9268 20804
rect 9100 20750 9102 20802
rect 9154 20750 9268 20802
rect 9100 20748 9268 20750
rect 9324 21588 9380 21598
rect 8652 20402 8708 20412
rect 8764 20690 8820 20702
rect 8764 20638 8766 20690
rect 8818 20638 8820 20690
rect 8764 20356 8820 20638
rect 8764 20290 8820 20300
rect 7980 19516 8372 19572
rect 7644 19070 7646 19122
rect 7698 19070 7700 19122
rect 7644 19058 7700 19070
rect 7756 19122 7812 19134
rect 7756 19070 7758 19122
rect 7810 19070 7812 19122
rect 7756 18900 7812 19070
rect 7980 18900 8036 19516
rect 9100 19460 9156 20748
rect 8428 19404 9156 19460
rect 8428 19234 8484 19404
rect 9324 19348 9380 21532
rect 9548 20804 9604 23324
rect 9660 23156 9716 23166
rect 9772 23156 9828 25228
rect 10892 24948 10948 26238
rect 10892 24882 10948 24892
rect 11004 26852 11172 26908
rect 11228 26852 11508 26908
rect 12236 26852 12516 26908
rect 12908 26852 13524 26908
rect 13580 26852 13860 26908
rect 9660 23154 9828 23156
rect 9660 23102 9662 23154
rect 9714 23102 9828 23154
rect 9660 23100 9828 23102
rect 9660 23090 9716 23100
rect 10332 23042 10388 23054
rect 10332 22990 10334 23042
rect 10386 22990 10388 23042
rect 10332 22258 10388 22990
rect 10668 22372 10724 22382
rect 10892 22372 10948 22382
rect 10668 22370 10892 22372
rect 10668 22318 10670 22370
rect 10722 22318 10892 22370
rect 10668 22316 10892 22318
rect 10668 22306 10724 22316
rect 10892 22306 10948 22316
rect 10332 22206 10334 22258
rect 10386 22206 10388 22258
rect 10332 22194 10388 22206
rect 10556 21700 10612 21710
rect 10892 21700 10948 21738
rect 10556 21698 10892 21700
rect 10556 21646 10558 21698
rect 10610 21646 10892 21698
rect 10556 21644 10892 21646
rect 10556 21634 10612 21644
rect 10892 21634 10948 21644
rect 11004 21476 11060 26852
rect 11116 21700 11172 21710
rect 11228 21700 11284 26852
rect 11676 26402 11732 26414
rect 11676 26350 11678 26402
rect 11730 26350 11732 26402
rect 11452 26292 11508 26302
rect 11452 26198 11508 26236
rect 11676 25620 11732 26350
rect 11676 25554 11732 25564
rect 12236 26290 12292 26852
rect 12908 26402 12964 26852
rect 12908 26350 12910 26402
rect 12962 26350 12964 26402
rect 12908 26338 12964 26350
rect 12236 26238 12238 26290
rect 12290 26238 12292 26290
rect 12236 25284 12292 26238
rect 12572 26292 12628 26302
rect 12236 25218 12292 25228
rect 12348 25620 12404 25630
rect 11676 24948 11732 24958
rect 11676 24854 11732 24892
rect 12012 24722 12068 24734
rect 12012 24670 12014 24722
rect 12066 24670 12068 24722
rect 12012 24388 12068 24670
rect 12348 24500 12404 25564
rect 12572 25396 12628 26236
rect 13580 25730 13636 26852
rect 13580 25678 13582 25730
rect 13634 25678 13636 25730
rect 13580 25666 13636 25678
rect 13916 26516 13972 27692
rect 15484 27074 15540 27086
rect 15484 27022 15486 27074
rect 15538 27022 15540 27074
rect 13916 25730 13972 26460
rect 15148 26852 15204 26862
rect 15484 26852 15540 27022
rect 15820 26908 15876 29262
rect 15932 28642 15988 29372
rect 15932 28590 15934 28642
rect 15986 28590 15988 28642
rect 15932 28578 15988 28590
rect 16156 28644 16212 30268
rect 16380 30258 16436 30268
rect 16716 30212 16772 33292
rect 17052 33234 17108 33740
rect 17052 33182 17054 33234
rect 17106 33182 17108 33234
rect 17052 33170 17108 33182
rect 16828 33124 16884 33134
rect 16828 32562 16884 33068
rect 16828 32510 16830 32562
rect 16882 32510 16884 32562
rect 16828 31892 16884 32510
rect 16828 31826 16884 31836
rect 17052 31668 17108 31678
rect 17052 31574 17108 31612
rect 16828 31556 16884 31566
rect 16828 31106 16884 31500
rect 16828 31054 16830 31106
rect 16882 31054 16884 31106
rect 16828 31042 16884 31054
rect 16828 30212 16884 30222
rect 16492 30210 16884 30212
rect 16492 30158 16830 30210
rect 16882 30158 16884 30210
rect 16492 30156 16884 30158
rect 17164 30212 17220 33964
rect 18508 33926 18564 33964
rect 17276 33572 17332 33582
rect 17276 32788 17332 33516
rect 18396 33348 18452 33358
rect 18396 33346 18564 33348
rect 18396 33294 18398 33346
rect 18450 33294 18564 33346
rect 18396 33292 18564 33294
rect 18396 33282 18452 33292
rect 17724 33124 17780 33134
rect 17724 33030 17780 33068
rect 17836 33122 17892 33134
rect 17836 33070 17838 33122
rect 17890 33070 17892 33122
rect 17836 32788 17892 33070
rect 17948 33124 18004 33134
rect 17948 33122 18340 33124
rect 17948 33070 17950 33122
rect 18002 33070 18340 33122
rect 17948 33068 18340 33070
rect 17948 33058 18004 33068
rect 17836 32732 18004 32788
rect 17276 32722 17332 32732
rect 17500 32562 17556 32574
rect 17500 32510 17502 32562
rect 17554 32510 17556 32562
rect 17500 32340 17556 32510
rect 17612 32562 17668 32574
rect 17612 32510 17614 32562
rect 17666 32510 17668 32562
rect 17612 32452 17668 32510
rect 17724 32564 17780 32574
rect 17724 32470 17780 32508
rect 17836 32562 17892 32574
rect 17836 32510 17838 32562
rect 17890 32510 17892 32562
rect 17612 32386 17668 32396
rect 17500 32274 17556 32284
rect 17836 32228 17892 32510
rect 17836 32162 17892 32172
rect 17388 31778 17444 31790
rect 17388 31726 17390 31778
rect 17442 31726 17444 31778
rect 17388 31556 17444 31726
rect 17388 31490 17444 31500
rect 17388 31220 17444 31230
rect 17388 31126 17444 31164
rect 17500 31108 17556 31118
rect 17500 31014 17556 31052
rect 17948 30996 18004 32732
rect 18060 32562 18116 32574
rect 18060 32510 18062 32562
rect 18114 32510 18116 32562
rect 18060 31556 18116 32510
rect 18060 31490 18116 31500
rect 18172 31668 18228 31678
rect 17948 30930 18004 30940
rect 18172 30994 18228 31612
rect 18172 30942 18174 30994
rect 18226 30942 18228 30994
rect 18172 30930 18228 30942
rect 18284 31106 18340 33068
rect 18508 32786 18564 33292
rect 18508 32734 18510 32786
rect 18562 32734 18564 32786
rect 18508 32722 18564 32734
rect 18396 32562 18452 32574
rect 18396 32510 18398 32562
rect 18450 32510 18452 32562
rect 18396 32004 18452 32510
rect 18620 32562 18676 32574
rect 18620 32510 18622 32562
rect 18674 32510 18676 32562
rect 18620 32452 18676 32510
rect 18620 32386 18676 32396
rect 18396 31938 18452 31948
rect 18732 32002 18788 35532
rect 18844 34468 18900 36988
rect 19068 36988 19236 37044
rect 19404 37044 19460 37054
rect 19068 36932 19124 36988
rect 18956 36820 19012 36830
rect 18956 36706 19012 36764
rect 18956 36654 18958 36706
rect 19010 36654 19012 36706
rect 18956 36642 19012 36654
rect 19068 36594 19124 36876
rect 19404 36820 19460 36988
rect 19068 36542 19070 36594
rect 19122 36542 19124 36594
rect 19068 36530 19124 36542
rect 19292 36764 19460 36820
rect 19292 36482 19348 36764
rect 19628 36594 19684 37324
rect 19628 36542 19630 36594
rect 19682 36542 19684 36594
rect 19628 36530 19684 36542
rect 19852 36706 19908 37436
rect 19852 36654 19854 36706
rect 19906 36654 19908 36706
rect 19292 36430 19294 36482
rect 19346 36430 19348 36482
rect 19292 36418 19348 36430
rect 19516 36484 19572 36494
rect 19068 36372 19124 36382
rect 19068 35026 19124 36316
rect 19068 34974 19070 35026
rect 19122 34974 19124 35026
rect 19068 34962 19124 34974
rect 19516 34914 19572 36428
rect 19852 36260 19908 36654
rect 20076 37378 20132 37390
rect 20076 37326 20078 37378
rect 20130 37326 20132 37378
rect 20076 36708 20132 37326
rect 20076 36642 20132 36652
rect 20188 37268 20244 37772
rect 20300 37734 20356 37772
rect 20076 36484 20132 36494
rect 20076 36390 20132 36428
rect 19516 34862 19518 34914
rect 19570 34862 19572 34914
rect 19516 34850 19572 34862
rect 19628 36204 19908 36260
rect 18956 34692 19012 34702
rect 18956 34598 19012 34636
rect 18844 34412 19236 34468
rect 18844 34244 18900 34254
rect 18844 34150 18900 34188
rect 19180 33572 19236 34412
rect 19292 34020 19348 34030
rect 19628 34020 19684 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20076 35700 20132 35710
rect 20188 35700 20244 37212
rect 20300 36482 20356 36494
rect 20300 36430 20302 36482
rect 20354 36430 20356 36482
rect 20300 36260 20356 36430
rect 20300 36194 20356 36204
rect 20524 35810 20580 38558
rect 20524 35758 20526 35810
rect 20578 35758 20580 35810
rect 20524 35746 20580 35758
rect 20076 35698 20244 35700
rect 20076 35646 20078 35698
rect 20130 35646 20244 35698
rect 20076 35644 20244 35646
rect 20076 35634 20132 35644
rect 19740 35588 19796 35598
rect 19740 35494 19796 35532
rect 19964 34916 20020 34926
rect 19964 34822 20020 34860
rect 20636 34916 20692 39004
rect 20748 36706 20804 39116
rect 20860 39106 20916 39116
rect 20972 38948 21028 38958
rect 21084 38948 21140 43596
rect 21196 43586 21252 43596
rect 21308 43204 21364 48076
rect 21196 43148 21364 43204
rect 21196 41972 21252 43148
rect 21308 42980 21364 42990
rect 21420 42980 21476 48748
rect 21644 46676 21700 49084
rect 21644 46610 21700 46620
rect 21756 45556 21812 50372
rect 21868 49252 21924 49262
rect 21868 49158 21924 49196
rect 21756 45490 21812 45500
rect 21756 45218 21812 45230
rect 21756 45166 21758 45218
rect 21810 45166 21812 45218
rect 21756 45108 21812 45166
rect 21532 44322 21588 44334
rect 21532 44270 21534 44322
rect 21586 44270 21588 44322
rect 21532 43876 21588 44270
rect 21756 44100 21812 45052
rect 21756 44044 21924 44100
rect 21532 43810 21588 43820
rect 21756 43876 21812 43886
rect 21756 43762 21812 43820
rect 21756 43710 21758 43762
rect 21810 43710 21812 43762
rect 21756 43698 21812 43710
rect 21532 43652 21588 43662
rect 21532 43092 21588 43596
rect 21644 43540 21700 43550
rect 21644 43446 21700 43484
rect 21868 43428 21924 44044
rect 21532 43026 21588 43036
rect 21756 43372 21924 43428
rect 21364 42924 21476 42980
rect 21308 42914 21364 42924
rect 21756 42868 21812 43372
rect 21532 42812 21812 42868
rect 21308 42756 21364 42766
rect 21308 42308 21364 42700
rect 21308 42242 21364 42252
rect 21196 41906 21252 41916
rect 21196 40628 21252 40638
rect 21532 40628 21588 42812
rect 21868 42756 21924 42766
rect 21756 42700 21868 42756
rect 21644 42196 21700 42206
rect 21644 41970 21700 42140
rect 21644 41918 21646 41970
rect 21698 41918 21700 41970
rect 21644 41906 21700 41918
rect 21196 40626 21588 40628
rect 21196 40574 21198 40626
rect 21250 40574 21588 40626
rect 21196 40572 21588 40574
rect 21196 40562 21252 40572
rect 21420 40404 21476 40414
rect 21308 40402 21476 40404
rect 21308 40350 21422 40402
rect 21474 40350 21476 40402
rect 21308 40348 21476 40350
rect 21028 38892 21140 38948
rect 21196 39844 21252 39854
rect 20972 38882 21028 38892
rect 20972 38724 21028 38734
rect 20972 38612 21140 38668
rect 20860 38164 20916 38174
rect 20860 37266 20916 38108
rect 20860 37214 20862 37266
rect 20914 37214 20916 37266
rect 20860 37202 20916 37214
rect 20748 36654 20750 36706
rect 20802 36654 20804 36706
rect 20748 36642 20804 36654
rect 21084 36372 21140 38612
rect 21196 38164 21252 39788
rect 21308 39060 21364 40348
rect 21420 40338 21476 40348
rect 21532 40404 21588 40414
rect 21532 40310 21588 40348
rect 21644 40402 21700 40414
rect 21644 40350 21646 40402
rect 21698 40350 21700 40402
rect 21644 39844 21700 40350
rect 21532 39788 21700 39844
rect 21532 39732 21588 39788
rect 21756 39732 21812 42700
rect 21868 42662 21924 42700
rect 21980 42084 22036 50988
rect 22204 50484 22260 50522
rect 22204 50418 22260 50428
rect 22316 49028 22372 52556
rect 22764 52500 22820 56028
rect 22876 54740 22932 59200
rect 23212 56308 23268 56318
rect 23212 56214 23268 56252
rect 23324 55412 23380 59200
rect 24220 56642 24276 59200
rect 24220 56590 24222 56642
rect 24274 56590 24276 56642
rect 24220 56578 24276 56590
rect 24668 56308 24724 59200
rect 24668 56242 24724 56252
rect 25004 56642 25060 56654
rect 25004 56590 25006 56642
rect 25058 56590 25060 56642
rect 23996 56084 24052 56094
rect 23996 56082 24164 56084
rect 23996 56030 23998 56082
rect 24050 56030 24164 56082
rect 23996 56028 24164 56030
rect 23996 56018 24052 56028
rect 24108 55972 24164 56028
rect 24556 55972 24612 55982
rect 24108 55970 24612 55972
rect 24108 55918 24558 55970
rect 24610 55918 24612 55970
rect 24108 55916 24612 55918
rect 23324 55356 23940 55412
rect 23100 55186 23156 55198
rect 23100 55134 23102 55186
rect 23154 55134 23156 55186
rect 22988 54740 23044 54750
rect 22876 54738 23044 54740
rect 22876 54686 22990 54738
rect 23042 54686 23044 54738
rect 22876 54684 23044 54686
rect 22988 54674 23044 54684
rect 22988 53844 23044 53854
rect 23100 53844 23156 55134
rect 23884 54738 23940 55356
rect 23884 54686 23886 54738
rect 23938 54686 23940 54738
rect 23884 54674 23940 54686
rect 22988 53842 23156 53844
rect 22988 53790 22990 53842
rect 23042 53790 23156 53842
rect 22988 53788 23156 53790
rect 23660 54516 23716 54526
rect 22988 53778 23044 53788
rect 23660 53730 23716 54460
rect 23660 53678 23662 53730
rect 23714 53678 23716 53730
rect 23660 53666 23716 53678
rect 23100 53620 23156 53630
rect 23436 53620 23492 53630
rect 23100 53526 23156 53564
rect 23212 53618 23492 53620
rect 23212 53566 23438 53618
rect 23490 53566 23492 53618
rect 23212 53564 23492 53566
rect 22876 53508 22932 53518
rect 22876 53414 22932 53452
rect 22764 52444 22932 52500
rect 22764 52276 22820 52286
rect 22764 52182 22820 52220
rect 22652 52164 22708 52174
rect 22540 52108 22652 52164
rect 22540 51602 22596 52108
rect 22652 52098 22708 52108
rect 22876 51716 22932 52444
rect 22876 51650 22932 51660
rect 22540 51550 22542 51602
rect 22594 51550 22596 51602
rect 22540 51538 22596 51550
rect 22652 51490 22708 51502
rect 22652 51438 22654 51490
rect 22706 51438 22708 51490
rect 22652 51380 22708 51438
rect 22540 51324 22652 51380
rect 22428 51156 22484 51166
rect 22428 51062 22484 51100
rect 22540 50932 22596 51324
rect 22652 51314 22708 51324
rect 23100 51380 23156 51390
rect 23100 51044 23156 51324
rect 23100 50978 23156 50988
rect 22428 50876 22596 50932
rect 22428 50484 22484 50876
rect 22540 50708 22596 50718
rect 22540 50706 23044 50708
rect 22540 50654 22542 50706
rect 22594 50654 23044 50706
rect 22540 50652 23044 50654
rect 22540 50642 22596 50652
rect 22988 50596 23044 50652
rect 23100 50596 23156 50606
rect 22988 50594 23156 50596
rect 22988 50542 23102 50594
rect 23154 50542 23156 50594
rect 22988 50540 23156 50542
rect 23100 50530 23156 50540
rect 22428 50370 22484 50428
rect 22876 50482 22932 50494
rect 22876 50430 22878 50482
rect 22930 50430 22932 50482
rect 22876 50428 22932 50430
rect 22876 50372 23044 50428
rect 22428 50318 22430 50370
rect 22482 50318 22484 50370
rect 22428 50306 22484 50318
rect 22876 49812 22932 49822
rect 22764 49810 22932 49812
rect 22764 49758 22878 49810
rect 22930 49758 22932 49810
rect 22764 49756 22932 49758
rect 22764 49138 22820 49756
rect 22876 49746 22932 49756
rect 22988 49252 23044 50372
rect 23212 50034 23268 53564
rect 23436 53554 23492 53564
rect 23772 53620 23828 53630
rect 23996 53620 24052 53630
rect 23772 53506 23828 53564
rect 23772 53454 23774 53506
rect 23826 53454 23828 53506
rect 23772 53442 23828 53454
rect 23884 53618 24052 53620
rect 23884 53566 23998 53618
rect 24050 53566 24052 53618
rect 23884 53564 24052 53566
rect 23884 53172 23940 53564
rect 23996 53554 24052 53564
rect 24108 53396 24164 55916
rect 24556 55906 24612 55916
rect 24668 55524 24724 55534
rect 24556 54516 24612 54526
rect 24556 54422 24612 54460
rect 24668 53954 24724 55468
rect 24668 53902 24670 53954
rect 24722 53902 24724 53954
rect 24668 53890 24724 53902
rect 24668 53730 24724 53742
rect 24668 53678 24670 53730
rect 24722 53678 24724 53730
rect 24332 53620 24388 53630
rect 23548 52948 23604 52958
rect 23772 52948 23828 52958
rect 23548 52854 23604 52892
rect 23660 52946 23828 52948
rect 23660 52894 23774 52946
rect 23826 52894 23828 52946
rect 23660 52892 23828 52894
rect 23324 52276 23380 52286
rect 23324 52162 23380 52220
rect 23324 52110 23326 52162
rect 23378 52110 23380 52162
rect 23324 52098 23380 52110
rect 23548 51940 23604 51950
rect 23436 51492 23492 51502
rect 23548 51492 23604 51884
rect 23436 51490 23604 51492
rect 23436 51438 23438 51490
rect 23490 51438 23604 51490
rect 23436 51436 23604 51438
rect 23436 51426 23492 51436
rect 23548 50706 23604 51436
rect 23548 50654 23550 50706
rect 23602 50654 23604 50706
rect 23548 50642 23604 50654
rect 23324 50596 23380 50606
rect 23324 50502 23380 50540
rect 23436 50484 23492 50494
rect 23660 50428 23716 52892
rect 23772 52882 23828 52892
rect 23884 51940 23940 53116
rect 23996 53340 24164 53396
rect 24220 53618 24388 53620
rect 24220 53566 24334 53618
rect 24386 53566 24388 53618
rect 24220 53564 24388 53566
rect 23996 53058 24052 53340
rect 24108 53172 24164 53182
rect 24108 53078 24164 53116
rect 23996 53006 23998 53058
rect 24050 53006 24052 53058
rect 23996 52994 24052 53006
rect 24108 52836 24164 52846
rect 24220 52836 24276 53564
rect 24332 53554 24388 53564
rect 24668 53508 24724 53678
rect 25004 53618 25060 56590
rect 25228 55410 25284 55422
rect 25228 55358 25230 55410
rect 25282 55358 25284 55410
rect 25228 54516 25284 55358
rect 25564 54738 25620 59200
rect 26012 56644 26068 59200
rect 26012 56588 26404 56644
rect 25788 55300 25844 55310
rect 25788 55206 25844 55244
rect 25564 54686 25566 54738
rect 25618 54686 25620 54738
rect 25564 54674 25620 54686
rect 26348 54740 26404 56588
rect 26684 55970 26740 55982
rect 26684 55918 26686 55970
rect 26738 55918 26740 55970
rect 26684 55524 26740 55918
rect 26684 55458 26740 55468
rect 26908 55468 26964 59200
rect 27356 57428 27412 59200
rect 27356 57372 28084 57428
rect 27356 56082 27412 56094
rect 27356 56030 27358 56082
rect 27410 56030 27412 56082
rect 26908 55412 27188 55468
rect 26460 55188 26516 55198
rect 26460 55186 26852 55188
rect 26460 55134 26462 55186
rect 26514 55134 26852 55186
rect 26460 55132 26852 55134
rect 26460 55122 26516 55132
rect 26460 54740 26516 54750
rect 26348 54738 26516 54740
rect 26348 54686 26462 54738
rect 26514 54686 26516 54738
rect 26348 54684 26516 54686
rect 26460 54674 26516 54684
rect 25228 54450 25284 54460
rect 25004 53566 25006 53618
rect 25058 53566 25060 53618
rect 25004 53554 25060 53566
rect 24668 53442 24724 53452
rect 25676 53508 25732 53518
rect 24108 52834 24276 52836
rect 24108 52782 24110 52834
rect 24162 52782 24276 52834
rect 24108 52780 24276 52782
rect 25452 53058 25508 53070
rect 25452 53006 25454 53058
rect 25506 53006 25508 53058
rect 25452 52948 25508 53006
rect 25676 52948 25732 53452
rect 26012 52948 26068 52958
rect 25452 52946 26068 52948
rect 25452 52894 26014 52946
rect 26066 52894 26068 52946
rect 25452 52892 26068 52894
rect 24108 52770 24164 52780
rect 24444 52724 24500 52734
rect 24332 52500 24388 52510
rect 23996 52164 24052 52174
rect 23996 52070 24052 52108
rect 24332 52052 24388 52444
rect 24444 52274 24500 52668
rect 25228 52724 25284 52734
rect 25228 52630 25284 52668
rect 25228 52500 25284 52510
rect 24444 52222 24446 52274
rect 24498 52222 24500 52274
rect 24444 52210 24500 52222
rect 24668 52276 24724 52286
rect 24444 52052 24500 52062
rect 24332 52050 24500 52052
rect 24332 51998 24446 52050
rect 24498 51998 24500 52050
rect 24332 51996 24500 51998
rect 24444 51986 24500 51996
rect 23884 51874 23940 51884
rect 24220 51938 24276 51950
rect 24220 51886 24222 51938
rect 24274 51886 24276 51938
rect 23772 51492 23828 51502
rect 23772 51398 23828 51436
rect 23996 51380 24052 51390
rect 23996 51286 24052 51324
rect 24108 51156 24164 51166
rect 23772 51100 24108 51156
rect 23772 50594 23828 51100
rect 24108 51090 24164 51100
rect 24108 50932 24164 50942
rect 24108 50706 24164 50876
rect 24108 50654 24110 50706
rect 24162 50654 24164 50706
rect 24108 50642 24164 50654
rect 23772 50542 23774 50594
rect 23826 50542 23828 50594
rect 23772 50530 23828 50542
rect 23884 50484 23940 50494
rect 23436 50372 23604 50428
rect 23660 50372 23828 50428
rect 23212 49982 23214 50034
rect 23266 49982 23268 50034
rect 23212 49970 23268 49982
rect 22764 49086 22766 49138
rect 22818 49086 22820 49138
rect 22764 49074 22820 49086
rect 22876 49196 23044 49252
rect 23212 49812 23268 49822
rect 23212 49252 23268 49756
rect 23548 49810 23604 50372
rect 23548 49758 23550 49810
rect 23602 49758 23604 49810
rect 23548 49746 23604 49758
rect 23324 49700 23380 49710
rect 23324 49606 23380 49644
rect 22316 48972 22708 49028
rect 22540 48802 22596 48814
rect 22540 48750 22542 48802
rect 22594 48750 22596 48802
rect 22540 48356 22596 48750
rect 22204 48300 22540 48356
rect 22092 47348 22148 47358
rect 22092 47254 22148 47292
rect 22204 47124 22260 48300
rect 22540 48262 22596 48300
rect 22652 48244 22708 48972
rect 22764 48916 22820 48926
rect 22764 48822 22820 48860
rect 22876 48468 22932 49196
rect 23100 49026 23156 49038
rect 23100 48974 23102 49026
rect 23154 48974 23156 49026
rect 23100 48804 23156 48974
rect 23212 49026 23268 49196
rect 23772 49138 23828 50372
rect 23884 50370 23940 50428
rect 23884 50318 23886 50370
rect 23938 50318 23940 50370
rect 23884 50306 23940 50318
rect 24108 50036 24164 50046
rect 24220 50036 24276 51886
rect 24556 51940 24612 51978
rect 24556 51874 24612 51884
rect 24556 51716 24612 51726
rect 24556 51490 24612 51660
rect 24556 51438 24558 51490
rect 24610 51438 24612 51490
rect 24444 51156 24500 51166
rect 24444 51062 24500 51100
rect 24556 50932 24612 51438
rect 24556 50866 24612 50876
rect 24108 50034 24276 50036
rect 24108 49982 24110 50034
rect 24162 49982 24276 50034
rect 24108 49980 24276 49982
rect 24332 50596 24388 50606
rect 24108 49970 24164 49980
rect 23996 49812 24052 49822
rect 23772 49086 23774 49138
rect 23826 49086 23828 49138
rect 23772 49074 23828 49086
rect 23884 49810 24052 49812
rect 23884 49758 23998 49810
rect 24050 49758 24052 49810
rect 23884 49756 24052 49758
rect 23212 48974 23214 49026
rect 23266 48974 23268 49026
rect 23212 48962 23268 48974
rect 23324 49028 23380 49038
rect 23100 48738 23156 48748
rect 22988 48468 23044 48478
rect 22876 48466 23044 48468
rect 22876 48414 22990 48466
rect 23042 48414 23044 48466
rect 22876 48412 23044 48414
rect 22988 48402 23044 48412
rect 23212 48468 23268 48478
rect 23324 48468 23380 48972
rect 23884 49028 23940 49756
rect 23996 49746 24052 49756
rect 24220 49810 24276 49822
rect 24220 49758 24222 49810
rect 24274 49758 24276 49810
rect 23884 48934 23940 48972
rect 23996 48916 24052 48926
rect 24220 48916 24276 49758
rect 24332 49252 24388 50540
rect 24668 50428 24724 52220
rect 25228 52274 25284 52444
rect 25228 52222 25230 52274
rect 25282 52222 25284 52274
rect 25228 52210 25284 52222
rect 25452 50428 25508 52892
rect 26012 52882 26068 52892
rect 25564 52724 25620 52734
rect 25564 52630 25620 52668
rect 26796 52164 26852 55132
rect 27132 53618 27188 55412
rect 27356 55300 27412 56030
rect 27412 55244 27748 55300
rect 27356 55234 27412 55244
rect 27692 54740 27748 55244
rect 27692 54738 27972 54740
rect 27692 54686 27694 54738
rect 27746 54686 27972 54738
rect 27692 54684 27972 54686
rect 27692 54674 27748 54684
rect 27132 53566 27134 53618
rect 27186 53566 27188 53618
rect 27132 53554 27188 53566
rect 27244 54514 27300 54526
rect 27244 54462 27246 54514
rect 27298 54462 27300 54514
rect 27244 52500 27300 54462
rect 27916 52948 27972 54684
rect 28028 54738 28084 57372
rect 28028 54686 28030 54738
rect 28082 54686 28084 54738
rect 28028 54674 28084 54686
rect 28252 54740 28308 59200
rect 28700 56642 28756 59200
rect 28700 56590 28702 56642
rect 28754 56590 28756 56642
rect 28700 56578 28756 56590
rect 29372 56642 29428 56654
rect 29372 56590 29374 56642
rect 29426 56590 29428 56642
rect 28700 56082 28756 56094
rect 28700 56030 28702 56082
rect 28754 56030 28756 56082
rect 28700 55468 28756 56030
rect 29372 55970 29428 56590
rect 29596 56420 29652 59200
rect 29596 56364 29876 56420
rect 29372 55918 29374 55970
rect 29426 55918 29428 55970
rect 29372 55906 29428 55918
rect 28588 55412 28756 55468
rect 28588 55410 28644 55412
rect 28588 55358 28590 55410
rect 28642 55358 28644 55410
rect 28588 55346 28644 55358
rect 29148 55300 29204 55310
rect 29148 55206 29204 55244
rect 28252 54674 28308 54684
rect 29148 54740 29204 54750
rect 29148 54646 29204 54684
rect 29820 54738 29876 56364
rect 30044 56308 30100 59200
rect 30044 56242 30100 56252
rect 30716 56308 30772 56318
rect 30716 56214 30772 56252
rect 30492 55970 30548 55982
rect 30492 55918 30494 55970
rect 30546 55918 30548 55970
rect 30492 55468 30548 55918
rect 30380 55412 30548 55468
rect 30940 55468 30996 59200
rect 31388 56308 31444 59200
rect 31388 56242 31444 56252
rect 31388 56082 31444 56094
rect 31388 56030 31390 56082
rect 31442 56030 31444 56082
rect 31388 55468 31444 56030
rect 32172 56082 32228 56094
rect 32172 56030 32174 56082
rect 32226 56030 32228 56082
rect 32172 55468 32228 56030
rect 30940 55412 31220 55468
rect 30380 55300 30436 55412
rect 29932 55188 29988 55198
rect 29932 55186 30324 55188
rect 29932 55134 29934 55186
rect 29986 55134 30324 55186
rect 29932 55132 30324 55134
rect 29932 55122 29988 55132
rect 29820 54686 29822 54738
rect 29874 54686 29876 54738
rect 29820 54674 29876 54686
rect 28812 54516 28868 54526
rect 28812 54514 28980 54516
rect 28812 54462 28814 54514
rect 28866 54462 28980 54514
rect 28812 54460 28980 54462
rect 28812 54450 28868 54460
rect 28812 53620 28868 53630
rect 28812 53058 28868 53564
rect 28924 53508 28980 54460
rect 29260 53508 29316 53518
rect 28924 53506 29316 53508
rect 28924 53454 29262 53506
rect 29314 53454 29316 53506
rect 28924 53452 29316 53454
rect 30268 53508 30324 55132
rect 30380 53732 30436 55244
rect 31164 54738 31220 55412
rect 31164 54686 31166 54738
rect 31218 54686 31220 54738
rect 31164 54674 31220 54686
rect 31276 55412 31444 55468
rect 32060 55412 32228 55468
rect 32284 55468 32340 59200
rect 32732 57092 32788 59200
rect 32732 57026 32788 57036
rect 32620 56308 32676 56318
rect 32620 55970 32676 56252
rect 33628 56308 33684 59200
rect 34076 56980 34132 59200
rect 34076 56914 34132 56924
rect 34188 57092 34244 57102
rect 33628 56242 33684 56252
rect 32620 55918 32622 55970
rect 32674 55918 32676 55970
rect 32620 55906 32676 55918
rect 33740 56082 33796 56094
rect 33740 56030 33742 56082
rect 33794 56030 33796 56082
rect 33740 55468 33796 56030
rect 34188 55970 34244 57036
rect 34188 55918 34190 55970
rect 34242 55918 34244 55970
rect 34188 55906 34244 55918
rect 32284 55412 32452 55468
rect 31276 54180 31332 55412
rect 32060 55410 32116 55412
rect 32060 55358 32062 55410
rect 32114 55358 32116 55410
rect 32060 55346 32116 55358
rect 32396 55186 32452 55412
rect 33404 55412 33796 55468
rect 34076 55860 34132 55870
rect 32396 55134 32398 55186
rect 32450 55134 32452 55186
rect 32396 55122 32452 55134
rect 32956 55298 33012 55310
rect 32956 55246 32958 55298
rect 33010 55246 33012 55298
rect 31052 54124 31332 54180
rect 32284 54402 32340 54414
rect 32284 54350 32286 54402
rect 32338 54350 32340 54402
rect 30436 53676 30548 53732
rect 30380 53666 30436 53676
rect 30380 53508 30436 53518
rect 30268 53506 30436 53508
rect 30268 53454 30382 53506
rect 30434 53454 30436 53506
rect 30268 53452 30436 53454
rect 28812 53006 28814 53058
rect 28866 53006 28868 53058
rect 28812 52994 28868 53006
rect 28028 52948 28084 52958
rect 27916 52946 28084 52948
rect 27916 52894 28030 52946
rect 28082 52894 28084 52946
rect 27916 52892 28084 52894
rect 27244 52434 27300 52444
rect 27356 52724 27412 52734
rect 27356 52274 27412 52668
rect 27356 52222 27358 52274
rect 27410 52222 27412 52274
rect 27356 52210 27412 52222
rect 28028 52276 28084 52892
rect 28588 52276 28644 52286
rect 28028 52274 29204 52276
rect 28028 52222 28590 52274
rect 28642 52222 29204 52274
rect 28028 52220 29204 52222
rect 28028 52164 28084 52220
rect 28588 52210 28644 52220
rect 26796 52108 26964 52164
rect 26908 51156 26964 52108
rect 26908 51090 26964 51100
rect 27468 52162 28084 52164
rect 27468 52110 28030 52162
rect 28082 52110 28084 52162
rect 27468 52108 28084 52110
rect 27468 50708 27524 52108
rect 28028 52098 28084 52108
rect 27020 50706 27524 50708
rect 27020 50654 27470 50706
rect 27522 50654 27524 50706
rect 27020 50652 27524 50654
rect 27020 50594 27076 50652
rect 27020 50542 27022 50594
rect 27074 50542 27076 50594
rect 27020 50530 27076 50542
rect 24332 49138 24388 49196
rect 24332 49086 24334 49138
rect 24386 49086 24388 49138
rect 24332 49074 24388 49086
rect 24444 50372 24724 50428
rect 25228 50372 25508 50428
rect 26236 50484 26292 50522
rect 26236 50418 26292 50428
rect 24052 48860 24276 48916
rect 23212 48466 23380 48468
rect 23212 48414 23214 48466
rect 23266 48414 23380 48466
rect 23212 48412 23380 48414
rect 23660 48804 23716 48814
rect 23212 48402 23268 48412
rect 23436 48356 23492 48366
rect 23436 48262 23492 48300
rect 22652 48188 22820 48244
rect 22428 48132 22484 48142
rect 22428 48038 22484 48076
rect 22652 48020 22708 48030
rect 22652 47926 22708 47964
rect 22316 47908 22372 47918
rect 22316 47458 22372 47852
rect 22316 47406 22318 47458
rect 22370 47406 22372 47458
rect 22316 47394 22372 47406
rect 22652 47460 22708 47470
rect 22652 47366 22708 47404
rect 22316 47236 22372 47246
rect 22764 47236 22820 48188
rect 23548 48242 23604 48254
rect 23548 48190 23550 48242
rect 23602 48190 23604 48242
rect 23548 48020 23604 48190
rect 22316 47234 22596 47236
rect 22316 47182 22318 47234
rect 22370 47182 22596 47234
rect 22316 47180 22596 47182
rect 22316 47170 22372 47180
rect 22092 47068 22260 47124
rect 22540 47068 22596 47180
rect 22092 45780 22148 47068
rect 22428 47012 22596 47068
rect 22652 47180 22820 47236
rect 23324 47348 23380 47358
rect 22316 46676 22372 46686
rect 22316 46582 22372 46620
rect 22204 46340 22260 46350
rect 22204 46002 22260 46284
rect 22428 46228 22484 47012
rect 22540 46788 22596 46798
rect 22540 46694 22596 46732
rect 22428 46162 22484 46172
rect 22540 46562 22596 46574
rect 22540 46510 22542 46562
rect 22594 46510 22596 46562
rect 22204 45950 22206 46002
rect 22258 45950 22260 46002
rect 22204 45938 22260 45950
rect 22428 46004 22484 46014
rect 22428 45890 22484 45948
rect 22428 45838 22430 45890
rect 22482 45838 22484 45890
rect 22428 45826 22484 45838
rect 22092 45724 22260 45780
rect 22092 45444 22148 45454
rect 22092 44436 22148 45388
rect 22092 44322 22148 44380
rect 22092 44270 22094 44322
rect 22146 44270 22148 44322
rect 22092 44258 22148 44270
rect 21980 42018 22036 42028
rect 22092 43428 22148 43438
rect 22092 41972 22148 43372
rect 22204 42194 22260 45724
rect 22540 45556 22596 46510
rect 22428 45500 22596 45556
rect 22316 44660 22372 44670
rect 22316 42756 22372 44604
rect 22316 42690 22372 42700
rect 22428 42644 22484 45500
rect 22540 44324 22596 44334
rect 22652 44324 22708 47180
rect 23212 46674 23268 46686
rect 23212 46622 23214 46674
rect 23266 46622 23268 46674
rect 22988 46562 23044 46574
rect 22988 46510 22990 46562
rect 23042 46510 23044 46562
rect 22988 45332 23044 46510
rect 23212 46340 23268 46622
rect 23212 46274 23268 46284
rect 22988 45266 23044 45276
rect 23100 46228 23156 46238
rect 22764 45218 22820 45230
rect 22764 45166 22766 45218
rect 22818 45166 22820 45218
rect 22764 44660 22820 45166
rect 22764 44594 22820 44604
rect 23100 44546 23156 46172
rect 23324 46116 23380 47292
rect 23548 47124 23604 47964
rect 23548 47058 23604 47068
rect 23100 44494 23102 44546
rect 23154 44494 23156 44546
rect 23100 44482 23156 44494
rect 23212 46060 23380 46116
rect 23212 44548 23268 46060
rect 23436 46004 23492 46014
rect 23324 44548 23380 44558
rect 23212 44546 23380 44548
rect 23212 44494 23326 44546
rect 23378 44494 23380 44546
rect 23212 44492 23380 44494
rect 23324 44482 23380 44492
rect 22540 44322 22708 44324
rect 22540 44270 22542 44322
rect 22594 44270 22708 44322
rect 22540 44268 22708 44270
rect 22540 43204 22596 44268
rect 22764 44100 22820 44110
rect 22764 44098 23044 44100
rect 22764 44046 22766 44098
rect 22818 44046 23044 44098
rect 22764 44044 23044 44046
rect 22764 44034 22820 44044
rect 22540 43138 22596 43148
rect 22876 43540 22932 43550
rect 22876 42754 22932 43484
rect 22988 43316 23044 44044
rect 23100 43652 23156 43662
rect 23100 43558 23156 43596
rect 23436 43538 23492 45948
rect 23548 45892 23604 45902
rect 23548 45798 23604 45836
rect 23548 44436 23604 44446
rect 23548 44342 23604 44380
rect 23436 43486 23438 43538
rect 23490 43486 23492 43538
rect 23436 43474 23492 43486
rect 23548 43652 23604 43662
rect 23324 43428 23380 43438
rect 23100 43316 23156 43326
rect 22988 43260 23100 43316
rect 22988 42980 23044 42990
rect 22988 42866 23044 42924
rect 22988 42814 22990 42866
rect 23042 42814 23044 42866
rect 22988 42802 23044 42814
rect 22876 42702 22878 42754
rect 22930 42702 22932 42754
rect 22876 42690 22932 42702
rect 23100 42754 23156 43260
rect 23100 42702 23102 42754
rect 23154 42702 23156 42754
rect 23100 42690 23156 42702
rect 23212 43204 23268 43214
rect 22428 42578 22484 42588
rect 22764 42644 22820 42654
rect 22204 42142 22206 42194
rect 22258 42142 22260 42194
rect 22204 42130 22260 42142
rect 22652 42530 22708 42542
rect 22652 42478 22654 42530
rect 22706 42478 22708 42530
rect 22652 42196 22708 42478
rect 22764 42196 22820 42588
rect 22988 42196 23044 42206
rect 22764 42194 23044 42196
rect 22764 42142 22990 42194
rect 23042 42142 23044 42194
rect 22764 42140 23044 42142
rect 22652 42130 22708 42140
rect 22092 41906 22148 41916
rect 22428 41970 22484 41982
rect 22764 41972 22820 41982
rect 22428 41918 22430 41970
rect 22482 41918 22484 41970
rect 21868 41746 21924 41758
rect 21868 41694 21870 41746
rect 21922 41694 21924 41746
rect 21868 40964 21924 41694
rect 22092 41524 22148 41534
rect 22092 41410 22148 41468
rect 22092 41358 22094 41410
rect 22146 41358 22148 41410
rect 22092 41346 22148 41358
rect 22204 41412 22260 41422
rect 22428 41412 22484 41918
rect 22260 41356 22484 41412
rect 22540 41970 22820 41972
rect 22540 41918 22766 41970
rect 22818 41918 22820 41970
rect 22540 41916 22820 41918
rect 22092 41188 22148 41198
rect 22092 41074 22148 41132
rect 22092 41022 22094 41074
rect 22146 41022 22148 41074
rect 22092 41010 22148 41022
rect 22204 41074 22260 41356
rect 22204 41022 22206 41074
rect 22258 41022 22260 41074
rect 21868 40898 21924 40908
rect 21980 40852 22036 40862
rect 21532 39666 21588 39676
rect 21644 39730 21812 39732
rect 21644 39678 21758 39730
rect 21810 39678 21812 39730
rect 21644 39676 21812 39678
rect 21308 38994 21364 39004
rect 21420 39508 21476 39518
rect 21420 38834 21476 39452
rect 21532 39506 21588 39518
rect 21532 39454 21534 39506
rect 21586 39454 21588 39506
rect 21532 39172 21588 39454
rect 21532 39106 21588 39116
rect 21420 38782 21422 38834
rect 21474 38782 21476 38834
rect 21308 38164 21364 38174
rect 21196 38162 21364 38164
rect 21196 38110 21310 38162
rect 21362 38110 21364 38162
rect 21196 38108 21364 38110
rect 21308 38098 21364 38108
rect 21420 37490 21476 38782
rect 21420 37438 21422 37490
rect 21474 37438 21476 37490
rect 21420 37426 21476 37438
rect 21532 36484 21588 36494
rect 21532 36390 21588 36428
rect 21308 36372 21364 36382
rect 21084 36370 21476 36372
rect 21084 36318 21310 36370
rect 21362 36318 21476 36370
rect 21084 36316 21476 36318
rect 21308 36306 21364 36316
rect 21420 36260 21476 36316
rect 21420 36204 21588 36260
rect 21420 35924 21476 35934
rect 21308 35922 21476 35924
rect 21308 35870 21422 35922
rect 21474 35870 21476 35922
rect 21308 35868 21476 35870
rect 20188 34802 20244 34814
rect 20188 34750 20190 34802
rect 20242 34750 20244 34802
rect 19852 34692 19908 34730
rect 19852 34626 19908 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19292 34018 19684 34020
rect 19292 33966 19294 34018
rect 19346 33966 19684 34018
rect 19292 33964 19684 33966
rect 20188 34132 20244 34750
rect 19292 33954 19348 33964
rect 18956 33348 19012 33358
rect 18956 33254 19012 33292
rect 19180 32788 19236 33516
rect 19628 33348 19684 33358
rect 19628 32900 19684 33292
rect 20188 33122 20244 34076
rect 20412 33684 20468 33694
rect 20468 33628 20580 33684
rect 20412 33618 20468 33628
rect 20188 33070 20190 33122
rect 20242 33070 20244 33122
rect 19516 32844 19628 32900
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19292 32788 19348 32798
rect 19180 32786 19348 32788
rect 19180 32734 19294 32786
rect 19346 32734 19348 32786
rect 19180 32732 19348 32734
rect 19292 32722 19348 32732
rect 18732 31950 18734 32002
rect 18786 31950 18788 32002
rect 18732 31938 18788 31950
rect 18844 32674 18900 32686
rect 18844 32622 18846 32674
rect 18898 32622 18900 32674
rect 18844 31780 18900 32622
rect 19516 32004 19572 32844
rect 19628 32834 19684 32844
rect 20076 32788 20132 32798
rect 19628 32676 19684 32686
rect 19628 32674 19796 32676
rect 19628 32622 19630 32674
rect 19682 32622 19796 32674
rect 19628 32620 19796 32622
rect 19628 32610 19684 32620
rect 19740 32340 19796 32620
rect 20076 32562 20132 32732
rect 20076 32510 20078 32562
rect 20130 32510 20132 32562
rect 20076 32498 20132 32510
rect 20188 32452 20244 33070
rect 20188 32386 20244 32396
rect 19740 32004 19796 32284
rect 19516 31948 19684 32004
rect 19516 31780 19572 31790
rect 18844 31686 18900 31724
rect 19292 31778 19572 31780
rect 19292 31726 19518 31778
rect 19570 31726 19572 31778
rect 19292 31724 19572 31726
rect 19180 31220 19236 31230
rect 19292 31220 19348 31724
rect 19516 31714 19572 31724
rect 19180 31218 19348 31220
rect 19180 31166 19182 31218
rect 19234 31166 19348 31218
rect 19180 31164 19348 31166
rect 19180 31154 19236 31164
rect 18284 31054 18286 31106
rect 18338 31054 18340 31106
rect 17500 30212 17556 30222
rect 17164 30210 17556 30212
rect 17164 30158 17502 30210
rect 17554 30158 17556 30210
rect 17164 30156 17556 30158
rect 16492 30100 16548 30156
rect 16268 30044 16548 30100
rect 16268 29650 16324 30044
rect 16268 29598 16270 29650
rect 16322 29598 16324 29650
rect 16268 29428 16324 29598
rect 16268 29362 16324 29372
rect 16156 28588 16548 28644
rect 16268 27972 16324 27982
rect 16044 27188 16100 27198
rect 15820 26852 15988 26908
rect 15148 26850 15540 26852
rect 15148 26798 15150 26850
rect 15202 26798 15540 26850
rect 15148 26796 15540 26798
rect 13916 25678 13918 25730
rect 13970 25678 13972 25730
rect 13916 25666 13972 25678
rect 15036 26178 15092 26190
rect 15036 26126 15038 26178
rect 15090 26126 15092 26178
rect 12012 24322 12068 24332
rect 12236 24444 12404 24500
rect 12460 24610 12516 24622
rect 12460 24558 12462 24610
rect 12514 24558 12516 24610
rect 11788 22596 11844 22606
rect 11676 22540 11788 22596
rect 11452 22372 11508 22382
rect 11452 22278 11508 22316
rect 11116 21698 11284 21700
rect 11116 21646 11118 21698
rect 11170 21646 11284 21698
rect 11116 21644 11284 21646
rect 11676 21698 11732 22540
rect 11788 22502 11844 22540
rect 11676 21646 11678 21698
rect 11730 21646 11732 21698
rect 11116 21634 11172 21644
rect 11676 21634 11732 21646
rect 12124 21700 12180 21710
rect 11004 21420 11284 21476
rect 10780 21362 10836 21374
rect 10780 21310 10782 21362
rect 10834 21310 10836 21362
rect 10108 21028 10164 21038
rect 10108 20934 10164 20972
rect 9660 20804 9716 20814
rect 9548 20802 9716 20804
rect 9548 20750 9662 20802
rect 9714 20750 9716 20802
rect 9548 20748 9716 20750
rect 9660 20738 9716 20748
rect 10220 20802 10276 20814
rect 10220 20750 10222 20802
rect 10274 20750 10276 20802
rect 8428 19182 8430 19234
rect 8482 19182 8484 19234
rect 8428 19170 8484 19182
rect 8876 19292 9380 19348
rect 9884 20690 9940 20702
rect 9884 20638 9886 20690
rect 9938 20638 9940 20690
rect 8092 19124 8148 19134
rect 8764 19124 8820 19134
rect 8876 19124 8932 19292
rect 9772 19234 9828 19246
rect 9772 19182 9774 19234
rect 9826 19182 9828 19234
rect 8092 19030 8148 19068
rect 8540 19122 8932 19124
rect 8540 19070 8766 19122
rect 8818 19070 8932 19122
rect 8540 19068 8932 19070
rect 9100 19124 9156 19134
rect 8204 19010 8260 19022
rect 8204 18958 8206 19010
rect 8258 18958 8260 19010
rect 7980 18844 8148 18900
rect 7756 18834 7812 18844
rect 6860 18562 6916 18574
rect 6860 18510 6862 18562
rect 6914 18510 6916 18562
rect 6860 18004 6916 18510
rect 7084 18452 7140 18732
rect 7532 18722 7588 18732
rect 7868 18788 7924 18798
rect 7924 18732 8036 18788
rect 7868 18722 7924 18732
rect 7308 18676 7364 18686
rect 6860 17938 6916 17948
rect 6972 18450 7140 18452
rect 6972 18398 7086 18450
rect 7138 18398 7140 18450
rect 6972 18396 7140 18398
rect 6748 17826 6804 17836
rect 6860 17668 6916 17678
rect 6972 17668 7028 18396
rect 7084 18386 7140 18396
rect 7196 18620 7308 18676
rect 6860 17666 7028 17668
rect 6860 17614 6862 17666
rect 6914 17614 7028 17666
rect 6860 17612 7028 17614
rect 6860 17602 6916 17612
rect 6300 17106 6468 17108
rect 6300 17054 6302 17106
rect 6354 17054 6468 17106
rect 6300 17052 6468 17054
rect 6748 17556 6804 17566
rect 6300 17042 6356 17052
rect 6412 16884 6468 16894
rect 6188 16772 6244 16782
rect 6076 16770 6244 16772
rect 6076 16718 6190 16770
rect 6242 16718 6244 16770
rect 6076 16716 6244 16718
rect 6076 16100 6132 16716
rect 6188 16706 6244 16716
rect 6076 16006 6132 16044
rect 5740 15876 5796 15886
rect 5740 15782 5796 15820
rect 6076 15540 6132 15550
rect 6076 15446 6132 15484
rect 6412 15316 6468 16828
rect 5628 15314 6468 15316
rect 5628 15262 6414 15314
rect 6466 15262 6468 15314
rect 5628 15260 6468 15262
rect 5628 15202 5684 15260
rect 6412 15250 6468 15260
rect 6748 15986 6804 17500
rect 7084 17108 7140 17118
rect 7196 17108 7252 18620
rect 7308 18610 7364 18620
rect 7532 18564 7588 18574
rect 7532 18470 7588 18508
rect 7756 18450 7812 18462
rect 7756 18398 7758 18450
rect 7810 18398 7812 18450
rect 7084 17106 7252 17108
rect 7084 17054 7086 17106
rect 7138 17054 7252 17106
rect 7084 17052 7252 17054
rect 7308 18004 7364 18014
rect 7084 17042 7140 17052
rect 7308 16996 7364 17948
rect 7756 17556 7812 18398
rect 7980 18450 8036 18732
rect 7980 18398 7982 18450
rect 8034 18398 8036 18450
rect 7980 18386 8036 18398
rect 8092 17556 8148 18844
rect 8204 18228 8260 18958
rect 8316 18788 8372 18798
rect 8316 18674 8372 18732
rect 8316 18622 8318 18674
rect 8370 18622 8372 18674
rect 8316 18610 8372 18622
rect 8316 18452 8372 18462
rect 8540 18452 8596 19068
rect 8764 19058 8820 19068
rect 9100 19030 9156 19068
rect 9772 19124 9828 19182
rect 9772 19058 9828 19068
rect 9548 18676 9604 18686
rect 8988 18564 9044 18574
rect 8988 18470 9044 18508
rect 9548 18562 9604 18620
rect 9548 18510 9550 18562
rect 9602 18510 9604 18562
rect 9548 18498 9604 18510
rect 9772 18564 9828 18574
rect 9884 18564 9940 20638
rect 10108 20578 10164 20590
rect 10108 20526 10110 20578
rect 10162 20526 10164 20578
rect 10108 19460 10164 20526
rect 10108 19394 10164 19404
rect 10220 20020 10276 20750
rect 10556 20690 10612 20702
rect 10556 20638 10558 20690
rect 10610 20638 10612 20690
rect 10556 20468 10612 20638
rect 10556 20412 10724 20468
rect 10668 20132 10724 20412
rect 10780 20244 10836 21310
rect 11004 20804 11060 20814
rect 10892 20802 11060 20804
rect 10892 20750 11006 20802
rect 11058 20750 11060 20802
rect 10892 20748 11060 20750
rect 10892 20690 10948 20748
rect 11004 20738 11060 20748
rect 10892 20638 10894 20690
rect 10946 20638 10948 20690
rect 10892 20626 10948 20638
rect 11228 20690 11284 21420
rect 12124 21140 12180 21644
rect 12236 21588 12292 24444
rect 12460 24388 12516 24558
rect 12460 24322 12516 24332
rect 12348 24164 12404 24174
rect 12572 24164 12628 25340
rect 14140 25396 14196 25406
rect 14140 25302 14196 25340
rect 14476 25396 14532 25406
rect 15036 25396 15092 26126
rect 15148 25508 15204 26796
rect 15372 26516 15428 26526
rect 15372 26422 15428 26460
rect 15708 26290 15764 26302
rect 15708 26238 15710 26290
rect 15762 26238 15764 26290
rect 15708 26068 15764 26238
rect 15708 26002 15764 26012
rect 15260 25508 15316 25518
rect 15148 25506 15316 25508
rect 15148 25454 15262 25506
rect 15314 25454 15316 25506
rect 15148 25452 15316 25454
rect 14476 25394 15092 25396
rect 14476 25342 14478 25394
rect 14530 25342 15092 25394
rect 14476 25340 15092 25342
rect 12796 25284 12852 25294
rect 12796 25190 12852 25228
rect 13916 25284 13972 25294
rect 12348 24162 12628 24164
rect 12348 24110 12350 24162
rect 12402 24110 12628 24162
rect 12348 24108 12628 24110
rect 12908 24948 12964 24958
rect 12348 24098 12404 24108
rect 12908 24050 12964 24892
rect 13580 24948 13636 24958
rect 13132 24612 13188 24622
rect 13132 24518 13188 24556
rect 13468 24612 13524 24622
rect 12908 23998 12910 24050
rect 12962 23998 12964 24050
rect 12684 23938 12740 23950
rect 12684 23886 12686 23938
rect 12738 23886 12740 23938
rect 12460 23042 12516 23054
rect 12460 22990 12462 23042
rect 12514 22990 12516 23042
rect 12460 22596 12516 22990
rect 12684 23044 12740 23886
rect 12908 23940 12964 23998
rect 12908 23874 12964 23884
rect 13244 24388 13300 24398
rect 13132 23044 13188 23054
rect 12684 23042 13188 23044
rect 12684 22990 13134 23042
rect 13186 22990 13188 23042
rect 12684 22988 13188 22990
rect 12460 22530 12516 22540
rect 13132 22596 13188 22988
rect 13132 22530 13188 22540
rect 12572 22370 12628 22382
rect 12572 22318 12574 22370
rect 12626 22318 12628 22370
rect 12460 22258 12516 22270
rect 12460 22206 12462 22258
rect 12514 22206 12516 22258
rect 12460 22148 12516 22206
rect 12572 22260 12628 22318
rect 13244 22260 13300 24332
rect 13468 23940 13524 24556
rect 12572 22194 12628 22204
rect 13132 22204 13300 22260
rect 13356 23938 13524 23940
rect 13356 23886 13470 23938
rect 13522 23886 13524 23938
rect 13356 23884 13524 23886
rect 12460 22082 12516 22092
rect 12348 21588 12404 21598
rect 12236 21586 12404 21588
rect 12236 21534 12350 21586
rect 12402 21534 12404 21586
rect 12236 21532 12404 21534
rect 12348 21522 12404 21532
rect 12684 21364 12740 21374
rect 12684 21270 12740 21308
rect 12124 21074 12180 21084
rect 11228 20638 11230 20690
rect 11282 20638 11284 20690
rect 11228 20626 11284 20638
rect 11340 20914 11396 20926
rect 11340 20862 11342 20914
rect 11394 20862 11396 20914
rect 11004 20244 11060 20254
rect 10780 20188 10948 20244
rect 10556 20020 10612 20030
rect 10220 19236 10276 19964
rect 9996 19180 10276 19236
rect 10332 20018 10612 20020
rect 10332 19966 10558 20018
rect 10610 19966 10612 20018
rect 10332 19964 10612 19966
rect 9996 19122 10052 19180
rect 9996 19070 9998 19122
rect 10050 19070 10052 19122
rect 9996 19058 10052 19070
rect 9828 18508 9940 18564
rect 9996 18674 10052 18686
rect 9996 18622 9998 18674
rect 10050 18622 10052 18674
rect 8316 18450 8596 18452
rect 8316 18398 8318 18450
rect 8370 18398 8596 18450
rect 8316 18396 8596 18398
rect 8764 18450 8820 18462
rect 8764 18398 8766 18450
rect 8818 18398 8820 18450
rect 8316 18386 8372 18396
rect 8204 18162 8260 18172
rect 8764 17780 8820 18398
rect 9772 18450 9828 18508
rect 9772 18398 9774 18450
rect 9826 18398 9828 18450
rect 9772 18386 9828 18398
rect 9884 18116 9940 18126
rect 9884 17780 9940 18060
rect 9996 18004 10052 18622
rect 10108 18450 10164 19180
rect 10108 18398 10110 18450
rect 10162 18398 10164 18450
rect 10108 18386 10164 18398
rect 10108 18228 10164 18238
rect 10108 18134 10164 18172
rect 9996 17948 10164 18004
rect 10108 17892 10164 17948
rect 10108 17826 10164 17836
rect 8764 17666 8820 17724
rect 8764 17614 8766 17666
rect 8818 17614 8820 17666
rect 8764 17602 8820 17614
rect 9436 17778 9940 17780
rect 9436 17726 9886 17778
rect 9938 17726 9940 17778
rect 9436 17724 9940 17726
rect 9436 17666 9492 17724
rect 9884 17714 9940 17724
rect 9436 17614 9438 17666
rect 9490 17614 9492 17666
rect 9436 17602 9492 17614
rect 8428 17556 8484 17566
rect 7756 17554 8484 17556
rect 7756 17502 8430 17554
rect 8482 17502 8484 17554
rect 7756 17500 8484 17502
rect 8428 17490 8484 17500
rect 9100 17556 9156 17566
rect 9100 17462 9156 17500
rect 9548 17556 9604 17566
rect 8092 17108 8148 17118
rect 8092 17014 8148 17052
rect 8540 17108 8596 17118
rect 8540 17014 8596 17052
rect 7756 16996 7812 17006
rect 7308 16994 7812 16996
rect 7308 16942 7758 16994
rect 7810 16942 7812 16994
rect 7308 16940 7812 16942
rect 6972 16884 7028 16894
rect 6972 16790 7028 16828
rect 6748 15934 6750 15986
rect 6802 15934 6804 15986
rect 5628 15150 5630 15202
rect 5682 15150 5684 15202
rect 5628 15138 5684 15150
rect 5068 14642 5124 15036
rect 5068 14590 5070 14642
rect 5122 14590 5124 14642
rect 4620 14578 4676 14588
rect 5068 14578 5124 14590
rect 5852 15092 5908 15102
rect 5852 14642 5908 15036
rect 5852 14590 5854 14642
rect 5906 14590 5908 14642
rect 5852 14578 5908 14590
rect 1820 14478 1822 14530
rect 1874 14478 1876 14530
rect 1820 14466 1876 14478
rect 6188 14084 6244 14094
rect 2604 13858 2660 13870
rect 2604 13806 2606 13858
rect 2658 13806 2660 13858
rect 2492 13076 2548 13086
rect 2604 13076 2660 13806
rect 6076 13858 6132 13870
rect 6076 13806 6078 13858
rect 6130 13806 6132 13858
rect 2940 13746 2996 13758
rect 2940 13694 2942 13746
rect 2994 13694 2996 13746
rect 2940 13188 2996 13694
rect 6076 13748 6132 13806
rect 6076 13682 6132 13692
rect 6188 13746 6244 14028
rect 6188 13694 6190 13746
rect 6242 13694 6244 13746
rect 5068 13522 5124 13534
rect 5068 13470 5070 13522
rect 5122 13470 5124 13522
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 2940 13122 2996 13132
rect 2492 13074 2660 13076
rect 2492 13022 2494 13074
rect 2546 13022 2660 13074
rect 2492 13020 2660 13022
rect 4620 13076 4676 13086
rect 2492 13010 2548 13020
rect 4620 12982 4676 13020
rect 1820 12962 1876 12974
rect 1820 12910 1822 12962
rect 1874 12910 1876 12962
rect 1820 12180 1876 12910
rect 3724 12964 3780 12974
rect 1820 12114 1876 12124
rect 2380 12180 2436 12190
rect 2380 12086 2436 12124
rect 3052 12068 3108 12078
rect 3052 12066 3332 12068
rect 3052 12014 3054 12066
rect 3106 12014 3332 12066
rect 3052 12012 3332 12014
rect 3052 12002 3108 12012
rect 3276 11284 3332 12012
rect 3724 11394 3780 12908
rect 5068 12964 5124 13470
rect 5404 13522 5460 13534
rect 5404 13470 5406 13522
rect 5458 13470 5460 13522
rect 5404 13300 5460 13470
rect 5068 12898 5124 12908
rect 5180 13244 5404 13300
rect 5068 12738 5124 12750
rect 5068 12686 5070 12738
rect 5122 12686 5124 12738
rect 5068 12180 5124 12686
rect 5068 12114 5124 12124
rect 5180 12066 5236 13244
rect 5404 13234 5460 13244
rect 5740 13188 5796 13198
rect 5740 13094 5796 13132
rect 6076 13076 6132 13086
rect 6076 12982 6132 13020
rect 6188 12852 6244 13694
rect 6300 12852 6356 12862
rect 6188 12850 6356 12852
rect 6188 12798 6302 12850
rect 6354 12798 6356 12850
rect 6188 12796 6356 12798
rect 6300 12786 6356 12796
rect 6748 12850 6804 15934
rect 6860 16100 6916 16110
rect 7196 16100 7252 16110
rect 6860 16098 7252 16100
rect 6860 16046 6862 16098
rect 6914 16046 7198 16098
rect 7250 16046 7252 16098
rect 6860 16044 7252 16046
rect 6860 15314 6916 16044
rect 7196 16034 7252 16044
rect 7196 15428 7252 15438
rect 7308 15428 7364 16940
rect 7756 16930 7812 16940
rect 8652 16996 8708 17006
rect 7420 16772 7476 16782
rect 7420 15986 7476 16716
rect 7868 16660 7924 16670
rect 7532 16100 7588 16110
rect 7868 16100 7924 16604
rect 7532 16098 7924 16100
rect 7532 16046 7534 16098
rect 7586 16046 7870 16098
rect 7922 16046 7924 16098
rect 7532 16044 7924 16046
rect 7532 16034 7588 16044
rect 7868 16034 7924 16044
rect 8540 16098 8596 16110
rect 8540 16046 8542 16098
rect 8594 16046 8596 16098
rect 7420 15934 7422 15986
rect 7474 15934 7476 15986
rect 7420 15876 7476 15934
rect 7420 15820 7924 15876
rect 7868 15764 7924 15820
rect 7868 15538 7924 15708
rect 7868 15486 7870 15538
rect 7922 15486 7924 15538
rect 7868 15474 7924 15486
rect 7980 15874 8036 15886
rect 7980 15822 7982 15874
rect 8034 15822 8036 15874
rect 6860 15262 6862 15314
rect 6914 15262 6916 15314
rect 6860 15250 6916 15262
rect 7084 15426 7364 15428
rect 7084 15374 7198 15426
rect 7250 15374 7364 15426
rect 7084 15372 7364 15374
rect 7980 15428 8036 15822
rect 6972 15092 7028 15102
rect 6972 14530 7028 15036
rect 6972 14478 6974 14530
rect 7026 14478 7028 14530
rect 6972 14466 7028 14478
rect 7084 13748 7140 15372
rect 7196 15362 7252 15372
rect 7980 15362 8036 15372
rect 8204 15874 8260 15886
rect 8204 15822 8206 15874
rect 8258 15822 8260 15874
rect 8204 15148 8260 15822
rect 8428 15428 8484 15438
rect 8428 15334 8484 15372
rect 7980 15092 8260 15148
rect 8540 15204 8596 16046
rect 8540 15138 8596 15148
rect 7980 14532 8036 15092
rect 7980 14476 8148 14532
rect 7644 14420 7700 14430
rect 7644 14418 8036 14420
rect 7644 14366 7646 14418
rect 7698 14366 8036 14418
rect 7644 14364 8036 14366
rect 7644 14354 7700 14364
rect 7980 13970 8036 14364
rect 7980 13918 7982 13970
rect 8034 13918 8036 13970
rect 7980 13906 8036 13918
rect 7084 13682 7140 13692
rect 7980 13748 8036 13758
rect 7532 12964 7588 12974
rect 6748 12798 6750 12850
rect 6802 12798 6804 12850
rect 5628 12180 5684 12190
rect 5628 12086 5684 12124
rect 6188 12180 6244 12190
rect 6188 12086 6244 12124
rect 5180 12014 5182 12066
rect 5234 12014 5236 12066
rect 5180 12002 5236 12014
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 3724 11342 3726 11394
rect 3778 11342 3780 11394
rect 3724 11330 3780 11342
rect 3388 11284 3444 11294
rect 3276 11282 3444 11284
rect 3276 11230 3390 11282
rect 3442 11230 3444 11282
rect 3276 11228 3444 11230
rect 3388 11218 3444 11228
rect 6748 11284 6804 12798
rect 7420 12962 7588 12964
rect 7420 12910 7534 12962
rect 7586 12910 7588 12962
rect 7420 12908 7588 12910
rect 7308 12740 7364 12750
rect 6860 12738 7364 12740
rect 6860 12686 7310 12738
rect 7362 12686 7364 12738
rect 6860 12684 7364 12686
rect 6860 12290 6916 12684
rect 7308 12674 7364 12684
rect 6860 12238 6862 12290
rect 6914 12238 6916 12290
rect 6860 12226 6916 12238
rect 7308 11620 7364 11630
rect 7420 11620 7476 12908
rect 7532 12898 7588 12908
rect 7308 11618 7476 11620
rect 7308 11566 7310 11618
rect 7362 11566 7476 11618
rect 7308 11564 7476 11566
rect 7644 11956 7700 11966
rect 7644 11618 7700 11900
rect 7644 11566 7646 11618
rect 7698 11566 7700 11618
rect 7308 11554 7364 11564
rect 7644 11554 7700 11566
rect 6748 11218 6804 11228
rect 7980 10722 8036 13692
rect 7980 10670 7982 10722
rect 8034 10670 8036 10722
rect 7980 10658 8036 10670
rect 8092 11394 8148 14476
rect 8316 13748 8372 13758
rect 8316 13654 8372 13692
rect 8652 13186 8708 16940
rect 9212 15988 9268 15998
rect 8988 15986 9268 15988
rect 8988 15934 9214 15986
rect 9266 15934 9268 15986
rect 8988 15932 9268 15934
rect 8988 15538 9044 15932
rect 9212 15922 9268 15932
rect 8988 15486 8990 15538
rect 9042 15486 9044 15538
rect 8988 15474 9044 15486
rect 8764 15314 8820 15326
rect 8764 15262 8766 15314
rect 8818 15262 8820 15314
rect 8764 14756 8820 15262
rect 8764 14690 8820 14700
rect 9100 15204 9156 15214
rect 9100 13970 9156 15148
rect 9100 13918 9102 13970
rect 9154 13918 9156 13970
rect 9100 13906 9156 13918
rect 9548 13748 9604 17500
rect 10332 17106 10388 19964
rect 10556 19954 10612 19964
rect 10668 19796 10724 20076
rect 10556 19740 10724 19796
rect 10780 20018 10836 20030
rect 10780 19966 10782 20018
rect 10834 19966 10836 20018
rect 10556 18676 10612 19740
rect 10556 18610 10612 18620
rect 10668 19124 10724 19134
rect 10780 19124 10836 19966
rect 10892 20020 10948 20188
rect 11004 20242 11284 20244
rect 11004 20190 11006 20242
rect 11058 20190 11284 20242
rect 11004 20188 11284 20190
rect 11004 20178 11060 20188
rect 11004 20020 11060 20030
rect 10892 20018 11060 20020
rect 10892 19966 11006 20018
rect 11058 19966 11060 20018
rect 10892 19964 11060 19966
rect 11004 19954 11060 19964
rect 11116 20020 11172 20030
rect 11116 19458 11172 19964
rect 11116 19406 11118 19458
rect 11170 19406 11172 19458
rect 11116 19394 11172 19406
rect 10668 19122 10836 19124
rect 10668 19070 10670 19122
rect 10722 19070 10836 19122
rect 10668 19068 10836 19070
rect 11004 19234 11060 19246
rect 11004 19182 11006 19234
rect 11058 19182 11060 19234
rect 10668 18564 10724 19068
rect 10668 18498 10724 18508
rect 10892 19010 10948 19022
rect 10892 18958 10894 19010
rect 10946 18958 10948 19010
rect 10892 18452 10948 18958
rect 10892 18386 10948 18396
rect 10332 17054 10334 17106
rect 10386 17054 10388 17106
rect 10332 17042 10388 17054
rect 11004 17106 11060 19182
rect 11228 18788 11284 20188
rect 11340 19234 11396 20862
rect 12796 20244 12852 20254
rect 12572 19460 12628 19470
rect 12572 19366 12628 19404
rect 12684 19236 12740 19246
rect 11340 19182 11342 19234
rect 11394 19182 11396 19234
rect 11340 19170 11396 19182
rect 12572 19234 12740 19236
rect 12572 19182 12686 19234
rect 12738 19182 12740 19234
rect 12572 19180 12740 19182
rect 12124 19124 12180 19134
rect 11900 19122 12180 19124
rect 11900 19070 12126 19122
rect 12178 19070 12180 19122
rect 11900 19068 12180 19070
rect 11228 18732 11508 18788
rect 11116 18676 11172 18686
rect 11172 18620 11284 18676
rect 11116 18610 11172 18620
rect 11004 17054 11006 17106
rect 11058 17054 11060 17106
rect 11004 17042 11060 17054
rect 11116 18450 11172 18462
rect 11116 18398 11118 18450
rect 11170 18398 11172 18450
rect 11116 16996 11172 18398
rect 11228 17556 11284 18620
rect 11340 18450 11396 18462
rect 11340 18398 11342 18450
rect 11394 18398 11396 18450
rect 11340 18228 11396 18398
rect 11452 18452 11508 18732
rect 11564 18676 11620 18686
rect 11564 18674 11844 18676
rect 11564 18622 11566 18674
rect 11618 18622 11844 18674
rect 11564 18620 11844 18622
rect 11564 18610 11620 18620
rect 11564 18452 11620 18462
rect 11452 18450 11620 18452
rect 11452 18398 11566 18450
rect 11618 18398 11620 18450
rect 11452 18396 11620 18398
rect 11564 18386 11620 18396
rect 11676 18450 11732 18462
rect 11676 18398 11678 18450
rect 11730 18398 11732 18450
rect 11676 18340 11732 18398
rect 11676 18274 11732 18284
rect 11452 18228 11508 18238
rect 11340 18172 11452 18228
rect 11452 18162 11508 18172
rect 11788 18004 11844 18620
rect 11788 17938 11844 17948
rect 11340 17556 11396 17566
rect 11228 17554 11396 17556
rect 11228 17502 11342 17554
rect 11394 17502 11396 17554
rect 11228 17500 11396 17502
rect 11340 17490 11396 17500
rect 11676 17444 11732 17454
rect 11676 17350 11732 17388
rect 11116 16930 11172 16940
rect 10220 16770 10276 16782
rect 10220 16718 10222 16770
rect 10274 16718 10276 16770
rect 9660 15876 9716 15886
rect 9660 14084 9716 15820
rect 9996 15316 10052 15326
rect 9996 15222 10052 15260
rect 10220 15148 10276 16718
rect 11116 16770 11172 16782
rect 11116 16718 11118 16770
rect 11170 16718 11172 16770
rect 11116 16212 11172 16718
rect 11564 16772 11620 16782
rect 11340 16212 11396 16222
rect 11116 16210 11508 16212
rect 11116 16158 11342 16210
rect 11394 16158 11508 16210
rect 11116 16156 11508 16158
rect 11340 16146 11396 16156
rect 10108 15092 10276 15148
rect 10108 14980 10164 15092
rect 9772 14924 10164 14980
rect 9772 14642 9828 14924
rect 9772 14590 9774 14642
rect 9826 14590 9828 14642
rect 9772 14578 9828 14590
rect 9660 14018 9716 14028
rect 9772 13748 9828 13758
rect 9548 13692 9716 13748
rect 9548 13524 9604 13534
rect 8652 13134 8654 13186
rect 8706 13134 8708 13186
rect 8652 13122 8708 13134
rect 8988 13300 9044 13310
rect 8988 13186 9044 13244
rect 8988 13134 8990 13186
rect 9042 13134 9044 13186
rect 8988 13122 9044 13134
rect 9548 12962 9604 13468
rect 9548 12910 9550 12962
rect 9602 12910 9604 12962
rect 9548 12898 9604 12910
rect 8988 12292 9044 12302
rect 8092 11342 8094 11394
rect 8146 11342 8148 11394
rect 8092 10610 8148 11342
rect 8428 12180 8484 12190
rect 8204 11284 8260 11294
rect 8204 11190 8260 11228
rect 8092 10558 8094 10610
rect 8146 10558 8148 10610
rect 8092 10546 8148 10558
rect 7084 10388 7140 10398
rect 6860 10386 7140 10388
rect 6860 10334 7086 10386
rect 7138 10334 7140 10386
rect 6860 10332 7140 10334
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 6860 9826 6916 10332
rect 7084 10322 7140 10332
rect 7420 10386 7476 10398
rect 7420 10334 7422 10386
rect 7474 10334 7476 10386
rect 6860 9774 6862 9826
rect 6914 9774 6916 9826
rect 6860 9762 6916 9774
rect 6524 9604 6580 9614
rect 6412 9602 6580 9604
rect 6412 9550 6526 9602
rect 6578 9550 6580 9602
rect 6412 9548 6580 9550
rect 6412 9154 6468 9548
rect 6524 9538 6580 9548
rect 6412 9102 6414 9154
rect 6466 9102 6468 9154
rect 6412 9090 6468 9102
rect 5740 9044 5796 9054
rect 5740 8950 5796 8988
rect 7420 8932 7476 10334
rect 8428 9826 8484 12124
rect 8988 12068 9044 12236
rect 8988 11974 9044 12012
rect 9212 12180 9268 12190
rect 9548 12180 9604 12190
rect 9268 12178 9604 12180
rect 9268 12126 9550 12178
rect 9602 12126 9604 12178
rect 9268 12124 9604 12126
rect 9212 11506 9268 12124
rect 9548 12114 9604 12124
rect 9660 11732 9716 13692
rect 9996 13748 10052 14924
rect 11116 14756 11172 14766
rect 11116 14662 11172 14700
rect 11452 14754 11508 16156
rect 11452 14702 11454 14754
rect 11506 14702 11508 14754
rect 11452 14690 11508 14702
rect 10444 14420 10500 14430
rect 10444 14418 11060 14420
rect 10444 14366 10446 14418
rect 10498 14366 11060 14418
rect 10444 14364 11060 14366
rect 10444 14354 10500 14364
rect 10108 14308 10164 14318
rect 10108 14306 10388 14308
rect 10108 14254 10110 14306
rect 10162 14254 10388 14306
rect 10108 14252 10388 14254
rect 10108 14242 10164 14252
rect 10108 13748 10164 13758
rect 9996 13746 10164 13748
rect 9996 13694 10110 13746
rect 10162 13694 10164 13746
rect 9996 13692 10164 13694
rect 9772 13654 9828 13692
rect 10108 13682 10164 13692
rect 9772 12852 9828 12862
rect 9772 12758 9828 12796
rect 10332 12290 10388 14252
rect 10892 14196 10948 14206
rect 10780 13860 10836 13870
rect 10780 13766 10836 13804
rect 10892 13746 10948 14140
rect 10892 13694 10894 13746
rect 10946 13694 10948 13746
rect 10892 13682 10948 13694
rect 10780 12964 10836 12974
rect 10780 12870 10836 12908
rect 11004 12740 11060 14364
rect 11452 13972 11508 13982
rect 11564 13972 11620 16716
rect 11788 16212 11844 16222
rect 11788 15204 11844 16156
rect 11788 15138 11844 15148
rect 11900 15148 11956 19068
rect 12124 19058 12180 19068
rect 12348 19122 12404 19134
rect 12348 19070 12350 19122
rect 12402 19070 12404 19122
rect 12236 18452 12292 18462
rect 12124 18450 12292 18452
rect 12124 18398 12238 18450
rect 12290 18398 12292 18450
rect 12124 18396 12292 18398
rect 12012 17556 12068 17566
rect 12012 17462 12068 17500
rect 12124 16772 12180 18396
rect 12236 18386 12292 18396
rect 12348 18452 12404 19070
rect 12460 18452 12516 18462
rect 12348 18450 12516 18452
rect 12348 18398 12462 18450
rect 12514 18398 12516 18450
rect 12348 18396 12516 18398
rect 12348 18228 12404 18396
rect 12460 18386 12516 18396
rect 12348 17666 12404 18172
rect 12572 18228 12628 19180
rect 12684 19170 12740 19180
rect 12684 18452 12740 18462
rect 12684 18358 12740 18396
rect 12796 18450 12852 20188
rect 12908 19348 12964 19358
rect 12908 19010 12964 19292
rect 12908 18958 12910 19010
rect 12962 18958 12964 19010
rect 12908 18946 12964 18958
rect 12796 18398 12798 18450
rect 12850 18398 12852 18450
rect 12796 18340 12852 18398
rect 13020 18674 13076 18686
rect 13020 18622 13022 18674
rect 13074 18622 13076 18674
rect 13020 18452 13076 18622
rect 13020 18386 13076 18396
rect 12796 18274 12852 18284
rect 12460 17892 12516 17902
rect 12460 17798 12516 17836
rect 12348 17614 12350 17666
rect 12402 17614 12404 17666
rect 12348 17556 12404 17614
rect 12572 17666 12628 18172
rect 12572 17614 12574 17666
rect 12626 17614 12628 17666
rect 12572 17602 12628 17614
rect 12796 17668 12852 17678
rect 12348 17490 12404 17500
rect 12796 17442 12852 17612
rect 12796 17390 12798 17442
rect 12850 17390 12852 17442
rect 12796 17378 12852 17390
rect 12124 16706 12180 16716
rect 12684 16324 12740 16334
rect 12236 15874 12292 15886
rect 12236 15822 12238 15874
rect 12290 15822 12292 15874
rect 12236 15764 12292 15822
rect 12236 15698 12292 15708
rect 12460 15874 12516 15886
rect 12460 15822 12462 15874
rect 12514 15822 12516 15874
rect 12460 15148 12516 15822
rect 12684 15874 12740 16268
rect 12796 16100 12852 16110
rect 12796 16006 12852 16044
rect 12684 15822 12686 15874
rect 12738 15822 12740 15874
rect 12684 15764 12740 15822
rect 12684 15698 12740 15708
rect 11900 15092 12180 15148
rect 12012 14418 12068 14430
rect 12012 14366 12014 14418
rect 12066 14366 12068 14418
rect 12012 14308 12068 14366
rect 12012 14242 12068 14252
rect 11452 13970 11620 13972
rect 11452 13918 11454 13970
rect 11506 13918 11620 13970
rect 11452 13916 11620 13918
rect 11452 13906 11508 13916
rect 11676 13860 11732 13870
rect 11564 12852 11620 12862
rect 11676 12852 11732 13804
rect 11788 13522 11844 13534
rect 11788 13470 11790 13522
rect 11842 13470 11844 13522
rect 11788 13076 11844 13470
rect 11788 13010 11844 13020
rect 12012 12852 12068 12862
rect 11676 12796 11844 12852
rect 11004 12684 11284 12740
rect 10332 12238 10334 12290
rect 10386 12238 10388 12290
rect 10332 12226 10388 12238
rect 9660 11666 9716 11676
rect 11228 11618 11284 12684
rect 11228 11566 11230 11618
rect 11282 11566 11284 11618
rect 11228 11554 11284 11566
rect 11564 12068 11620 12796
rect 11564 11618 11620 12012
rect 11564 11566 11566 11618
rect 11618 11566 11620 11618
rect 11564 11554 11620 11566
rect 11676 11732 11732 11742
rect 9212 11454 9214 11506
rect 9266 11454 9268 11506
rect 9212 11442 9268 11454
rect 11564 10836 11620 10846
rect 11564 10742 11620 10780
rect 8428 9774 8430 9826
rect 8482 9774 8484 9826
rect 8428 9044 8484 9774
rect 10892 10612 10948 10622
rect 8428 8978 8484 8988
rect 8540 9716 8596 9726
rect 7420 8866 7476 8876
rect 8540 8932 8596 9660
rect 9100 9716 9156 9726
rect 9100 9714 9604 9716
rect 9100 9662 9102 9714
rect 9154 9662 9604 9714
rect 9100 9660 9604 9662
rect 9100 9650 9156 9660
rect 9548 9266 9604 9660
rect 9548 9214 9550 9266
rect 9602 9214 9604 9266
rect 9548 9202 9604 9214
rect 8540 8838 8596 8876
rect 8988 9044 9044 9054
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 8988 8428 9044 8988
rect 9884 9044 9940 9054
rect 9884 8950 9940 8988
rect 10444 9044 10500 9054
rect 10444 8950 10500 8988
rect 10780 9044 10836 9054
rect 10892 9044 10948 10556
rect 10780 9042 10948 9044
rect 10780 8990 10782 9042
rect 10834 8990 10948 9042
rect 10780 8988 10948 8990
rect 10780 8978 10836 8988
rect 8988 8372 9380 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 9324 6692 9380 8372
rect 10892 7924 10948 8988
rect 11004 10500 11060 10510
rect 11004 8428 11060 10444
rect 11676 10050 11732 11676
rect 11788 11172 11844 12796
rect 12012 11394 12068 12796
rect 12124 11844 12180 15092
rect 12348 15092 12516 15148
rect 12572 15316 12628 15326
rect 12572 15202 12628 15260
rect 12572 15150 12574 15202
rect 12626 15150 12628 15202
rect 12236 14532 12292 14542
rect 12348 14532 12404 15092
rect 12236 14530 12404 14532
rect 12236 14478 12238 14530
rect 12290 14478 12404 14530
rect 12236 14476 12404 14478
rect 12572 14532 12628 15150
rect 13132 15148 13188 22204
rect 13244 21474 13300 21486
rect 13244 21422 13246 21474
rect 13298 21422 13300 21474
rect 13244 21140 13300 21422
rect 13244 21074 13300 21084
rect 13356 20020 13412 23884
rect 13468 23874 13524 23884
rect 13580 23378 13636 24892
rect 13804 24722 13860 24734
rect 13804 24670 13806 24722
rect 13858 24670 13860 24722
rect 13804 23548 13860 24670
rect 13580 23326 13582 23378
rect 13634 23326 13636 23378
rect 13580 23314 13636 23326
rect 13692 23492 13860 23548
rect 13692 23380 13748 23492
rect 13692 23314 13748 23324
rect 13692 23154 13748 23166
rect 13692 23102 13694 23154
rect 13746 23102 13748 23154
rect 13580 22930 13636 22942
rect 13580 22878 13582 22930
rect 13634 22878 13636 22930
rect 13580 22260 13636 22878
rect 13692 22820 13748 23102
rect 13692 22754 13748 22764
rect 13692 22484 13748 22494
rect 13916 22484 13972 25228
rect 14028 24836 14084 24846
rect 14028 24834 14308 24836
rect 14028 24782 14030 24834
rect 14082 24782 14308 24834
rect 14028 24780 14308 24782
rect 14028 24770 14084 24780
rect 14252 24050 14308 24780
rect 14252 23998 14254 24050
rect 14306 23998 14308 24050
rect 14252 23986 14308 23998
rect 14364 23492 14420 23502
rect 14028 23380 14084 23390
rect 14028 22594 14084 23324
rect 14028 22542 14030 22594
rect 14082 22542 14084 22594
rect 14028 22530 14084 22542
rect 14140 22930 14196 22942
rect 14140 22878 14142 22930
rect 14194 22878 14196 22930
rect 13692 22482 13972 22484
rect 13692 22430 13694 22482
rect 13746 22430 13972 22482
rect 13692 22428 13972 22430
rect 13692 22418 13748 22428
rect 14140 22260 14196 22878
rect 14364 22594 14420 23436
rect 14476 23154 14532 25340
rect 14924 24612 14980 24622
rect 15260 24612 15316 25452
rect 14980 24556 15316 24612
rect 14924 24518 14980 24556
rect 15260 23492 15316 23502
rect 15260 23266 15316 23436
rect 15596 23268 15652 23278
rect 15260 23214 15262 23266
rect 15314 23214 15316 23266
rect 15260 23202 15316 23214
rect 15484 23212 15596 23268
rect 14476 23102 14478 23154
rect 14530 23102 14532 23154
rect 14476 23090 14532 23102
rect 15148 23154 15204 23166
rect 15148 23102 15150 23154
rect 15202 23102 15204 23154
rect 14588 22820 14644 22830
rect 14364 22542 14366 22594
rect 14418 22542 14420 22594
rect 14364 22530 14420 22542
rect 14476 22764 14588 22820
rect 13580 22194 13636 22204
rect 13804 22204 14196 22260
rect 13804 21698 13860 22204
rect 13804 21646 13806 21698
rect 13858 21646 13860 21698
rect 13804 21634 13860 21646
rect 14252 21812 14308 21822
rect 14028 21588 14084 21598
rect 13916 21586 14084 21588
rect 13916 21534 14030 21586
rect 14082 21534 14084 21586
rect 13916 21532 14084 21534
rect 13916 21476 13972 21532
rect 14028 21522 14084 21532
rect 14252 21586 14308 21756
rect 14252 21534 14254 21586
rect 14306 21534 14308 21586
rect 14252 21522 14308 21534
rect 14364 21588 14420 21598
rect 13692 21420 13972 21476
rect 13468 21364 13524 21374
rect 13468 20802 13524 21308
rect 13468 20750 13470 20802
rect 13522 20750 13524 20802
rect 13468 20738 13524 20750
rect 13692 20802 13748 21420
rect 13916 21252 13972 21262
rect 13916 21026 13972 21196
rect 13916 20974 13918 21026
rect 13970 20974 13972 21026
rect 13916 20962 13972 20974
rect 13692 20750 13694 20802
rect 13746 20750 13748 20802
rect 13244 19964 13412 20020
rect 13580 20578 13636 20590
rect 13580 20526 13582 20578
rect 13634 20526 13636 20578
rect 13244 16212 13300 19964
rect 13356 19796 13412 19806
rect 13356 19702 13412 19740
rect 13468 19794 13524 19806
rect 13468 19742 13470 19794
rect 13522 19742 13524 19794
rect 13468 19348 13524 19742
rect 13580 19796 13636 20526
rect 13692 20020 13748 20750
rect 13804 20804 13860 20814
rect 13804 20130 13860 20748
rect 14028 20804 14084 20814
rect 14364 20804 14420 21532
rect 14028 20802 14420 20804
rect 14028 20750 14030 20802
rect 14082 20750 14420 20802
rect 14028 20748 14420 20750
rect 14028 20244 14084 20748
rect 14028 20178 14084 20188
rect 14364 20580 14420 20590
rect 13804 20078 13806 20130
rect 13858 20078 13860 20130
rect 13804 20066 13860 20078
rect 13916 20132 13972 20142
rect 13692 19954 13748 19964
rect 13580 19730 13636 19740
rect 13692 19794 13748 19806
rect 13692 19742 13694 19794
rect 13746 19742 13748 19794
rect 13468 19282 13524 19292
rect 13580 19236 13636 19246
rect 13356 17556 13412 17566
rect 13356 17106 13412 17500
rect 13356 17054 13358 17106
rect 13410 17054 13412 17106
rect 13356 17042 13412 17054
rect 13244 15316 13300 16156
rect 13580 16100 13636 19180
rect 13692 19012 13748 19742
rect 13916 19012 13972 20076
rect 13692 18946 13748 18956
rect 13804 18956 13972 19012
rect 14028 20020 14084 20030
rect 14028 19122 14084 19964
rect 14028 19070 14030 19122
rect 14082 19070 14084 19122
rect 13692 18676 13748 18686
rect 13692 18450 13748 18620
rect 13692 18398 13694 18450
rect 13746 18398 13748 18450
rect 13692 18228 13748 18398
rect 13692 18162 13748 18172
rect 13804 18004 13860 18956
rect 13916 18788 13972 18798
rect 13916 18226 13972 18732
rect 14028 18452 14084 19070
rect 14140 20018 14196 20030
rect 14140 19966 14142 20018
rect 14194 19966 14196 20018
rect 14140 18676 14196 19966
rect 14364 19794 14420 20524
rect 14364 19742 14366 19794
rect 14418 19742 14420 19794
rect 14364 19730 14420 19742
rect 14140 18610 14196 18620
rect 14252 19234 14308 19246
rect 14252 19182 14254 19234
rect 14306 19182 14308 19234
rect 14252 18900 14308 19182
rect 14476 19236 14532 22764
rect 14588 22754 14644 22764
rect 14924 22708 14980 22718
rect 14588 22260 14644 22270
rect 14588 22166 14644 22204
rect 14924 22260 14980 22652
rect 14924 22258 15092 22260
rect 14924 22206 14926 22258
rect 14978 22206 15092 22258
rect 14924 22204 15092 22206
rect 14924 22194 14980 22204
rect 15036 21924 15092 22204
rect 15148 22036 15204 23102
rect 15260 22036 15316 22046
rect 15148 21980 15260 22036
rect 15260 21970 15316 21980
rect 15036 21858 15092 21868
rect 14588 21810 14644 21822
rect 14588 21758 14590 21810
rect 14642 21758 14644 21810
rect 14588 19236 14644 21758
rect 15148 20804 15204 20814
rect 15148 20710 15204 20748
rect 15372 20802 15428 20814
rect 15372 20750 15374 20802
rect 15426 20750 15428 20802
rect 15372 20244 15428 20750
rect 15372 20178 15428 20188
rect 14700 20020 14756 20030
rect 14700 19926 14756 19964
rect 14924 20020 14980 20030
rect 15484 20020 15540 23212
rect 15596 23202 15652 23212
rect 15820 23042 15876 23054
rect 15820 22990 15822 23042
rect 15874 22990 15876 23042
rect 15820 22820 15876 22990
rect 15820 22754 15876 22764
rect 15708 22146 15764 22158
rect 15708 22094 15710 22146
rect 15762 22094 15764 22146
rect 15708 22036 15764 22094
rect 15708 21970 15764 21980
rect 15932 21924 15988 26852
rect 16044 25618 16100 27132
rect 16268 27186 16324 27916
rect 16268 27134 16270 27186
rect 16322 27134 16324 27186
rect 16268 27122 16324 27134
rect 16156 26178 16212 26190
rect 16156 26126 16158 26178
rect 16210 26126 16212 26178
rect 16156 26068 16212 26126
rect 16156 26002 16212 26012
rect 16044 25566 16046 25618
rect 16098 25566 16100 25618
rect 16044 25554 16100 25566
rect 16380 24050 16436 24062
rect 16380 23998 16382 24050
rect 16434 23998 16436 24050
rect 16380 23492 16436 23998
rect 16380 23426 16436 23436
rect 16380 23268 16436 23278
rect 16380 23174 16436 23212
rect 16156 22484 16212 22494
rect 16044 22428 16156 22484
rect 16044 22146 16100 22428
rect 16156 22418 16212 22428
rect 16044 22094 16046 22146
rect 16098 22094 16100 22146
rect 16044 22082 16100 22094
rect 16380 22148 16436 22158
rect 16380 22054 16436 22092
rect 15932 21868 16212 21924
rect 15932 21700 15988 21710
rect 15932 21606 15988 21644
rect 15596 21588 15652 21598
rect 15596 21028 15652 21532
rect 16156 21586 16212 21868
rect 16156 21534 16158 21586
rect 16210 21534 16212 21586
rect 16156 21364 16212 21534
rect 16156 21298 16212 21308
rect 16156 21140 16212 21150
rect 15596 20972 16100 21028
rect 15596 20802 15652 20972
rect 15596 20750 15598 20802
rect 15650 20750 15652 20802
rect 15596 20738 15652 20750
rect 15932 20804 15988 20814
rect 15932 20242 15988 20748
rect 15932 20190 15934 20242
rect 15986 20190 15988 20242
rect 15932 20178 15988 20190
rect 15820 20020 15876 20030
rect 14924 19926 14980 19964
rect 15148 19964 15540 20020
rect 15708 20018 15876 20020
rect 15708 19966 15822 20018
rect 15874 19966 15876 20018
rect 15708 19964 15876 19966
rect 14812 19906 14868 19918
rect 14812 19854 14814 19906
rect 14866 19854 14868 19906
rect 14812 19460 14868 19854
rect 14924 19460 14980 19470
rect 15148 19460 15204 19964
rect 15596 19908 15652 19918
rect 14812 19458 14980 19460
rect 14812 19406 14926 19458
rect 14978 19406 14980 19458
rect 14812 19404 14980 19406
rect 14924 19394 14980 19404
rect 15036 19404 15204 19460
rect 15260 19906 15652 19908
rect 15260 19854 15598 19906
rect 15650 19854 15652 19906
rect 15260 19852 15652 19854
rect 15260 19458 15316 19852
rect 15596 19842 15652 19852
rect 15260 19406 15262 19458
rect 15314 19406 15316 19458
rect 14700 19236 14756 19246
rect 14588 19234 14756 19236
rect 14588 19182 14702 19234
rect 14754 19182 14756 19234
rect 14588 19180 14756 19182
rect 14476 19170 14532 19180
rect 14700 19170 14756 19180
rect 14140 18452 14196 18462
rect 14028 18450 14196 18452
rect 14028 18398 14142 18450
rect 14194 18398 14196 18450
rect 14028 18396 14196 18398
rect 14140 18386 14196 18396
rect 14252 18228 14308 18844
rect 15036 18788 15092 19404
rect 15260 19394 15316 19406
rect 15148 19234 15204 19246
rect 15148 19182 15150 19234
rect 15202 19182 15204 19234
rect 15148 19012 15204 19182
rect 15708 19124 15764 19964
rect 15820 19954 15876 19964
rect 16044 20018 16100 20972
rect 16044 19966 16046 20018
rect 16098 19966 16100 20018
rect 16044 19954 16100 19966
rect 16156 19796 16212 21084
rect 16380 20578 16436 20590
rect 16380 20526 16382 20578
rect 16434 20526 16436 20578
rect 16380 20244 16436 20526
rect 16380 20178 16436 20188
rect 15148 18946 15204 18956
rect 15372 19068 15764 19124
rect 15932 19740 16212 19796
rect 14364 18732 14644 18788
rect 15036 18732 15204 18788
rect 14364 18674 14420 18732
rect 14364 18622 14366 18674
rect 14418 18622 14420 18674
rect 14364 18610 14420 18622
rect 14588 18676 14644 18732
rect 14588 18620 14868 18676
rect 14476 18564 14532 18574
rect 14476 18562 14756 18564
rect 14476 18510 14478 18562
rect 14530 18510 14756 18562
rect 14476 18508 14756 18510
rect 14476 18498 14532 18508
rect 13916 18174 13918 18226
rect 13970 18174 13972 18226
rect 13916 18162 13972 18174
rect 14140 18172 14308 18228
rect 14028 18004 14084 18014
rect 13804 17948 13972 18004
rect 13804 17668 13860 17678
rect 13804 17574 13860 17612
rect 13916 17442 13972 17948
rect 14028 17890 14084 17948
rect 14028 17838 14030 17890
rect 14082 17838 14084 17890
rect 14028 17826 14084 17838
rect 13916 17390 13918 17442
rect 13970 17390 13972 17442
rect 13916 17378 13972 17390
rect 13692 17108 13748 17118
rect 14140 17108 14196 18172
rect 14252 17892 14308 17902
rect 14252 17798 14308 17836
rect 13692 17106 14196 17108
rect 13692 17054 13694 17106
rect 13746 17054 14196 17106
rect 13692 17052 14196 17054
rect 14252 17444 14308 17454
rect 13692 17042 13748 17052
rect 13468 16044 13636 16100
rect 13692 16100 13748 16110
rect 13468 15540 13524 16044
rect 13580 15876 13636 15886
rect 13580 15782 13636 15820
rect 13580 15540 13636 15550
rect 13468 15538 13636 15540
rect 13468 15486 13582 15538
rect 13634 15486 13636 15538
rect 13468 15484 13636 15486
rect 13580 15428 13636 15484
rect 13580 15362 13636 15372
rect 13692 15426 13748 16044
rect 14140 16100 14196 16110
rect 14140 16006 14196 16044
rect 13804 15986 13860 15998
rect 13804 15934 13806 15986
rect 13858 15934 13860 15986
rect 13804 15540 13860 15934
rect 13804 15474 13860 15484
rect 13916 15988 13972 15998
rect 13692 15374 13694 15426
rect 13746 15374 13748 15426
rect 13692 15362 13748 15374
rect 13244 15250 13300 15260
rect 13132 15092 13300 15148
rect 12236 14196 12292 14476
rect 12572 14466 12628 14476
rect 13132 14532 13188 14542
rect 12236 14130 12292 14140
rect 12684 14420 12740 14430
rect 12460 13858 12516 13870
rect 12460 13806 12462 13858
rect 12514 13806 12516 13858
rect 12460 13188 12516 13806
rect 12572 13748 12628 13758
rect 12684 13748 12740 14364
rect 12572 13746 12740 13748
rect 12572 13694 12574 13746
rect 12626 13694 12740 13746
rect 12572 13692 12740 13694
rect 12572 13682 12628 13692
rect 12460 13122 12516 13132
rect 12684 13524 12740 13692
rect 12572 13076 12628 13086
rect 12236 12068 12292 12078
rect 12460 12068 12516 12078
rect 12292 12066 12516 12068
rect 12292 12014 12462 12066
rect 12514 12014 12516 12066
rect 12292 12012 12516 12014
rect 12236 12002 12292 12012
rect 12460 12002 12516 12012
rect 12572 12068 12628 13020
rect 12124 11788 12404 11844
rect 12012 11342 12014 11394
rect 12066 11342 12068 11394
rect 12012 11330 12068 11342
rect 12236 11620 12292 11630
rect 12124 11282 12180 11294
rect 12124 11230 12126 11282
rect 12178 11230 12180 11282
rect 12124 11172 12180 11230
rect 11788 11116 12180 11172
rect 12124 10836 12180 10846
rect 12236 10836 12292 11564
rect 12180 10780 12292 10836
rect 12124 10742 12180 10780
rect 11788 10722 11844 10734
rect 11788 10670 11790 10722
rect 11842 10670 11844 10722
rect 11788 10612 11844 10670
rect 11788 10546 11844 10556
rect 11676 9998 11678 10050
rect 11730 9998 11732 10050
rect 11676 9986 11732 9998
rect 11228 9940 11284 9950
rect 12012 9940 12068 9950
rect 11284 9884 11396 9940
rect 11228 9846 11284 9884
rect 11340 9154 11396 9884
rect 12012 9846 12068 9884
rect 11340 9102 11342 9154
rect 11394 9102 11396 9154
rect 11340 9090 11396 9102
rect 11564 9604 11620 9614
rect 11564 9042 11620 9548
rect 12236 9268 12292 9278
rect 12348 9268 12404 11788
rect 12460 10612 12516 10622
rect 12572 10612 12628 12012
rect 12460 10610 12628 10612
rect 12460 10558 12462 10610
rect 12514 10558 12628 10610
rect 12460 10556 12628 10558
rect 12460 10500 12516 10556
rect 12460 10434 12516 10444
rect 12684 9828 12740 13468
rect 12908 14306 12964 14318
rect 12908 14254 12910 14306
rect 12962 14254 12964 14306
rect 12908 13748 12964 14254
rect 12908 13076 12964 13692
rect 13020 13634 13076 13646
rect 13020 13582 13022 13634
rect 13074 13582 13076 13634
rect 13020 13188 13076 13582
rect 13020 13122 13076 13132
rect 12908 13010 12964 13020
rect 13132 12964 13188 14476
rect 13132 12402 13188 12908
rect 13132 12350 13134 12402
rect 13186 12350 13188 12402
rect 13132 12338 13188 12350
rect 13244 11620 13300 15092
rect 13580 15092 13636 15102
rect 13580 15090 13748 15092
rect 13580 15038 13582 15090
rect 13634 15038 13748 15090
rect 13580 15036 13748 15038
rect 13580 15026 13636 15036
rect 13468 14420 13524 14430
rect 13468 14326 13524 14364
rect 13692 12852 13748 15036
rect 13916 14308 13972 15932
rect 14252 15148 14308 17388
rect 14700 16884 14756 18508
rect 14812 18450 14868 18620
rect 14812 18398 14814 18450
rect 14866 18398 14868 18450
rect 14812 18386 14868 18398
rect 15036 18452 15092 18462
rect 15036 18358 15092 18396
rect 15148 18004 15204 18732
rect 15372 18562 15428 19068
rect 15820 19010 15876 19022
rect 15820 18958 15822 19010
rect 15874 18958 15876 19010
rect 15820 18564 15876 18958
rect 15372 18510 15374 18562
rect 15426 18510 15428 18562
rect 15372 18498 15428 18510
rect 15484 18508 15876 18564
rect 15148 17556 15204 17948
rect 15260 18228 15316 18238
rect 15484 18228 15540 18508
rect 15932 18452 15988 19740
rect 15260 18226 15540 18228
rect 15260 18174 15262 18226
rect 15314 18174 15540 18226
rect 15260 18172 15540 18174
rect 15708 18396 15988 18452
rect 16044 19236 16100 19246
rect 15260 17892 15316 18172
rect 15260 17826 15316 17836
rect 15596 18116 15652 18126
rect 14812 17500 15204 17556
rect 14812 17106 14868 17500
rect 14812 17054 14814 17106
rect 14866 17054 14868 17106
rect 14812 17042 14868 17054
rect 15148 17108 15204 17500
rect 15596 17554 15652 18060
rect 15596 17502 15598 17554
rect 15650 17502 15652 17554
rect 15596 17490 15652 17502
rect 15372 17108 15428 17118
rect 15148 17106 15428 17108
rect 15148 17054 15374 17106
rect 15426 17054 15428 17106
rect 15148 17052 15428 17054
rect 15372 17042 15428 17052
rect 15036 16996 15092 17006
rect 15036 16902 15092 16940
rect 15148 16884 15204 16894
rect 14700 16828 14868 16884
rect 14700 16660 14756 16670
rect 14700 16324 14756 16604
rect 14812 16548 14868 16828
rect 14812 16492 15092 16548
rect 14924 16324 14980 16334
rect 14700 16322 14980 16324
rect 14700 16270 14926 16322
rect 14978 16270 14980 16322
rect 14700 16268 14980 16270
rect 14924 16258 14980 16268
rect 14588 15874 14644 15886
rect 14588 15822 14590 15874
rect 14642 15822 14644 15874
rect 14476 15540 14532 15550
rect 14476 15446 14532 15484
rect 14028 15092 14308 15148
rect 14028 14530 14084 15092
rect 14588 14756 14644 15822
rect 14924 15428 14980 15438
rect 14924 15334 14980 15372
rect 14028 14478 14030 14530
rect 14082 14478 14084 14530
rect 14028 14466 14084 14478
rect 14252 14700 14644 14756
rect 13692 12786 13748 12796
rect 13804 12852 13860 12862
rect 13916 12852 13972 14252
rect 13804 12850 13972 12852
rect 13804 12798 13806 12850
rect 13858 12798 13972 12850
rect 13804 12796 13972 12798
rect 14028 12852 14084 12862
rect 13804 12786 13860 12796
rect 14028 12758 14084 12796
rect 14028 12292 14084 12302
rect 14028 12198 14084 12236
rect 13468 12068 13524 12078
rect 13468 11974 13524 12012
rect 13244 11554 13300 11564
rect 13692 11394 13748 11406
rect 13692 11342 13694 11394
rect 13746 11342 13748 11394
rect 13468 11172 13524 11182
rect 13244 11170 13524 11172
rect 13244 11118 13470 11170
rect 13522 11118 13524 11170
rect 13244 11116 13524 11118
rect 13244 10722 13300 11116
rect 13468 11106 13524 11116
rect 13244 10670 13246 10722
rect 13298 10670 13300 10722
rect 13244 10658 13300 10670
rect 13692 10050 13748 11342
rect 13692 9998 13694 10050
rect 13746 9998 13748 10050
rect 13692 9986 13748 9998
rect 12796 9828 12852 9838
rect 12684 9826 12852 9828
rect 12684 9774 12798 9826
rect 12850 9774 12852 9826
rect 12684 9772 12852 9774
rect 12572 9716 12628 9726
rect 12572 9622 12628 9660
rect 12236 9266 12404 9268
rect 12236 9214 12238 9266
rect 12290 9214 12404 9266
rect 12236 9212 12404 9214
rect 12236 9202 12292 9212
rect 12796 9154 12852 9772
rect 14028 9828 14084 9838
rect 12796 9102 12798 9154
rect 12850 9102 12852 9154
rect 12796 9090 12852 9102
rect 13356 9156 13412 9166
rect 13356 9062 13412 9100
rect 11564 8990 11566 9042
rect 11618 8990 11620 9042
rect 11564 8978 11620 8990
rect 12572 8818 12628 8830
rect 12572 8766 12574 8818
rect 12626 8766 12628 8818
rect 12572 8428 12628 8766
rect 14028 8428 14084 9772
rect 14252 9714 14308 14700
rect 14476 14532 14532 14542
rect 14476 14530 14644 14532
rect 14476 14478 14478 14530
rect 14530 14478 14644 14530
rect 14476 14476 14644 14478
rect 14476 14466 14532 14476
rect 14364 13188 14420 13198
rect 14588 13188 14644 14476
rect 14700 14308 14756 14318
rect 14700 14214 14756 14252
rect 14700 13188 14756 13198
rect 14588 13186 14756 13188
rect 14588 13134 14702 13186
rect 14754 13134 14756 13186
rect 14588 13132 14756 13134
rect 14364 13094 14420 13132
rect 14700 13122 14756 13132
rect 14476 12404 14532 12414
rect 14476 12290 14532 12348
rect 15036 12402 15092 16492
rect 15148 16098 15204 16828
rect 15148 16046 15150 16098
rect 15202 16046 15204 16098
rect 15148 15540 15204 16046
rect 15484 15876 15540 15886
rect 15484 15874 15652 15876
rect 15484 15822 15486 15874
rect 15538 15822 15652 15874
rect 15484 15820 15652 15822
rect 15484 15810 15540 15820
rect 15484 15540 15540 15550
rect 15148 15538 15540 15540
rect 15148 15486 15486 15538
rect 15538 15486 15540 15538
rect 15148 15484 15540 15486
rect 15484 15474 15540 15484
rect 15148 14308 15204 14318
rect 15148 13858 15204 14252
rect 15148 13806 15150 13858
rect 15202 13806 15204 13858
rect 15148 13794 15204 13806
rect 15596 13860 15652 15820
rect 15708 15148 15764 18396
rect 16044 17780 16100 19180
rect 16156 19236 16212 19246
rect 16492 19236 16548 28588
rect 16604 26514 16660 30156
rect 16828 30146 16884 30156
rect 17500 30146 17556 30156
rect 17948 30212 18004 30222
rect 17948 30098 18004 30156
rect 17948 30046 17950 30098
rect 18002 30046 18004 30098
rect 17948 30034 18004 30046
rect 18172 29652 18228 29662
rect 18284 29652 18340 31054
rect 19068 30996 19124 31006
rect 19628 30996 19684 31948
rect 19740 31938 19796 31948
rect 20076 31666 20132 31678
rect 20076 31614 20078 31666
rect 20130 31614 20132 31666
rect 20076 31556 20132 31614
rect 20076 31490 20132 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19068 30902 19124 30940
rect 19292 30994 19684 30996
rect 19292 30942 19630 30994
rect 19682 30942 19684 30994
rect 19292 30940 19684 30942
rect 19292 30324 19348 30940
rect 19628 30930 19684 30940
rect 20412 30882 20468 30894
rect 20412 30830 20414 30882
rect 20466 30830 20468 30882
rect 19516 30548 19572 30558
rect 19292 30322 19460 30324
rect 19292 30270 19294 30322
rect 19346 30270 19460 30322
rect 19292 30268 19460 30270
rect 19292 30258 19348 30268
rect 18620 30210 18676 30222
rect 18620 30158 18622 30210
rect 18674 30158 18676 30210
rect 18172 29650 18340 29652
rect 18172 29598 18174 29650
rect 18226 29598 18340 29650
rect 18172 29596 18340 29598
rect 18396 29986 18452 29998
rect 18396 29934 18398 29986
rect 18450 29934 18452 29986
rect 18172 29586 18228 29596
rect 18396 29540 18452 29934
rect 18396 29474 18452 29484
rect 18060 29316 18116 29326
rect 16716 28756 16772 28766
rect 16716 28662 16772 28700
rect 16604 26462 16606 26514
rect 16658 26462 16660 26514
rect 16604 26450 16660 26462
rect 17948 26292 18004 26302
rect 17836 26180 17892 26190
rect 17836 26086 17892 26124
rect 17948 24722 18004 26236
rect 17948 24670 17950 24722
rect 18002 24670 18004 24722
rect 17500 24612 17556 24622
rect 17500 24518 17556 24556
rect 17948 23492 18004 24670
rect 17948 23426 18004 23436
rect 18060 23826 18116 29260
rect 18284 29316 18340 29326
rect 18620 29316 18676 30158
rect 18284 29314 18452 29316
rect 18284 29262 18286 29314
rect 18338 29262 18452 29314
rect 18284 29260 18452 29262
rect 18284 29250 18340 29260
rect 18396 27186 18452 29260
rect 18620 29250 18676 29260
rect 18956 29316 19012 29326
rect 18956 29222 19012 29260
rect 19404 28756 19460 30268
rect 19516 29652 19572 30492
rect 20412 30434 20468 30830
rect 20412 30382 20414 30434
rect 20466 30382 20468 30434
rect 20412 30370 20468 30382
rect 19740 30212 19796 30222
rect 19740 30118 19796 30156
rect 20524 30098 20580 33628
rect 20636 33460 20692 34860
rect 20748 34916 20804 34926
rect 20972 34916 21028 34926
rect 20748 34914 20972 34916
rect 20748 34862 20750 34914
rect 20802 34862 20972 34914
rect 20748 34860 20972 34862
rect 20748 34356 20804 34860
rect 20972 34850 21028 34860
rect 20748 34290 20804 34300
rect 20748 33460 20804 33470
rect 20636 33458 20804 33460
rect 20636 33406 20750 33458
rect 20802 33406 20804 33458
rect 20636 33404 20804 33406
rect 20748 33394 20804 33404
rect 21308 33348 21364 35868
rect 21420 35858 21476 35868
rect 21532 35026 21588 36204
rect 21644 35924 21700 39676
rect 21756 39666 21812 39676
rect 21868 40628 21924 40638
rect 21756 39060 21812 39070
rect 21868 39060 21924 40572
rect 21756 39058 21924 39060
rect 21756 39006 21758 39058
rect 21810 39006 21924 39058
rect 21756 39004 21924 39006
rect 21980 40402 22036 40796
rect 22204 40628 22260 41022
rect 22540 41300 22596 41916
rect 22764 41906 22820 41916
rect 22876 41412 22932 41422
rect 22540 41244 22820 41300
rect 22316 40964 22372 40974
rect 22372 40908 22484 40964
rect 22316 40898 22372 40908
rect 22316 40628 22372 40638
rect 22204 40626 22372 40628
rect 22204 40574 22318 40626
rect 22370 40574 22372 40626
rect 22204 40572 22372 40574
rect 22316 40562 22372 40572
rect 21980 40350 21982 40402
rect 22034 40350 22036 40402
rect 21756 38994 21812 39004
rect 21980 38668 22036 40350
rect 22092 40514 22148 40526
rect 22092 40462 22094 40514
rect 22146 40462 22148 40514
rect 22092 40292 22148 40462
rect 22092 40226 22148 40236
rect 22428 39508 22484 40908
rect 22540 40628 22596 41244
rect 22764 41186 22820 41244
rect 22764 41134 22766 41186
rect 22818 41134 22820 41186
rect 22764 41122 22820 41134
rect 22876 41186 22932 41356
rect 22876 41134 22878 41186
rect 22930 41134 22932 41186
rect 22876 41122 22932 41134
rect 22652 41074 22708 41086
rect 22652 41022 22654 41074
rect 22706 41022 22708 41074
rect 22652 40964 22708 41022
rect 22988 40964 23044 42140
rect 23100 41748 23156 41758
rect 23100 41654 23156 41692
rect 22652 40908 23044 40964
rect 23100 41188 23156 41198
rect 23100 40852 23156 41132
rect 22764 40796 23156 40852
rect 22652 40628 22708 40638
rect 22540 40626 22708 40628
rect 22540 40574 22654 40626
rect 22706 40574 22708 40626
rect 22540 40572 22708 40574
rect 22652 40562 22708 40572
rect 22540 40404 22596 40414
rect 22540 40310 22596 40348
rect 22540 39508 22596 39518
rect 22428 39506 22596 39508
rect 22428 39454 22542 39506
rect 22594 39454 22596 39506
rect 22428 39452 22596 39454
rect 22092 39396 22148 39406
rect 22092 38834 22148 39340
rect 22204 39394 22260 39406
rect 22204 39342 22206 39394
rect 22258 39342 22260 39394
rect 22204 39060 22260 39342
rect 22204 38994 22260 39004
rect 22092 38782 22094 38834
rect 22146 38782 22148 38834
rect 22092 38770 22148 38782
rect 22428 38834 22484 39452
rect 22540 39442 22596 39452
rect 22428 38782 22430 38834
rect 22482 38782 22484 38834
rect 22428 38770 22484 38782
rect 22764 38724 22820 40796
rect 23100 40628 23156 40638
rect 22988 39620 23044 39630
rect 21980 38612 22260 38668
rect 22764 38658 22820 38668
rect 22876 38836 22932 38846
rect 21868 37828 21924 37838
rect 21868 37826 22036 37828
rect 21868 37774 21870 37826
rect 21922 37774 22036 37826
rect 21868 37772 22036 37774
rect 21868 37762 21924 37772
rect 21868 37492 21924 37502
rect 21868 36372 21924 37436
rect 21980 37044 22036 37772
rect 21980 36950 22036 36988
rect 22092 37154 22148 37166
rect 22092 37102 22094 37154
rect 22146 37102 22148 37154
rect 21868 36306 21924 36316
rect 21980 36596 22036 36606
rect 21868 35924 21924 35934
rect 21644 35922 21924 35924
rect 21644 35870 21870 35922
rect 21922 35870 21924 35922
rect 21644 35868 21924 35870
rect 21532 34974 21534 35026
rect 21586 34974 21588 35026
rect 21532 34962 21588 34974
rect 21420 34692 21476 34702
rect 21420 34242 21476 34636
rect 21420 34190 21422 34242
rect 21474 34190 21476 34242
rect 21420 34178 21476 34190
rect 21644 33348 21700 33358
rect 21756 33348 21812 35868
rect 21868 35858 21924 35868
rect 21980 35812 22036 36540
rect 22092 36484 22148 37102
rect 22204 36820 22260 38612
rect 22652 38052 22708 38062
rect 22652 37958 22708 37996
rect 22204 36754 22260 36764
rect 22876 37154 22932 38780
rect 22988 38834 23044 39564
rect 22988 38782 22990 38834
rect 23042 38782 23044 38834
rect 22988 38770 23044 38782
rect 22876 37102 22878 37154
rect 22930 37102 22932 37154
rect 22876 36596 22932 37102
rect 22540 36540 22932 36596
rect 22988 37044 23044 37054
rect 22092 36418 22148 36428
rect 22204 36482 22260 36494
rect 22204 36430 22206 36482
rect 22258 36430 22260 36482
rect 22204 35924 22260 36430
rect 22540 36036 22596 36540
rect 22652 36372 22708 36382
rect 22652 36278 22708 36316
rect 22764 36258 22820 36270
rect 22764 36206 22766 36258
rect 22818 36206 22820 36258
rect 22764 36036 22820 36206
rect 22876 36260 22932 36270
rect 22988 36260 23044 36988
rect 22876 36258 23044 36260
rect 22876 36206 22878 36258
rect 22930 36206 23044 36258
rect 22876 36204 23044 36206
rect 22876 36194 22932 36204
rect 22540 35980 22708 36036
rect 22764 35980 23044 36036
rect 22204 35858 22260 35868
rect 21980 35746 22036 35756
rect 22316 35812 22372 35822
rect 22204 35588 22260 35598
rect 21980 35532 22204 35588
rect 21980 34914 22036 35532
rect 22204 35522 22260 35532
rect 22316 35308 22372 35756
rect 22428 35700 22484 35710
rect 22652 35700 22708 35980
rect 22876 35812 22932 35822
rect 22876 35718 22932 35756
rect 22428 35606 22484 35644
rect 22540 35644 22708 35700
rect 22764 35700 22820 35710
rect 21980 34862 21982 34914
rect 22034 34862 22036 34914
rect 21980 34850 22036 34862
rect 22204 35252 22372 35308
rect 21308 33346 21476 33348
rect 21308 33294 21310 33346
rect 21362 33294 21476 33346
rect 21308 33292 21476 33294
rect 21308 33282 21364 33292
rect 20748 32452 20804 32462
rect 20748 32450 21364 32452
rect 20748 32398 20750 32450
rect 20802 32398 21364 32450
rect 20748 32396 21364 32398
rect 20748 32386 20804 32396
rect 20748 32228 20804 32238
rect 20748 30434 20804 32172
rect 20748 30382 20750 30434
rect 20802 30382 20804 30434
rect 20748 30370 20804 30382
rect 21196 30660 21252 30670
rect 21196 30212 21252 30604
rect 21308 30434 21364 32396
rect 21420 30548 21476 33292
rect 21644 33346 21812 33348
rect 21644 33294 21646 33346
rect 21698 33294 21812 33346
rect 21644 33292 21812 33294
rect 21980 34692 22036 34702
rect 21980 34244 22036 34636
rect 21980 33346 22036 34188
rect 21980 33294 21982 33346
rect 22034 33294 22036 33346
rect 21644 33282 21700 33292
rect 21980 33282 22036 33294
rect 22092 34130 22148 34142
rect 22092 34078 22094 34130
rect 22146 34078 22148 34130
rect 22092 33348 22148 34078
rect 22092 33282 22148 33292
rect 21756 33122 21812 33134
rect 21756 33070 21758 33122
rect 21810 33070 21812 33122
rect 21756 32340 21812 33070
rect 22204 32340 22260 35252
rect 21756 32274 21812 32284
rect 22092 32284 22260 32340
rect 22428 35026 22484 35038
rect 22428 34974 22430 35026
rect 22482 34974 22484 35026
rect 21868 31892 21924 31902
rect 21420 30482 21476 30492
rect 21644 31890 21924 31892
rect 21644 31838 21870 31890
rect 21922 31838 21924 31890
rect 21644 31836 21924 31838
rect 21644 30772 21700 31836
rect 21868 31826 21924 31836
rect 21868 31668 21924 31678
rect 21868 31574 21924 31612
rect 21980 31556 22036 31566
rect 21980 31462 22036 31500
rect 21308 30382 21310 30434
rect 21362 30382 21364 30434
rect 21308 30370 21364 30382
rect 21644 30434 21700 30716
rect 21644 30382 21646 30434
rect 21698 30382 21700 30434
rect 21644 30370 21700 30382
rect 21308 30212 21364 30222
rect 21196 30210 21364 30212
rect 21196 30158 21310 30210
rect 21362 30158 21364 30210
rect 21196 30156 21364 30158
rect 22092 30212 22148 32284
rect 22204 32116 22260 32126
rect 22204 31778 22260 32060
rect 22428 31892 22484 34974
rect 22540 34132 22596 35644
rect 22652 34916 22708 34926
rect 22652 34822 22708 34860
rect 22652 34356 22708 34366
rect 22764 34356 22820 35644
rect 22988 34468 23044 35980
rect 23100 34692 23156 40572
rect 23212 38050 23268 43148
rect 23324 42420 23380 43372
rect 23436 42420 23492 42430
rect 23324 42364 23436 42420
rect 23436 42354 23492 42364
rect 23436 41972 23492 41982
rect 23324 41524 23380 41534
rect 23324 41410 23380 41468
rect 23324 41358 23326 41410
rect 23378 41358 23380 41410
rect 23324 41346 23380 41358
rect 23436 40964 23492 41916
rect 23548 41076 23604 43596
rect 23660 41300 23716 48748
rect 23884 47796 23940 47806
rect 23772 47572 23828 47582
rect 23772 46564 23828 47516
rect 23884 47570 23940 47740
rect 23884 47518 23886 47570
rect 23938 47518 23940 47570
rect 23884 47506 23940 47518
rect 23884 46788 23940 46798
rect 23884 46694 23940 46732
rect 23772 46498 23828 46508
rect 23996 45444 24052 48860
rect 24332 48244 24388 48254
rect 24220 48188 24332 48244
rect 24108 47684 24164 47694
rect 24108 47458 24164 47628
rect 24108 47406 24110 47458
rect 24162 47406 24164 47458
rect 24108 47394 24164 47406
rect 24220 47460 24276 48188
rect 24332 48150 24388 48188
rect 24220 47394 24276 47404
rect 24332 48018 24388 48030
rect 24332 47966 24334 48018
rect 24386 47966 24388 48018
rect 24332 47236 24388 47966
rect 24444 47460 24500 50372
rect 24556 49812 24612 49822
rect 24556 49718 24612 49756
rect 24668 48356 24724 48366
rect 24668 48262 24724 48300
rect 24444 47404 24612 47460
rect 24332 47170 24388 47180
rect 24444 47234 24500 47246
rect 24444 47182 24446 47234
rect 24498 47182 24500 47234
rect 24220 47124 24276 47134
rect 24108 46676 24164 46686
rect 24108 45890 24164 46620
rect 24108 45838 24110 45890
rect 24162 45838 24164 45890
rect 24108 45826 24164 45838
rect 23996 45388 24164 45444
rect 23996 45220 24052 45230
rect 23884 44660 23940 44670
rect 23884 44434 23940 44604
rect 23884 44382 23886 44434
rect 23938 44382 23940 44434
rect 23884 44370 23940 44382
rect 23996 44436 24052 45164
rect 23996 44322 24052 44380
rect 23996 44270 23998 44322
rect 24050 44270 24052 44322
rect 23996 44258 24052 44270
rect 23772 44098 23828 44110
rect 23772 44046 23774 44098
rect 23826 44046 23828 44098
rect 23772 43708 23828 44046
rect 24108 43764 24164 45388
rect 24220 44884 24276 47068
rect 24444 46788 24500 47182
rect 24332 46732 24500 46788
rect 24332 46452 24388 46732
rect 24444 46564 24500 46574
rect 24444 46470 24500 46508
rect 24332 46386 24388 46396
rect 24444 46116 24500 46126
rect 24556 46116 24612 47404
rect 24668 47234 24724 47246
rect 24668 47182 24670 47234
rect 24722 47182 24724 47234
rect 24668 47124 24724 47182
rect 24668 47058 24724 47068
rect 24780 47234 24836 47246
rect 24780 47182 24782 47234
rect 24834 47182 24836 47234
rect 24556 46060 24724 46116
rect 24332 46002 24388 46014
rect 24332 45950 24334 46002
rect 24386 45950 24388 46002
rect 24332 45106 24388 45950
rect 24444 45892 24500 46060
rect 24556 45892 24612 45902
rect 24444 45890 24612 45892
rect 24444 45838 24558 45890
rect 24610 45838 24612 45890
rect 24444 45836 24612 45838
rect 24556 45780 24612 45836
rect 24556 45714 24612 45724
rect 24556 45220 24612 45230
rect 24556 45126 24612 45164
rect 24332 45054 24334 45106
rect 24386 45054 24388 45106
rect 24332 45042 24388 45054
rect 24220 44828 24388 44884
rect 23996 43708 24164 43764
rect 24332 43762 24388 44828
rect 24444 44324 24500 44334
rect 24444 44230 24500 44268
rect 24332 43710 24334 43762
rect 24386 43710 24388 43762
rect 23772 43652 23940 43708
rect 23772 43538 23828 43550
rect 23772 43486 23774 43538
rect 23826 43486 23828 43538
rect 23772 42980 23828 43486
rect 23884 43428 23940 43652
rect 23884 43362 23940 43372
rect 23772 42914 23828 42924
rect 23884 42756 23940 42766
rect 23884 42662 23940 42700
rect 23996 42194 24052 43708
rect 24332 43698 24388 43710
rect 24220 43652 24276 43662
rect 24220 43558 24276 43596
rect 24444 43540 24500 43550
rect 24444 43538 24612 43540
rect 24444 43486 24446 43538
rect 24498 43486 24612 43538
rect 24444 43484 24612 43486
rect 24444 43474 24500 43484
rect 24444 43316 24500 43326
rect 24332 43260 24444 43316
rect 24332 42754 24388 43260
rect 24444 43250 24500 43260
rect 24332 42702 24334 42754
rect 24386 42702 24388 42754
rect 24332 42690 24388 42702
rect 24444 42644 24500 42654
rect 24444 42550 24500 42588
rect 23996 42142 23998 42194
rect 24050 42142 24052 42194
rect 23996 42130 24052 42142
rect 24108 42196 24164 42206
rect 24556 42196 24612 43484
rect 24668 42756 24724 46060
rect 24780 44324 24836 47182
rect 25004 47236 25060 47246
rect 25004 47142 25060 47180
rect 25228 45556 25284 50372
rect 27468 49810 27524 50652
rect 27916 50540 28420 50596
rect 27468 49758 27470 49810
rect 27522 49758 27524 49810
rect 27468 49746 27524 49758
rect 27804 50482 27860 50494
rect 27804 50430 27806 50482
rect 27858 50430 27860 50482
rect 26796 49700 26852 49710
rect 26460 49588 26516 49598
rect 26348 49532 26460 49588
rect 26012 49140 26068 49150
rect 26012 49046 26068 49084
rect 25564 49028 25620 49038
rect 25564 48802 25620 48972
rect 25564 48750 25566 48802
rect 25618 48750 25620 48802
rect 25452 48018 25508 48030
rect 25452 47966 25454 48018
rect 25506 47966 25508 48018
rect 25452 47348 25508 47966
rect 25564 47460 25620 48750
rect 26348 48468 26404 49532
rect 26460 49522 26516 49532
rect 26796 49138 26852 49644
rect 26796 49086 26798 49138
rect 26850 49086 26852 49138
rect 26796 49074 26852 49086
rect 27020 49698 27076 49710
rect 27020 49646 27022 49698
rect 27074 49646 27076 49698
rect 27020 49140 27076 49646
rect 27804 49476 27860 50430
rect 27916 50482 27972 50540
rect 27916 50430 27918 50482
rect 27970 50430 27972 50482
rect 27916 50418 27972 50430
rect 28364 50484 28420 50540
rect 29148 50594 29204 52220
rect 29260 51268 29316 53452
rect 30380 53442 30436 53452
rect 30492 52162 30548 53676
rect 30716 53618 30772 53630
rect 30716 53566 30718 53618
rect 30770 53566 30772 53618
rect 30716 53172 30772 53566
rect 30716 53106 30772 53116
rect 30940 52836 30996 52846
rect 31052 52836 31108 54124
rect 31164 53732 31220 53742
rect 32284 53732 32340 54350
rect 32956 54404 33012 55246
rect 33180 54404 33236 54414
rect 32956 54348 33180 54404
rect 31220 53676 31444 53732
rect 31164 53638 31220 53676
rect 31388 53170 31444 53676
rect 33180 53732 33236 54348
rect 33292 53732 33348 53742
rect 33180 53676 33292 53732
rect 32284 53666 32340 53676
rect 31948 53620 32004 53630
rect 31948 53618 32228 53620
rect 31948 53566 31950 53618
rect 32002 53566 32228 53618
rect 31948 53564 32228 53566
rect 31948 53554 32004 53564
rect 31388 53118 31390 53170
rect 31442 53118 31444 53170
rect 31388 53106 31444 53118
rect 32172 53170 32228 53564
rect 32172 53118 32174 53170
rect 32226 53118 32228 53170
rect 32172 53106 32228 53118
rect 32508 53060 32564 53070
rect 32508 52966 32564 53004
rect 30940 52834 31108 52836
rect 30940 52782 30942 52834
rect 30994 52782 31108 52834
rect 30940 52780 31108 52782
rect 30940 52770 30996 52780
rect 30492 52110 30494 52162
rect 30546 52110 30548 52162
rect 30492 52098 30548 52110
rect 31276 52052 31332 52062
rect 31276 51958 31332 51996
rect 33292 52052 33348 53676
rect 33404 52274 33460 55412
rect 33628 55186 33684 55198
rect 33628 55134 33630 55186
rect 33682 55134 33684 55186
rect 33628 53172 33684 55134
rect 34076 53842 34132 55804
rect 34972 55188 35028 59200
rect 35420 57092 35476 59200
rect 35420 57026 35476 57036
rect 35308 56308 35364 56318
rect 35308 56214 35364 56252
rect 36316 56308 36372 59200
rect 36316 56242 36372 56252
rect 36428 56980 36484 56990
rect 35756 56084 35812 56094
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35756 55410 35812 56028
rect 35980 56082 36036 56094
rect 35980 56030 35982 56082
rect 36034 56030 36036 56082
rect 35980 55860 36036 56030
rect 36428 55970 36484 56924
rect 36764 56084 36820 59200
rect 37548 56084 37604 56094
rect 36764 56028 36932 56084
rect 36428 55918 36430 55970
rect 36482 55918 36484 55970
rect 36428 55906 36484 55918
rect 35980 55794 36036 55804
rect 36876 55468 36932 56028
rect 37548 55990 37604 56028
rect 37660 55468 37716 59200
rect 37996 57092 38052 57102
rect 37996 55970 38052 57036
rect 38108 56644 38164 59200
rect 38108 56578 38164 56588
rect 37996 55918 37998 55970
rect 38050 55918 38052 55970
rect 37996 55906 38052 55918
rect 39004 55468 39060 59200
rect 39452 56980 39508 59200
rect 39452 56914 39508 56924
rect 39116 56308 39172 56318
rect 39116 56214 39172 56252
rect 39788 56082 39844 56094
rect 39788 56030 39790 56082
rect 39842 56030 39844 56082
rect 39788 55468 39844 56030
rect 36876 55412 37492 55468
rect 37660 55412 38612 55468
rect 39004 55412 39284 55468
rect 35756 55358 35758 55410
rect 35810 55358 35812 55410
rect 35756 55346 35812 55358
rect 37436 55410 37492 55412
rect 37436 55358 37438 55410
rect 37490 55358 37492 55410
rect 37436 55346 37492 55358
rect 38108 55298 38164 55310
rect 38108 55246 38110 55298
rect 38162 55246 38164 55298
rect 34972 55122 35028 55132
rect 36092 55188 36148 55198
rect 36092 55094 36148 55132
rect 35308 54514 35364 54526
rect 35308 54462 35310 54514
rect 35362 54462 35364 54514
rect 34300 54404 34356 54414
rect 34300 54310 34356 54348
rect 34860 54404 34916 54414
rect 34860 54310 34916 54348
rect 35308 54404 35364 54462
rect 35980 54404 36036 54414
rect 35308 54338 35364 54348
rect 35868 54402 36036 54404
rect 35868 54350 35982 54402
rect 36034 54350 36036 54402
rect 35868 54348 36036 54350
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35196 53844 35252 53854
rect 34076 53790 34078 53842
rect 34130 53790 34132 53842
rect 34076 53778 34132 53790
rect 34300 53842 35252 53844
rect 34300 53790 35198 53842
rect 35250 53790 35252 53842
rect 34300 53788 35252 53790
rect 33852 53172 33908 53182
rect 33628 53170 33908 53172
rect 33628 53118 33854 53170
rect 33906 53118 33908 53170
rect 33628 53116 33908 53118
rect 33852 53106 33908 53116
rect 33964 53058 34020 53070
rect 33964 53006 33966 53058
rect 34018 53006 34020 53058
rect 33852 52388 33908 52398
rect 33964 52388 34020 53006
rect 33852 52386 34020 52388
rect 33852 52334 33854 52386
rect 33906 52334 34020 52386
rect 33852 52332 34020 52334
rect 34188 52948 34244 52958
rect 34300 52948 34356 53788
rect 35196 53778 35252 53788
rect 34636 53620 34692 53630
rect 34524 53618 34692 53620
rect 34524 53566 34638 53618
rect 34690 53566 34692 53618
rect 34524 53564 34692 53566
rect 34188 52946 34356 52948
rect 34188 52894 34190 52946
rect 34242 52894 34356 52946
rect 34188 52892 34356 52894
rect 34412 52948 34468 52958
rect 34524 52948 34580 53564
rect 34636 53554 34692 53564
rect 35532 53620 35588 53630
rect 35532 53618 35812 53620
rect 35532 53566 35534 53618
rect 35586 53566 35812 53618
rect 35532 53564 35812 53566
rect 35532 53554 35588 53564
rect 34748 53506 34804 53518
rect 34748 53454 34750 53506
rect 34802 53454 34804 53506
rect 34748 53284 34804 53454
rect 34972 53508 35028 53518
rect 35308 53508 35364 53518
rect 34972 53506 35252 53508
rect 34972 53454 34974 53506
rect 35026 53454 35252 53506
rect 34972 53452 35252 53454
rect 34972 53442 35028 53452
rect 34748 53218 34804 53228
rect 34636 53172 34692 53182
rect 34636 53078 34692 53116
rect 35196 53060 35252 53452
rect 35308 53414 35364 53452
rect 35196 53004 35588 53060
rect 34412 52946 34580 52948
rect 34412 52894 34414 52946
rect 34466 52894 34580 52946
rect 34412 52892 34580 52894
rect 35532 52948 35588 53004
rect 35756 52948 35812 53564
rect 35868 53618 35924 54348
rect 35980 54338 36036 54348
rect 38108 54402 38164 55246
rect 38556 55186 38612 55412
rect 38556 55134 38558 55186
rect 38610 55134 38612 55186
rect 38556 55122 38612 55134
rect 39228 54738 39284 55412
rect 39340 55412 39844 55468
rect 39900 55468 39956 59200
rect 40348 56868 40404 59200
rect 40348 56802 40404 56812
rect 40348 56644 40404 56654
rect 40348 55970 40404 56588
rect 40348 55918 40350 55970
rect 40402 55918 40404 55970
rect 40348 55906 40404 55918
rect 40796 55468 40852 59200
rect 41692 57092 41748 59200
rect 41692 57026 41748 57036
rect 42028 56980 42084 56990
rect 42028 55970 42084 56924
rect 42140 56308 42196 59200
rect 42140 56242 42196 56252
rect 42924 56868 42980 56878
rect 42028 55918 42030 55970
rect 42082 55918 42084 55970
rect 42028 55906 42084 55918
rect 42476 56082 42532 56094
rect 42476 56030 42478 56082
rect 42530 56030 42532 56082
rect 39900 55412 40516 55468
rect 40796 55412 41636 55468
rect 39340 55410 39396 55412
rect 39340 55358 39342 55410
rect 39394 55358 39396 55410
rect 39340 55346 39396 55358
rect 39228 54686 39230 54738
rect 39282 54686 39284 54738
rect 39228 54674 39284 54686
rect 40460 54740 40516 55412
rect 41468 55188 41524 55198
rect 41468 55094 41524 55132
rect 40460 54738 40964 54740
rect 40460 54686 40462 54738
rect 40514 54686 40964 54738
rect 40460 54684 40964 54686
rect 40460 54674 40516 54684
rect 40908 54626 40964 54684
rect 41580 54738 41636 55412
rect 41580 54686 41582 54738
rect 41634 54686 41636 54738
rect 41580 54674 41636 54686
rect 42140 55298 42196 55310
rect 42140 55246 42142 55298
rect 42194 55246 42196 55298
rect 40908 54574 40910 54626
rect 40962 54574 40964 54626
rect 40908 54562 40964 54574
rect 41244 54626 41300 54638
rect 41244 54574 41246 54626
rect 41298 54574 41300 54626
rect 38108 54350 38110 54402
rect 38162 54350 38164 54402
rect 38108 54338 38164 54350
rect 38668 53844 38724 53854
rect 38668 53750 38724 53788
rect 38892 53730 38948 53742
rect 38892 53678 38894 53730
rect 38946 53678 38948 53730
rect 35868 53566 35870 53618
rect 35922 53566 35924 53618
rect 35868 53554 35924 53566
rect 36204 53620 36260 53630
rect 36204 53618 36820 53620
rect 36204 53566 36206 53618
rect 36258 53566 36820 53618
rect 36204 53564 36820 53566
rect 36204 53554 36260 53564
rect 36764 53170 36820 53564
rect 38668 53618 38724 53630
rect 38668 53566 38670 53618
rect 38722 53566 38724 53618
rect 36764 53118 36766 53170
rect 36818 53118 36820 53170
rect 36764 53106 36820 53118
rect 38108 53508 38164 53518
rect 38444 53508 38500 53518
rect 37212 53060 37268 53070
rect 37212 52966 37268 53004
rect 35868 52948 35924 52958
rect 35756 52946 35924 52948
rect 35756 52894 35870 52946
rect 35922 52894 35924 52946
rect 35756 52892 35924 52894
rect 33852 52322 33908 52332
rect 34188 52276 34244 52892
rect 33404 52222 33406 52274
rect 33458 52222 33460 52274
rect 33404 52210 33460 52222
rect 33964 52220 34244 52276
rect 34300 52386 34356 52398
rect 34300 52334 34302 52386
rect 34354 52334 34356 52386
rect 33852 52164 33908 52174
rect 33516 52162 33908 52164
rect 33516 52110 33854 52162
rect 33906 52110 33908 52162
rect 33516 52108 33908 52110
rect 33516 52052 33572 52108
rect 33852 52098 33908 52108
rect 33292 51996 33572 52052
rect 29260 51202 29316 51212
rect 32060 50708 32116 50718
rect 29148 50542 29150 50594
rect 29202 50542 29204 50594
rect 29148 50530 29204 50542
rect 31836 50706 32116 50708
rect 31836 50654 32062 50706
rect 32114 50654 32116 50706
rect 31836 50652 32116 50654
rect 28476 50484 28532 50494
rect 28364 50482 28532 50484
rect 28364 50430 28478 50482
rect 28530 50430 28532 50482
rect 28364 50428 28532 50430
rect 28140 50370 28196 50382
rect 28140 50318 28142 50370
rect 28194 50318 28196 50370
rect 28140 49924 28196 50318
rect 28140 49858 28196 49868
rect 28252 50370 28308 50382
rect 28252 50318 28254 50370
rect 28306 50318 28308 50370
rect 28140 49700 28196 49710
rect 28140 49606 28196 49644
rect 26684 48916 26740 48926
rect 26684 48822 26740 48860
rect 25788 48466 26404 48468
rect 25788 48414 26350 48466
rect 26402 48414 26404 48466
rect 25788 48412 26404 48414
rect 25788 48356 25844 48412
rect 26348 48402 26404 48412
rect 26460 48802 26516 48814
rect 26460 48750 26462 48802
rect 26514 48750 26516 48802
rect 25788 48242 25844 48300
rect 25788 48190 25790 48242
rect 25842 48190 25844 48242
rect 25788 48178 25844 48190
rect 26012 48244 26068 48254
rect 26012 48150 26068 48188
rect 26460 47684 26516 48750
rect 26908 48802 26964 48814
rect 26908 48750 26910 48802
rect 26962 48750 26964 48802
rect 26684 48354 26740 48366
rect 26684 48302 26686 48354
rect 26738 48302 26740 48354
rect 26460 47618 26516 47628
rect 26572 47796 26628 47806
rect 25564 47404 25956 47460
rect 25452 47292 25844 47348
rect 25340 47236 25396 47246
rect 25340 47234 25508 47236
rect 25340 47182 25342 47234
rect 25394 47182 25508 47234
rect 25340 47180 25508 47182
rect 25340 47170 25396 47180
rect 25452 47124 25508 47180
rect 25340 47012 25508 47068
rect 25788 47234 25844 47292
rect 25788 47182 25790 47234
rect 25842 47182 25844 47234
rect 25676 47012 25732 47022
rect 25340 46788 25396 47012
rect 25340 46722 25396 46732
rect 25676 46674 25732 46956
rect 25676 46622 25678 46674
rect 25730 46622 25732 46674
rect 25676 46610 25732 46622
rect 25788 46676 25844 47182
rect 25788 46610 25844 46620
rect 25340 46562 25396 46574
rect 25340 46510 25342 46562
rect 25394 46510 25396 46562
rect 25340 46452 25396 46510
rect 25340 46386 25396 46396
rect 25900 45892 25956 47404
rect 26124 47234 26180 47246
rect 26572 47236 26628 47740
rect 26684 47348 26740 48302
rect 26908 48244 26964 48750
rect 27020 48356 27076 49084
rect 27468 49420 27860 49476
rect 27356 49028 27412 49038
rect 27356 48934 27412 48972
rect 27244 48916 27300 48926
rect 27244 48822 27300 48860
rect 27468 48692 27524 49420
rect 28252 49364 28308 50318
rect 27692 49308 28308 49364
rect 27580 49140 27636 49150
rect 27580 49026 27636 49084
rect 27580 48974 27582 49026
rect 27634 48974 27636 49026
rect 27580 48962 27636 48974
rect 27468 48626 27524 48636
rect 27468 48468 27524 48478
rect 27244 48466 27524 48468
rect 27244 48414 27470 48466
rect 27522 48414 27524 48466
rect 27244 48412 27524 48414
rect 27132 48356 27188 48366
rect 27020 48354 27188 48356
rect 27020 48302 27134 48354
rect 27186 48302 27188 48354
rect 27020 48300 27188 48302
rect 27132 48290 27188 48300
rect 26908 48188 27076 48244
rect 27020 48132 27076 48188
rect 27244 48132 27300 48412
rect 27468 48402 27524 48412
rect 27580 48468 27636 48478
rect 27692 48468 27748 49308
rect 28364 49028 28420 50428
rect 28476 50418 28532 50428
rect 28588 50484 28644 50494
rect 29932 50484 29988 50494
rect 28588 50482 28980 50484
rect 28588 50430 28590 50482
rect 28642 50430 28980 50482
rect 28588 50428 28980 50430
rect 29596 50482 29988 50484
rect 29596 50430 29934 50482
rect 29986 50430 29988 50482
rect 29596 50428 29988 50430
rect 28588 50418 28644 50428
rect 28924 50372 29316 50428
rect 29036 49924 29092 49934
rect 27580 48466 27748 48468
rect 27580 48414 27582 48466
rect 27634 48414 27748 48466
rect 27580 48412 27748 48414
rect 27804 48692 27860 48702
rect 27580 48402 27636 48412
rect 27020 48076 27300 48132
rect 27356 48242 27412 48254
rect 27356 48190 27358 48242
rect 27410 48190 27412 48242
rect 26684 47282 26740 47292
rect 26124 47182 26126 47234
rect 26178 47182 26180 47234
rect 26124 46788 26180 47182
rect 26124 46722 26180 46732
rect 26348 47234 26628 47236
rect 26348 47182 26574 47234
rect 26626 47182 26628 47234
rect 26348 47180 26628 47182
rect 26348 47012 26404 47180
rect 26572 47170 26628 47180
rect 27132 47234 27188 47246
rect 27132 47182 27134 47234
rect 27186 47182 27188 47234
rect 26236 46562 26292 46574
rect 26236 46510 26238 46562
rect 26290 46510 26292 46562
rect 26124 46452 26180 46462
rect 26124 46114 26180 46396
rect 26124 46062 26126 46114
rect 26178 46062 26180 46114
rect 26124 46050 26180 46062
rect 25900 45836 26180 45892
rect 25228 45490 25284 45500
rect 25228 45218 25284 45230
rect 25228 45166 25230 45218
rect 25282 45166 25284 45218
rect 24780 44258 24836 44268
rect 25004 44436 25060 44446
rect 25228 44436 25284 45166
rect 25060 44380 25284 44436
rect 25564 45106 25620 45118
rect 25564 45054 25566 45106
rect 25618 45054 25620 45106
rect 25004 44322 25060 44380
rect 25004 44270 25006 44322
rect 25058 44270 25060 44322
rect 25004 44258 25060 44270
rect 25452 44210 25508 44222
rect 25452 44158 25454 44210
rect 25506 44158 25508 44210
rect 24780 44098 24836 44110
rect 24780 44046 24782 44098
rect 24834 44046 24836 44098
rect 24780 43540 24836 44046
rect 24892 44098 24948 44110
rect 24892 44046 24894 44098
rect 24946 44046 24948 44098
rect 24892 43652 24948 44046
rect 25452 43876 25508 44158
rect 25452 43810 25508 43820
rect 24892 43586 24948 43596
rect 25340 43650 25396 43662
rect 25340 43598 25342 43650
rect 25394 43598 25396 43650
rect 24780 43474 24836 43484
rect 25116 43092 25172 43102
rect 25116 42756 25172 43036
rect 25340 42980 25396 43598
rect 25564 43316 25620 45054
rect 26012 45106 26068 45118
rect 26012 45054 26014 45106
rect 26066 45054 26068 45106
rect 26012 44884 26068 45054
rect 26124 44884 26180 45836
rect 26236 45108 26292 46510
rect 26348 45778 26404 46956
rect 26796 47124 26852 47134
rect 26796 46898 26852 47068
rect 26796 46846 26798 46898
rect 26850 46846 26852 46898
rect 26796 46834 26852 46846
rect 27132 47012 27188 47182
rect 27356 47124 27412 48190
rect 27692 48242 27748 48254
rect 27692 48190 27694 48242
rect 27746 48190 27748 48242
rect 27356 47058 27412 47068
rect 27580 47458 27636 47470
rect 27580 47406 27582 47458
rect 27634 47406 27636 47458
rect 26572 46788 26628 46798
rect 26460 46674 26516 46686
rect 26460 46622 26462 46674
rect 26514 46622 26516 46674
rect 26460 46002 26516 46622
rect 26572 46452 26628 46732
rect 27020 46786 27076 46798
rect 27020 46734 27022 46786
rect 27074 46734 27076 46786
rect 26572 46386 26628 46396
rect 26684 46564 26740 46574
rect 26460 45950 26462 46002
rect 26514 45950 26516 46002
rect 26460 45892 26516 45950
rect 26460 45826 26516 45836
rect 26684 45890 26740 46508
rect 27020 46564 27076 46734
rect 27132 46676 27188 46956
rect 27580 46898 27636 47406
rect 27692 47124 27748 48190
rect 27804 47684 27860 48636
rect 28140 48130 28196 48142
rect 28140 48078 28142 48130
rect 28194 48078 28196 48130
rect 28140 48020 28196 48078
rect 28252 48132 28308 48142
rect 28252 48038 28308 48076
rect 27804 47628 28084 47684
rect 27916 47458 27972 47470
rect 27916 47406 27918 47458
rect 27970 47406 27972 47458
rect 27692 47058 27748 47068
rect 27804 47234 27860 47246
rect 27804 47182 27806 47234
rect 27858 47182 27860 47234
rect 27580 46846 27582 46898
rect 27634 46846 27636 46898
rect 27580 46834 27636 46846
rect 27356 46676 27412 46686
rect 27132 46674 27412 46676
rect 27132 46622 27358 46674
rect 27410 46622 27412 46674
rect 27132 46620 27412 46622
rect 27356 46610 27412 46620
rect 27020 46498 27076 46508
rect 27132 46450 27188 46462
rect 27132 46398 27134 46450
rect 27186 46398 27188 46450
rect 27132 46116 27188 46398
rect 27132 46050 27188 46060
rect 27244 46452 27300 46462
rect 27132 45892 27188 45902
rect 27244 45892 27300 46396
rect 27692 46452 27748 46462
rect 27692 46358 27748 46396
rect 27804 46228 27860 47182
rect 27804 46162 27860 46172
rect 26684 45838 26686 45890
rect 26738 45838 26740 45890
rect 26348 45726 26350 45778
rect 26402 45726 26404 45778
rect 26348 45714 26404 45726
rect 26236 45042 26292 45052
rect 26348 44994 26404 45006
rect 26348 44942 26350 44994
rect 26402 44942 26404 44994
rect 26348 44884 26404 44942
rect 26124 44828 26404 44884
rect 26012 44818 26068 44828
rect 25788 44436 25844 44446
rect 25788 44322 25844 44380
rect 25788 44270 25790 44322
rect 25842 44270 25844 44322
rect 25788 44258 25844 44270
rect 26348 44100 26404 44828
rect 26236 44044 26404 44100
rect 26572 44322 26628 44334
rect 26572 44270 26574 44322
rect 26626 44270 26628 44322
rect 26572 44100 26628 44270
rect 26012 43876 26068 43886
rect 25676 43540 25732 43550
rect 25676 43446 25732 43484
rect 25620 43260 25732 43316
rect 25564 43250 25620 43260
rect 25340 42924 25508 42980
rect 25340 42756 25396 42766
rect 25116 42700 25284 42756
rect 24668 42690 24724 42700
rect 25228 42642 25284 42700
rect 25228 42590 25230 42642
rect 25282 42590 25284 42642
rect 25228 42578 25284 42590
rect 25452 42756 25508 42924
rect 25564 42756 25620 42766
rect 25452 42754 25620 42756
rect 25452 42702 25566 42754
rect 25618 42702 25620 42754
rect 25452 42700 25620 42702
rect 25340 42642 25396 42700
rect 25564 42690 25620 42700
rect 25340 42590 25342 42642
rect 25394 42590 25396 42642
rect 25340 42578 25396 42590
rect 25676 42644 25732 43260
rect 26012 42980 26068 43820
rect 26012 42914 26068 42924
rect 26124 43538 26180 43550
rect 26124 43486 26126 43538
rect 26178 43486 26180 43538
rect 25788 42644 25844 42654
rect 25676 42642 25844 42644
rect 25676 42590 25790 42642
rect 25842 42590 25844 42642
rect 25676 42588 25844 42590
rect 25788 42578 25844 42588
rect 26124 42644 26180 43486
rect 26236 42868 26292 44044
rect 26572 44034 26628 44044
rect 26348 43876 26404 43886
rect 26348 43650 26404 43820
rect 26348 43598 26350 43650
rect 26402 43598 26404 43650
rect 26348 43586 26404 43598
rect 26684 43540 26740 45838
rect 26796 45890 27300 45892
rect 26796 45838 27134 45890
rect 27186 45838 27300 45890
rect 26796 45836 27300 45838
rect 27356 45892 27412 45902
rect 26796 45220 26852 45836
rect 27132 45826 27188 45836
rect 27356 45798 27412 45836
rect 27804 45892 27860 45902
rect 27804 45798 27860 45836
rect 27916 45780 27972 47406
rect 28028 47236 28084 47628
rect 28140 47572 28196 47964
rect 28140 47506 28196 47516
rect 28252 47460 28308 47470
rect 28364 47460 28420 48972
rect 28252 47458 28420 47460
rect 28252 47406 28254 47458
rect 28306 47406 28420 47458
rect 28252 47404 28420 47406
rect 28476 49026 28532 49038
rect 28476 48974 28478 49026
rect 28530 48974 28532 49026
rect 28476 47908 28532 48974
rect 29036 49026 29092 49868
rect 29036 48974 29038 49026
rect 29090 48974 29092 49026
rect 29036 48962 29092 48974
rect 29148 49252 29204 49262
rect 28924 48916 28980 48926
rect 28700 48580 28756 48590
rect 28700 48466 28756 48524
rect 28700 48414 28702 48466
rect 28754 48414 28756 48466
rect 28700 48356 28756 48414
rect 28812 48468 28868 48478
rect 28924 48468 28980 48860
rect 28812 48466 28980 48468
rect 28812 48414 28814 48466
rect 28866 48414 28980 48466
rect 28812 48412 28980 48414
rect 28812 48402 28868 48412
rect 28700 48290 28756 48300
rect 28924 48242 28980 48254
rect 28924 48190 28926 48242
rect 28978 48190 28980 48242
rect 28924 47908 28980 48190
rect 29036 48242 29092 48254
rect 29036 48190 29038 48242
rect 29090 48190 29092 48242
rect 29036 48132 29092 48190
rect 29036 48066 29092 48076
rect 28476 47852 28980 47908
rect 28252 47394 28308 47404
rect 28140 47236 28196 47246
rect 28028 47180 28140 47236
rect 28140 46564 28196 47180
rect 28252 46900 28308 46910
rect 28476 46900 28532 47852
rect 28812 47572 28868 47582
rect 29148 47572 29204 49196
rect 29260 47908 29316 50372
rect 29596 49138 29652 50428
rect 29932 50418 29988 50428
rect 31836 50148 31892 50652
rect 32060 50642 32116 50652
rect 31164 50092 31892 50148
rect 31164 49922 31220 50092
rect 31164 49870 31166 49922
rect 31218 49870 31220 49922
rect 31164 49858 31220 49870
rect 31500 49922 31556 49934
rect 31500 49870 31502 49922
rect 31554 49870 31556 49922
rect 30940 49812 30996 49822
rect 30492 49810 30996 49812
rect 30492 49758 30942 49810
rect 30994 49758 30996 49810
rect 30492 49756 30996 49758
rect 29596 49086 29598 49138
rect 29650 49086 29652 49138
rect 29596 49074 29652 49086
rect 30268 49700 30324 49710
rect 30492 49700 30548 49756
rect 30940 49746 30996 49756
rect 30268 49698 30548 49700
rect 30268 49646 30270 49698
rect 30322 49646 30548 49698
rect 30268 49644 30548 49646
rect 29484 49028 29540 49038
rect 29484 48934 29540 48972
rect 30044 49028 30100 49038
rect 30044 48914 30100 48972
rect 30044 48862 30046 48914
rect 30098 48862 30100 48914
rect 30044 48850 30100 48862
rect 29372 48804 29428 48814
rect 29372 48242 29428 48748
rect 29708 48804 29764 48814
rect 29708 48710 29764 48748
rect 30268 48356 30324 49644
rect 30604 49588 30660 49598
rect 30604 49494 30660 49532
rect 31500 49364 31556 49870
rect 31836 49922 31892 50092
rect 31836 49870 31838 49922
rect 31890 49870 31892 49922
rect 31836 49858 31892 49870
rect 32508 50370 32564 50382
rect 32508 50318 32510 50370
rect 32562 50318 32564 50370
rect 30604 49308 31556 49364
rect 32284 49700 32340 49710
rect 32508 49700 32564 50318
rect 32284 49698 32564 49700
rect 32284 49646 32286 49698
rect 32338 49646 32564 49698
rect 32284 49644 32564 49646
rect 33180 49700 33236 49710
rect 33292 49700 33348 51996
rect 33628 51828 33684 51838
rect 33516 51492 33572 51502
rect 33516 50594 33572 51436
rect 33628 50818 33684 51772
rect 33852 51492 33908 51502
rect 33852 51398 33908 51436
rect 33740 51268 33796 51278
rect 33740 51174 33796 51212
rect 33964 51156 34020 52220
rect 34300 51940 34356 52334
rect 34300 51874 34356 51884
rect 34412 51604 34468 52892
rect 35532 52854 35588 52892
rect 35084 52836 35140 52846
rect 35084 52742 35140 52780
rect 34860 52724 34916 52734
rect 34412 51538 34468 51548
rect 34524 52274 34580 52286
rect 34524 52222 34526 52274
rect 34578 52222 34580 52274
rect 34524 51490 34580 52222
rect 34860 52162 34916 52668
rect 35308 52724 35364 52762
rect 35308 52658 35364 52668
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35644 52500 35700 52510
rect 34860 52110 34862 52162
rect 34914 52110 34916 52162
rect 34524 51438 34526 51490
rect 34578 51438 34580 51490
rect 34524 51426 34580 51438
rect 34636 51938 34692 51950
rect 34636 51886 34638 51938
rect 34690 51886 34692 51938
rect 33628 50766 33630 50818
rect 33682 50766 33684 50818
rect 33628 50754 33684 50766
rect 33852 51100 34020 51156
rect 34076 51378 34132 51390
rect 34076 51326 34078 51378
rect 34130 51326 34132 51378
rect 33516 50542 33518 50594
rect 33570 50542 33572 50594
rect 33516 50530 33572 50542
rect 33740 50596 33796 50606
rect 33852 50596 33908 51100
rect 34076 50708 34132 51326
rect 34300 51378 34356 51390
rect 34300 51326 34302 51378
rect 34354 51326 34356 51378
rect 34300 51268 34356 51326
rect 33740 50594 33908 50596
rect 33740 50542 33742 50594
rect 33794 50542 33908 50594
rect 33740 50540 33908 50542
rect 33964 50652 34132 50708
rect 34188 51212 34300 51268
rect 33740 50530 33796 50540
rect 33964 50484 34020 50652
rect 34188 50594 34244 51212
rect 34300 51202 34356 51212
rect 34636 50820 34692 51886
rect 34860 51602 34916 52110
rect 35532 51940 35588 51950
rect 35644 51940 35700 52444
rect 35868 52274 35924 52892
rect 36092 52948 36148 52958
rect 36092 52854 36148 52892
rect 38108 52948 38164 53452
rect 38332 53506 38500 53508
rect 38332 53454 38446 53506
rect 38498 53454 38500 53506
rect 38332 53452 38500 53454
rect 38668 53508 38724 53566
rect 38780 53508 38836 53518
rect 38668 53452 38780 53508
rect 38108 52946 38276 52948
rect 38108 52894 38110 52946
rect 38162 52894 38276 52946
rect 38108 52892 38276 52894
rect 38108 52882 38164 52892
rect 36316 52722 36372 52734
rect 36316 52670 36318 52722
rect 36370 52670 36372 52722
rect 35868 52222 35870 52274
rect 35922 52222 35924 52274
rect 35868 52210 35924 52222
rect 35980 52388 36036 52398
rect 35980 52050 36036 52332
rect 35980 51998 35982 52050
rect 36034 51998 36036 52050
rect 35980 51986 36036 51998
rect 35532 51938 35700 51940
rect 35532 51886 35534 51938
rect 35586 51886 35700 51938
rect 35532 51884 35700 51886
rect 35532 51874 35588 51884
rect 34860 51550 34862 51602
rect 34914 51550 34916 51602
rect 34860 51538 34916 51550
rect 35532 51716 35588 51726
rect 35532 51490 35588 51660
rect 35532 51438 35534 51490
rect 35586 51438 35588 51490
rect 35532 51426 35588 51438
rect 35644 51492 35700 51884
rect 35756 51938 35812 51950
rect 35756 51886 35758 51938
rect 35810 51886 35812 51938
rect 35756 51716 35812 51886
rect 36316 51940 36372 52670
rect 37660 52724 37716 52734
rect 37660 52630 37716 52668
rect 37884 52722 37940 52734
rect 37884 52670 37886 52722
rect 37938 52670 37940 52722
rect 37660 52388 37716 52398
rect 37660 52162 37716 52332
rect 37884 52276 37940 52670
rect 37884 52210 37940 52220
rect 37660 52110 37662 52162
rect 37714 52110 37716 52162
rect 37660 52098 37716 52110
rect 37996 52052 38052 52062
rect 37996 51958 38052 51996
rect 36316 51884 37044 51940
rect 35756 51650 35812 51660
rect 36092 51828 36148 51838
rect 35980 51604 36036 51614
rect 35980 51510 36036 51548
rect 36092 51602 36148 51772
rect 36092 51550 36094 51602
rect 36146 51550 36148 51602
rect 35756 51492 35812 51502
rect 35644 51490 35812 51492
rect 35644 51438 35758 51490
rect 35810 51438 35812 51490
rect 35644 51436 35812 51438
rect 35756 51426 35812 51436
rect 34860 51380 34916 51390
rect 34860 50932 34916 51324
rect 35196 51380 35252 51390
rect 36092 51380 36148 51550
rect 34972 51156 35028 51166
rect 35196 51156 35252 51324
rect 35868 51324 36148 51380
rect 36316 51380 36372 51418
rect 35868 51268 35924 51324
rect 36316 51314 36372 51324
rect 36540 51378 36596 51390
rect 36764 51380 36820 51390
rect 36540 51326 36542 51378
rect 36594 51326 36596 51378
rect 34972 51062 35028 51100
rect 35084 51154 35252 51156
rect 35084 51102 35198 51154
rect 35250 51102 35252 51154
rect 35084 51100 35252 51102
rect 34860 50876 35028 50932
rect 34636 50754 34692 50764
rect 34188 50542 34190 50594
rect 34242 50542 34244 50594
rect 34188 50530 34244 50542
rect 34748 50596 34804 50606
rect 34748 50502 34804 50540
rect 34412 50484 34468 50494
rect 33964 50482 34132 50484
rect 33964 50430 33966 50482
rect 34018 50430 34132 50482
rect 33964 50428 34132 50430
rect 34300 50482 34468 50484
rect 34300 50430 34414 50482
rect 34466 50430 34468 50482
rect 34300 50428 34468 50430
rect 33964 50418 34020 50428
rect 34076 50372 34356 50428
rect 34412 50418 34468 50428
rect 33180 49698 33348 49700
rect 33180 49646 33182 49698
rect 33234 49646 33348 49698
rect 33180 49644 33348 49646
rect 29372 48190 29374 48242
rect 29426 48190 29428 48242
rect 29372 48178 29428 48190
rect 30044 48244 30100 48254
rect 30268 48244 30324 48300
rect 30044 48242 30324 48244
rect 30044 48190 30046 48242
rect 30098 48190 30324 48242
rect 30044 48188 30324 48190
rect 30380 48804 30436 48814
rect 30604 48804 30660 49308
rect 31164 49138 31220 49150
rect 31164 49086 31166 49138
rect 31218 49086 31220 49138
rect 30828 48914 30884 48926
rect 30828 48862 30830 48914
rect 30882 48862 30884 48914
rect 30380 48802 30660 48804
rect 30380 48750 30382 48802
rect 30434 48750 30660 48802
rect 30380 48748 30660 48750
rect 30716 48802 30772 48814
rect 30716 48750 30718 48802
rect 30770 48750 30772 48802
rect 30380 48242 30436 48748
rect 30716 48580 30772 48750
rect 30716 48514 30772 48524
rect 30604 48356 30660 48366
rect 30828 48356 30884 48862
rect 30604 48354 31108 48356
rect 30604 48302 30606 48354
rect 30658 48302 31108 48354
rect 30604 48300 31108 48302
rect 30604 48290 30660 48300
rect 30380 48190 30382 48242
rect 30434 48190 30436 48242
rect 29596 48018 29652 48030
rect 29596 47966 29598 48018
rect 29650 47966 29652 48018
rect 29260 47852 29428 47908
rect 29260 47684 29316 47694
rect 29260 47590 29316 47628
rect 28252 46898 28532 46900
rect 28252 46846 28254 46898
rect 28306 46846 28532 46898
rect 28252 46844 28532 46846
rect 28700 46900 28756 46910
rect 28252 46834 28308 46844
rect 28700 46806 28756 46844
rect 28812 46786 28868 47516
rect 28812 46734 28814 46786
rect 28866 46734 28868 46786
rect 28812 46722 28868 46734
rect 28924 47516 29204 47572
rect 28028 46562 28196 46564
rect 28028 46510 28142 46562
rect 28194 46510 28196 46562
rect 28028 46508 28196 46510
rect 28028 46004 28084 46508
rect 28140 46498 28196 46508
rect 28476 46674 28532 46686
rect 28476 46622 28478 46674
rect 28530 46622 28532 46674
rect 28028 45938 28084 45948
rect 28140 46116 28196 46126
rect 27916 45714 27972 45724
rect 27132 45668 27188 45678
rect 27020 45444 27076 45454
rect 26796 45126 26852 45164
rect 26908 45388 27020 45444
rect 26908 44322 26964 45388
rect 27020 45378 27076 45388
rect 27132 45106 27188 45612
rect 27244 45668 27300 45678
rect 27692 45668 27748 45678
rect 27244 45666 27412 45668
rect 27244 45614 27246 45666
rect 27298 45614 27412 45666
rect 27244 45612 27412 45614
rect 27244 45602 27300 45612
rect 27132 45054 27134 45106
rect 27186 45054 27188 45106
rect 27132 45042 27188 45054
rect 27244 44996 27300 45006
rect 27244 44902 27300 44940
rect 27356 44436 27412 45612
rect 27468 45666 27748 45668
rect 27468 45614 27694 45666
rect 27746 45614 27748 45666
rect 27468 45612 27748 45614
rect 27468 45106 27524 45612
rect 27692 45602 27748 45612
rect 28140 45444 28196 46060
rect 28476 45892 28532 46622
rect 28476 45826 28532 45836
rect 28364 45668 28420 45678
rect 28364 45666 28532 45668
rect 28364 45614 28366 45666
rect 28418 45614 28532 45666
rect 28364 45612 28532 45614
rect 28364 45602 28420 45612
rect 28364 45444 28420 45454
rect 28140 45388 28308 45444
rect 27916 45220 27972 45230
rect 27468 45054 27470 45106
rect 27522 45054 27524 45106
rect 27468 45042 27524 45054
rect 27692 45108 27748 45118
rect 27692 45014 27748 45052
rect 27916 45106 27972 45164
rect 27916 45054 27918 45106
rect 27970 45054 27972 45106
rect 27916 45042 27972 45054
rect 28140 45220 28196 45230
rect 27356 44370 27412 44380
rect 28140 44994 28196 45164
rect 28140 44942 28142 44994
rect 28194 44942 28196 44994
rect 26908 44270 26910 44322
rect 26962 44270 26964 44322
rect 26908 44258 26964 44270
rect 26684 43474 26740 43484
rect 27020 44212 27076 44222
rect 27020 43538 27076 44156
rect 27356 44212 27412 44222
rect 27356 44118 27412 44156
rect 27020 43486 27022 43538
rect 27074 43486 27076 43538
rect 27020 43474 27076 43486
rect 27132 44098 27188 44110
rect 27804 44100 27860 44110
rect 27132 44046 27134 44098
rect 27186 44046 27188 44098
rect 26796 42980 26852 42990
rect 26348 42868 26404 42878
rect 26236 42812 26348 42868
rect 26348 42802 26404 42812
rect 26124 42578 26180 42588
rect 25900 42530 25956 42542
rect 25900 42478 25902 42530
rect 25954 42478 25956 42530
rect 24108 42102 24164 42140
rect 24444 42140 24612 42196
rect 25228 42420 25284 42430
rect 24332 42084 24388 42094
rect 23884 41970 23940 41982
rect 23884 41918 23886 41970
rect 23938 41918 23940 41970
rect 23884 41860 23940 41918
rect 23884 41794 23940 41804
rect 23772 41300 23828 41310
rect 23660 41298 23828 41300
rect 23660 41246 23774 41298
rect 23826 41246 23828 41298
rect 23660 41244 23828 41246
rect 23772 41234 23828 41244
rect 23884 41300 23940 41310
rect 23660 41076 23716 41086
rect 23548 41074 23828 41076
rect 23548 41022 23662 41074
rect 23714 41022 23828 41074
rect 23548 41020 23828 41022
rect 23660 41010 23716 41020
rect 23436 40898 23492 40908
rect 23212 37998 23214 38050
rect 23266 37998 23268 38050
rect 23212 37986 23268 37998
rect 23324 40292 23380 40302
rect 23324 37266 23380 40236
rect 23436 39394 23492 39406
rect 23436 39342 23438 39394
rect 23490 39342 23492 39394
rect 23436 38836 23492 39342
rect 23660 38836 23716 38874
rect 23436 38780 23660 38836
rect 23660 38770 23716 38780
rect 23772 38668 23828 41020
rect 23884 40068 23940 41244
rect 23996 41188 24052 41198
rect 23996 41094 24052 41132
rect 24108 41186 24164 41198
rect 24108 41134 24110 41186
rect 24162 41134 24164 41186
rect 24108 40626 24164 41134
rect 24108 40574 24110 40626
rect 24162 40574 24164 40626
rect 24108 40562 24164 40574
rect 24332 40402 24388 42028
rect 24444 41972 24500 42140
rect 25116 42084 25172 42094
rect 24444 41906 24500 41916
rect 24556 42082 25172 42084
rect 24556 42030 25118 42082
rect 25170 42030 25172 42082
rect 24556 42028 25172 42030
rect 24556 41970 24612 42028
rect 25116 42018 25172 42028
rect 24556 41918 24558 41970
rect 24610 41918 24612 41970
rect 24556 41906 24612 41918
rect 24332 40350 24334 40402
rect 24386 40350 24388 40402
rect 23884 40002 23940 40012
rect 23996 40180 24052 40190
rect 23996 39058 24052 40124
rect 23996 39006 23998 39058
rect 24050 39006 24052 39058
rect 23996 38994 24052 39006
rect 23324 37214 23326 37266
rect 23378 37214 23380 37266
rect 23324 37202 23380 37214
rect 23436 38612 23492 38622
rect 23324 37044 23380 37054
rect 23324 36482 23380 36988
rect 23324 36430 23326 36482
rect 23378 36430 23380 36482
rect 23324 36418 23380 36430
rect 23436 35698 23492 38556
rect 23436 35646 23438 35698
rect 23490 35646 23492 35698
rect 23436 35588 23492 35646
rect 23436 35522 23492 35532
rect 23548 38612 23828 38668
rect 24332 38668 24388 40350
rect 24556 41412 24612 41422
rect 24556 41298 24612 41356
rect 25228 41412 25284 42364
rect 25452 42420 25508 42430
rect 25340 42084 25396 42094
rect 25340 41990 25396 42028
rect 25452 42082 25508 42364
rect 25900 42420 25956 42478
rect 25900 42308 25956 42364
rect 25452 42030 25454 42082
rect 25506 42030 25508 42082
rect 25452 42018 25508 42030
rect 25676 42252 25956 42308
rect 25676 41748 25732 42252
rect 26796 42196 26852 42924
rect 25900 42084 25956 42094
rect 26348 42084 26404 42094
rect 25900 42082 26404 42084
rect 25900 42030 25902 42082
rect 25954 42030 26350 42082
rect 26402 42030 26404 42082
rect 25900 42028 26404 42030
rect 25900 42018 25956 42028
rect 26348 42018 26404 42028
rect 26796 42082 26852 42140
rect 26908 42420 26964 42430
rect 26908 42194 26964 42364
rect 27132 42420 27188 44046
rect 27692 44098 27860 44100
rect 27692 44046 27806 44098
rect 27858 44046 27860 44098
rect 27692 44044 27860 44046
rect 27580 43762 27636 43774
rect 27580 43710 27582 43762
rect 27634 43710 27636 43762
rect 27580 43092 27636 43710
rect 27692 43540 27748 44044
rect 27804 44034 27860 44044
rect 28140 43988 28196 44942
rect 28140 43922 28196 43932
rect 28028 43652 28084 43662
rect 28252 43652 28308 45388
rect 28364 45330 28420 45388
rect 28364 45278 28366 45330
rect 28418 45278 28420 45330
rect 28364 45266 28420 45278
rect 28476 45220 28532 45612
rect 28476 45154 28532 45164
rect 28588 45108 28644 45118
rect 28588 45014 28644 45052
rect 28476 44994 28532 45006
rect 28476 44942 28478 44994
rect 28530 44942 28532 44994
rect 28476 43764 28532 44942
rect 28924 44884 28980 47516
rect 29148 47346 29204 47358
rect 29148 47294 29150 47346
rect 29202 47294 29204 47346
rect 29148 47236 29204 47294
rect 29260 47348 29316 47358
rect 29372 47348 29428 47852
rect 29260 47346 29428 47348
rect 29260 47294 29262 47346
rect 29314 47294 29428 47346
rect 29260 47292 29428 47294
rect 29260 47282 29316 47292
rect 29148 47170 29204 47180
rect 29036 47124 29092 47134
rect 29036 47012 29092 47068
rect 29036 46956 29204 47012
rect 29148 46340 29204 46956
rect 29260 46900 29316 46910
rect 29260 46674 29316 46844
rect 29260 46622 29262 46674
rect 29314 46622 29316 46674
rect 29260 46610 29316 46622
rect 29372 46564 29428 47292
rect 29596 47012 29652 47966
rect 30044 47572 30100 48188
rect 30268 48020 30324 48030
rect 30380 48020 30436 48190
rect 31052 48244 31108 48300
rect 31164 48244 31220 49086
rect 31836 48356 31892 48366
rect 31500 48354 31892 48356
rect 31500 48302 31838 48354
rect 31890 48302 31892 48354
rect 31500 48300 31892 48302
rect 31388 48244 31444 48254
rect 31052 48242 31444 48244
rect 31052 48190 31390 48242
rect 31442 48190 31444 48242
rect 31052 48188 31444 48190
rect 31388 48178 31444 48188
rect 30940 48130 30996 48142
rect 30940 48078 30942 48130
rect 30994 48078 30996 48130
rect 30380 47964 30772 48020
rect 30268 47926 30324 47964
rect 30044 47506 30100 47516
rect 29596 46946 29652 46956
rect 29484 46788 29540 46798
rect 30044 46788 30100 46798
rect 29484 46786 30100 46788
rect 29484 46734 29486 46786
rect 29538 46734 30046 46786
rect 30098 46734 30100 46786
rect 29484 46732 30100 46734
rect 29484 46722 29540 46732
rect 29820 46564 29876 46574
rect 29372 46508 29820 46564
rect 29820 46470 29876 46508
rect 29148 46284 29540 46340
rect 29372 46002 29428 46014
rect 29372 45950 29374 46002
rect 29426 45950 29428 46002
rect 29260 45892 29316 45902
rect 29260 45106 29316 45836
rect 29372 45444 29428 45950
rect 29372 45378 29428 45388
rect 29484 45890 29540 46284
rect 29484 45838 29486 45890
rect 29538 45838 29540 45890
rect 29260 45054 29262 45106
rect 29314 45054 29316 45106
rect 29260 45042 29316 45054
rect 29372 45108 29428 45118
rect 29372 44994 29428 45052
rect 29372 44942 29374 44994
rect 29426 44942 29428 44994
rect 29372 44930 29428 44942
rect 28700 44828 28980 44884
rect 28588 44098 28644 44110
rect 28588 44046 28590 44098
rect 28642 44046 28644 44098
rect 28588 43988 28644 44046
rect 28588 43922 28644 43932
rect 28476 43698 28532 43708
rect 28028 43558 28084 43596
rect 28140 43650 28308 43652
rect 28140 43598 28254 43650
rect 28306 43598 28308 43650
rect 28140 43596 28308 43598
rect 27692 43474 27748 43484
rect 27804 43538 27860 43550
rect 27804 43486 27806 43538
rect 27858 43486 27860 43538
rect 27580 43026 27636 43036
rect 27804 42978 27860 43486
rect 27804 42926 27806 42978
rect 27858 42926 27860 42978
rect 27804 42914 27860 42926
rect 27916 43428 27972 43438
rect 27356 42868 27412 42878
rect 27412 42812 27748 42868
rect 27356 42774 27412 42812
rect 27692 42644 27748 42812
rect 27916 42754 27972 43372
rect 27916 42702 27918 42754
rect 27970 42702 27972 42754
rect 27916 42690 27972 42702
rect 28028 43204 28084 43214
rect 27804 42644 27860 42654
rect 27692 42642 27860 42644
rect 27692 42590 27806 42642
rect 27858 42590 27860 42642
rect 27692 42588 27860 42590
rect 27804 42578 27860 42588
rect 27132 42354 27188 42364
rect 26908 42142 26910 42194
rect 26962 42142 26964 42194
rect 26908 42130 26964 42142
rect 27132 42196 27188 42206
rect 27916 42196 27972 42206
rect 27132 42194 27972 42196
rect 27132 42142 27134 42194
rect 27186 42142 27918 42194
rect 27970 42142 27972 42194
rect 27132 42140 27972 42142
rect 27132 42130 27188 42140
rect 27916 42130 27972 42140
rect 26796 42030 26798 42082
rect 26850 42030 26852 42082
rect 26796 42018 26852 42030
rect 25228 41346 25284 41356
rect 25452 41692 25732 41748
rect 25788 41972 25844 41982
rect 25788 41748 25844 41916
rect 26460 41972 26516 41982
rect 26908 41972 26964 41982
rect 26460 41970 26628 41972
rect 26460 41918 26462 41970
rect 26514 41918 26628 41970
rect 26460 41916 26628 41918
rect 26460 41906 26516 41916
rect 26348 41860 26404 41870
rect 25788 41692 26068 41748
rect 24556 41246 24558 41298
rect 24610 41246 24612 41298
rect 24556 40292 24612 41246
rect 24668 41188 24724 41198
rect 24668 41094 24724 41132
rect 25452 41186 25508 41692
rect 25900 41412 25956 41422
rect 25900 41298 25956 41356
rect 25900 41246 25902 41298
rect 25954 41246 25956 41298
rect 25452 41134 25454 41186
rect 25506 41134 25508 41186
rect 25452 41122 25508 41134
rect 25676 41188 25732 41198
rect 25676 41094 25732 41132
rect 24556 40226 24612 40236
rect 24668 40964 24724 40974
rect 24444 38836 24500 38846
rect 24444 38742 24500 38780
rect 24332 38612 24612 38668
rect 23548 36596 23604 38612
rect 23884 38164 23940 38174
rect 23884 38162 24500 38164
rect 23884 38110 23886 38162
rect 23938 38110 24500 38162
rect 23884 38108 24500 38110
rect 23884 38098 23940 38108
rect 23660 38052 23716 38062
rect 23660 37958 23716 37996
rect 24220 37940 24276 37950
rect 23772 37938 24276 37940
rect 23772 37886 24222 37938
rect 24274 37886 24276 37938
rect 23772 37884 24276 37886
rect 23772 37378 23828 37884
rect 24220 37874 24276 37884
rect 24332 37940 24388 37950
rect 24332 37846 24388 37884
rect 24444 37938 24500 38108
rect 24444 37886 24446 37938
rect 24498 37886 24500 37938
rect 24444 37874 24500 37886
rect 23772 37326 23774 37378
rect 23826 37326 23828 37378
rect 23772 37314 23828 37326
rect 24444 37492 24500 37502
rect 24556 37492 24612 38612
rect 24668 37716 24724 40908
rect 25788 40628 25844 40638
rect 25788 40534 25844 40572
rect 25564 40514 25620 40526
rect 25564 40462 25566 40514
rect 25618 40462 25620 40514
rect 25004 40404 25060 40414
rect 25004 38500 25060 40348
rect 25452 40402 25508 40414
rect 25452 40350 25454 40402
rect 25506 40350 25508 40402
rect 25452 40180 25508 40350
rect 25452 40114 25508 40124
rect 25564 40404 25620 40462
rect 25900 40404 25956 41246
rect 26012 41300 26068 41692
rect 26348 41746 26404 41804
rect 26348 41694 26350 41746
rect 26402 41694 26404 41746
rect 26012 40514 26068 41244
rect 26012 40462 26014 40514
rect 26066 40462 26068 40514
rect 26012 40450 26068 40462
rect 26124 41636 26180 41646
rect 25452 39844 25508 39854
rect 25228 39620 25284 39630
rect 25228 39526 25284 39564
rect 25452 39506 25508 39788
rect 25452 39454 25454 39506
rect 25506 39454 25508 39506
rect 25452 39442 25508 39454
rect 25564 39058 25620 40348
rect 25564 39006 25566 39058
rect 25618 39006 25620 39058
rect 25564 38994 25620 39006
rect 25788 40348 25956 40404
rect 25004 38434 25060 38444
rect 25228 38834 25284 38846
rect 25228 38782 25230 38834
rect 25282 38782 25284 38834
rect 25228 38612 25284 38782
rect 25004 38052 25060 38062
rect 25228 38052 25284 38556
rect 25340 38164 25396 38174
rect 25340 38070 25396 38108
rect 25060 37996 25284 38052
rect 24724 37660 24836 37716
rect 24668 37650 24724 37660
rect 24444 37490 24612 37492
rect 24444 37438 24446 37490
rect 24498 37438 24612 37490
rect 24444 37436 24612 37438
rect 24108 37266 24164 37278
rect 24108 37214 24110 37266
rect 24162 37214 24164 37266
rect 23660 36596 23716 36606
rect 23548 36594 23716 36596
rect 23548 36542 23662 36594
rect 23714 36542 23716 36594
rect 23548 36540 23716 36542
rect 23548 35586 23604 36540
rect 23660 36530 23716 36540
rect 24108 36594 24164 37214
rect 24444 37044 24500 37436
rect 24444 36978 24500 36988
rect 24108 36542 24110 36594
rect 24162 36542 24164 36594
rect 24108 36484 24164 36542
rect 24108 36418 24164 36428
rect 24780 35922 24836 37660
rect 25004 37604 25060 37996
rect 25340 37940 25396 37950
rect 25116 37884 25340 37940
rect 25116 37826 25172 37884
rect 25340 37874 25396 37884
rect 25564 37940 25620 37950
rect 25116 37774 25118 37826
rect 25170 37774 25172 37826
rect 25116 37762 25172 37774
rect 25228 37716 25284 37726
rect 25284 37660 25396 37716
rect 25228 37650 25284 37660
rect 25004 37548 25172 37604
rect 24780 35870 24782 35922
rect 24834 35870 24836 35922
rect 24780 35858 24836 35870
rect 23884 35700 23940 35710
rect 23884 35606 23940 35644
rect 23548 35534 23550 35586
rect 23602 35534 23604 35586
rect 23548 35522 23604 35534
rect 23100 34626 23156 34636
rect 23212 34692 23268 34702
rect 23548 34692 23604 34702
rect 23996 34692 24052 34702
rect 23212 34690 23380 34692
rect 23212 34638 23214 34690
rect 23266 34638 23380 34690
rect 23212 34636 23380 34638
rect 23212 34626 23268 34636
rect 22988 34412 23268 34468
rect 22652 34354 22932 34356
rect 22652 34302 22654 34354
rect 22706 34302 22932 34354
rect 22652 34300 22932 34302
rect 22652 34290 22708 34300
rect 22540 34076 22708 34132
rect 22204 31726 22206 31778
rect 22258 31726 22260 31778
rect 22204 31714 22260 31726
rect 22316 31836 22484 31892
rect 22092 30156 22260 30212
rect 20524 30046 20526 30098
rect 20578 30046 20580 30098
rect 20524 30034 20580 30046
rect 21308 29876 21364 30156
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 21308 29810 21364 29820
rect 22092 29986 22148 29998
rect 22092 29934 22094 29986
rect 22146 29934 22148 29986
rect 22092 29876 22148 29934
rect 22092 29810 22148 29820
rect 19836 29754 20100 29764
rect 19516 29650 19684 29652
rect 19516 29598 19518 29650
rect 19570 29598 19684 29650
rect 19516 29596 19684 29598
rect 19516 29586 19572 29596
rect 19516 28756 19572 28766
rect 19404 28754 19572 28756
rect 19404 28702 19518 28754
rect 19570 28702 19572 28754
rect 19404 28700 19572 28702
rect 19516 28690 19572 28700
rect 19628 28532 19684 29596
rect 21308 29426 21364 29438
rect 21308 29374 21310 29426
rect 21362 29374 21364 29426
rect 21308 29316 21364 29374
rect 21308 29250 21364 29260
rect 21980 29314 22036 29326
rect 21980 29262 21982 29314
rect 22034 29262 22036 29314
rect 21980 28866 22036 29262
rect 22204 29204 22260 30156
rect 21980 28814 21982 28866
rect 22034 28814 22036 28866
rect 21980 28802 22036 28814
rect 22092 29148 22260 29204
rect 21308 28532 21364 28542
rect 19068 28476 19684 28532
rect 18956 28420 19012 28430
rect 18956 28326 19012 28364
rect 18844 28084 18900 28094
rect 18732 27748 18788 27758
rect 18396 27134 18398 27186
rect 18450 27134 18452 27186
rect 18284 26290 18340 26302
rect 18284 26238 18286 26290
rect 18338 26238 18340 26290
rect 18172 25620 18228 25630
rect 18284 25620 18340 26238
rect 18396 26292 18452 27134
rect 18620 27746 18788 27748
rect 18620 27694 18734 27746
rect 18786 27694 18788 27746
rect 18620 27692 18788 27694
rect 18620 26964 18676 27692
rect 18732 27682 18788 27692
rect 18732 27188 18788 27198
rect 18732 27094 18788 27132
rect 18620 26898 18676 26908
rect 18844 26962 18900 28028
rect 19068 27858 19124 28476
rect 19292 27972 19348 27982
rect 19068 27806 19070 27858
rect 19122 27806 19124 27858
rect 19068 27794 19124 27806
rect 19180 27970 19348 27972
rect 19180 27918 19294 27970
rect 19346 27918 19348 27970
rect 19180 27916 19348 27918
rect 18844 26910 18846 26962
rect 18898 26910 18900 26962
rect 18844 26898 18900 26910
rect 19068 26962 19124 26974
rect 19068 26910 19070 26962
rect 19122 26910 19124 26962
rect 19068 26740 19124 26910
rect 19068 26674 19124 26684
rect 19180 26404 19236 27916
rect 19292 27906 19348 27916
rect 19628 27860 19684 28476
rect 21084 28476 21308 28532
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19740 28084 19796 28094
rect 19740 27990 19796 28028
rect 19852 28084 19908 28094
rect 19852 28082 20132 28084
rect 19852 28030 19854 28082
rect 19906 28030 20132 28082
rect 19852 28028 20132 28030
rect 19852 28018 19908 28028
rect 20076 27972 20132 28028
rect 20188 27972 20244 27982
rect 20076 27916 20188 27972
rect 20188 27906 20244 27916
rect 20524 27972 20580 27982
rect 20524 27878 20580 27916
rect 20748 27860 20804 27870
rect 19628 27804 20132 27860
rect 19964 27636 20020 27646
rect 19404 27634 20020 27636
rect 19404 27582 19966 27634
rect 20018 27582 20020 27634
rect 19404 27580 20020 27582
rect 19404 27186 19460 27580
rect 19964 27570 20020 27580
rect 20076 27300 20132 27804
rect 20748 27766 20804 27804
rect 21084 27858 21140 28476
rect 21084 27806 21086 27858
rect 21138 27806 21140 27858
rect 21084 27794 21140 27806
rect 20412 27636 20468 27646
rect 19404 27134 19406 27186
rect 19458 27134 19460 27186
rect 19404 27122 19460 27134
rect 19852 27244 20132 27300
rect 20300 27634 20468 27636
rect 20300 27582 20414 27634
rect 20466 27582 20468 27634
rect 20300 27580 20468 27582
rect 19068 26348 19236 26404
rect 19292 26852 19348 26862
rect 18620 26292 18676 26302
rect 18396 26236 18620 26292
rect 18620 26198 18676 26236
rect 18844 26292 18900 26302
rect 18172 25618 18340 25620
rect 18172 25566 18174 25618
rect 18226 25566 18340 25618
rect 18172 25564 18340 25566
rect 18172 25554 18228 25564
rect 18284 25508 18340 25564
rect 18284 25442 18340 25452
rect 18620 25956 18676 25966
rect 18508 25396 18564 25406
rect 18396 25394 18564 25396
rect 18396 25342 18510 25394
rect 18562 25342 18564 25394
rect 18396 25340 18564 25342
rect 18284 25172 18340 25182
rect 18396 25172 18452 25340
rect 18508 25330 18564 25340
rect 18340 25116 18452 25172
rect 18284 25106 18340 25116
rect 18396 24948 18452 24958
rect 18396 24854 18452 24892
rect 18060 23774 18062 23826
rect 18114 23774 18116 23826
rect 16716 23266 16772 23278
rect 16716 23214 16718 23266
rect 16770 23214 16772 23266
rect 16716 22708 16772 23214
rect 17500 23268 17556 23278
rect 17500 23174 17556 23212
rect 16716 22642 16772 22652
rect 18060 23154 18116 23774
rect 18060 23102 18062 23154
rect 18114 23102 18116 23154
rect 16940 22484 16996 22494
rect 16716 22260 16772 22270
rect 16156 19234 16548 19236
rect 16156 19182 16158 19234
rect 16210 19182 16494 19234
rect 16546 19182 16548 19234
rect 16156 19180 16548 19182
rect 16156 19170 16212 19180
rect 16492 19170 16548 19180
rect 16604 22204 16716 22260
rect 16604 19236 16660 22204
rect 16716 22166 16772 22204
rect 16940 21700 16996 22428
rect 17948 22372 18004 22382
rect 17948 22278 18004 22316
rect 17164 22260 17220 22270
rect 17164 22166 17220 22204
rect 18060 22258 18116 23102
rect 18396 23940 18452 23950
rect 18060 22206 18062 22258
rect 18114 22206 18116 22258
rect 18060 22194 18116 22206
rect 18284 22930 18340 22942
rect 18284 22878 18286 22930
rect 18338 22878 18340 22930
rect 17500 22148 17556 22158
rect 16604 19170 16660 19180
rect 16716 21644 16996 21700
rect 17276 22146 17556 22148
rect 17276 22094 17502 22146
rect 17554 22094 17556 22146
rect 17276 22092 17556 22094
rect 16716 21586 16772 21644
rect 16716 21534 16718 21586
rect 16770 21534 16772 21586
rect 16604 19012 16660 19022
rect 16604 18676 16660 18956
rect 16604 18610 16660 18620
rect 16716 18228 16772 21534
rect 16940 20802 16996 20814
rect 16940 20750 16942 20802
rect 16994 20750 16996 20802
rect 16940 18452 16996 20750
rect 16940 18386 16996 18396
rect 16716 18172 17220 18228
rect 15820 17724 16100 17780
rect 16716 17892 16772 17902
rect 15820 17108 15876 17724
rect 16604 17666 16660 17678
rect 16604 17614 16606 17666
rect 16658 17614 16660 17666
rect 15932 17556 15988 17566
rect 16380 17556 16436 17566
rect 15932 17554 16100 17556
rect 15932 17502 15934 17554
rect 15986 17502 16100 17554
rect 15932 17500 16100 17502
rect 15932 17490 15988 17500
rect 15820 16100 15876 17052
rect 15932 16996 15988 17006
rect 15932 16882 15988 16940
rect 15932 16830 15934 16882
rect 15986 16830 15988 16882
rect 15932 16818 15988 16830
rect 16044 16324 16100 17500
rect 16380 17462 16436 17500
rect 16604 17444 16660 17614
rect 16492 17108 16548 17118
rect 16492 17014 16548 17052
rect 16156 16994 16212 17006
rect 16156 16942 16158 16994
rect 16210 16942 16212 16994
rect 16156 16772 16212 16942
rect 16156 16706 16212 16716
rect 16604 16772 16660 17388
rect 16716 17108 16772 17836
rect 16716 17042 16772 17052
rect 17164 17778 17220 18172
rect 17164 17726 17166 17778
rect 17218 17726 17220 17778
rect 16604 16706 16660 16716
rect 16828 16994 16884 17006
rect 17164 16996 17220 17726
rect 16828 16942 16830 16994
rect 16882 16942 16884 16994
rect 16716 16548 16772 16558
rect 16156 16324 16212 16334
rect 16044 16322 16660 16324
rect 16044 16270 16158 16322
rect 16210 16270 16660 16322
rect 16044 16268 16660 16270
rect 16156 16258 16212 16268
rect 16604 16100 16660 16268
rect 15820 16098 16212 16100
rect 15820 16046 15822 16098
rect 15874 16046 16212 16098
rect 15820 16044 16212 16046
rect 15820 16034 15876 16044
rect 16156 15538 16212 16044
rect 16492 16044 16660 16100
rect 16268 15986 16324 15998
rect 16268 15934 16270 15986
rect 16322 15934 16324 15986
rect 16268 15876 16324 15934
rect 16268 15810 16324 15820
rect 16156 15486 16158 15538
rect 16210 15486 16212 15538
rect 16156 15474 16212 15486
rect 16492 15538 16548 16044
rect 16716 15988 16772 16492
rect 16828 16436 16884 16942
rect 16828 16370 16884 16380
rect 17052 16940 17164 16996
rect 17052 16098 17108 16940
rect 17164 16930 17220 16940
rect 17276 16660 17332 22092
rect 17500 22082 17556 22092
rect 18172 21364 18228 21374
rect 17836 21362 18228 21364
rect 17836 21310 18174 21362
rect 18226 21310 18228 21362
rect 17836 21308 18228 21310
rect 17612 20690 17668 20702
rect 17612 20638 17614 20690
rect 17666 20638 17668 20690
rect 17500 20244 17556 20254
rect 17612 20244 17668 20638
rect 17500 20242 17668 20244
rect 17500 20190 17502 20242
rect 17554 20190 17668 20242
rect 17500 20188 17668 20190
rect 17500 20178 17556 20188
rect 17836 20130 17892 21308
rect 18172 21298 18228 21308
rect 17836 20078 17838 20130
rect 17890 20078 17892 20130
rect 17836 20066 17892 20078
rect 18172 19908 18228 19918
rect 18172 19814 18228 19852
rect 17500 18452 17556 18462
rect 17500 16882 17556 18396
rect 18284 17892 18340 22878
rect 18396 22258 18452 23884
rect 18508 23828 18564 23838
rect 18508 22482 18564 23772
rect 18508 22430 18510 22482
rect 18562 22430 18564 22482
rect 18508 22418 18564 22430
rect 18396 22206 18398 22258
rect 18450 22206 18452 22258
rect 18396 22194 18452 22206
rect 18620 21588 18676 25900
rect 18844 25620 18900 26236
rect 18620 21522 18676 21532
rect 18732 25506 18788 25518
rect 18732 25454 18734 25506
rect 18786 25454 18788 25506
rect 18732 25396 18788 25454
rect 18844 25506 18900 25564
rect 18844 25454 18846 25506
rect 18898 25454 18900 25506
rect 18844 25442 18900 25454
rect 18732 24050 18788 25340
rect 18732 23998 18734 24050
rect 18786 23998 18788 24050
rect 18508 21362 18564 21374
rect 18508 21310 18510 21362
rect 18562 21310 18564 21362
rect 18508 20132 18564 21310
rect 18508 20066 18564 20076
rect 18732 19906 18788 23998
rect 18844 24834 18900 24846
rect 18844 24782 18846 24834
rect 18898 24782 18900 24834
rect 18844 22372 18900 24782
rect 19068 24052 19124 26348
rect 19180 26180 19236 26190
rect 19292 26180 19348 26796
rect 19852 26852 19908 27244
rect 20300 27186 20356 27580
rect 20412 27570 20468 27580
rect 20300 27134 20302 27186
rect 20354 27134 20356 27186
rect 20300 27122 20356 27134
rect 20076 27076 20132 27086
rect 20076 26982 20132 27020
rect 21308 27074 21364 28476
rect 22092 28530 22148 29148
rect 22316 28756 22372 31836
rect 22428 31668 22484 31678
rect 22428 31574 22484 31612
rect 22540 30884 22596 30894
rect 22092 28478 22094 28530
rect 22146 28478 22148 28530
rect 21644 28420 21700 28430
rect 21644 28326 21700 28364
rect 22092 28084 22148 28478
rect 22204 28700 22372 28756
rect 22428 30882 22596 30884
rect 22428 30830 22542 30882
rect 22594 30830 22596 30882
rect 22428 30828 22596 30830
rect 22652 30884 22708 34076
rect 22764 33348 22820 33358
rect 22764 33254 22820 33292
rect 22876 32676 22932 34300
rect 23212 34242 23268 34412
rect 23212 34190 23214 34242
rect 23266 34190 23268 34242
rect 23212 34178 23268 34190
rect 23212 33684 23268 33694
rect 23324 33684 23380 34636
rect 23548 34690 24052 34692
rect 23548 34638 23550 34690
rect 23602 34638 23998 34690
rect 24050 34638 24052 34690
rect 23548 34636 24052 34638
rect 23548 34626 23604 34636
rect 23996 34356 24052 34636
rect 23996 34290 24052 34300
rect 24444 34468 24500 34478
rect 23548 34130 23604 34142
rect 23548 34078 23550 34130
rect 23602 34078 23604 34130
rect 23268 33628 23380 33684
rect 23436 34018 23492 34030
rect 23436 33966 23438 34018
rect 23490 33966 23492 34018
rect 23212 33618 23268 33628
rect 22764 32620 22932 32676
rect 23100 33122 23156 33134
rect 23100 33070 23102 33122
rect 23154 33070 23156 33122
rect 22764 31332 22820 32620
rect 22876 32450 22932 32462
rect 22876 32398 22878 32450
rect 22930 32398 22932 32450
rect 22876 31668 22932 32398
rect 23100 32116 23156 33070
rect 23436 33124 23492 33966
rect 23548 33572 23604 34078
rect 24444 34130 24500 34412
rect 24444 34078 24446 34130
rect 24498 34078 24500 34130
rect 24444 34066 24500 34078
rect 23548 33506 23604 33516
rect 24108 33906 24164 33918
rect 24108 33854 24110 33906
rect 24162 33854 24164 33906
rect 23772 33348 23828 33358
rect 23772 33254 23828 33292
rect 23436 33030 23492 33068
rect 24108 32788 24164 33854
rect 24444 33908 24500 33918
rect 24444 33906 24612 33908
rect 24444 33854 24446 33906
rect 24498 33854 24612 33906
rect 24444 33852 24612 33854
rect 24444 33842 24500 33852
rect 24556 33458 24612 33852
rect 24556 33406 24558 33458
rect 24610 33406 24612 33458
rect 24556 33394 24612 33406
rect 24892 33460 24948 33470
rect 23660 32732 24164 32788
rect 23100 32050 23156 32060
rect 23324 32562 23380 32574
rect 23324 32510 23326 32562
rect 23378 32510 23380 32562
rect 23324 32004 23380 32510
rect 23548 32564 23604 32574
rect 23548 32470 23604 32508
rect 23660 32450 23716 32732
rect 23660 32398 23662 32450
rect 23714 32398 23716 32450
rect 23548 32228 23604 32238
rect 23660 32228 23716 32398
rect 23604 32172 23716 32228
rect 23772 32562 23828 32574
rect 23772 32510 23774 32562
rect 23826 32510 23828 32562
rect 23548 32162 23604 32172
rect 23772 32116 23828 32510
rect 23996 32564 24052 32574
rect 24332 32564 24388 32574
rect 23996 32562 24388 32564
rect 23996 32510 23998 32562
rect 24050 32510 24334 32562
rect 24386 32510 24388 32562
rect 23996 32508 24388 32510
rect 23996 32498 24052 32508
rect 24332 32498 24388 32508
rect 24892 32564 24948 33404
rect 23772 32050 23828 32060
rect 24444 32450 24500 32462
rect 24444 32398 24446 32450
rect 24498 32398 24500 32450
rect 23324 31938 23380 31948
rect 23548 32002 23604 32014
rect 23548 31950 23550 32002
rect 23602 31950 23604 32002
rect 23100 31778 23156 31790
rect 23100 31726 23102 31778
rect 23154 31726 23156 31778
rect 23100 31668 23156 31726
rect 22876 31612 23156 31668
rect 22876 31556 22932 31612
rect 22876 31490 22932 31500
rect 22764 31276 22932 31332
rect 22652 30828 22820 30884
rect 22204 28532 22260 28700
rect 22204 28466 22260 28476
rect 22316 28530 22372 28542
rect 22316 28478 22318 28530
rect 22370 28478 22372 28530
rect 21644 27972 21700 27982
rect 21532 27860 21588 27870
rect 21308 27022 21310 27074
rect 21362 27022 21364 27074
rect 21308 27010 21364 27022
rect 21420 27746 21476 27758
rect 21420 27694 21422 27746
rect 21474 27694 21476 27746
rect 21196 26962 21252 26974
rect 21196 26910 21198 26962
rect 21250 26910 21252 26962
rect 21196 26908 21252 26910
rect 19852 26786 19908 26796
rect 20412 26852 21252 26908
rect 19404 26740 19460 26750
rect 19460 26684 19572 26740
rect 19404 26674 19460 26684
rect 19516 26402 19572 26684
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19516 26350 19518 26402
rect 19570 26350 19572 26402
rect 19516 26338 19572 26350
rect 19964 26290 20020 26302
rect 19964 26238 19966 26290
rect 20018 26238 20020 26290
rect 19180 26178 19348 26180
rect 19180 26126 19182 26178
rect 19234 26126 19348 26178
rect 19180 26124 19348 26126
rect 19180 26114 19236 26124
rect 19068 23996 19236 24052
rect 19068 23828 19124 23838
rect 19068 23734 19124 23772
rect 18844 22278 18900 22316
rect 19068 23492 19124 23502
rect 19068 22258 19124 23436
rect 19180 22372 19236 23996
rect 19292 23044 19348 26124
rect 19628 26180 19684 26190
rect 19628 24500 19684 26124
rect 19964 26180 20020 26238
rect 20412 26290 20468 26852
rect 21420 26404 21476 27694
rect 21532 26964 21588 27804
rect 21644 27860 21700 27916
rect 21644 27858 21812 27860
rect 21644 27806 21646 27858
rect 21698 27806 21812 27858
rect 21644 27804 21812 27806
rect 21644 27794 21700 27804
rect 21532 26898 21588 26908
rect 21644 27636 21700 27646
rect 21420 26338 21476 26348
rect 20412 26238 20414 26290
rect 20466 26238 20468 26290
rect 20412 26226 20468 26238
rect 21532 26292 21588 26302
rect 21644 26292 21700 27580
rect 21532 26290 21700 26292
rect 21532 26238 21534 26290
rect 21586 26238 21700 26290
rect 21532 26236 21700 26238
rect 21756 27076 21812 27804
rect 22092 27412 22148 28028
rect 22316 27970 22372 28478
rect 22316 27918 22318 27970
rect 22370 27918 22372 27970
rect 22316 27906 22372 27918
rect 22092 27346 22148 27356
rect 21868 27076 21924 27086
rect 21756 27074 21924 27076
rect 21756 27022 21870 27074
rect 21922 27022 21924 27074
rect 21756 27020 21924 27022
rect 21084 26180 21140 26190
rect 21532 26180 21588 26236
rect 19964 26114 20020 26124
rect 20636 26178 21140 26180
rect 20636 26126 21086 26178
rect 21138 26126 21140 26178
rect 20636 26124 21140 26126
rect 19740 25396 19796 25406
rect 19740 25302 19796 25340
rect 20188 25394 20244 25406
rect 20188 25342 20190 25394
rect 20242 25342 20244 25394
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20076 24836 20132 24846
rect 19852 24780 20076 24836
rect 19852 24722 19908 24780
rect 20076 24770 20132 24780
rect 19852 24670 19854 24722
rect 19906 24670 19908 24722
rect 19852 24658 19908 24670
rect 20076 24610 20132 24622
rect 20076 24558 20078 24610
rect 20130 24558 20132 24610
rect 20076 24500 20132 24558
rect 19628 24444 20132 24500
rect 19628 23828 19684 24444
rect 20188 23940 20244 25342
rect 20636 24836 20692 26124
rect 21084 26114 21140 26124
rect 21308 26124 21588 26180
rect 20748 25508 20804 25518
rect 21308 25508 21364 26124
rect 20748 25506 21364 25508
rect 20748 25454 20750 25506
rect 20802 25454 21364 25506
rect 20748 25452 21364 25454
rect 21420 25508 21476 25518
rect 20748 25442 20804 25452
rect 20188 23874 20244 23884
rect 20524 24780 20636 24836
rect 19628 23380 19684 23772
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23324 19908 23380
rect 19852 23266 19908 23324
rect 19852 23214 19854 23266
rect 19906 23214 19908 23266
rect 19852 23202 19908 23214
rect 19740 23156 19796 23166
rect 19628 23044 19684 23054
rect 19292 22988 19628 23044
rect 19628 22950 19684 22988
rect 19740 22930 19796 23100
rect 20524 23156 20580 24780
rect 20636 24770 20692 24780
rect 20748 25060 20804 25070
rect 21420 25060 21476 25452
rect 21532 25284 21588 25294
rect 21532 25190 21588 25228
rect 20524 23062 20580 23100
rect 20748 24612 20804 25004
rect 20748 23938 20804 24556
rect 21308 25004 21476 25060
rect 20748 23886 20750 23938
rect 20802 23886 20804 23938
rect 20636 22932 20692 22942
rect 19740 22878 19742 22930
rect 19794 22878 19796 22930
rect 19740 22866 19796 22878
rect 20300 22876 20636 22932
rect 20300 22594 20356 22876
rect 20300 22542 20302 22594
rect 20354 22542 20356 22594
rect 20300 22530 20356 22542
rect 19180 22278 19236 22316
rect 20188 22372 20244 22382
rect 19740 22260 19796 22270
rect 19068 22206 19070 22258
rect 19122 22206 19124 22258
rect 19068 22194 19124 22206
rect 19628 22258 19796 22260
rect 19628 22206 19742 22258
rect 19794 22206 19796 22258
rect 19628 22204 19796 22206
rect 19292 22148 19348 22158
rect 19068 21700 19124 21710
rect 19068 21606 19124 21644
rect 19180 21586 19236 21598
rect 19180 21534 19182 21586
rect 19234 21534 19236 21586
rect 19180 20692 19236 21534
rect 19180 20018 19236 20636
rect 19292 20130 19348 22092
rect 19292 20078 19294 20130
rect 19346 20078 19348 20130
rect 19292 20066 19348 20078
rect 19180 19966 19182 20018
rect 19234 19966 19236 20018
rect 19180 19954 19236 19966
rect 18732 19854 18734 19906
rect 18786 19854 18788 19906
rect 18508 19794 18564 19806
rect 18508 19742 18510 19794
rect 18562 19742 18564 19794
rect 18508 19572 18564 19742
rect 18508 19506 18564 19516
rect 18732 19236 18788 19854
rect 18732 19170 18788 19180
rect 19180 19796 19236 19806
rect 19180 19234 19236 19740
rect 19180 19182 19182 19234
rect 19234 19182 19236 19234
rect 19180 19170 19236 19182
rect 19404 19012 19460 19022
rect 19404 19010 19572 19012
rect 19404 18958 19406 19010
rect 19458 18958 19572 19010
rect 19404 18956 19572 18958
rect 19404 18946 19460 18956
rect 19516 18562 19572 18956
rect 19516 18510 19518 18562
rect 19570 18510 19572 18562
rect 19516 18498 19572 18510
rect 18732 18452 18788 18462
rect 18732 18358 18788 18396
rect 19628 18340 19684 22204
rect 19740 22194 19796 22204
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21698 20244 22316
rect 20300 21812 20356 21822
rect 20300 21718 20356 21756
rect 20188 21646 20190 21698
rect 20242 21646 20244 21698
rect 20188 21634 20244 21646
rect 20412 21588 20468 22876
rect 20636 22866 20692 22876
rect 20636 22596 20692 22606
rect 20748 22596 20804 23886
rect 20636 22594 20804 22596
rect 20636 22542 20638 22594
rect 20690 22542 20804 22594
rect 20636 22540 20804 22542
rect 20860 23940 20916 23950
rect 20636 22530 20692 22540
rect 20524 22370 20580 22382
rect 20524 22318 20526 22370
rect 20578 22318 20580 22370
rect 20524 21812 20580 22318
rect 20748 21812 20804 21822
rect 20524 21810 20804 21812
rect 20524 21758 20750 21810
rect 20802 21758 20804 21810
rect 20524 21756 20804 21758
rect 20748 21746 20804 21756
rect 20860 21698 20916 23884
rect 21196 23380 21252 23390
rect 21084 23324 21196 23380
rect 20972 23266 21028 23278
rect 20972 23214 20974 23266
rect 21026 23214 21028 23266
rect 20972 22932 21028 23214
rect 20972 22866 21028 22876
rect 20860 21646 20862 21698
rect 20914 21646 20916 21698
rect 20860 21634 20916 21646
rect 21084 21924 21140 23324
rect 21196 23314 21252 23324
rect 20524 21588 20580 21598
rect 20412 21586 20580 21588
rect 20412 21534 20526 21586
rect 20578 21534 20580 21586
rect 20412 21532 20580 21534
rect 20524 21522 20580 21532
rect 21084 21364 21140 21868
rect 21308 21812 21364 25004
rect 21756 24276 21812 27020
rect 21868 27010 21924 27020
rect 22428 26908 22484 30828
rect 22540 30818 22596 30828
rect 22652 27972 22708 27982
rect 22652 27878 22708 27916
rect 22540 27076 22596 27086
rect 22540 26982 22596 27020
rect 22764 26908 22820 30828
rect 22876 30212 22932 31276
rect 22988 31220 23044 31230
rect 22988 31126 23044 31164
rect 23100 31106 23156 31612
rect 23100 31054 23102 31106
rect 23154 31054 23156 31106
rect 23100 31042 23156 31054
rect 23548 31668 23604 31950
rect 23660 31780 23716 31790
rect 23660 31778 23828 31780
rect 23660 31726 23662 31778
rect 23714 31726 23828 31778
rect 23660 31724 23828 31726
rect 23660 31714 23716 31724
rect 22876 30146 22932 30156
rect 22988 30212 23044 30222
rect 22988 30210 23268 30212
rect 22988 30158 22990 30210
rect 23042 30158 23268 30210
rect 22988 30156 23268 30158
rect 22988 30146 23044 30156
rect 23212 28754 23268 30156
rect 23212 28702 23214 28754
rect 23266 28702 23268 28754
rect 23212 28690 23268 28702
rect 23548 28754 23604 31612
rect 23772 31332 23828 31724
rect 24444 31556 24500 32398
rect 24444 31490 24500 31500
rect 24556 31890 24612 31902
rect 24556 31838 24558 31890
rect 24610 31838 24612 31890
rect 24556 31668 24612 31838
rect 24892 31668 24948 32508
rect 23772 31276 24276 31332
rect 24220 31218 24276 31276
rect 24220 31166 24222 31218
rect 24274 31166 24276 31218
rect 24220 31154 24276 31166
rect 23884 31106 23940 31118
rect 23884 31054 23886 31106
rect 23938 31054 23940 31106
rect 23884 30772 23940 31054
rect 24444 31106 24500 31118
rect 24444 31054 24446 31106
rect 24498 31054 24500 31106
rect 23996 30996 24052 31006
rect 23996 30902 24052 30940
rect 24444 30772 24500 31054
rect 24556 30996 24612 31612
rect 24556 30902 24612 30940
rect 24668 31666 24948 31668
rect 24668 31614 24894 31666
rect 24946 31614 24948 31666
rect 24668 31612 24948 31614
rect 24668 30772 24724 31612
rect 24892 31602 24948 31612
rect 25004 32340 25060 32350
rect 23884 30716 24724 30772
rect 24332 30212 24388 30222
rect 24332 30118 24388 30156
rect 23548 28702 23550 28754
rect 23602 28702 23604 28754
rect 23548 28690 23604 28702
rect 24108 29314 24164 29326
rect 24108 29262 24110 29314
rect 24162 29262 24164 29314
rect 23660 28644 23716 28654
rect 24108 28644 24164 29262
rect 23660 28642 24164 28644
rect 23660 28590 23662 28642
rect 23714 28590 24164 28642
rect 23660 28588 24164 28590
rect 24668 29316 24724 29326
rect 22876 27858 22932 27870
rect 22876 27806 22878 27858
rect 22930 27806 22932 27858
rect 22876 27636 22932 27806
rect 22876 27570 22932 27580
rect 23660 27636 23716 28588
rect 23996 28420 24052 28430
rect 23996 27972 24052 28364
rect 24668 28196 24724 29260
rect 25004 28868 25060 32284
rect 25004 28802 25060 28812
rect 24668 28140 24948 28196
rect 23996 27858 24052 27916
rect 24668 27972 24724 27982
rect 23996 27806 23998 27858
rect 24050 27806 24052 27858
rect 23996 27794 24052 27806
rect 24444 27860 24500 27870
rect 24444 27766 24500 27804
rect 24556 27858 24612 27870
rect 24556 27806 24558 27858
rect 24610 27806 24612 27858
rect 23660 27570 23716 27580
rect 24220 27746 24276 27758
rect 24220 27694 24222 27746
rect 24274 27694 24276 27746
rect 23660 27412 23716 27422
rect 21980 26852 22036 26862
rect 22316 26852 22484 26908
rect 22652 26852 22820 26908
rect 22876 26964 22932 26974
rect 22036 26796 22148 26852
rect 21980 26786 22036 26796
rect 21980 26402 22036 26414
rect 21980 26350 21982 26402
rect 22034 26350 22036 26402
rect 21308 21746 21364 21756
rect 21420 24220 21812 24276
rect 21868 26066 21924 26078
rect 21868 26014 21870 26066
rect 21922 26014 21924 26066
rect 21420 21810 21476 24220
rect 21868 23604 21924 26014
rect 21980 25508 22036 26350
rect 21980 25442 22036 25452
rect 22092 25506 22148 26796
rect 22092 25454 22094 25506
rect 22146 25454 22148 25506
rect 22092 25442 22148 25454
rect 22204 26290 22260 26302
rect 22204 26238 22206 26290
rect 22258 26238 22260 26290
rect 22204 25060 22260 26238
rect 22204 24994 22260 25004
rect 22204 24834 22260 24846
rect 22204 24782 22206 24834
rect 22258 24782 22260 24834
rect 22204 24612 22260 24782
rect 22204 24546 22260 24556
rect 21756 23548 21924 23604
rect 21532 23156 21588 23166
rect 21532 22482 21588 23100
rect 21756 22596 21812 23548
rect 21868 23380 21924 23390
rect 21868 23286 21924 23324
rect 22316 23268 22372 26852
rect 22652 26516 22708 26852
rect 22652 26460 22820 26516
rect 22540 26404 22596 26414
rect 22596 26348 22708 26404
rect 22540 26338 22596 26348
rect 22428 26290 22484 26302
rect 22428 26238 22430 26290
rect 22482 26238 22484 26290
rect 22428 25396 22484 26238
rect 22652 25508 22708 26348
rect 22764 26068 22820 26460
rect 22876 26292 22932 26908
rect 23436 26852 23492 26862
rect 23324 26850 23492 26852
rect 23324 26798 23438 26850
rect 23490 26798 23492 26850
rect 23324 26796 23492 26798
rect 22876 26290 23044 26292
rect 22876 26238 22878 26290
rect 22930 26238 23044 26290
rect 22876 26236 23044 26238
rect 22876 26226 22932 26236
rect 22764 26012 22932 26068
rect 22764 25508 22820 25518
rect 22652 25506 22820 25508
rect 22652 25454 22766 25506
rect 22818 25454 22820 25506
rect 22652 25452 22820 25454
rect 22764 25442 22820 25452
rect 22540 25396 22596 25406
rect 22428 25394 22596 25396
rect 22428 25342 22542 25394
rect 22594 25342 22596 25394
rect 22428 25340 22596 25342
rect 21532 22430 21534 22482
rect 21586 22430 21588 22482
rect 21532 22418 21588 22430
rect 21644 22594 21812 22596
rect 21644 22542 21758 22594
rect 21810 22542 21812 22594
rect 21644 22540 21812 22542
rect 21420 21758 21422 21810
rect 21474 21758 21476 21810
rect 21420 21746 21476 21758
rect 21644 21698 21700 22540
rect 21756 22530 21812 22540
rect 22092 23212 22372 23268
rect 22428 24610 22484 24622
rect 22428 24558 22430 24610
rect 22482 24558 22484 24610
rect 22092 22372 22148 23212
rect 22204 23044 22260 23054
rect 22204 22950 22260 22988
rect 22092 22316 22260 22372
rect 22092 22148 22148 22158
rect 22092 22054 22148 22092
rect 21644 21646 21646 21698
rect 21698 21646 21700 21698
rect 21644 21634 21700 21646
rect 22092 21700 22148 21710
rect 21532 21476 21588 21486
rect 21532 21474 21812 21476
rect 21532 21422 21534 21474
rect 21586 21422 21812 21474
rect 21532 21420 21812 21422
rect 21532 21410 21588 21420
rect 20636 21308 21140 21364
rect 19740 20914 19796 20926
rect 19740 20862 19742 20914
rect 19794 20862 19796 20914
rect 19740 20580 19796 20862
rect 20636 20802 20692 21308
rect 20636 20750 20638 20802
rect 20690 20750 20692 20802
rect 20636 20738 20692 20750
rect 20300 20692 20356 20702
rect 20300 20598 20356 20636
rect 20524 20580 20580 20590
rect 19740 20524 20244 20580
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20132 20244 20524
rect 20524 20486 20580 20524
rect 21420 20580 21476 20590
rect 21420 20486 21476 20524
rect 20188 20066 20244 20076
rect 21084 20468 21140 20478
rect 20860 19906 20916 19918
rect 20860 19854 20862 19906
rect 20914 19854 20916 19906
rect 19964 19794 20020 19806
rect 19964 19742 19966 19794
rect 20018 19742 20020 19794
rect 19852 19236 19908 19246
rect 19852 19142 19908 19180
rect 19964 19012 20020 19742
rect 20300 19796 20356 19806
rect 20300 19702 20356 19740
rect 19964 18956 20244 19012
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 18060 17836 18340 17892
rect 19292 18284 19684 18340
rect 17500 16830 17502 16882
rect 17554 16830 17556 16882
rect 17500 16818 17556 16830
rect 17612 16996 17668 17006
rect 17276 16594 17332 16604
rect 17388 16772 17444 16782
rect 17052 16046 17054 16098
rect 17106 16046 17108 16098
rect 17052 16034 17108 16046
rect 16492 15486 16494 15538
rect 16546 15486 16548 15538
rect 16492 15474 16548 15486
rect 16604 15986 16772 15988
rect 16604 15934 16718 15986
rect 16770 15934 16772 15986
rect 16604 15932 16772 15934
rect 15708 15092 16100 15148
rect 15596 13794 15652 13804
rect 16044 14418 16100 15092
rect 16604 14530 16660 15932
rect 16716 15922 16772 15932
rect 17388 15538 17444 16716
rect 17500 16212 17556 16222
rect 17612 16212 17668 16940
rect 17500 16210 17668 16212
rect 17500 16158 17502 16210
rect 17554 16158 17668 16210
rect 17500 16156 17668 16158
rect 17500 16146 17556 16156
rect 18060 16100 18116 17836
rect 18172 16772 18228 16782
rect 18172 16770 18340 16772
rect 18172 16718 18174 16770
rect 18226 16718 18340 16770
rect 18172 16716 18340 16718
rect 18172 16706 18228 16716
rect 18060 16034 18116 16044
rect 18284 15986 18340 16716
rect 18284 15934 18286 15986
rect 18338 15934 18340 15986
rect 18284 15922 18340 15934
rect 18620 15988 18676 15998
rect 19180 15988 19236 15998
rect 18620 15986 19236 15988
rect 18620 15934 18622 15986
rect 18674 15934 19182 15986
rect 19234 15934 19236 15986
rect 18620 15932 19236 15934
rect 18620 15922 18676 15932
rect 19180 15922 19236 15932
rect 17388 15486 17390 15538
rect 17442 15486 17444 15538
rect 17388 15474 17444 15486
rect 16828 15426 16884 15438
rect 16828 15374 16830 15426
rect 16882 15374 16884 15426
rect 16604 14478 16606 14530
rect 16658 14478 16660 14530
rect 16604 14466 16660 14478
rect 16716 15316 16772 15326
rect 16716 14532 16772 15260
rect 16828 14756 16884 15374
rect 17724 15428 17780 15438
rect 17724 15334 17780 15372
rect 16828 14690 16884 14700
rect 16940 14532 16996 14542
rect 16716 14530 16996 14532
rect 16716 14478 16942 14530
rect 16994 14478 16996 14530
rect 16716 14476 16996 14478
rect 16044 14366 16046 14418
rect 16098 14366 16100 14418
rect 15820 13748 15876 13758
rect 15820 13654 15876 13692
rect 15036 12350 15038 12402
rect 15090 12350 15092 12402
rect 15036 12338 15092 12350
rect 15596 12404 15652 12414
rect 14476 12238 14478 12290
rect 14530 12238 14532 12290
rect 14476 12226 14532 12238
rect 15596 12066 15652 12348
rect 16044 12404 16100 14366
rect 16716 13970 16772 14476
rect 16940 14466 16996 14476
rect 17724 14420 17780 14430
rect 17724 14418 18004 14420
rect 17724 14366 17726 14418
rect 17778 14366 18004 14418
rect 17724 14364 18004 14366
rect 17724 14354 17780 14364
rect 16716 13918 16718 13970
rect 16770 13918 16772 13970
rect 16716 13906 16772 13918
rect 17948 12850 18004 14364
rect 19068 13748 19124 13758
rect 18620 13524 18676 13534
rect 18284 13522 18676 13524
rect 18284 13470 18622 13522
rect 18674 13470 18676 13522
rect 18284 13468 18676 13470
rect 18284 12962 18340 13468
rect 18620 13458 18676 13468
rect 18956 13522 19012 13534
rect 18956 13470 18958 13522
rect 19010 13470 19012 13522
rect 18956 13412 19012 13470
rect 18956 13346 19012 13356
rect 19068 13186 19124 13692
rect 19068 13134 19070 13186
rect 19122 13134 19124 13186
rect 19068 13122 19124 13134
rect 18284 12910 18286 12962
rect 18338 12910 18340 12962
rect 18284 12898 18340 12910
rect 18956 12852 19012 12862
rect 17948 12798 17950 12850
rect 18002 12798 18004 12850
rect 17948 12786 18004 12798
rect 18508 12850 19012 12852
rect 18508 12798 18958 12850
rect 19010 12798 19012 12850
rect 18508 12796 19012 12798
rect 16044 12338 16100 12348
rect 15596 12014 15598 12066
rect 15650 12014 15652 12066
rect 14252 9662 14254 9714
rect 14306 9662 14308 9714
rect 14252 9604 14308 9662
rect 14700 11954 14756 11966
rect 14700 11902 14702 11954
rect 14754 11902 14756 11954
rect 14700 10724 14756 11902
rect 15596 11620 15652 12014
rect 15596 11564 15876 11620
rect 14700 9714 14756 10668
rect 14700 9662 14702 9714
rect 14754 9662 14756 9714
rect 14700 9650 14756 9662
rect 15260 11396 15316 11406
rect 15596 11396 15652 11406
rect 15260 11394 15652 11396
rect 15260 11342 15262 11394
rect 15314 11342 15598 11394
rect 15650 11342 15652 11394
rect 15260 11340 15652 11342
rect 15260 10500 15316 11340
rect 15596 11330 15652 11340
rect 14252 9538 14308 9548
rect 11004 8372 11508 8428
rect 11452 8370 11508 8372
rect 11452 8318 11454 8370
rect 11506 8318 11508 8370
rect 11452 8306 11508 8318
rect 12236 8372 12628 8428
rect 13356 8372 14084 8428
rect 15260 8372 15316 10444
rect 15372 10724 15428 10734
rect 15372 10498 15428 10668
rect 15372 10446 15374 10498
rect 15426 10446 15428 10498
rect 15372 10434 15428 10446
rect 15708 10722 15764 10734
rect 15708 10670 15710 10722
rect 15762 10670 15764 10722
rect 15708 10388 15764 10670
rect 15708 9828 15764 10332
rect 15708 9762 15764 9772
rect 15820 9604 15876 11564
rect 18508 11506 18564 12796
rect 18956 12786 19012 12796
rect 19292 12404 19348 18284
rect 20188 18228 20244 18956
rect 20188 18162 20244 18172
rect 20748 18452 20804 18462
rect 20860 18452 20916 19854
rect 20804 18396 20916 18452
rect 19292 12338 19348 12348
rect 19404 18116 19460 18126
rect 18508 11454 18510 11506
rect 18562 11454 18564 11506
rect 16380 11282 16436 11294
rect 18508 11284 18564 11454
rect 16380 11230 16382 11282
rect 16434 11230 16436 11282
rect 16380 10834 16436 11230
rect 16380 10782 16382 10834
rect 16434 10782 16436 10834
rect 16380 10770 16436 10782
rect 18396 11228 18564 11284
rect 19180 11282 19236 11294
rect 19180 11230 19182 11282
rect 19234 11230 19236 11282
rect 18396 10722 18452 11228
rect 18844 11172 18900 11182
rect 18396 10670 18398 10722
rect 18450 10670 18452 10722
rect 18396 10658 18452 10670
rect 18508 11170 18900 11172
rect 18508 11118 18846 11170
rect 18898 11118 18900 11170
rect 18508 11116 18900 11118
rect 16044 10610 16100 10622
rect 16044 10558 16046 10610
rect 16098 10558 16100 10610
rect 16044 10276 16100 10558
rect 16716 10612 16772 10622
rect 16716 10518 16772 10556
rect 17500 10612 17556 10622
rect 17500 10518 17556 10556
rect 17724 10500 17780 10510
rect 16044 9940 16100 10220
rect 17164 10388 17220 10398
rect 16380 9940 16436 9950
rect 16044 9938 16436 9940
rect 16044 9886 16382 9938
rect 16434 9886 16436 9938
rect 16044 9884 16436 9886
rect 16380 9874 16436 9884
rect 15708 9548 15876 9604
rect 10892 7868 11508 7924
rect 10220 7586 10276 7598
rect 10220 7534 10222 7586
rect 10274 7534 10276 7586
rect 10108 6804 10164 6814
rect 10220 6804 10276 7534
rect 10556 7476 10612 7486
rect 11116 7476 11172 7486
rect 10556 7474 11172 7476
rect 10556 7422 10558 7474
rect 10610 7422 11118 7474
rect 11170 7422 11172 7474
rect 10556 7420 11172 7422
rect 10556 7410 10612 7420
rect 11116 7410 11172 7420
rect 11452 7474 11508 7868
rect 11452 7422 11454 7474
rect 11506 7422 11508 7474
rect 11452 7410 11508 7422
rect 12124 7812 12180 7822
rect 12124 7474 12180 7756
rect 12124 7422 12126 7474
rect 12178 7422 12180 7474
rect 12124 7410 12180 7422
rect 12236 7586 12292 8372
rect 12236 7534 12238 7586
rect 12290 7534 12292 7586
rect 10108 6802 10276 6804
rect 10108 6750 10110 6802
rect 10162 6750 10276 6802
rect 10108 6748 10276 6750
rect 12236 6802 12292 7534
rect 13356 7474 13412 8372
rect 15260 8370 15652 8372
rect 15260 8318 15262 8370
rect 15314 8318 15652 8370
rect 15260 8316 15652 8318
rect 14140 7812 14196 7822
rect 13356 7422 13358 7474
rect 13410 7422 13412 7474
rect 13356 7410 13412 7422
rect 14028 7756 14140 7812
rect 14028 7474 14084 7756
rect 14140 7746 14196 7756
rect 14700 7700 14756 7710
rect 14700 7606 14756 7644
rect 14028 7422 14030 7474
rect 14082 7422 14084 7474
rect 14028 7410 14084 7422
rect 14140 7586 14196 7598
rect 14140 7534 14142 7586
rect 14194 7534 14196 7586
rect 13020 7252 13076 7262
rect 14140 7252 14196 7534
rect 15036 7252 15092 7262
rect 13020 7250 13412 7252
rect 13020 7198 13022 7250
rect 13074 7198 13412 7250
rect 13020 7196 13412 7198
rect 14140 7250 15092 7252
rect 14140 7198 15038 7250
rect 15090 7198 15092 7250
rect 14140 7196 15092 7198
rect 13020 7186 13076 7196
rect 12236 6750 12238 6802
rect 12290 6750 12292 6802
rect 10108 6738 10164 6748
rect 12236 6738 12292 6750
rect 9324 6598 9380 6636
rect 11788 6692 11844 6702
rect 11788 6132 11844 6636
rect 12684 6692 12740 6702
rect 13356 6692 13412 7196
rect 13692 6692 13748 6702
rect 13356 6690 13748 6692
rect 13356 6638 13694 6690
rect 13746 6638 13748 6690
rect 13356 6636 13748 6638
rect 12684 6598 12740 6636
rect 13692 6626 13748 6636
rect 13468 6468 13524 6478
rect 12908 6466 13524 6468
rect 12908 6414 13470 6466
rect 13522 6414 13524 6466
rect 12908 6412 13524 6414
rect 11788 6130 12180 6132
rect 11788 6078 11790 6130
rect 11842 6078 12180 6130
rect 11788 6076 12180 6078
rect 11788 6066 11844 6076
rect 12124 5906 12180 6076
rect 12908 6018 12964 6412
rect 13468 6402 13524 6412
rect 12908 5966 12910 6018
rect 12962 5966 12964 6018
rect 12908 5954 12964 5966
rect 12124 5854 12126 5906
rect 12178 5854 12180 5906
rect 12124 5842 12180 5854
rect 15036 5794 15092 7196
rect 15036 5742 15038 5794
rect 15090 5742 15092 5794
rect 15036 5730 15092 5742
rect 15260 6692 15316 8316
rect 15596 8258 15652 8316
rect 15596 8206 15598 8258
rect 15650 8206 15652 8258
rect 15596 8194 15652 8206
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 15260 5236 15316 6636
rect 15708 7474 15764 9548
rect 16380 8146 16436 8158
rect 16380 8094 16382 8146
rect 16434 8094 16436 8146
rect 16380 7698 16436 8094
rect 16380 7646 16382 7698
rect 16434 7646 16436 7698
rect 16380 7634 16436 7646
rect 15708 7422 15710 7474
rect 15762 7422 15764 7474
rect 15708 6356 15764 7422
rect 15820 7586 15876 7598
rect 15820 7534 15822 7586
rect 15874 7534 15876 7586
rect 15820 6580 15876 7534
rect 16716 7476 16772 7486
rect 16716 7382 16772 7420
rect 17164 6914 17220 10332
rect 17724 10052 17780 10444
rect 17836 10388 17892 10398
rect 18508 10388 18564 11116
rect 18844 11106 18900 11116
rect 19180 10834 19236 11230
rect 19180 10782 19182 10834
rect 19234 10782 19236 10834
rect 19180 10770 19236 10782
rect 18620 10612 18676 10622
rect 18620 10518 18676 10556
rect 17836 10294 17892 10332
rect 18396 10332 18564 10388
rect 17724 9996 17892 10052
rect 17724 9828 17780 9838
rect 17724 9734 17780 9772
rect 17500 7476 17556 7486
rect 17500 7382 17556 7420
rect 17836 7474 17892 9996
rect 18396 9938 18452 10332
rect 18396 9886 18398 9938
rect 18450 9886 18452 9938
rect 18396 9874 18452 9886
rect 19292 10052 19348 10062
rect 19292 9266 19348 9996
rect 19292 9214 19294 9266
rect 19346 9214 19348 9266
rect 18508 9156 18564 9166
rect 18060 8930 18116 8942
rect 18060 8878 18062 8930
rect 18114 8878 18116 8930
rect 18060 7812 18116 8878
rect 18396 8932 18452 8942
rect 18396 8838 18452 8876
rect 18060 7746 18116 7756
rect 18508 8370 18564 9100
rect 18620 9044 18676 9054
rect 18620 9042 19124 9044
rect 18620 8990 18622 9042
rect 18674 8990 19124 9042
rect 18620 8988 19124 8990
rect 18620 8978 18676 8988
rect 19068 8818 19124 8988
rect 19292 8932 19348 9214
rect 19292 8866 19348 8876
rect 19068 8766 19070 8818
rect 19122 8766 19124 8818
rect 19068 8754 19124 8766
rect 19404 8818 19460 18060
rect 19628 17668 19684 17678
rect 19628 16436 19684 17612
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20748 17106 20804 18396
rect 20748 17054 20750 17106
rect 20802 17054 20804 17106
rect 20748 17042 20804 17054
rect 19628 16370 19684 16380
rect 20300 16770 20356 16782
rect 20300 16718 20302 16770
rect 20354 16718 20356 16770
rect 19516 16324 19572 16334
rect 19516 16230 19572 16268
rect 20300 16324 20356 16718
rect 20300 16258 20356 16268
rect 21084 16212 21140 20412
rect 21420 20132 21476 20142
rect 21420 20038 21476 20076
rect 21532 20130 21588 20142
rect 21532 20078 21534 20130
rect 21586 20078 21588 20130
rect 21308 20020 21364 20030
rect 21308 19236 21364 19964
rect 21420 19908 21476 19918
rect 21532 19908 21588 20078
rect 21644 20132 21700 20142
rect 21644 20038 21700 20076
rect 21756 20132 21812 21420
rect 22092 20580 22148 21644
rect 22204 21476 22260 22316
rect 22428 22370 22484 24558
rect 22540 24612 22596 25340
rect 22540 24546 22596 24556
rect 22764 24722 22820 24734
rect 22764 24670 22766 24722
rect 22818 24670 22820 24722
rect 22764 24052 22820 24670
rect 22652 23996 22764 24052
rect 22652 22932 22708 23996
rect 22764 23986 22820 23996
rect 22764 23828 22820 23838
rect 22764 23734 22820 23772
rect 22876 23716 22932 26012
rect 22988 25732 23044 26236
rect 23324 26180 23380 26796
rect 23436 26786 23492 26796
rect 23660 26290 23716 27356
rect 23772 27076 23828 27086
rect 23772 26982 23828 27020
rect 24220 26908 24276 27694
rect 24444 26962 24500 26974
rect 24444 26910 24446 26962
rect 24498 26910 24500 26962
rect 24444 26908 24500 26910
rect 23660 26238 23662 26290
rect 23714 26238 23716 26290
rect 23660 26226 23716 26238
rect 23996 26852 24276 26908
rect 24332 26852 24500 26908
rect 23996 26290 24052 26852
rect 24220 26516 24276 26526
rect 24332 26516 24388 26852
rect 24556 26628 24612 27806
rect 24556 26562 24612 26572
rect 24220 26514 24388 26516
rect 24220 26462 24222 26514
rect 24274 26462 24388 26514
rect 24220 26460 24388 26462
rect 24220 26450 24276 26460
rect 24444 26404 24500 26414
rect 24668 26404 24724 27916
rect 24892 27076 24948 28140
rect 24892 27010 24948 27020
rect 25116 26908 25172 37548
rect 25340 37490 25396 37660
rect 25340 37438 25342 37490
rect 25394 37438 25396 37490
rect 25340 37426 25396 37438
rect 25564 37266 25620 37884
rect 25788 37490 25844 40348
rect 26124 40292 26180 41580
rect 26348 41188 26404 41694
rect 26348 41122 26404 41132
rect 26572 41186 26628 41916
rect 26796 41412 26852 41422
rect 26796 41318 26852 41356
rect 26572 41134 26574 41186
rect 26626 41134 26628 41186
rect 26572 40628 26628 41134
rect 26572 40562 26628 40572
rect 26908 41186 26964 41916
rect 27692 41972 27748 41982
rect 27692 41878 27748 41916
rect 26908 41134 26910 41186
rect 26962 41134 26964 41186
rect 26348 40404 26404 40414
rect 26348 40310 26404 40348
rect 26012 40236 26180 40292
rect 26236 40290 26292 40302
rect 26236 40238 26238 40290
rect 26290 40238 26292 40290
rect 25900 39394 25956 39406
rect 25900 39342 25902 39394
rect 25954 39342 25956 39394
rect 25900 38612 25956 39342
rect 26012 38946 26068 40236
rect 26236 40180 26292 40238
rect 26236 40114 26292 40124
rect 26796 40180 26852 40190
rect 26348 39732 26404 39742
rect 26124 39676 26348 39732
rect 26124 39058 26180 39676
rect 26348 39638 26404 39676
rect 26796 39506 26852 40124
rect 26908 39844 26964 41134
rect 27804 41746 27860 41758
rect 27804 41694 27806 41746
rect 27858 41694 27860 41746
rect 27804 41188 27860 41694
rect 27916 41188 27972 41198
rect 27804 41186 27972 41188
rect 27804 41134 27918 41186
rect 27970 41134 27972 41186
rect 27804 41132 27972 41134
rect 27916 41122 27972 41132
rect 27580 40852 27636 40862
rect 27244 40740 27300 40750
rect 27020 39844 27076 39854
rect 26908 39788 27020 39844
rect 27020 39750 27076 39788
rect 26908 39620 26964 39630
rect 26908 39526 26964 39564
rect 26796 39454 26798 39506
rect 26850 39454 26852 39506
rect 26796 39442 26852 39454
rect 26124 39006 26126 39058
rect 26178 39006 26180 39058
rect 26124 38994 26180 39006
rect 26908 39172 26964 39182
rect 26908 39058 26964 39116
rect 26908 39006 26910 39058
rect 26962 39006 26964 39058
rect 26908 38994 26964 39006
rect 26012 38894 26014 38946
rect 26066 38894 26068 38946
rect 26012 38882 26068 38894
rect 27244 38834 27300 40684
rect 27356 40514 27412 40526
rect 27356 40462 27358 40514
rect 27410 40462 27412 40514
rect 27356 40292 27412 40462
rect 27580 40514 27636 40796
rect 28028 40740 28084 43148
rect 28140 42194 28196 43596
rect 28252 43586 28308 43596
rect 28476 43540 28532 43550
rect 28476 43446 28532 43484
rect 28364 43316 28420 43326
rect 28364 43222 28420 43260
rect 28140 42142 28142 42194
rect 28194 42142 28196 42194
rect 28140 42130 28196 42142
rect 28364 42084 28420 42094
rect 28364 41970 28420 42028
rect 28364 41918 28366 41970
rect 28418 41918 28420 41970
rect 28364 41906 28420 41918
rect 28588 41748 28644 41758
rect 28588 41300 28644 41692
rect 28588 41186 28644 41244
rect 28588 41134 28590 41186
rect 28642 41134 28644 41186
rect 28588 41122 28644 41134
rect 28476 41076 28532 41086
rect 28476 40982 28532 41020
rect 28364 40964 28420 40974
rect 28028 40674 28084 40684
rect 28252 40908 28364 40964
rect 27580 40462 27582 40514
rect 27634 40462 27636 40514
rect 27580 40450 27636 40462
rect 27916 40516 27972 40526
rect 27916 40422 27972 40460
rect 27356 39956 27412 40236
rect 27468 40404 27524 40414
rect 27468 40290 27524 40348
rect 27468 40238 27470 40290
rect 27522 40238 27524 40290
rect 27468 40226 27524 40238
rect 28140 40402 28196 40414
rect 28140 40350 28142 40402
rect 28194 40350 28196 40402
rect 27356 39900 27748 39956
rect 27580 39620 27636 39630
rect 27580 39526 27636 39564
rect 27692 39506 27748 39900
rect 27916 39620 27972 39630
rect 28140 39620 28196 40350
rect 28252 40068 28308 40908
rect 28364 40870 28420 40908
rect 28364 40628 28420 40638
rect 28700 40628 28756 44828
rect 29484 44772 29540 45838
rect 29820 46228 29876 46238
rect 29708 45780 29764 45790
rect 29596 45218 29652 45230
rect 29596 45166 29598 45218
rect 29650 45166 29652 45218
rect 29596 44884 29652 45166
rect 29596 44818 29652 44828
rect 29372 44716 29540 44772
rect 28364 40534 28420 40572
rect 28588 40572 28756 40628
rect 28812 44660 28868 44670
rect 28812 40628 28868 44604
rect 29372 44322 29428 44716
rect 29596 44660 29652 44670
rect 29372 44270 29374 44322
rect 29426 44270 29428 44322
rect 29372 44258 29428 44270
rect 29484 44604 29596 44660
rect 29036 44098 29092 44110
rect 29036 44046 29038 44098
rect 29090 44046 29092 44098
rect 28924 42082 28980 42094
rect 28924 42030 28926 42082
rect 28978 42030 28980 42082
rect 28924 41860 28980 42030
rect 29036 42084 29092 44046
rect 29148 44100 29204 44110
rect 29148 44006 29204 44044
rect 29260 43988 29316 43998
rect 29260 43762 29316 43932
rect 29260 43710 29262 43762
rect 29314 43710 29316 43762
rect 29260 43698 29316 43710
rect 29036 42018 29092 42028
rect 29148 43540 29204 43550
rect 29148 42754 29204 43484
rect 29484 42868 29540 44604
rect 29596 44594 29652 44604
rect 29708 44322 29764 45724
rect 29708 44270 29710 44322
rect 29762 44270 29764 44322
rect 29708 44258 29764 44270
rect 29596 43988 29652 43998
rect 29596 43650 29652 43932
rect 29596 43598 29598 43650
rect 29650 43598 29652 43650
rect 29596 43586 29652 43598
rect 29708 43764 29764 43774
rect 29596 42868 29652 42878
rect 29484 42866 29652 42868
rect 29484 42814 29598 42866
rect 29650 42814 29652 42866
rect 29484 42812 29652 42814
rect 29596 42802 29652 42812
rect 29148 42702 29150 42754
rect 29202 42702 29204 42754
rect 29148 41860 29204 42702
rect 29708 42754 29764 43708
rect 29820 43538 29876 46172
rect 30044 45892 30100 46732
rect 30716 46788 30772 47964
rect 30716 46694 30772 46732
rect 30828 47012 30884 47022
rect 30828 46898 30884 46956
rect 30828 46846 30830 46898
rect 30882 46846 30884 46898
rect 30604 46674 30660 46686
rect 30604 46622 30606 46674
rect 30658 46622 30660 46674
rect 30044 45798 30100 45836
rect 30156 46450 30212 46462
rect 30156 46398 30158 46450
rect 30210 46398 30212 46450
rect 30044 44996 30100 45006
rect 30044 44546 30100 44940
rect 30156 44660 30212 46398
rect 30380 45890 30436 45902
rect 30380 45838 30382 45890
rect 30434 45838 30436 45890
rect 30380 44884 30436 45838
rect 30604 45892 30660 46622
rect 30604 45218 30660 45836
rect 30828 45780 30884 46846
rect 30940 46900 30996 48078
rect 31388 46900 31444 46910
rect 31500 46900 31556 48300
rect 31836 48290 31892 48300
rect 32060 48356 32116 48366
rect 32060 48242 32116 48300
rect 32060 48190 32062 48242
rect 32114 48190 32116 48242
rect 32060 48178 32116 48190
rect 32284 47572 32340 49644
rect 33180 48244 33236 49644
rect 34076 49026 34132 49038
rect 34076 48974 34078 49026
rect 34130 48974 34132 49026
rect 33292 48916 33348 48926
rect 33292 48822 33348 48860
rect 34076 48804 34132 48974
rect 34524 48804 34580 48814
rect 34076 48802 34580 48804
rect 34076 48750 34526 48802
rect 34578 48750 34580 48802
rect 34076 48748 34580 48750
rect 33740 48468 33796 48478
rect 33404 48244 33460 48254
rect 33180 48242 33460 48244
rect 33180 48190 33406 48242
rect 33458 48190 33460 48242
rect 33180 48188 33460 48190
rect 32396 47572 32452 47582
rect 32284 47516 32396 47572
rect 32396 47478 32452 47516
rect 33404 47572 33460 48188
rect 33404 47506 33460 47516
rect 30940 46834 30996 46844
rect 31164 46898 31556 46900
rect 31164 46846 31390 46898
rect 31442 46846 31556 46898
rect 31164 46844 31556 46846
rect 33180 47458 33236 47470
rect 33180 47406 33182 47458
rect 33234 47406 33236 47458
rect 31164 46674 31220 46844
rect 31164 46622 31166 46674
rect 31218 46622 31220 46674
rect 31164 46610 31220 46622
rect 31276 46116 31332 46844
rect 31388 46834 31444 46844
rect 31724 46786 31780 46798
rect 31724 46734 31726 46786
rect 31778 46734 31780 46786
rect 31612 46676 31668 46686
rect 31500 46620 31612 46676
rect 31276 46114 31444 46116
rect 31276 46062 31278 46114
rect 31330 46062 31444 46114
rect 31276 46060 31444 46062
rect 31276 46050 31332 46060
rect 30828 45714 30884 45724
rect 30604 45166 30606 45218
rect 30658 45166 30660 45218
rect 30604 45154 30660 45166
rect 30828 45108 30884 45118
rect 30380 44818 30436 44828
rect 30716 44884 30772 44894
rect 30156 44604 30660 44660
rect 30044 44494 30046 44546
rect 30098 44494 30100 44546
rect 30044 44482 30100 44494
rect 29932 44322 29988 44334
rect 29932 44270 29934 44322
rect 29986 44270 29988 44322
rect 29932 43988 29988 44270
rect 30604 44322 30660 44604
rect 30604 44270 30606 44322
rect 30658 44270 30660 44322
rect 30604 44258 30660 44270
rect 30156 44100 30212 44110
rect 30212 44044 30324 44100
rect 30156 44034 30212 44044
rect 29932 43922 29988 43932
rect 29820 43486 29822 43538
rect 29874 43486 29876 43538
rect 29820 43474 29876 43486
rect 30156 43764 30212 43774
rect 30156 43316 30212 43708
rect 30268 43428 30324 44044
rect 30380 44098 30436 44110
rect 30380 44046 30382 44098
rect 30434 44046 30436 44098
rect 30380 43540 30436 44046
rect 30716 43988 30772 44828
rect 30828 44436 30884 45052
rect 31052 45106 31108 45118
rect 31052 45054 31054 45106
rect 31106 45054 31108 45106
rect 31052 44884 31108 45054
rect 31388 45106 31444 46060
rect 31500 45778 31556 46620
rect 31612 46610 31668 46620
rect 31724 46564 31780 46734
rect 32060 46788 32116 46798
rect 32060 46694 32116 46732
rect 32172 46676 32228 46686
rect 32172 46582 32228 46620
rect 33068 46676 33124 46686
rect 33068 46582 33124 46620
rect 31780 46508 31892 46564
rect 31724 46498 31780 46508
rect 31500 45726 31502 45778
rect 31554 45726 31556 45778
rect 31500 45714 31556 45726
rect 31612 46002 31668 46014
rect 31612 45950 31614 46002
rect 31666 45950 31668 46002
rect 31612 45220 31668 45950
rect 31612 45154 31668 45164
rect 31388 45054 31390 45106
rect 31442 45054 31444 45106
rect 31388 45042 31444 45054
rect 31164 44996 31220 45006
rect 31164 44994 31332 44996
rect 31164 44942 31166 44994
rect 31218 44942 31332 44994
rect 31164 44940 31332 44942
rect 31164 44930 31220 44940
rect 31052 44818 31108 44828
rect 30828 44322 30884 44380
rect 30828 44270 30830 44322
rect 30882 44270 30884 44322
rect 30828 44258 30884 44270
rect 30940 44434 30996 44446
rect 30940 44382 30942 44434
rect 30994 44382 30996 44434
rect 30940 44324 30996 44382
rect 31164 44324 31220 44334
rect 30940 44258 30996 44268
rect 31052 44322 31220 44324
rect 31052 44270 31166 44322
rect 31218 44270 31220 44322
rect 31052 44268 31220 44270
rect 30604 43932 30772 43988
rect 30604 43764 30660 43932
rect 31052 43876 31108 44268
rect 31164 44258 31220 44268
rect 30604 43698 30660 43708
rect 30716 43820 31108 43876
rect 30604 43540 30660 43550
rect 30380 43538 30660 43540
rect 30380 43486 30606 43538
rect 30658 43486 30660 43538
rect 30380 43484 30660 43486
rect 30268 43372 30548 43428
rect 30156 43260 30436 43316
rect 29708 42702 29710 42754
rect 29762 42702 29764 42754
rect 29708 42690 29764 42702
rect 29820 43092 29876 43102
rect 29484 42532 29540 42542
rect 29260 42530 29540 42532
rect 29260 42478 29486 42530
rect 29538 42478 29540 42530
rect 29260 42476 29540 42478
rect 29260 42196 29316 42476
rect 29484 42466 29540 42476
rect 29820 42308 29876 43036
rect 29484 42252 29876 42308
rect 29932 42756 29988 42766
rect 29260 42140 29428 42196
rect 28924 41804 29204 41860
rect 29260 41970 29316 41982
rect 29260 41918 29262 41970
rect 29314 41918 29316 41970
rect 28924 40628 28980 40638
rect 28812 40626 28980 40628
rect 28812 40574 28926 40626
rect 28978 40574 28980 40626
rect 28812 40572 28980 40574
rect 28476 40180 28532 40190
rect 28476 40086 28532 40124
rect 28252 40012 28420 40068
rect 27916 39618 28196 39620
rect 27916 39566 27918 39618
rect 27970 39566 28196 39618
rect 27916 39564 28196 39566
rect 28252 39844 28308 39854
rect 28252 39618 28308 39788
rect 28252 39566 28254 39618
rect 28306 39566 28308 39618
rect 27916 39554 27972 39564
rect 28252 39554 28308 39566
rect 27692 39454 27694 39506
rect 27746 39454 27748 39506
rect 27692 39442 27748 39454
rect 28364 39508 28420 40012
rect 28476 39508 28532 39518
rect 28364 39506 28532 39508
rect 28364 39454 28478 39506
rect 28530 39454 28532 39506
rect 28364 39452 28532 39454
rect 28476 39442 28532 39452
rect 28364 39172 28420 39182
rect 28364 39058 28420 39116
rect 28364 39006 28366 39058
rect 28418 39006 28420 39058
rect 28364 38994 28420 39006
rect 28588 39060 28644 40572
rect 28924 40562 28980 40572
rect 29036 40628 29092 41804
rect 29148 41524 29204 41534
rect 29260 41524 29316 41918
rect 29204 41468 29316 41524
rect 29372 41972 29428 42140
rect 29148 41458 29204 41468
rect 29372 41412 29428 41916
rect 29372 41346 29428 41356
rect 29148 41188 29204 41198
rect 29148 41094 29204 41132
rect 29484 41074 29540 42252
rect 29820 42082 29876 42094
rect 29820 42030 29822 42082
rect 29874 42030 29876 42082
rect 29596 41748 29652 41758
rect 29596 41654 29652 41692
rect 29820 41412 29876 42030
rect 29932 41858 29988 42700
rect 30380 42754 30436 43260
rect 30380 42702 30382 42754
rect 30434 42702 30436 42754
rect 30380 42690 30436 42702
rect 30492 42642 30548 43372
rect 30492 42590 30494 42642
rect 30546 42590 30548 42642
rect 30492 42578 30548 42590
rect 30604 41972 30660 43484
rect 30716 42754 30772 43820
rect 31276 43538 31332 44940
rect 31612 44436 31668 44446
rect 31668 44380 31780 44436
rect 31612 44370 31668 44380
rect 31388 44324 31444 44334
rect 31444 44268 31556 44324
rect 31388 44258 31444 44268
rect 31276 43486 31278 43538
rect 31330 43486 31332 43538
rect 31276 43428 31332 43486
rect 31276 43362 31332 43372
rect 31388 44098 31444 44110
rect 31388 44046 31390 44098
rect 31442 44046 31444 44098
rect 30716 42702 30718 42754
rect 30770 42702 30772 42754
rect 30716 42690 30772 42702
rect 30940 43314 30996 43326
rect 30940 43262 30942 43314
rect 30994 43262 30996 43314
rect 30828 41972 30884 41982
rect 30604 41970 30884 41972
rect 30604 41918 30830 41970
rect 30882 41918 30884 41970
rect 30604 41916 30884 41918
rect 29932 41806 29934 41858
rect 29986 41806 29988 41858
rect 29932 41794 29988 41806
rect 29484 41022 29486 41074
rect 29538 41022 29540 41074
rect 29484 41010 29540 41022
rect 29596 41356 29876 41412
rect 30268 41524 30324 41534
rect 29372 40964 29428 40974
rect 29372 40852 29428 40908
rect 29596 40852 29652 41356
rect 29932 41298 29988 41310
rect 29932 41246 29934 41298
rect 29986 41246 29988 41298
rect 29820 41188 29876 41198
rect 29820 41094 29876 41132
rect 29372 40796 29652 40852
rect 29148 40628 29204 40638
rect 29092 40626 29204 40628
rect 29092 40574 29150 40626
rect 29202 40574 29204 40626
rect 29092 40572 29204 40574
rect 29036 40534 29092 40572
rect 29148 40562 29204 40572
rect 29820 40628 29876 40638
rect 29820 40534 29876 40572
rect 28700 40404 28756 40414
rect 28700 40310 28756 40348
rect 28812 40290 28868 40302
rect 28812 40238 28814 40290
rect 28866 40238 28868 40290
rect 28700 39060 28756 39070
rect 28588 39058 28756 39060
rect 28588 39006 28702 39058
rect 28754 39006 28756 39058
rect 28588 39004 28756 39006
rect 27244 38782 27246 38834
rect 27298 38782 27300 38834
rect 27244 38770 27300 38782
rect 27692 38834 27748 38846
rect 27692 38782 27694 38834
rect 27746 38782 27748 38834
rect 25900 38546 25956 38556
rect 26124 38612 26180 38622
rect 26124 38518 26180 38556
rect 27468 38612 27524 38622
rect 27468 38162 27524 38556
rect 27468 38110 27470 38162
rect 27522 38110 27524 38162
rect 27468 38098 27524 38110
rect 27692 38164 27748 38782
rect 27692 38098 27748 38108
rect 28140 38050 28196 38062
rect 28140 37998 28142 38050
rect 28194 37998 28196 38050
rect 25788 37438 25790 37490
rect 25842 37438 25844 37490
rect 25788 37426 25844 37438
rect 26796 37492 26852 37502
rect 26796 37378 26852 37436
rect 26796 37326 26798 37378
rect 26850 37326 26852 37378
rect 26796 37314 26852 37326
rect 27020 37490 27076 37502
rect 27020 37438 27022 37490
rect 27074 37438 27076 37490
rect 27020 37380 27076 37438
rect 27132 37380 27188 37390
rect 27020 37324 27132 37380
rect 25564 37214 25566 37266
rect 25618 37214 25620 37266
rect 25452 35924 25508 35934
rect 25452 34468 25508 35868
rect 25564 35252 25620 37214
rect 25676 37156 25732 37166
rect 26460 37156 26516 37166
rect 27020 37156 27076 37324
rect 27132 37314 27188 37324
rect 27580 37266 27636 37278
rect 27580 37214 27582 37266
rect 27634 37214 27636 37266
rect 25676 37154 26292 37156
rect 25676 37102 25678 37154
rect 25730 37102 26292 37154
rect 25676 37100 26292 37102
rect 25676 37090 25732 37100
rect 26236 36594 26292 37100
rect 26460 37154 27076 37156
rect 26460 37102 26462 37154
rect 26514 37102 27076 37154
rect 26460 37100 27076 37102
rect 27132 37156 27188 37166
rect 26460 37090 26516 37100
rect 26236 36542 26238 36594
rect 26290 36542 26292 36594
rect 26236 36530 26292 36542
rect 26236 36372 26292 36382
rect 25788 35812 25844 35822
rect 25788 35718 25844 35756
rect 26124 35810 26180 35822
rect 26124 35758 26126 35810
rect 26178 35758 26180 35810
rect 26124 35252 26180 35758
rect 25564 35196 26180 35252
rect 25788 34692 25844 35196
rect 25900 35028 25956 35038
rect 26236 35028 26292 36316
rect 26908 36148 26964 37100
rect 27132 37062 27188 37100
rect 27580 36932 27636 37214
rect 28140 36932 28196 37998
rect 28252 37156 28308 37166
rect 28252 37062 28308 37100
rect 28252 36932 28308 36942
rect 28140 36876 28252 36932
rect 27580 36596 27636 36876
rect 28252 36866 28308 36876
rect 28588 36932 28644 36942
rect 27020 36594 27636 36596
rect 27020 36542 27582 36594
rect 27634 36542 27636 36594
rect 27020 36540 27636 36542
rect 27020 36482 27076 36540
rect 27580 36530 27636 36540
rect 28588 36594 28644 36876
rect 28588 36542 28590 36594
rect 28642 36542 28644 36594
rect 28588 36530 28644 36542
rect 27020 36430 27022 36482
rect 27074 36430 27076 36482
rect 27020 36418 27076 36430
rect 26908 36092 27188 36148
rect 26460 35812 26516 35822
rect 26460 35718 26516 35756
rect 25900 35026 26292 35028
rect 25900 34974 25902 35026
rect 25954 34974 26238 35026
rect 26290 34974 26292 35026
rect 25900 34972 26292 34974
rect 25900 34916 25956 34972
rect 26236 34962 26292 34972
rect 27132 35026 27188 36092
rect 27244 35700 27300 35710
rect 27300 35644 27636 35700
rect 27244 35606 27300 35644
rect 27132 34974 27134 35026
rect 27186 34974 27188 35026
rect 25900 34850 25956 34860
rect 26796 34914 26852 34926
rect 26796 34862 26798 34914
rect 26850 34862 26852 34914
rect 26348 34692 26404 34702
rect 25788 34636 25956 34692
rect 25452 34354 25508 34412
rect 25452 34302 25454 34354
rect 25506 34302 25508 34354
rect 25452 34290 25508 34302
rect 25564 33572 25620 33582
rect 25564 32674 25620 33516
rect 25564 32622 25566 32674
rect 25618 32622 25620 32674
rect 25564 32610 25620 32622
rect 25676 32452 25732 32462
rect 25676 32358 25732 32396
rect 25452 31556 25508 31566
rect 25676 31556 25732 31566
rect 25508 31554 25732 31556
rect 25508 31502 25678 31554
rect 25730 31502 25732 31554
rect 25508 31500 25732 31502
rect 25228 31444 25284 31454
rect 25228 30322 25284 31388
rect 25228 30270 25230 30322
rect 25282 30270 25284 30322
rect 25228 30258 25284 30270
rect 25340 30212 25396 30222
rect 25340 29538 25396 30156
rect 25340 29486 25342 29538
rect 25394 29486 25396 29538
rect 25340 29474 25396 29486
rect 25452 30210 25508 31500
rect 25676 31490 25732 31500
rect 25452 30158 25454 30210
rect 25506 30158 25508 30210
rect 25452 29426 25508 30158
rect 25788 30098 25844 30110
rect 25788 30046 25790 30098
rect 25842 30046 25844 30098
rect 25452 29374 25454 29426
rect 25506 29374 25508 29426
rect 25452 29362 25508 29374
rect 25676 29428 25732 29438
rect 25788 29428 25844 30046
rect 25900 29876 25956 34636
rect 26348 34690 26516 34692
rect 26348 34638 26350 34690
rect 26402 34638 26516 34690
rect 26348 34636 26516 34638
rect 26348 34626 26404 34636
rect 26012 33124 26068 33134
rect 26012 32674 26068 33068
rect 26012 32622 26014 32674
rect 26066 32622 26068 32674
rect 26012 32610 26068 32622
rect 26348 32788 26404 32798
rect 26124 32564 26180 32574
rect 26124 32470 26180 32508
rect 26348 32562 26404 32732
rect 26348 32510 26350 32562
rect 26402 32510 26404 32562
rect 26348 32498 26404 32510
rect 26348 31668 26404 31678
rect 26348 31574 26404 31612
rect 26460 31332 26516 34636
rect 26796 34356 26852 34862
rect 26796 34290 26852 34300
rect 27132 33796 27188 34974
rect 27580 34914 27636 35644
rect 27580 34862 27582 34914
rect 27634 34862 27636 34914
rect 27580 34850 27636 34862
rect 28140 34916 28196 34926
rect 28140 34822 28196 34860
rect 28588 34692 28644 34702
rect 28700 34692 28756 39004
rect 28812 38836 28868 40238
rect 28812 38770 28868 38780
rect 29148 39172 29204 39182
rect 29148 39058 29204 39116
rect 29148 39006 29150 39058
rect 29202 39006 29204 39058
rect 29148 38668 29204 39006
rect 29148 38612 29540 38668
rect 29484 38050 29540 38612
rect 29484 37998 29486 38050
rect 29538 37998 29540 38050
rect 29484 37986 29540 37998
rect 29820 37940 29876 37950
rect 29820 37846 29876 37884
rect 29932 35698 29988 41246
rect 30268 41186 30324 41468
rect 30268 41134 30270 41186
rect 30322 41134 30324 41186
rect 30268 40628 30324 41134
rect 30604 41188 30660 41198
rect 30828 41188 30884 41916
rect 30660 41132 30884 41188
rect 30604 41074 30660 41132
rect 30604 41022 30606 41074
rect 30658 41022 30660 41074
rect 30604 41010 30660 41022
rect 30940 40740 30996 43262
rect 31164 42420 31220 42430
rect 31388 42420 31444 44046
rect 31164 42194 31220 42364
rect 31164 42142 31166 42194
rect 31218 42142 31220 42194
rect 31164 42130 31220 42142
rect 31276 42364 31444 42420
rect 30268 40562 30324 40572
rect 30828 40684 30996 40740
rect 30156 40514 30212 40526
rect 30156 40462 30158 40514
rect 30210 40462 30212 40514
rect 30156 38052 30212 40462
rect 30828 40292 30884 40684
rect 30940 40516 30996 40526
rect 31276 40516 31332 42364
rect 30940 40514 31332 40516
rect 30940 40462 30942 40514
rect 30994 40462 31332 40514
rect 30940 40460 31332 40462
rect 31388 42196 31444 42206
rect 30940 40450 30996 40460
rect 31388 40402 31444 42140
rect 31500 41970 31556 44268
rect 31612 44212 31668 44222
rect 31612 44118 31668 44156
rect 31724 43538 31780 44380
rect 31836 44322 31892 46508
rect 33068 45892 33124 45902
rect 33180 45892 33236 47406
rect 33740 47458 33796 48412
rect 34524 48356 34580 48748
rect 34524 48290 34580 48300
rect 34188 48132 34244 48142
rect 34188 48130 34916 48132
rect 34188 48078 34190 48130
rect 34242 48078 34916 48130
rect 34188 48076 34916 48078
rect 34188 48066 34244 48076
rect 33964 47572 34020 47582
rect 34748 47572 34804 47582
rect 33964 47570 34804 47572
rect 33964 47518 33966 47570
rect 34018 47518 34750 47570
rect 34802 47518 34804 47570
rect 33964 47516 34804 47518
rect 33964 47506 34020 47516
rect 34748 47506 34804 47516
rect 34860 47570 34916 48076
rect 34860 47518 34862 47570
rect 34914 47518 34916 47570
rect 34860 47506 34916 47518
rect 33740 47406 33742 47458
rect 33794 47406 33796 47458
rect 33740 47394 33796 47406
rect 34188 47348 34244 47358
rect 34076 47346 34244 47348
rect 34076 47294 34190 47346
rect 34242 47294 34244 47346
rect 34076 47292 34244 47294
rect 33124 45836 33236 45892
rect 33516 46562 33572 46574
rect 33516 46510 33518 46562
rect 33570 46510 33572 46562
rect 33068 45798 33124 45836
rect 33516 45332 33572 46510
rect 34076 46562 34132 47292
rect 34188 47282 34244 47292
rect 34412 47348 34468 47358
rect 34972 47348 35028 50876
rect 35084 50596 35140 51100
rect 35196 51090 35252 51100
rect 35756 51212 35924 51268
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 50596 35252 50606
rect 35084 50594 35476 50596
rect 35084 50542 35198 50594
rect 35250 50542 35476 50594
rect 35084 50540 35476 50542
rect 35196 50530 35252 50540
rect 35420 49922 35476 50540
rect 35756 50594 35812 51212
rect 36316 51156 36372 51166
rect 35756 50542 35758 50594
rect 35810 50542 35812 50594
rect 35756 50530 35812 50542
rect 35980 50820 36036 50830
rect 35868 50484 35924 50494
rect 35868 50390 35924 50428
rect 35980 50034 36036 50764
rect 36316 50818 36372 51100
rect 36540 50932 36596 51326
rect 36316 50766 36318 50818
rect 36370 50766 36372 50818
rect 36316 50754 36372 50766
rect 36428 50876 36540 50932
rect 35980 49982 35982 50034
rect 36034 49982 36036 50034
rect 35980 49970 36036 49982
rect 36092 50708 36148 50718
rect 36092 50034 36148 50652
rect 36428 50706 36484 50876
rect 36540 50866 36596 50876
rect 36652 51378 36820 51380
rect 36652 51326 36766 51378
rect 36818 51326 36820 51378
rect 36652 51324 36820 51326
rect 36428 50654 36430 50706
rect 36482 50654 36484 50706
rect 36428 50596 36484 50654
rect 36428 50530 36484 50540
rect 36652 50428 36708 51324
rect 36764 51314 36820 51324
rect 36988 51266 37044 51884
rect 37884 51938 37940 51950
rect 37884 51886 37886 51938
rect 37938 51886 37940 51938
rect 37324 51490 37380 51502
rect 37324 51438 37326 51490
rect 37378 51438 37380 51490
rect 36988 51214 36990 51266
rect 37042 51214 37044 51266
rect 36988 51202 37044 51214
rect 37100 51378 37156 51390
rect 37100 51326 37102 51378
rect 37154 51326 37156 51378
rect 37100 51268 37156 51326
rect 37100 51044 37156 51212
rect 37100 50978 37156 50988
rect 37324 50820 37380 51438
rect 37100 50764 37380 50820
rect 36092 49982 36094 50034
rect 36146 49982 36148 50034
rect 36092 49970 36148 49982
rect 36204 50372 36708 50428
rect 36988 50596 37044 50606
rect 37100 50596 37156 50764
rect 37548 50596 37604 50606
rect 36988 50594 37156 50596
rect 36988 50542 36990 50594
rect 37042 50542 37156 50594
rect 36988 50540 37156 50542
rect 37324 50594 37604 50596
rect 37324 50542 37550 50594
rect 37602 50542 37604 50594
rect 37324 50540 37604 50542
rect 36988 50372 37044 50540
rect 37324 50428 37380 50540
rect 37548 50530 37604 50540
rect 35420 49870 35422 49922
rect 35474 49870 35476 49922
rect 35420 49588 35476 49870
rect 35644 49812 35700 49822
rect 35644 49718 35700 49756
rect 36204 49588 36260 50372
rect 36988 50306 37044 50316
rect 37212 50372 37380 50428
rect 37660 50484 37716 50494
rect 36540 50148 36596 50158
rect 36316 50036 36372 50046
rect 36316 49942 36372 49980
rect 36540 49922 36596 50092
rect 37212 50036 37268 50372
rect 36540 49870 36542 49922
rect 36594 49870 36596 49922
rect 36540 49858 36596 49870
rect 36876 49922 36932 49934
rect 36876 49870 36878 49922
rect 36930 49870 36932 49922
rect 36876 49700 36932 49870
rect 37100 49924 37156 49934
rect 37100 49830 37156 49868
rect 36876 49634 36932 49644
rect 37212 49698 37268 49980
rect 37212 49646 37214 49698
rect 37266 49646 37268 49698
rect 37212 49634 37268 49646
rect 37436 50260 37492 50270
rect 37436 49810 37492 50204
rect 37660 50260 37716 50428
rect 37884 50484 37940 51886
rect 38108 51604 38164 51614
rect 38108 51510 38164 51548
rect 37884 50418 37940 50428
rect 37996 51380 38052 51390
rect 37996 50260 38052 51324
rect 38108 51156 38164 51166
rect 38108 51062 38164 51100
rect 38220 50818 38276 52892
rect 38332 52388 38388 53452
rect 38444 53442 38500 53452
rect 38780 53442 38836 53452
rect 38332 52322 38388 52332
rect 38444 53284 38500 53294
rect 38444 52946 38500 53228
rect 38668 53060 38724 53098
rect 38668 52994 38724 53004
rect 38444 52894 38446 52946
rect 38498 52894 38500 52946
rect 38444 52164 38500 52894
rect 38780 52948 38836 52958
rect 38780 52854 38836 52892
rect 38668 52836 38724 52846
rect 38556 52276 38612 52286
rect 38668 52276 38724 52780
rect 38556 52274 38724 52276
rect 38556 52222 38558 52274
rect 38610 52222 38724 52274
rect 38556 52220 38724 52222
rect 38780 52724 38836 52734
rect 38556 52210 38612 52220
rect 38220 50766 38222 50818
rect 38274 50766 38276 50818
rect 38220 50754 38276 50766
rect 38332 52108 38500 52164
rect 38332 50708 38388 52108
rect 38444 51940 38500 51950
rect 38444 51268 38500 51884
rect 38668 51938 38724 51950
rect 38668 51886 38670 51938
rect 38722 51886 38724 51938
rect 38444 51202 38500 51212
rect 38556 51378 38612 51390
rect 38556 51326 38558 51378
rect 38610 51326 38612 51378
rect 38332 50594 38388 50652
rect 38332 50542 38334 50594
rect 38386 50542 38388 50594
rect 38332 50530 38388 50542
rect 37660 50204 38052 50260
rect 38444 50482 38500 50494
rect 38444 50430 38446 50482
rect 38498 50430 38500 50482
rect 37660 50034 37716 50204
rect 38444 50148 38500 50430
rect 38444 50082 38500 50092
rect 37660 49982 37662 50034
rect 37714 49982 37716 50034
rect 37660 49970 37716 49982
rect 37996 49924 38052 49934
rect 37996 49830 38052 49868
rect 37436 49758 37438 49810
rect 37490 49758 37492 49810
rect 35420 49532 35924 49588
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35868 48916 35924 49532
rect 35980 49532 36260 49588
rect 35980 49250 36036 49532
rect 35980 49198 35982 49250
rect 36034 49198 36036 49250
rect 35980 49186 36036 49198
rect 36092 49028 36148 49038
rect 36092 48934 36148 48972
rect 37436 49028 37492 49758
rect 38556 49476 38612 51326
rect 38668 51380 38724 51886
rect 38780 51602 38836 52668
rect 38892 52388 38948 53678
rect 39228 53732 39284 53742
rect 39900 53732 39956 53742
rect 39228 53730 39508 53732
rect 39228 53678 39230 53730
rect 39282 53678 39508 53730
rect 39228 53676 39508 53678
rect 39228 53666 39284 53676
rect 39452 53170 39508 53676
rect 39900 53730 40404 53732
rect 39900 53678 39902 53730
rect 39954 53678 40404 53730
rect 39900 53676 40404 53678
rect 39900 53666 39956 53676
rect 40348 53618 40404 53676
rect 40348 53566 40350 53618
rect 40402 53566 40404 53618
rect 39452 53118 39454 53170
rect 39506 53118 39508 53170
rect 39452 53106 39508 53118
rect 39564 53506 39620 53518
rect 39564 53454 39566 53506
rect 39618 53454 39620 53506
rect 39116 53060 39172 53070
rect 39116 52500 39172 53004
rect 39228 52946 39284 52958
rect 39228 52894 39230 52946
rect 39282 52894 39284 52946
rect 39228 52612 39284 52894
rect 39564 52948 39620 53454
rect 40124 53508 40180 53518
rect 40236 53508 40292 53518
rect 40180 53506 40292 53508
rect 40180 53454 40238 53506
rect 40290 53454 40292 53506
rect 40180 53452 40292 53454
rect 39676 53172 39732 53182
rect 39676 53078 39732 53116
rect 39564 52892 39956 52948
rect 39228 52556 39844 52612
rect 38892 52332 39060 52388
rect 38892 52164 38948 52174
rect 38892 52070 38948 52108
rect 39004 51940 39060 52332
rect 39116 52386 39172 52444
rect 39116 52334 39118 52386
rect 39170 52334 39172 52386
rect 39116 52322 39172 52334
rect 39452 52388 39508 52398
rect 39452 52162 39508 52332
rect 39564 52276 39620 52286
rect 39564 52182 39620 52220
rect 39452 52110 39454 52162
rect 39506 52110 39508 52162
rect 39452 52098 39508 52110
rect 39676 52106 39732 52118
rect 39004 51874 39060 51884
rect 39340 52052 39396 52062
rect 38780 51550 38782 51602
rect 38834 51550 38836 51602
rect 38780 51538 38836 51550
rect 39116 51604 39172 51614
rect 38668 51314 38724 51324
rect 38892 51378 38948 51390
rect 38892 51326 38894 51378
rect 38946 51326 38948 51378
rect 38892 51268 38948 51326
rect 38892 51202 38948 51212
rect 38668 51044 38724 51054
rect 38668 50594 38724 50988
rect 38668 50542 38670 50594
rect 38722 50542 38724 50594
rect 38668 50530 38724 50542
rect 38892 50708 38948 50718
rect 38780 50484 38836 50494
rect 38780 49810 38836 50428
rect 38892 50482 38948 50652
rect 39004 50596 39060 50606
rect 39004 50502 39060 50540
rect 38892 50430 38894 50482
rect 38946 50430 38948 50482
rect 38892 50418 38948 50430
rect 39116 50428 39172 51548
rect 39228 51492 39284 51502
rect 39228 51044 39284 51436
rect 39340 51380 39396 51996
rect 39676 52054 39678 52106
rect 39730 52054 39732 52106
rect 39676 52052 39732 52054
rect 39676 51986 39732 51996
rect 39788 52050 39844 52556
rect 39788 51998 39790 52050
rect 39842 51998 39844 52050
rect 39340 51314 39396 51324
rect 39564 51492 39620 51502
rect 39564 51378 39620 51436
rect 39564 51326 39566 51378
rect 39618 51326 39620 51378
rect 39564 51314 39620 51326
rect 39452 51156 39508 51166
rect 39452 51062 39508 51100
rect 39228 50978 39284 50988
rect 39564 51044 39620 51054
rect 39340 50820 39396 50830
rect 39116 50372 39284 50428
rect 39228 50036 39284 50372
rect 39228 49970 39284 49980
rect 39228 49812 39284 49822
rect 38780 49758 38782 49810
rect 38834 49758 38836 49810
rect 38780 49746 38836 49758
rect 39116 49810 39284 49812
rect 39116 49758 39230 49810
rect 39282 49758 39284 49810
rect 39116 49756 39284 49758
rect 39116 49700 39172 49756
rect 39228 49746 39284 49756
rect 38556 49420 38724 49476
rect 37436 48962 37492 48972
rect 35980 48916 36036 48926
rect 35868 48914 36036 48916
rect 35868 48862 35982 48914
rect 36034 48862 36036 48914
rect 35868 48860 36036 48862
rect 35980 48850 36036 48860
rect 38668 48916 38724 49420
rect 38668 48850 38724 48860
rect 39004 48804 39060 48814
rect 39116 48804 39172 49644
rect 39340 49026 39396 50764
rect 39452 50372 39508 50382
rect 39452 50278 39508 50316
rect 39340 48974 39342 49026
rect 39394 48974 39396 49026
rect 39340 48962 39396 48974
rect 39452 49252 39508 49262
rect 39060 48748 39172 48804
rect 39228 48916 39284 48926
rect 39004 48710 39060 48748
rect 39228 48466 39284 48860
rect 39452 48692 39508 49196
rect 39564 49138 39620 50988
rect 39676 50484 39732 50494
rect 39676 49700 39732 50428
rect 39676 49634 39732 49644
rect 39788 49586 39844 51998
rect 39900 51604 39956 52892
rect 39900 51538 39956 51548
rect 40012 52722 40068 52734
rect 40012 52670 40014 52722
rect 40066 52670 40068 52722
rect 40012 51492 40068 52670
rect 40124 51828 40180 53452
rect 40236 53442 40292 53452
rect 40236 52948 40292 52958
rect 40348 52948 40404 53566
rect 41020 53060 41076 53070
rect 41244 53060 41300 54574
rect 42140 54402 42196 55246
rect 42140 54350 42142 54402
rect 42194 54350 42196 54402
rect 42140 53732 42196 54350
rect 42476 54402 42532 56030
rect 42924 55970 42980 56812
rect 42924 55918 42926 55970
rect 42978 55918 42980 55970
rect 42924 55906 42980 55918
rect 43036 55972 43092 59200
rect 43036 55906 43092 55916
rect 43484 55412 43540 59200
rect 43596 57092 43652 57102
rect 43596 55970 43652 57036
rect 44380 56642 44436 59200
rect 44828 57764 44884 59200
rect 44828 57708 45332 57764
rect 44380 56590 44382 56642
rect 44434 56590 44436 56642
rect 44380 56578 44436 56590
rect 44940 56642 44996 56654
rect 44940 56590 44942 56642
rect 44994 56590 44996 56642
rect 44044 56308 44100 56318
rect 44044 56214 44100 56252
rect 43596 55918 43598 55970
rect 43650 55918 43652 55970
rect 43596 55906 43652 55918
rect 44492 55972 44548 55982
rect 44492 55878 44548 55916
rect 44940 55970 44996 56590
rect 45276 56308 45332 57708
rect 45388 56308 45444 56318
rect 45276 56306 45444 56308
rect 45276 56254 45390 56306
rect 45442 56254 45444 56306
rect 45276 56252 45444 56254
rect 45388 56242 45444 56252
rect 44940 55918 44942 55970
rect 44994 55918 44996 55970
rect 44940 55906 44996 55918
rect 45724 55972 45780 59200
rect 46172 56308 46228 59200
rect 46396 56308 46452 56318
rect 46172 56306 46452 56308
rect 46172 56254 46398 56306
rect 46450 56254 46452 56306
rect 46172 56252 46452 56254
rect 46396 56242 46452 56252
rect 45948 55972 46004 55982
rect 45724 55970 46004 55972
rect 45724 55918 45950 55970
rect 46002 55918 46004 55970
rect 45724 55916 46004 55918
rect 47068 55972 47124 59200
rect 47516 57764 47572 59200
rect 47516 57708 47908 57764
rect 47852 56306 47908 57708
rect 47852 56254 47854 56306
rect 47906 56254 47908 56306
rect 47852 56242 47908 56254
rect 47404 55972 47460 55982
rect 47068 55970 47460 55972
rect 47068 55918 47406 55970
rect 47458 55918 47460 55970
rect 47068 55916 47460 55918
rect 48412 55972 48468 59200
rect 48860 56308 48916 59200
rect 49084 56308 49140 56318
rect 48860 56306 49140 56308
rect 48860 56254 49086 56306
rect 49138 56254 49140 56306
rect 48860 56252 49140 56254
rect 49084 56242 49140 56252
rect 48636 55972 48692 55982
rect 48412 55970 48692 55972
rect 48412 55918 48638 55970
rect 48690 55918 48692 55970
rect 48412 55916 48692 55918
rect 49756 55972 49812 59200
rect 50204 56308 50260 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 50428 56308 50484 56318
rect 50204 56306 50484 56308
rect 50204 56254 50430 56306
rect 50482 56254 50484 56306
rect 50204 56252 50484 56254
rect 50428 56242 50484 56252
rect 49980 55972 50036 55982
rect 49756 55970 50036 55972
rect 49756 55918 49982 55970
rect 50034 55918 50036 55970
rect 49756 55916 50036 55918
rect 51100 55972 51156 59200
rect 51548 56308 51604 59200
rect 51772 56308 51828 56318
rect 51548 56306 51828 56308
rect 51548 56254 51774 56306
rect 51826 56254 51828 56306
rect 51548 56252 51828 56254
rect 51772 56242 51828 56252
rect 51324 55972 51380 55982
rect 51100 55970 51380 55972
rect 51100 55918 51326 55970
rect 51378 55918 51380 55970
rect 51100 55916 51380 55918
rect 52444 55972 52500 59200
rect 52892 56308 52948 59200
rect 53116 56308 53172 56318
rect 52892 56306 53172 56308
rect 52892 56254 53118 56306
rect 53170 56254 53172 56306
rect 52892 56252 53172 56254
rect 53116 56242 53172 56252
rect 52668 55972 52724 55982
rect 52444 55970 52724 55972
rect 52444 55918 52670 55970
rect 52722 55918 52724 55970
rect 52444 55916 52724 55918
rect 53788 55972 53844 59200
rect 54236 56866 54292 59200
rect 54236 56814 54238 56866
rect 54290 56814 54292 56866
rect 54236 56802 54292 56814
rect 55020 56866 55076 56878
rect 55020 56814 55022 56866
rect 55074 56814 55076 56866
rect 55020 56306 55076 56814
rect 55020 56254 55022 56306
rect 55074 56254 55076 56306
rect 55020 56242 55076 56254
rect 55132 56196 55188 59200
rect 55580 57316 55636 59200
rect 55580 57260 55972 57316
rect 55916 56306 55972 57260
rect 55916 56254 55918 56306
rect 55970 56254 55972 56306
rect 55916 56242 55972 56254
rect 55132 56140 55412 56196
rect 54012 55972 54068 55982
rect 53788 55970 54068 55972
rect 53788 55918 54014 55970
rect 54066 55918 54068 55970
rect 53788 55916 54068 55918
rect 55356 55972 55412 56140
rect 55468 55972 55524 55982
rect 55356 55970 55524 55972
rect 55356 55918 55470 55970
rect 55522 55918 55524 55970
rect 55356 55916 55524 55918
rect 45948 55906 46004 55916
rect 47404 55906 47460 55916
rect 48636 55906 48692 55916
rect 49980 55906 50036 55916
rect 51324 55906 51380 55916
rect 52668 55906 52724 55916
rect 54012 55906 54068 55916
rect 55468 55906 55524 55916
rect 43484 55356 43988 55412
rect 42588 55188 42644 55198
rect 42588 55094 42644 55132
rect 42700 55186 42756 55198
rect 43260 55188 43316 55198
rect 42700 55134 42702 55186
rect 42754 55134 42756 55186
rect 42700 55076 42756 55134
rect 42700 55010 42756 55020
rect 42924 55186 43316 55188
rect 42924 55134 43262 55186
rect 43314 55134 43316 55186
rect 42924 55132 43316 55134
rect 42476 54350 42478 54402
rect 42530 54350 42532 54402
rect 42476 54338 42532 54350
rect 42924 53842 42980 55132
rect 43260 55122 43316 55132
rect 43932 55186 43988 55356
rect 43932 55134 43934 55186
rect 43986 55134 43988 55186
rect 43932 55122 43988 55134
rect 43596 55076 43652 55086
rect 43596 54982 43652 55020
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 44604 54628 44660 54638
rect 44604 54534 44660 54572
rect 45388 54514 45444 54526
rect 45388 54462 45390 54514
rect 45442 54462 45444 54514
rect 45388 54404 45444 54462
rect 45836 54404 45892 54414
rect 45388 54348 45836 54404
rect 42924 53790 42926 53842
rect 42978 53790 42980 53842
rect 42924 53778 42980 53790
rect 43260 53842 43316 53854
rect 43260 53790 43262 53842
rect 43314 53790 43316 53842
rect 42140 53666 42196 53676
rect 42028 53284 42084 53294
rect 42084 53228 42196 53284
rect 42028 53218 42084 53228
rect 41916 53060 41972 53070
rect 41020 53058 41188 53060
rect 41020 53006 41022 53058
rect 41074 53006 41188 53058
rect 41020 53004 41188 53006
rect 41020 52994 41076 53004
rect 40908 52948 40964 52958
rect 40292 52892 40404 52948
rect 40460 52946 40964 52948
rect 40460 52894 40910 52946
rect 40962 52894 40964 52946
rect 40460 52892 40964 52894
rect 40236 52854 40292 52892
rect 40236 52388 40292 52398
rect 40236 52162 40292 52332
rect 40236 52110 40238 52162
rect 40290 52110 40292 52162
rect 40236 52098 40292 52110
rect 40348 52164 40404 52174
rect 40460 52164 40516 52892
rect 40908 52882 40964 52892
rect 41020 52722 41076 52734
rect 41020 52670 41022 52722
rect 41074 52670 41076 52722
rect 40404 52108 40516 52164
rect 40684 52500 40740 52510
rect 40684 52162 40740 52444
rect 41020 52388 41076 52670
rect 41020 52322 41076 52332
rect 41132 52276 41188 53004
rect 41300 53004 41524 53060
rect 41244 52994 41300 53004
rect 41356 52276 41412 52286
rect 41132 52274 41412 52276
rect 41132 52222 41358 52274
rect 41410 52222 41412 52274
rect 41132 52220 41412 52222
rect 40684 52110 40686 52162
rect 40738 52110 40740 52162
rect 40348 51940 40404 52108
rect 40684 52098 40740 52110
rect 41020 52164 41076 52174
rect 41132 52164 41188 52220
rect 41020 52162 41188 52164
rect 41020 52110 41022 52162
rect 41074 52110 41188 52162
rect 41020 52108 41188 52110
rect 41020 52098 41076 52108
rect 40124 51762 40180 51772
rect 40236 51884 40404 51940
rect 40796 51940 40852 51950
rect 40012 51426 40068 51436
rect 40124 51490 40180 51502
rect 40124 51438 40126 51490
rect 40178 51438 40180 51490
rect 40124 51380 40180 51438
rect 39900 51156 39956 51166
rect 39900 51154 40068 51156
rect 39900 51102 39902 51154
rect 39954 51102 40068 51154
rect 39900 51100 40068 51102
rect 39900 51090 39956 51100
rect 39900 50482 39956 50494
rect 39900 50430 39902 50482
rect 39954 50430 39956 50482
rect 39900 50372 39956 50430
rect 39900 50306 39956 50316
rect 39900 50036 39956 50046
rect 39900 49810 39956 49980
rect 39900 49758 39902 49810
rect 39954 49758 39956 49810
rect 39900 49746 39956 49758
rect 40012 49924 40068 51100
rect 40124 50820 40180 51324
rect 40236 51266 40292 51884
rect 40236 51214 40238 51266
rect 40290 51214 40292 51266
rect 40236 51202 40292 51214
rect 40124 50754 40180 50764
rect 40236 51044 40292 51054
rect 40124 50484 40180 50494
rect 40124 50390 40180 50428
rect 40012 49588 40068 49868
rect 39788 49534 39790 49586
rect 39842 49534 39844 49586
rect 39788 49522 39844 49534
rect 39900 49532 40068 49588
rect 40236 50372 40292 50988
rect 40796 50706 40852 51884
rect 40908 51938 40964 51950
rect 40908 51886 40910 51938
rect 40962 51886 40964 51938
rect 40908 51604 40964 51886
rect 40908 51538 40964 51548
rect 41020 51828 41076 51838
rect 41356 51828 41412 52220
rect 41468 52050 41524 53004
rect 41916 52966 41972 53004
rect 42028 52162 42084 52174
rect 42028 52110 42030 52162
rect 42082 52110 42084 52162
rect 41468 51998 41470 52050
rect 41522 51998 41524 52050
rect 41468 51986 41524 51998
rect 41692 52052 41748 52062
rect 41692 51958 41748 51996
rect 41356 51772 41636 51828
rect 40796 50654 40798 50706
rect 40850 50654 40852 50706
rect 40796 50642 40852 50654
rect 40460 50594 40516 50606
rect 40460 50542 40462 50594
rect 40514 50542 40516 50594
rect 40460 50484 40516 50542
rect 40460 50418 40516 50428
rect 41020 50482 41076 51772
rect 41356 51604 41412 51614
rect 41356 51378 41412 51548
rect 41356 51326 41358 51378
rect 41410 51326 41412 51378
rect 41356 51314 41412 51326
rect 41580 51378 41636 51772
rect 42028 51492 42084 52110
rect 42140 51938 42196 53228
rect 42252 53058 42308 53070
rect 42252 53006 42254 53058
rect 42306 53006 42308 53058
rect 42252 52948 42308 53006
rect 42588 53060 42644 53070
rect 42588 52966 42644 53004
rect 42252 52882 42308 52892
rect 43036 52834 43092 52846
rect 43036 52782 43038 52834
rect 43090 52782 43092 52834
rect 43036 52612 43092 52782
rect 43260 52836 43316 53790
rect 43484 53730 43540 53742
rect 43484 53678 43486 53730
rect 43538 53678 43540 53730
rect 43372 52836 43428 52846
rect 43260 52780 43372 52836
rect 43372 52770 43428 52780
rect 43484 52612 43540 53678
rect 44828 53732 44884 53742
rect 44828 53638 44884 53676
rect 45276 53732 45332 53742
rect 45388 53732 45444 54348
rect 45836 54310 45892 54348
rect 48076 54404 48132 54414
rect 48132 54348 48468 54404
rect 45332 53676 45444 53732
rect 45276 53666 45332 53676
rect 43036 52556 43540 52612
rect 43596 52948 43652 52958
rect 43036 52276 43092 52556
rect 42700 52220 43092 52276
rect 43484 52276 43540 52286
rect 42364 52052 42420 52062
rect 42140 51886 42142 51938
rect 42194 51886 42196 51938
rect 42140 51874 42196 51886
rect 42252 51996 42364 52052
rect 42140 51492 42196 51502
rect 42084 51490 42196 51492
rect 42084 51438 42142 51490
rect 42194 51438 42196 51490
rect 42084 51436 42196 51438
rect 42028 51398 42084 51436
rect 42140 51426 42196 51436
rect 41580 51326 41582 51378
rect 41634 51326 41636 51378
rect 41580 51314 41636 51326
rect 41916 51154 41972 51166
rect 41916 51102 41918 51154
rect 41970 51102 41972 51154
rect 41020 50430 41022 50482
rect 41074 50430 41076 50482
rect 41020 50418 41076 50430
rect 41132 50932 41188 50942
rect 41132 50594 41188 50876
rect 41132 50542 41134 50594
rect 41186 50542 41188 50594
rect 39564 49086 39566 49138
rect 39618 49086 39620 49138
rect 39564 49074 39620 49086
rect 39228 48414 39230 48466
rect 39282 48414 39284 48466
rect 39228 48402 39284 48414
rect 39340 48636 39508 48692
rect 39340 48354 39396 48636
rect 39676 48468 39732 48478
rect 39900 48468 39956 49532
rect 39676 48466 39956 48468
rect 39676 48414 39678 48466
rect 39730 48414 39956 48466
rect 39676 48412 39956 48414
rect 40012 49252 40068 49262
rect 40012 48466 40068 49196
rect 40124 48916 40180 48926
rect 40236 48916 40292 50316
rect 40124 48914 40292 48916
rect 40124 48862 40126 48914
rect 40178 48862 40292 48914
rect 40124 48860 40292 48862
rect 40684 49924 40740 49934
rect 40684 48914 40740 49868
rect 40908 49700 40964 49710
rect 40796 49028 40852 49038
rect 40908 49028 40964 49644
rect 40796 49026 40964 49028
rect 40796 48974 40798 49026
rect 40850 48974 40964 49026
rect 40796 48972 40964 48974
rect 40796 48962 40852 48972
rect 40684 48862 40686 48914
rect 40738 48862 40740 48914
rect 40124 48850 40180 48860
rect 40684 48850 40740 48862
rect 41132 48914 41188 50542
rect 41916 50596 41972 51102
rect 41916 50530 41972 50540
rect 42140 50708 42196 50718
rect 41580 50484 41636 50494
rect 41580 50390 41636 50428
rect 42028 50484 42084 50494
rect 41356 50370 41412 50382
rect 41356 50318 41358 50370
rect 41410 50318 41412 50370
rect 41356 49924 41412 50318
rect 42028 49924 42084 50428
rect 42140 50148 42196 50652
rect 42252 50594 42308 51996
rect 42364 51986 42420 51996
rect 42476 52052 42532 52062
rect 42700 52052 42756 52220
rect 42476 52050 42756 52052
rect 42476 51998 42478 52050
rect 42530 51998 42756 52050
rect 42476 51996 42756 51998
rect 42812 52052 42868 52062
rect 42364 51044 42420 51054
rect 42476 51044 42532 51996
rect 42812 51490 42868 51996
rect 43372 51940 43428 51950
rect 42812 51438 42814 51490
rect 42866 51438 42868 51490
rect 42812 51426 42868 51438
rect 42924 51938 43428 51940
rect 42924 51886 43374 51938
rect 43426 51886 43428 51938
rect 42924 51884 43428 51886
rect 42924 51156 42980 51884
rect 43372 51874 43428 51884
rect 43372 51604 43428 51614
rect 43036 51490 43092 51502
rect 43036 51438 43038 51490
rect 43090 51438 43092 51490
rect 43036 51380 43092 51438
rect 43372 51380 43428 51548
rect 43036 51314 43092 51324
rect 43148 51378 43428 51380
rect 43148 51326 43374 51378
rect 43426 51326 43428 51378
rect 43148 51324 43428 51326
rect 42420 50988 42532 51044
rect 42588 51100 42980 51156
rect 42364 50978 42420 50988
rect 42252 50542 42254 50594
rect 42306 50542 42308 50594
rect 42252 50484 42308 50542
rect 42252 50418 42308 50428
rect 42476 50820 42532 50830
rect 42476 50706 42532 50764
rect 42588 50818 42644 51100
rect 43148 51044 43204 51324
rect 43372 51314 43428 51324
rect 42588 50766 42590 50818
rect 42642 50766 42644 50818
rect 42588 50754 42644 50766
rect 42924 50988 43204 51044
rect 42476 50654 42478 50706
rect 42530 50654 42532 50706
rect 42476 50260 42532 50654
rect 42924 50482 42980 50988
rect 43484 50708 43540 52220
rect 43596 52050 43652 52892
rect 44044 52836 44100 52846
rect 45388 52836 45444 53676
rect 47740 53842 47796 53854
rect 47740 53790 47742 53842
rect 47794 53790 47796 53842
rect 45612 53618 45668 53630
rect 45612 53566 45614 53618
rect 45666 53566 45668 53618
rect 45612 53170 45668 53566
rect 45612 53118 45614 53170
rect 45666 53118 45668 53170
rect 45612 53106 45668 53118
rect 45500 53058 45556 53070
rect 45500 53006 45502 53058
rect 45554 53006 45556 53058
rect 45500 52948 45556 53006
rect 46060 52948 46116 52958
rect 45500 52946 46116 52948
rect 45500 52894 46062 52946
rect 46114 52894 46116 52946
rect 45500 52892 46116 52894
rect 45388 52780 45556 52836
rect 43596 51998 43598 52050
rect 43650 51998 43652 52050
rect 43596 51986 43652 51998
rect 43708 52050 43764 52062
rect 43708 51998 43710 52050
rect 43762 51998 43764 52050
rect 43708 51604 43764 51998
rect 43932 51604 43988 51614
rect 43708 51538 43764 51548
rect 43820 51548 43932 51604
rect 43820 51490 43876 51548
rect 43820 51438 43822 51490
rect 43874 51438 43876 51490
rect 43820 51426 43876 51438
rect 43708 51380 43764 51390
rect 43596 51378 43764 51380
rect 43596 51326 43710 51378
rect 43762 51326 43764 51378
rect 43596 51324 43764 51326
rect 43596 50932 43652 51324
rect 43708 51314 43764 51324
rect 43820 51156 43876 51166
rect 43820 51062 43876 51100
rect 43596 50866 43652 50876
rect 43708 51044 43764 51054
rect 43260 50652 43540 50708
rect 43260 50596 43316 50652
rect 42924 50430 42926 50482
rect 42978 50430 42980 50482
rect 42924 50418 42980 50430
rect 43036 50594 43316 50596
rect 43036 50542 43262 50594
rect 43314 50542 43316 50594
rect 43036 50540 43316 50542
rect 42476 50194 42532 50204
rect 42140 50092 42420 50148
rect 42028 49868 42308 49924
rect 41356 49858 41412 49868
rect 41468 49812 41524 49822
rect 41468 49026 41524 49756
rect 42140 49252 42196 49262
rect 42252 49252 42308 49868
rect 42364 49810 42420 50092
rect 42476 50034 42532 50046
rect 42476 49982 42478 50034
rect 42530 49982 42532 50034
rect 42476 49924 42532 49982
rect 42476 49858 42532 49868
rect 43036 49922 43092 50540
rect 43260 50530 43316 50540
rect 43596 50484 43652 50494
rect 43372 50482 43652 50484
rect 43372 50430 43598 50482
rect 43650 50430 43652 50482
rect 43372 50428 43652 50430
rect 43372 50372 43428 50428
rect 43596 50418 43652 50428
rect 43372 50306 43428 50316
rect 43596 50148 43652 50158
rect 43036 49870 43038 49922
rect 43090 49870 43092 49922
rect 43036 49858 43092 49870
rect 43372 50036 43428 50046
rect 42364 49758 42366 49810
rect 42418 49758 42420 49810
rect 42364 49746 42420 49758
rect 42588 49812 42644 49822
rect 43148 49812 43204 49822
rect 42588 49810 42980 49812
rect 42588 49758 42590 49810
rect 42642 49758 42980 49810
rect 42588 49756 42980 49758
rect 42588 49746 42644 49756
rect 42140 49250 42308 49252
rect 42140 49198 42142 49250
rect 42194 49198 42308 49250
rect 42140 49196 42308 49198
rect 42924 49252 42980 49756
rect 43148 49718 43204 49756
rect 43372 49810 43428 49980
rect 43596 50034 43652 50092
rect 43596 49982 43598 50034
rect 43650 49982 43652 50034
rect 43596 49970 43652 49982
rect 43372 49758 43374 49810
rect 43426 49758 43428 49810
rect 43372 49746 43428 49758
rect 42140 49186 42196 49196
rect 42924 49158 42980 49196
rect 43596 49476 43652 49486
rect 41468 48974 41470 49026
rect 41522 48974 41524 49026
rect 41468 48962 41524 48974
rect 43260 49028 43316 49038
rect 43260 48934 43316 48972
rect 41132 48862 41134 48914
rect 41186 48862 41188 48914
rect 41132 48850 41188 48862
rect 41804 48916 41860 48926
rect 41804 48822 41860 48860
rect 42028 48804 42084 48814
rect 42028 48710 42084 48748
rect 40012 48414 40014 48466
rect 40066 48414 40068 48466
rect 39676 48402 39732 48412
rect 40012 48402 40068 48414
rect 39340 48302 39342 48354
rect 39394 48302 39396 48354
rect 39340 48290 39396 48302
rect 41356 48356 41412 48366
rect 36316 48132 36372 48142
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 34412 47254 34468 47292
rect 34860 47292 35028 47348
rect 35084 47458 35140 47470
rect 35084 47406 35086 47458
rect 35138 47406 35140 47458
rect 34076 46510 34078 46562
rect 34130 46510 34132 46562
rect 33852 45892 33908 45902
rect 33516 45276 33684 45332
rect 31948 45220 32004 45230
rect 31948 45126 32004 45164
rect 32284 45108 32340 45146
rect 33180 45108 33236 45118
rect 33516 45108 33572 45118
rect 32284 45042 32340 45052
rect 32396 45106 33572 45108
rect 32396 45054 33182 45106
rect 33234 45054 33518 45106
rect 33570 45054 33572 45106
rect 32396 45052 33572 45054
rect 31836 44270 31838 44322
rect 31890 44270 31892 44322
rect 31836 44258 31892 44270
rect 32060 44994 32116 45006
rect 32060 44942 32062 44994
rect 32114 44942 32116 44994
rect 32060 43876 32116 44942
rect 32396 44772 32452 45052
rect 33180 45042 33236 45052
rect 33516 45042 33572 45052
rect 32060 43810 32116 43820
rect 32172 44716 32452 44772
rect 33516 44884 33572 44894
rect 33628 44884 33684 45276
rect 33572 44828 33684 44884
rect 33740 45106 33796 45118
rect 33740 45054 33742 45106
rect 33794 45054 33796 45106
rect 31724 43486 31726 43538
rect 31778 43486 31780 43538
rect 31724 43474 31780 43486
rect 32172 42644 32228 44716
rect 32396 44548 32452 44558
rect 32284 44212 32340 44222
rect 32284 44118 32340 44156
rect 32396 42868 32452 44492
rect 32620 44436 32676 44446
rect 32620 44434 33460 44436
rect 32620 44382 32622 44434
rect 32674 44382 33460 44434
rect 32620 44380 33460 44382
rect 32620 44370 32676 44380
rect 33404 44322 33460 44380
rect 33404 44270 33406 44322
rect 33458 44270 33460 44322
rect 33404 44258 33460 44270
rect 33180 44210 33236 44222
rect 33180 44158 33182 44210
rect 33234 44158 33236 44210
rect 32396 42802 32452 42812
rect 32508 44098 32564 44110
rect 32508 44046 32510 44098
rect 32562 44046 32564 44098
rect 32508 43540 32564 44046
rect 33180 44100 33236 44158
rect 33516 44100 33572 44828
rect 33740 44660 33796 45054
rect 33740 44594 33796 44604
rect 33628 44548 33684 44558
rect 33628 44434 33684 44492
rect 33628 44382 33630 44434
rect 33682 44382 33684 44434
rect 33628 44370 33684 44382
rect 33628 44212 33684 44222
rect 33628 44118 33684 44156
rect 33180 44044 33572 44100
rect 33740 44098 33796 44110
rect 33740 44046 33742 44098
rect 33794 44046 33796 44098
rect 33740 43988 33796 44046
rect 33516 43932 33796 43988
rect 33404 43652 33460 43662
rect 33516 43652 33572 43932
rect 33852 43876 33908 45836
rect 33964 45220 34020 45230
rect 33964 45126 34020 45164
rect 33404 43650 33572 43652
rect 33404 43598 33406 43650
rect 33458 43598 33572 43650
rect 33404 43596 33572 43598
rect 33628 43820 33908 43876
rect 33068 43540 33124 43550
rect 32508 43538 33124 43540
rect 32508 43486 33070 43538
rect 33122 43486 33124 43538
rect 32508 43484 33124 43486
rect 31948 42588 32228 42644
rect 31948 42420 32004 42588
rect 31836 42364 32004 42420
rect 32172 42420 32228 42430
rect 31500 41918 31502 41970
rect 31554 41918 31556 41970
rect 31500 41906 31556 41918
rect 31724 41972 31780 41982
rect 31724 41878 31780 41916
rect 31836 41860 31892 42364
rect 31948 42196 32004 42206
rect 31948 42102 32004 42140
rect 32172 42194 32228 42364
rect 32172 42142 32174 42194
rect 32226 42142 32228 42194
rect 32172 42130 32228 42142
rect 32060 41972 32116 41982
rect 32508 41972 32564 43484
rect 33068 43474 33124 43484
rect 33404 43540 33460 43596
rect 32620 42530 32676 42542
rect 32620 42478 32622 42530
rect 32674 42478 32676 42530
rect 32620 42196 32676 42478
rect 32620 42130 32676 42140
rect 33292 42084 33348 42094
rect 33292 41990 33348 42028
rect 32060 41970 32452 41972
rect 32060 41918 32062 41970
rect 32114 41918 32452 41970
rect 32060 41916 32452 41918
rect 32060 41906 32116 41916
rect 31836 41804 32004 41860
rect 31948 41412 32004 41804
rect 32396 41748 32452 41916
rect 32508 41906 32564 41916
rect 33180 41858 33236 41870
rect 33180 41806 33182 41858
rect 33234 41806 33236 41858
rect 33068 41748 33124 41758
rect 32396 41746 33124 41748
rect 32396 41694 33070 41746
rect 33122 41694 33124 41746
rect 32396 41692 33124 41694
rect 33068 41682 33124 41692
rect 33180 41412 33236 41806
rect 31948 41356 32116 41412
rect 31948 41188 32004 41198
rect 31388 40350 31390 40402
rect 31442 40350 31444 40402
rect 31388 40338 31444 40350
rect 31612 41186 32004 41188
rect 31612 41134 31950 41186
rect 32002 41134 32004 41186
rect 31612 41132 32004 41134
rect 31612 40628 31668 41132
rect 31948 41122 32004 41132
rect 31836 40964 31892 40974
rect 30828 40236 30996 40292
rect 30492 39956 30548 39966
rect 30492 39060 30548 39900
rect 30492 38722 30548 39004
rect 30492 38670 30494 38722
rect 30546 38670 30548 38722
rect 30492 38658 30548 38670
rect 30828 38834 30884 38846
rect 30828 38782 30830 38834
rect 30882 38782 30884 38834
rect 30828 38668 30884 38782
rect 30716 38612 30884 38668
rect 30940 38668 30996 40236
rect 31500 39620 31556 39630
rect 31612 39620 31668 40572
rect 31724 40852 31780 40862
rect 31724 39732 31780 40796
rect 31836 40626 31892 40908
rect 31836 40574 31838 40626
rect 31890 40574 31892 40626
rect 31836 40562 31892 40574
rect 31724 39666 31780 39676
rect 31948 40402 32004 40414
rect 31948 40350 31950 40402
rect 32002 40350 32004 40402
rect 31500 39618 31668 39620
rect 31500 39566 31502 39618
rect 31554 39566 31668 39618
rect 31500 39564 31668 39566
rect 31948 39620 32004 40350
rect 30940 38612 31220 38668
rect 30212 37996 30324 38052
rect 30156 37986 30212 37996
rect 30156 36372 30212 36382
rect 30156 36278 30212 36316
rect 30268 35924 30324 37996
rect 30380 37940 30436 37950
rect 30380 37846 30436 37884
rect 30716 37938 30772 38612
rect 31052 38050 31108 38062
rect 31052 37998 31054 38050
rect 31106 37998 31108 38050
rect 31052 37940 31108 37998
rect 30716 37886 30718 37938
rect 30770 37886 30772 37938
rect 30380 37154 30436 37166
rect 30380 37102 30382 37154
rect 30434 37102 30436 37154
rect 30380 37044 30436 37102
rect 30604 37044 30660 37054
rect 30380 37042 30660 37044
rect 30380 36990 30606 37042
rect 30658 36990 30660 37042
rect 30380 36988 30660 36990
rect 30604 36978 30660 36988
rect 30716 36708 30772 37886
rect 30940 37884 31108 37940
rect 30828 37604 30884 37614
rect 30828 37490 30884 37548
rect 30828 37438 30830 37490
rect 30882 37438 30884 37490
rect 30828 36932 30884 37438
rect 30940 37042 30996 37884
rect 31164 37828 31220 38612
rect 30940 36990 30942 37042
rect 30994 36990 30996 37042
rect 30940 36978 30996 36990
rect 31052 37772 31220 37828
rect 31276 38050 31332 38062
rect 31276 37998 31278 38050
rect 31330 37998 31332 38050
rect 31276 37940 31332 37998
rect 30828 36866 30884 36876
rect 30716 36652 30884 36708
rect 30716 36482 30772 36494
rect 30716 36430 30718 36482
rect 30770 36430 30772 36482
rect 30492 36260 30548 36270
rect 30716 36260 30772 36430
rect 30492 36258 30660 36260
rect 30492 36206 30494 36258
rect 30546 36206 30660 36258
rect 30492 36204 30660 36206
rect 30492 36194 30548 36204
rect 30492 35924 30548 35934
rect 30268 35922 30548 35924
rect 30268 35870 30494 35922
rect 30546 35870 30548 35922
rect 30268 35868 30548 35870
rect 30492 35858 30548 35868
rect 29932 35646 29934 35698
rect 29986 35646 29988 35698
rect 29932 35634 29988 35646
rect 30268 35698 30324 35710
rect 30268 35646 30270 35698
rect 30322 35646 30324 35698
rect 30268 35364 30324 35646
rect 30268 35298 30324 35308
rect 30380 35586 30436 35598
rect 30380 35534 30382 35586
rect 30434 35534 30436 35586
rect 29708 35140 29764 35150
rect 29708 35026 29764 35084
rect 30380 35138 30436 35534
rect 30380 35086 30382 35138
rect 30434 35086 30436 35138
rect 30380 35074 30436 35086
rect 30044 35028 30100 35038
rect 29708 34974 29710 35026
rect 29762 34974 29764 35026
rect 29708 34962 29764 34974
rect 29820 35026 30100 35028
rect 29820 34974 30046 35026
rect 30098 34974 30100 35026
rect 29820 34972 30100 34974
rect 29148 34692 29204 34702
rect 28588 34690 29204 34692
rect 28588 34638 28590 34690
rect 28642 34638 29150 34690
rect 29202 34638 29204 34690
rect 28588 34636 29204 34638
rect 27580 34356 27636 34366
rect 27580 34262 27636 34300
rect 28588 34356 28644 34636
rect 29148 34626 29204 34636
rect 29820 34356 29876 34972
rect 30044 34962 30100 34972
rect 28588 34290 28644 34300
rect 29372 34300 29876 34356
rect 30156 34692 30212 34702
rect 29372 34242 29428 34300
rect 29372 34190 29374 34242
rect 29426 34190 29428 34242
rect 29372 34178 29428 34190
rect 27132 33730 27188 33740
rect 28700 34130 28756 34142
rect 28700 34078 28702 34130
rect 28754 34078 28756 34130
rect 28700 33572 28756 34078
rect 28700 33506 28756 33516
rect 30044 33572 30100 33582
rect 26684 33460 26740 33470
rect 26684 33366 26740 33404
rect 27468 33346 27524 33358
rect 27468 33294 27470 33346
rect 27522 33294 27524 33346
rect 27020 33234 27076 33246
rect 27020 33182 27022 33234
rect 27074 33182 27076 33234
rect 26684 32452 26740 32462
rect 26572 32450 26740 32452
rect 26572 32398 26686 32450
rect 26738 32398 26740 32450
rect 26572 32396 26740 32398
rect 26572 31668 26628 32396
rect 26684 32386 26740 32396
rect 27020 32452 27076 33182
rect 27020 31778 27076 32396
rect 27020 31726 27022 31778
rect 27074 31726 27076 31778
rect 27020 31714 27076 31726
rect 27244 33234 27300 33246
rect 27244 33182 27246 33234
rect 27298 33182 27300 33234
rect 27244 32788 27300 33182
rect 27244 31778 27300 32732
rect 27468 32564 27524 33294
rect 27468 32002 27524 32508
rect 27468 31950 27470 32002
rect 27522 31950 27524 32002
rect 27468 31938 27524 31950
rect 27580 33346 27636 33358
rect 27580 33294 27582 33346
rect 27634 33294 27636 33346
rect 27580 32900 27636 33294
rect 27804 33124 27860 33134
rect 27804 33030 27860 33068
rect 28812 33124 28868 33134
rect 27244 31726 27246 31778
rect 27298 31726 27300 31778
rect 26572 31602 26628 31612
rect 26684 31556 26740 31566
rect 26684 31554 27076 31556
rect 26684 31502 26686 31554
rect 26738 31502 27076 31554
rect 26684 31500 27076 31502
rect 26684 31490 26740 31500
rect 25900 29810 25956 29820
rect 26348 31276 26516 31332
rect 27020 31332 27076 31500
rect 27244 31332 27300 31726
rect 27020 31276 27300 31332
rect 25676 29426 25844 29428
rect 25676 29374 25678 29426
rect 25730 29374 25844 29426
rect 25676 29372 25844 29374
rect 25452 28644 25508 28654
rect 25452 28082 25508 28588
rect 25452 28030 25454 28082
rect 25506 28030 25508 28082
rect 25452 28018 25508 28030
rect 25340 27972 25396 27982
rect 25340 27878 25396 27916
rect 25564 27970 25620 27982
rect 25564 27918 25566 27970
rect 25618 27918 25620 27970
rect 24332 26402 24724 26404
rect 24332 26350 24446 26402
rect 24498 26350 24724 26402
rect 24332 26348 24724 26350
rect 24780 26852 25172 26908
rect 25452 27860 25508 27870
rect 25564 27860 25620 27918
rect 25508 27804 25620 27860
rect 25452 26964 25508 27804
rect 25452 26898 25508 26908
rect 25564 27188 25620 27198
rect 25676 27188 25732 29372
rect 26348 28530 26404 31276
rect 26572 30210 26628 30222
rect 26572 30158 26574 30210
rect 26626 30158 26628 30210
rect 26460 30098 26516 30110
rect 26460 30046 26462 30098
rect 26514 30046 26516 30098
rect 26460 29426 26516 30046
rect 26460 29374 26462 29426
rect 26514 29374 26516 29426
rect 26460 29362 26516 29374
rect 26572 28756 26628 30158
rect 27020 30210 27076 31276
rect 27580 30884 27636 32844
rect 28812 32674 28868 33068
rect 30044 32788 30100 33516
rect 28812 32622 28814 32674
rect 28866 32622 28868 32674
rect 28812 32610 28868 32622
rect 29596 32786 30100 32788
rect 29596 32734 30046 32786
rect 30098 32734 30100 32786
rect 29596 32732 30100 32734
rect 29596 32562 29652 32732
rect 30044 32722 30100 32732
rect 29596 32510 29598 32562
rect 29650 32510 29652 32562
rect 29596 32498 29652 32510
rect 29932 32340 29988 32350
rect 27804 31892 27860 31902
rect 27804 31778 27860 31836
rect 28364 31892 28420 31902
rect 28364 31798 28420 31836
rect 27804 31726 27806 31778
rect 27858 31726 27860 31778
rect 27804 31714 27860 31726
rect 29932 31668 29988 32284
rect 29708 31666 29988 31668
rect 29708 31614 29934 31666
rect 29986 31614 29988 31666
rect 29708 31612 29988 31614
rect 27804 31556 27860 31566
rect 27804 31554 28308 31556
rect 27804 31502 27806 31554
rect 27858 31502 28308 31554
rect 27804 31500 28308 31502
rect 27804 31490 27860 31500
rect 27020 30158 27022 30210
rect 27074 30158 27076 30210
rect 27020 30146 27076 30158
rect 27468 30828 27636 30884
rect 26348 28478 26350 28530
rect 26402 28478 26404 28530
rect 26348 28466 26404 28478
rect 26460 28700 26628 28756
rect 26460 28308 26516 28700
rect 25620 27132 25732 27188
rect 26012 28252 26516 28308
rect 26684 28642 26740 28654
rect 26684 28590 26686 28642
rect 26738 28590 26740 28642
rect 26012 27746 26068 28252
rect 26012 27694 26014 27746
rect 26066 27694 26068 27746
rect 23996 26238 23998 26290
rect 24050 26238 24052 26290
rect 23996 26226 24052 26238
rect 24108 26290 24164 26302
rect 24108 26238 24110 26290
rect 24162 26238 24164 26290
rect 23324 26086 23380 26124
rect 24108 26180 24164 26238
rect 23436 25732 23492 25742
rect 22988 25730 23492 25732
rect 22988 25678 23438 25730
rect 23490 25678 23492 25730
rect 22988 25676 23492 25678
rect 22988 25394 23044 25676
rect 23436 25666 23492 25676
rect 23100 25508 23156 25518
rect 23100 25414 23156 25452
rect 23772 25506 23828 25518
rect 23772 25454 23774 25506
rect 23826 25454 23828 25506
rect 22988 25342 22990 25394
rect 23042 25342 23044 25394
rect 22988 25330 23044 25342
rect 23772 25396 23828 25454
rect 23772 25330 23828 25340
rect 23996 25506 24052 25518
rect 23996 25454 23998 25506
rect 24050 25454 24052 25506
rect 23660 25172 23716 25182
rect 23548 25116 23660 25172
rect 22988 25060 23044 25070
rect 22988 23938 23044 25004
rect 23436 25060 23492 25070
rect 23436 24722 23492 25004
rect 23436 24670 23438 24722
rect 23490 24670 23492 24722
rect 23436 24658 23492 24670
rect 23436 24052 23492 24062
rect 22988 23886 22990 23938
rect 23042 23886 23044 23938
rect 22988 23874 23044 23886
rect 23212 23940 23268 23950
rect 23212 23846 23268 23884
rect 22876 23660 23268 23716
rect 23100 23492 23156 23502
rect 22652 22876 22932 22932
rect 22428 22318 22430 22370
rect 22482 22318 22484 22370
rect 22316 21700 22372 21710
rect 22316 21606 22372 21644
rect 22204 21420 22372 21476
rect 22204 20580 22260 20590
rect 22092 20524 22204 20580
rect 22204 20242 22260 20524
rect 22204 20190 22206 20242
rect 22258 20190 22260 20242
rect 22204 20178 22260 20190
rect 22092 20132 22148 20142
rect 21756 20130 22148 20132
rect 21756 20078 22094 20130
rect 22146 20078 22148 20130
rect 21756 20076 22148 20078
rect 21476 19852 21588 19908
rect 21420 19842 21476 19852
rect 21084 16146 21140 16156
rect 21196 17442 21252 17454
rect 21196 17390 21198 17442
rect 21250 17390 21252 17442
rect 20300 16100 20356 16110
rect 19516 15988 19572 15998
rect 19516 13858 19572 15932
rect 20076 15988 20132 15998
rect 20076 15894 20132 15932
rect 20188 15876 20244 15886
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15314 20244 15820
rect 20188 15262 20190 15314
rect 20242 15262 20244 15314
rect 20188 15250 20244 15262
rect 20300 15148 20356 16044
rect 21196 16100 21252 17390
rect 21196 16034 21252 16044
rect 21308 15428 21364 19180
rect 21644 19012 21700 19022
rect 21644 18918 21700 18956
rect 21644 18338 21700 18350
rect 21644 18286 21646 18338
rect 21698 18286 21700 18338
rect 21644 18228 21700 18286
rect 21644 18162 21700 18172
rect 21532 17668 21588 17678
rect 21756 17668 21812 20076
rect 22092 20066 22148 20076
rect 21980 19236 22036 19246
rect 22316 19236 22372 21420
rect 22428 21028 22484 22318
rect 22540 22596 22596 22606
rect 22540 21140 22596 22540
rect 22876 22370 22932 22876
rect 22876 22318 22878 22370
rect 22930 22318 22932 22370
rect 22876 22306 22932 22318
rect 23100 22370 23156 23436
rect 23100 22318 23102 22370
rect 23154 22318 23156 22370
rect 23100 22306 23156 22318
rect 22988 22146 23044 22158
rect 22988 22094 22990 22146
rect 23042 22094 23044 22146
rect 22652 21812 22708 21822
rect 22988 21812 23044 22094
rect 22652 21810 23044 21812
rect 22652 21758 22654 21810
rect 22706 21758 23044 21810
rect 22652 21756 23044 21758
rect 22652 21746 22708 21756
rect 22988 21698 23044 21756
rect 22988 21646 22990 21698
rect 23042 21646 23044 21698
rect 22988 21634 23044 21646
rect 23100 21362 23156 21374
rect 23100 21310 23102 21362
rect 23154 21310 23156 21362
rect 22540 21084 22932 21140
rect 22428 20972 22708 21028
rect 22428 20132 22484 20142
rect 22428 20038 22484 20076
rect 21980 19234 22372 19236
rect 21980 19182 21982 19234
rect 22034 19182 22318 19234
rect 22370 19182 22372 19234
rect 21980 19180 22372 19182
rect 21980 19170 22036 19180
rect 22316 19170 22372 19180
rect 22540 19012 22596 20972
rect 22652 20914 22708 20972
rect 22652 20862 22654 20914
rect 22706 20862 22708 20914
rect 22652 20850 22708 20862
rect 22764 20580 22820 20590
rect 22764 20242 22820 20524
rect 22764 20190 22766 20242
rect 22818 20190 22820 20242
rect 22764 20178 22820 20190
rect 22876 19796 22932 21084
rect 22988 20804 23044 20814
rect 22988 20710 23044 20748
rect 23100 20468 23156 21310
rect 23212 20916 23268 23660
rect 23436 23378 23492 23996
rect 23436 23326 23438 23378
rect 23490 23326 23492 23378
rect 23324 23154 23380 23166
rect 23324 23102 23326 23154
rect 23378 23102 23380 23154
rect 23324 22372 23380 23102
rect 23324 22258 23380 22316
rect 23324 22206 23326 22258
rect 23378 22206 23380 22258
rect 23324 22194 23380 22206
rect 23436 21812 23492 23326
rect 23436 21746 23492 21756
rect 23436 20916 23492 20926
rect 23212 20914 23492 20916
rect 23212 20862 23438 20914
rect 23490 20862 23492 20914
rect 23212 20860 23492 20862
rect 23436 20850 23492 20860
rect 23100 20412 23268 20468
rect 23100 20244 23156 20254
rect 23100 20018 23156 20188
rect 23100 19966 23102 20018
rect 23154 19966 23156 20018
rect 23100 19954 23156 19966
rect 22876 19730 22932 19740
rect 23212 19684 23268 20412
rect 23548 19906 23604 25116
rect 23660 25106 23716 25116
rect 23884 25060 23940 25070
rect 23884 23268 23940 25004
rect 23996 24948 24052 25454
rect 24108 25284 24164 26124
rect 24108 25218 24164 25228
rect 24220 25620 24276 25630
rect 23996 24882 24052 24892
rect 23996 24612 24052 24622
rect 23996 23826 24052 24556
rect 24220 24388 24276 25564
rect 24332 25508 24388 26348
rect 24444 26338 24500 26348
rect 24332 25442 24388 25452
rect 24444 26180 24500 26190
rect 24444 25618 24500 26124
rect 24444 25566 24446 25618
rect 24498 25566 24500 25618
rect 24444 25060 24500 25566
rect 24780 25172 24836 26852
rect 25564 26514 25620 27132
rect 26012 26908 26068 27694
rect 26572 27212 26628 27224
rect 26460 27188 26516 27198
rect 26572 27188 26574 27212
rect 26516 27160 26574 27188
rect 26626 27160 26628 27212
rect 26516 27132 26628 27160
rect 26460 27122 26516 27132
rect 26684 26964 26740 28590
rect 26796 28644 26852 28654
rect 26796 28550 26852 28588
rect 27132 28644 27188 28654
rect 27468 28644 27524 30828
rect 28252 30436 28308 31500
rect 29148 30882 29204 30894
rect 29148 30830 29150 30882
rect 29202 30830 29204 30882
rect 28252 30380 28420 30436
rect 28252 30212 28308 30222
rect 28252 30118 28308 30156
rect 27804 29428 27860 29438
rect 27580 28868 27636 28878
rect 27580 28774 27636 28812
rect 27132 28642 27524 28644
rect 27132 28590 27134 28642
rect 27186 28590 27524 28642
rect 27132 28588 27524 28590
rect 27132 28578 27188 28588
rect 27804 28530 27860 29372
rect 28364 29316 28420 30380
rect 28588 30100 28644 30110
rect 29148 30100 29204 30830
rect 29484 30100 29540 30110
rect 28588 30098 29652 30100
rect 28588 30046 28590 30098
rect 28642 30046 29486 30098
rect 29538 30046 29652 30098
rect 28588 30044 29652 30046
rect 28588 30034 28644 30044
rect 29484 30034 29540 30044
rect 28476 29986 28532 29998
rect 28476 29934 28478 29986
rect 28530 29934 28532 29986
rect 28476 29428 28532 29934
rect 29596 29988 29652 30044
rect 29596 29922 29652 29932
rect 29036 29652 29092 29662
rect 29708 29652 29764 31612
rect 29932 31602 29988 31612
rect 29820 30884 29876 30894
rect 29820 30434 29876 30828
rect 29820 30382 29822 30434
rect 29874 30382 29876 30434
rect 29820 30370 29876 30382
rect 29820 30212 29876 30222
rect 30156 30212 30212 34636
rect 30492 34692 30548 34702
rect 30604 34692 30660 36204
rect 30716 35812 30772 36204
rect 30716 35746 30772 35756
rect 30548 34636 30660 34692
rect 30492 34626 30548 34636
rect 30828 33236 30884 36652
rect 31052 35924 31108 37772
rect 31164 37266 31220 37278
rect 31164 37214 31166 37266
rect 31218 37214 31220 37266
rect 31164 36596 31220 37214
rect 31276 37268 31332 37884
rect 31500 37716 31556 39564
rect 31948 39554 32004 39564
rect 31724 39508 31780 39518
rect 31612 39060 31668 39070
rect 31612 38966 31668 39004
rect 31612 38276 31668 38286
rect 31724 38276 31780 39452
rect 32060 39060 32116 41356
rect 32732 41356 33236 41412
rect 32732 41298 32788 41356
rect 32732 41246 32734 41298
rect 32786 41246 32788 41298
rect 32732 41234 32788 41246
rect 32508 40516 32564 40526
rect 33404 40516 33460 43484
rect 32508 40514 33460 40516
rect 32508 40462 32510 40514
rect 32562 40462 33460 40514
rect 32508 40460 33460 40462
rect 33516 42084 33572 42094
rect 32508 40450 32564 40460
rect 33068 40068 33124 40078
rect 32172 39506 32228 39518
rect 32172 39454 32174 39506
rect 32226 39454 32228 39506
rect 32172 39060 32228 39454
rect 32284 39060 32340 39070
rect 32172 39058 32340 39060
rect 32172 39006 32286 39058
rect 32338 39006 32340 39058
rect 32172 39004 32340 39006
rect 32060 38834 32116 39004
rect 32284 38994 32340 39004
rect 32060 38782 32062 38834
rect 32114 38782 32116 38834
rect 32060 38770 32116 38782
rect 32172 38836 32228 38846
rect 32172 38742 32228 38780
rect 32620 38836 32676 38846
rect 32956 38836 33012 38846
rect 32620 38834 33012 38836
rect 32620 38782 32622 38834
rect 32674 38782 32958 38834
rect 33010 38782 33012 38834
rect 32620 38780 33012 38782
rect 32620 38770 32676 38780
rect 32956 38770 33012 38780
rect 33068 38668 33124 40012
rect 33180 39060 33236 39070
rect 33180 38966 33236 39004
rect 33292 38946 33348 40460
rect 33292 38894 33294 38946
rect 33346 38894 33348 38946
rect 33292 38882 33348 38894
rect 33292 38724 33348 38734
rect 33068 38612 33236 38668
rect 31612 38274 31780 38276
rect 31612 38222 31614 38274
rect 31666 38222 31780 38274
rect 31612 38220 31780 38222
rect 31612 38210 31668 38220
rect 31500 37650 31556 37660
rect 31612 38052 31668 38062
rect 31500 37492 31556 37502
rect 31500 37398 31556 37436
rect 31276 37202 31332 37212
rect 31500 36708 31556 36718
rect 31500 36614 31556 36652
rect 31164 36540 31332 36596
rect 31164 36372 31220 36382
rect 31164 36278 31220 36316
rect 31276 36260 31332 36540
rect 31276 36194 31332 36204
rect 31388 36258 31444 36270
rect 31388 36206 31390 36258
rect 31442 36206 31444 36258
rect 31164 35924 31220 35934
rect 31388 35924 31444 36206
rect 31052 35922 31220 35924
rect 31052 35870 31166 35922
rect 31218 35870 31220 35922
rect 31052 35868 31220 35870
rect 31164 35858 31220 35868
rect 31276 35868 31444 35924
rect 31612 35922 31668 37996
rect 33068 37716 33124 37726
rect 32172 37378 32228 37390
rect 32172 37326 32174 37378
rect 32226 37326 32228 37378
rect 31948 37268 32004 37278
rect 31948 36484 32004 37212
rect 32060 36484 32116 36494
rect 31948 36482 32116 36484
rect 31948 36430 32062 36482
rect 32114 36430 32116 36482
rect 31948 36428 32116 36430
rect 32060 36418 32116 36428
rect 32172 36484 32228 37326
rect 33068 37266 33124 37660
rect 33068 37214 33070 37266
rect 33122 37214 33124 37266
rect 33068 37202 33124 37214
rect 31836 36260 31892 36270
rect 31836 36166 31892 36204
rect 31612 35870 31614 35922
rect 31666 35870 31668 35922
rect 30940 35364 30996 35374
rect 30940 34468 30996 35308
rect 31052 34916 31108 34926
rect 31276 34916 31332 35868
rect 31612 35858 31668 35870
rect 31388 35700 31444 35710
rect 31388 35606 31444 35644
rect 31500 35586 31556 35598
rect 31500 35534 31502 35586
rect 31554 35534 31556 35586
rect 31388 35140 31444 35150
rect 31500 35140 31556 35534
rect 31388 35138 31556 35140
rect 31388 35086 31390 35138
rect 31442 35086 31556 35138
rect 31388 35084 31556 35086
rect 31388 35074 31444 35084
rect 31052 34914 31332 34916
rect 31052 34862 31054 34914
rect 31106 34862 31332 34914
rect 31052 34860 31332 34862
rect 31052 34692 31108 34860
rect 31052 34626 31108 34636
rect 31276 34692 31332 34702
rect 31276 34690 31780 34692
rect 31276 34638 31278 34690
rect 31330 34638 31780 34690
rect 31276 34636 31780 34638
rect 31276 34626 31332 34636
rect 30940 34412 31556 34468
rect 31500 34018 31556 34412
rect 31500 33966 31502 34018
rect 31554 33966 31556 34018
rect 31500 33954 31556 33966
rect 31052 33572 31108 33582
rect 31052 33346 31108 33516
rect 31724 33458 31780 34636
rect 32060 34020 32116 34030
rect 31724 33406 31726 33458
rect 31778 33406 31780 33458
rect 31724 33394 31780 33406
rect 31948 34018 32116 34020
rect 31948 33966 32062 34018
rect 32114 33966 32116 34018
rect 31948 33964 32116 33966
rect 31948 33572 32004 33964
rect 32060 33954 32116 33964
rect 31052 33294 31054 33346
rect 31106 33294 31108 33346
rect 31052 33282 31108 33294
rect 30604 33180 30884 33236
rect 30604 32564 30660 33180
rect 30268 32562 30660 32564
rect 30268 32510 30606 32562
rect 30658 32510 30660 32562
rect 30268 32508 30660 32510
rect 30268 31780 30324 32508
rect 30604 32498 30660 32508
rect 30828 32676 30884 32686
rect 30828 31892 30884 32620
rect 30828 31826 30884 31836
rect 30268 31686 30324 31724
rect 31500 31780 31556 31790
rect 31500 31686 31556 31724
rect 31948 30996 32004 33516
rect 32172 32788 32228 36428
rect 33068 34130 33124 34142
rect 33068 34078 33070 34130
rect 33122 34078 33124 34130
rect 33068 33572 33124 34078
rect 33068 33506 33124 33516
rect 32172 32694 32228 32732
rect 32508 32900 32564 32910
rect 32508 32786 32564 32844
rect 32508 32734 32510 32786
rect 32562 32734 32564 32786
rect 32508 32722 32564 32734
rect 33180 32452 33236 38612
rect 33292 36708 33348 38668
rect 33292 36642 33348 36652
rect 33404 38500 33460 38510
rect 33404 37156 33460 38444
rect 33516 37492 33572 42028
rect 33516 37426 33572 37436
rect 33628 37828 33684 43820
rect 33964 43652 34020 43662
rect 33964 43558 34020 43596
rect 33852 43540 33908 43550
rect 33852 43446 33908 43484
rect 33964 43204 34020 43214
rect 34076 43204 34132 46510
rect 34524 46562 34580 46574
rect 34524 46510 34526 46562
rect 34578 46510 34580 46562
rect 34524 45892 34580 46510
rect 34524 45826 34580 45836
rect 34748 46004 34804 46014
rect 34188 45106 34244 45118
rect 34188 45054 34190 45106
rect 34242 45054 34244 45106
rect 34188 43762 34244 45054
rect 34524 45108 34580 45118
rect 34748 45108 34804 45948
rect 34524 45106 34804 45108
rect 34524 45054 34526 45106
rect 34578 45054 34804 45106
rect 34524 45052 34804 45054
rect 34524 45042 34580 45052
rect 34412 44548 34468 44558
rect 34412 44454 34468 44492
rect 34188 43710 34190 43762
rect 34242 43710 34244 43762
rect 34188 43698 34244 43710
rect 34412 44268 34692 44324
rect 34020 43148 34132 43204
rect 34300 43316 34356 43326
rect 33964 43138 34020 43148
rect 34300 42978 34356 43260
rect 34300 42926 34302 42978
rect 34354 42926 34356 42978
rect 34300 42914 34356 42926
rect 34188 42868 34244 42878
rect 33964 42530 34020 42542
rect 33964 42478 33966 42530
rect 34018 42478 34020 42530
rect 33964 42308 34020 42478
rect 33964 42242 34020 42252
rect 34188 41970 34244 42812
rect 34412 42532 34468 44268
rect 34636 44210 34692 44268
rect 34636 44158 34638 44210
rect 34690 44158 34692 44210
rect 34636 44146 34692 44158
rect 34524 44098 34580 44110
rect 34524 44046 34526 44098
rect 34578 44046 34580 44098
rect 34524 43652 34580 44046
rect 34524 43586 34580 43596
rect 34524 43428 34580 43438
rect 34748 43428 34804 45052
rect 34860 44436 34916 47292
rect 35084 47236 35140 47406
rect 36316 47348 36372 48076
rect 41356 47460 41412 48300
rect 43596 48132 43652 49420
rect 43708 49026 43764 50988
rect 43820 50820 43876 50830
rect 43820 50148 43876 50764
rect 43932 50708 43988 51548
rect 44044 51044 44100 52780
rect 45276 52388 45332 52398
rect 45276 52164 45332 52332
rect 44940 51604 44996 51614
rect 44940 51510 44996 51548
rect 45276 51378 45332 52108
rect 45276 51326 45278 51378
rect 45330 51326 45332 51378
rect 45276 51314 45332 51326
rect 44044 50978 44100 50988
rect 45500 50708 45556 52780
rect 45612 52500 45668 52892
rect 46060 52882 46116 52892
rect 46620 52946 46676 52958
rect 46620 52894 46622 52946
rect 46674 52894 46676 52946
rect 45724 52724 45780 52734
rect 45948 52724 46004 52734
rect 45724 52722 45948 52724
rect 45724 52670 45726 52722
rect 45778 52670 45948 52722
rect 45724 52668 45948 52670
rect 45724 52658 45780 52668
rect 45836 52500 45892 52510
rect 45612 52444 45780 52500
rect 45612 52164 45668 52174
rect 45612 52070 45668 52108
rect 45612 51492 45668 51502
rect 45724 51492 45780 52444
rect 45836 52386 45892 52444
rect 45836 52334 45838 52386
rect 45890 52334 45892 52386
rect 45836 52322 45892 52334
rect 45612 51490 45780 51492
rect 45612 51438 45614 51490
rect 45666 51438 45780 51490
rect 45612 51436 45780 51438
rect 45612 51044 45668 51436
rect 45612 50978 45668 50988
rect 43932 50642 43988 50652
rect 45052 50706 45556 50708
rect 45052 50654 45502 50706
rect 45554 50654 45556 50706
rect 45052 50652 45556 50654
rect 43932 50482 43988 50494
rect 43932 50430 43934 50482
rect 43986 50430 43988 50482
rect 43932 50428 43988 50430
rect 43932 50372 44100 50428
rect 43820 50092 43988 50148
rect 43820 49924 43876 49934
rect 43820 49830 43876 49868
rect 43932 49922 43988 50092
rect 44044 50036 44100 50372
rect 44044 49970 44100 49980
rect 44940 50370 44996 50382
rect 44940 50318 44942 50370
rect 44994 50318 44996 50370
rect 43932 49870 43934 49922
rect 43986 49870 43988 49922
rect 43932 49858 43988 49870
rect 44940 49812 44996 50318
rect 43708 48974 43710 49026
rect 43762 48974 43764 49026
rect 43708 48962 43764 48974
rect 44604 49700 44660 49710
rect 44940 49700 44996 49756
rect 44604 49698 44996 49700
rect 44604 49646 44606 49698
rect 44658 49646 44996 49698
rect 44604 49644 44996 49646
rect 44044 48916 44100 48926
rect 44044 48914 44324 48916
rect 44044 48862 44046 48914
rect 44098 48862 44324 48914
rect 44044 48860 44324 48862
rect 44044 48850 44100 48860
rect 43596 48066 43652 48076
rect 44268 47572 44324 48860
rect 44492 48356 44548 48366
rect 44492 48262 44548 48300
rect 44268 47478 44324 47516
rect 41356 47458 41636 47460
rect 41356 47406 41358 47458
rect 41410 47406 41636 47458
rect 41356 47404 41636 47406
rect 41356 47394 41412 47404
rect 36316 47282 36372 47292
rect 35084 47170 35140 47180
rect 35644 47236 35700 47246
rect 35644 47142 35700 47180
rect 40348 47236 40404 47246
rect 37660 47124 37716 47134
rect 35532 46676 35588 46686
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35532 45892 35588 46620
rect 35868 46674 35924 46686
rect 35868 46622 35870 46674
rect 35922 46622 35924 46674
rect 35644 46564 35700 46574
rect 35868 46564 35924 46622
rect 35644 46562 35924 46564
rect 35644 46510 35646 46562
rect 35698 46510 35924 46562
rect 35644 46508 35924 46510
rect 36652 46562 36708 46574
rect 36652 46510 36654 46562
rect 36706 46510 36708 46562
rect 35644 46004 35700 46508
rect 35644 45938 35700 45948
rect 35532 45798 35588 45836
rect 34972 45220 35028 45230
rect 35196 45220 35252 45230
rect 35028 45218 35252 45220
rect 35028 45166 35198 45218
rect 35250 45166 35252 45218
rect 35028 45164 35252 45166
rect 34972 45154 35028 45164
rect 35196 45154 35252 45164
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34972 44436 35028 44446
rect 34860 44380 34972 44436
rect 34972 44370 35028 44380
rect 36428 43764 36484 43774
rect 35644 43652 35700 43662
rect 35644 43558 35700 43596
rect 34860 43538 34916 43550
rect 34860 43486 34862 43538
rect 34914 43486 34916 43538
rect 34860 43428 34916 43486
rect 34524 43426 34916 43428
rect 34524 43374 34526 43426
rect 34578 43374 34916 43426
rect 34524 43372 34916 43374
rect 34524 43362 34580 43372
rect 34524 42756 34580 42766
rect 34524 42662 34580 42700
rect 34300 42084 34356 42094
rect 34412 42084 34468 42476
rect 34356 42028 34468 42084
rect 34524 42084 34580 42094
rect 34636 42084 34692 43372
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35420 42868 35476 42878
rect 35420 42774 35476 42812
rect 35868 42754 35924 42766
rect 35868 42702 35870 42754
rect 35922 42702 35924 42754
rect 34860 42644 34916 42654
rect 34860 42550 34916 42588
rect 34748 42530 34804 42542
rect 34748 42478 34750 42530
rect 34802 42478 34804 42530
rect 34748 42196 34804 42478
rect 34972 42532 35028 42542
rect 34972 42530 35140 42532
rect 34972 42478 34974 42530
rect 35026 42478 35140 42530
rect 34972 42476 35140 42478
rect 34972 42466 35028 42476
rect 35084 42420 35140 42476
rect 34972 42196 35028 42206
rect 34748 42140 34916 42196
rect 34580 42028 34692 42084
rect 34300 42018 34356 42028
rect 34188 41918 34190 41970
rect 34242 41918 34244 41970
rect 34188 41746 34244 41918
rect 34188 41694 34190 41746
rect 34242 41694 34244 41746
rect 34188 41682 34244 41694
rect 34524 41858 34580 42028
rect 34524 41806 34526 41858
rect 34578 41806 34580 41858
rect 34524 40628 34580 41806
rect 34748 41970 34804 41982
rect 34748 41918 34750 41970
rect 34802 41918 34804 41970
rect 34636 41748 34692 41758
rect 34748 41748 34804 41918
rect 34636 41746 34804 41748
rect 34636 41694 34638 41746
rect 34690 41694 34804 41746
rect 34636 41692 34804 41694
rect 34860 41748 34916 42140
rect 34636 41682 34692 41692
rect 34860 41682 34916 41692
rect 35084 42196 35140 42364
rect 35868 42308 35924 42702
rect 35868 42242 35924 42252
rect 36428 42530 36484 43708
rect 36428 42478 36430 42530
rect 36482 42478 36484 42530
rect 35420 42196 35476 42206
rect 35084 42140 35420 42196
rect 34860 41300 34916 41310
rect 34972 41300 35028 42140
rect 35420 42102 35476 42140
rect 35756 42084 35812 42094
rect 35196 41972 35252 41982
rect 35196 41878 35252 41916
rect 35756 41972 35812 42028
rect 36428 41972 36484 42478
rect 35756 41970 36484 41972
rect 35756 41918 35758 41970
rect 35810 41918 36484 41970
rect 35756 41916 36484 41918
rect 36540 42308 36596 42318
rect 36540 41970 36596 42252
rect 36540 41918 36542 41970
rect 36594 41918 36596 41970
rect 35756 41906 35812 41916
rect 35308 41858 35364 41870
rect 35308 41806 35310 41858
rect 35362 41806 35364 41858
rect 35308 41748 35364 41806
rect 34916 41244 35028 41300
rect 35084 41692 35364 41748
rect 34860 41206 34916 41244
rect 35084 41188 35140 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 41188 35252 41198
rect 35084 41186 35252 41188
rect 35084 41134 35198 41186
rect 35250 41134 35252 41186
rect 35084 41132 35252 41134
rect 35196 41122 35252 41132
rect 35532 41186 35588 41198
rect 35532 41134 35534 41186
rect 35586 41134 35588 41186
rect 34580 40572 34804 40628
rect 34524 40534 34580 40572
rect 34748 40404 34804 40572
rect 34860 40404 34916 40414
rect 34748 40402 34916 40404
rect 34748 40350 34862 40402
rect 34914 40350 34916 40402
rect 34748 40348 34916 40350
rect 33740 40180 33796 40190
rect 33740 37938 33796 40124
rect 34300 39730 34356 39742
rect 34300 39678 34302 39730
rect 34354 39678 34356 39730
rect 34300 39060 34356 39678
rect 34748 39730 34804 40348
rect 34860 40338 34916 40348
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34748 39678 34750 39730
rect 34802 39678 34804 39730
rect 34748 39666 34804 39678
rect 34300 38668 34356 39004
rect 34300 38612 34916 38668
rect 34076 38052 34132 38062
rect 34524 38052 34580 38062
rect 34076 38050 34580 38052
rect 34076 37998 34078 38050
rect 34130 37998 34526 38050
rect 34578 37998 34580 38050
rect 34076 37996 34580 37998
rect 34076 37986 34132 37996
rect 34524 37986 34580 37996
rect 33740 37886 33742 37938
rect 33794 37886 33796 37938
rect 33740 37874 33796 37886
rect 33404 36594 33460 37100
rect 33404 36542 33406 36594
rect 33458 36542 33460 36594
rect 33404 36530 33460 36542
rect 33516 34916 33572 34926
rect 33516 34822 33572 34860
rect 33516 32788 33572 32798
rect 33516 32562 33572 32732
rect 33516 32510 33518 32562
rect 33570 32510 33572 32562
rect 33516 32498 33572 32510
rect 33180 32450 33460 32452
rect 33180 32398 33182 32450
rect 33234 32398 33460 32450
rect 33180 32396 33460 32398
rect 33180 32386 33236 32396
rect 33404 31892 33460 32396
rect 33516 31892 33572 31902
rect 33404 31890 33572 31892
rect 33404 31838 33518 31890
rect 33570 31838 33572 31890
rect 33404 31836 33572 31838
rect 32060 31780 32116 31790
rect 32060 31778 32340 31780
rect 32060 31726 32062 31778
rect 32114 31726 32340 31778
rect 32060 31724 32340 31726
rect 32060 31714 32116 31724
rect 32060 30996 32116 31006
rect 31948 30940 32060 30996
rect 31276 30884 31332 30894
rect 31276 30790 31332 30828
rect 29820 30210 30212 30212
rect 29820 30158 29822 30210
rect 29874 30158 30212 30210
rect 29820 30156 30212 30158
rect 30268 30212 30324 30222
rect 29820 30146 29876 30156
rect 30268 30118 30324 30156
rect 29036 29650 29540 29652
rect 29036 29598 29038 29650
rect 29090 29598 29540 29650
rect 29036 29596 29540 29598
rect 29036 29586 29092 29596
rect 28812 29540 28868 29550
rect 28868 29484 28980 29540
rect 28812 29446 28868 29484
rect 28700 29428 28756 29438
rect 28476 29372 28700 29428
rect 28700 29334 28756 29372
rect 28364 29260 28644 29316
rect 28588 29204 28644 29260
rect 28924 29204 28980 29484
rect 29484 29538 29540 29596
rect 29708 29540 29764 29596
rect 29484 29486 29486 29538
rect 29538 29486 29540 29538
rect 29484 29474 29540 29486
rect 29596 29484 29764 29540
rect 30156 29988 30212 29998
rect 30156 29538 30212 29932
rect 31276 29652 31332 29662
rect 31276 29558 31332 29596
rect 30156 29486 30158 29538
rect 30210 29486 30212 29538
rect 29372 29426 29428 29438
rect 29372 29374 29374 29426
rect 29426 29374 29428 29426
rect 29372 29316 29428 29374
rect 29596 29316 29652 29484
rect 30156 29474 30212 29486
rect 30268 29540 30324 29550
rect 30828 29540 30884 29550
rect 30268 29538 30436 29540
rect 30268 29486 30270 29538
rect 30322 29486 30436 29538
rect 30268 29484 30436 29486
rect 30268 29474 30324 29484
rect 29932 29426 29988 29438
rect 29932 29374 29934 29426
rect 29986 29374 29988 29426
rect 29372 29260 29652 29316
rect 29708 29314 29764 29326
rect 29708 29262 29710 29314
rect 29762 29262 29764 29314
rect 28588 29148 28756 29204
rect 28924 29148 29204 29204
rect 28252 28868 28308 28878
rect 28252 28774 28308 28812
rect 27916 28756 27972 28766
rect 27916 28754 28084 28756
rect 27916 28702 27918 28754
rect 27970 28702 28084 28754
rect 27916 28700 28084 28702
rect 27916 28690 27972 28700
rect 27804 28478 27806 28530
rect 27858 28478 27860 28530
rect 27804 28466 27860 28478
rect 27132 28418 27188 28430
rect 27132 28366 27134 28418
rect 27186 28366 27188 28418
rect 27132 27972 27188 28366
rect 28028 28196 28084 28700
rect 28588 28754 28644 28766
rect 28588 28702 28590 28754
rect 28642 28702 28644 28754
rect 28476 28644 28532 28654
rect 28476 28530 28532 28588
rect 28476 28478 28478 28530
rect 28530 28478 28532 28530
rect 28476 28466 28532 28478
rect 28028 28140 28308 28196
rect 28140 27972 28196 27982
rect 27132 27970 28196 27972
rect 27132 27918 28142 27970
rect 28194 27918 28196 27970
rect 27132 27916 28196 27918
rect 28140 27906 28196 27916
rect 27020 27076 27076 27086
rect 27020 26982 27076 27020
rect 26012 26852 26180 26908
rect 26684 26898 26740 26908
rect 25564 26462 25566 26514
rect 25618 26462 25620 26514
rect 25564 26450 25620 26462
rect 25228 26402 25284 26414
rect 25228 26350 25230 26402
rect 25282 26350 25284 26402
rect 24780 25106 24836 25116
rect 24892 25284 24948 25294
rect 25228 25284 25284 26350
rect 26124 26292 26180 26852
rect 26460 26852 26516 26862
rect 26460 26402 26516 26796
rect 26460 26350 26462 26402
rect 26514 26350 26516 26402
rect 26236 26292 26292 26302
rect 26124 26290 26292 26292
rect 26124 26238 26238 26290
rect 26290 26238 26292 26290
rect 26124 26236 26292 26238
rect 24892 25282 25284 25284
rect 24892 25230 24894 25282
rect 24946 25230 25284 25282
rect 24892 25228 25284 25230
rect 25676 25396 25732 25406
rect 24444 24994 24500 25004
rect 24556 24948 24612 24958
rect 24892 24948 24948 25228
rect 24612 24892 24948 24948
rect 25116 25060 25172 25070
rect 24556 24834 24612 24892
rect 24556 24782 24558 24834
rect 24610 24782 24612 24834
rect 24444 24722 24500 24734
rect 24444 24670 24446 24722
rect 24498 24670 24500 24722
rect 24444 24612 24500 24670
rect 24444 24546 24500 24556
rect 24220 24332 24500 24388
rect 24332 24050 24388 24062
rect 24332 23998 24334 24050
rect 24386 23998 24388 24050
rect 23996 23774 23998 23826
rect 24050 23774 24052 23826
rect 23996 23762 24052 23774
rect 24220 23940 24276 23950
rect 24220 23492 24276 23884
rect 24332 23716 24388 23998
rect 24332 23650 24388 23660
rect 24220 23436 24388 23492
rect 23884 23266 24276 23268
rect 23884 23214 23886 23266
rect 23938 23214 24276 23266
rect 23884 23212 24276 23214
rect 23884 23202 23940 23212
rect 23660 23154 23716 23166
rect 23660 23102 23662 23154
rect 23714 23102 23716 23154
rect 23660 23044 23716 23102
rect 24108 23044 24164 23054
rect 23660 23042 24164 23044
rect 23660 22990 24110 23042
rect 24162 22990 24164 23042
rect 23660 22988 24164 22990
rect 23660 22372 23716 22988
rect 24108 22978 24164 22988
rect 23772 22372 23828 22382
rect 23660 22370 23828 22372
rect 23660 22318 23774 22370
rect 23826 22318 23828 22370
rect 23660 22316 23828 22318
rect 23772 22306 23828 22316
rect 24220 22370 24276 23212
rect 24220 22318 24222 22370
rect 24274 22318 24276 22370
rect 24220 22306 24276 22318
rect 23884 22146 23940 22158
rect 23884 22094 23886 22146
rect 23938 22094 23940 22146
rect 23660 21924 23716 21934
rect 23716 21868 23828 21924
rect 23660 21858 23716 21868
rect 23660 21588 23716 21598
rect 23660 20690 23716 21532
rect 23660 20638 23662 20690
rect 23714 20638 23716 20690
rect 23660 20580 23716 20638
rect 23660 20514 23716 20524
rect 23548 19854 23550 19906
rect 23602 19854 23604 19906
rect 23548 19842 23604 19854
rect 23100 19628 23268 19684
rect 23324 19796 23380 19806
rect 23100 19572 23156 19628
rect 22652 19124 22708 19134
rect 22652 19030 22708 19068
rect 22204 18956 22596 19012
rect 22876 19012 22932 19022
rect 22092 18452 22148 18462
rect 22092 18358 22148 18396
rect 21532 17666 21812 17668
rect 21532 17614 21534 17666
rect 21586 17614 21812 17666
rect 21532 17612 21812 17614
rect 21980 18116 22036 18126
rect 21532 17602 21588 17612
rect 21420 17444 21476 17454
rect 21980 17444 22036 18060
rect 21420 17442 22036 17444
rect 21420 17390 21422 17442
rect 21474 17390 21982 17442
rect 22034 17390 22036 17442
rect 21420 17388 22036 17390
rect 21420 16884 21476 17388
rect 21980 17378 22036 17388
rect 21420 16818 21476 16828
rect 21308 15362 21364 15372
rect 20860 15202 20916 15214
rect 20860 15150 20862 15202
rect 20914 15150 20916 15202
rect 20860 15148 20916 15150
rect 21532 15204 21588 15214
rect 22204 15148 22260 18956
rect 22540 17666 22596 17678
rect 22540 17614 22542 17666
rect 22594 17614 22596 17666
rect 22540 17556 22596 17614
rect 22540 17490 22596 17500
rect 20300 15092 20580 15148
rect 19852 14644 19908 14654
rect 19516 13806 19518 13858
rect 19570 13806 19572 13858
rect 19516 13794 19572 13806
rect 19628 14642 19908 14644
rect 19628 14590 19854 14642
rect 19906 14590 19908 14642
rect 19628 14588 19908 14590
rect 19516 13636 19572 13646
rect 19516 12850 19572 13580
rect 19628 13412 19684 14588
rect 19852 14578 19908 14588
rect 20412 14530 20468 14542
rect 20412 14478 20414 14530
rect 20466 14478 20468 14530
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20412 14084 20468 14478
rect 20412 14018 20468 14028
rect 20300 13858 20356 13870
rect 20300 13806 20302 13858
rect 20354 13806 20356 13858
rect 19628 13346 19684 13356
rect 19740 13746 19796 13758
rect 19740 13694 19742 13746
rect 19794 13694 19796 13746
rect 19740 13076 19796 13694
rect 20300 13636 20356 13806
rect 20524 13746 20580 15092
rect 20636 15092 20916 15148
rect 21084 15092 21588 15148
rect 22092 15092 22260 15148
rect 22316 17442 22372 17454
rect 22316 17390 22318 17442
rect 22370 17390 22372 17442
rect 22316 16884 22372 17390
rect 20636 14418 20692 15092
rect 20636 14366 20638 14418
rect 20690 14366 20692 14418
rect 20636 14354 20692 14366
rect 20524 13694 20526 13746
rect 20578 13694 20580 13746
rect 20524 13682 20580 13694
rect 21084 13746 21140 15092
rect 21196 14084 21252 14094
rect 21252 14028 21476 14084
rect 21196 14018 21252 14028
rect 21420 13970 21476 14028
rect 21420 13918 21422 13970
rect 21474 13918 21476 13970
rect 21420 13906 21476 13918
rect 21084 13694 21086 13746
rect 21138 13694 21140 13746
rect 21084 13682 21140 13694
rect 21868 13748 21924 13758
rect 21868 13654 21924 13692
rect 20300 13570 20356 13580
rect 19740 12962 19796 13020
rect 19740 12910 19742 12962
rect 19794 12910 19796 12962
rect 19740 12898 19796 12910
rect 20300 13188 20356 13198
rect 19516 12798 19518 12850
rect 19570 12798 19572 12850
rect 19516 12786 19572 12798
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19964 12404 20020 12414
rect 19964 11620 20020 12348
rect 20188 12068 20244 12078
rect 20300 12068 20356 13132
rect 21308 13076 21364 13086
rect 21308 12982 21364 13020
rect 21644 12962 21700 12974
rect 21644 12910 21646 12962
rect 21698 12910 21700 12962
rect 20188 12066 20356 12068
rect 20188 12014 20190 12066
rect 20242 12014 20356 12066
rect 20188 12012 20356 12014
rect 20636 12738 20692 12750
rect 20636 12686 20638 12738
rect 20690 12686 20692 12738
rect 20188 12002 20244 12012
rect 19964 11506 20020 11564
rect 19964 11454 19966 11506
rect 20018 11454 20020 11506
rect 19964 11442 20020 11454
rect 20076 11508 20132 11518
rect 20076 11394 20132 11452
rect 20076 11342 20078 11394
rect 20130 11342 20132 11394
rect 20076 11330 20132 11342
rect 20636 11396 20692 12686
rect 21532 12180 21588 12190
rect 20636 11330 20692 11340
rect 20748 11620 20804 11630
rect 20748 11506 20804 11564
rect 20748 11454 20750 11506
rect 20802 11454 20804 11506
rect 19516 11282 19572 11294
rect 19516 11230 19518 11282
rect 19570 11230 19572 11282
rect 19516 10724 19572 11230
rect 20300 11284 20356 11294
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19740 10724 19796 10734
rect 19516 10722 19796 10724
rect 19516 10670 19742 10722
rect 19794 10670 19796 10722
rect 19516 10668 19796 10670
rect 19740 10612 19796 10668
rect 20300 10724 20356 11228
rect 20300 10722 20580 10724
rect 20300 10670 20302 10722
rect 20354 10670 20580 10722
rect 20300 10668 20580 10670
rect 20300 10658 20356 10668
rect 19740 10546 19796 10556
rect 19516 10500 19572 10510
rect 19516 10406 19572 10444
rect 20524 9938 20580 10668
rect 20524 9886 20526 9938
rect 20578 9886 20580 9938
rect 20524 9874 20580 9886
rect 19740 9828 19796 9838
rect 19404 8766 19406 8818
rect 19458 8766 19460 8818
rect 18508 8318 18510 8370
rect 18562 8318 18564 8370
rect 18060 7588 18116 7598
rect 17836 7422 17838 7474
rect 17890 7422 17892 7474
rect 17836 7410 17892 7422
rect 17948 7532 18060 7588
rect 17164 6862 17166 6914
rect 17218 6862 17220 6914
rect 17164 6850 17220 6862
rect 17948 6690 18004 7532
rect 18060 7494 18116 7532
rect 18508 7586 18564 8318
rect 19404 8258 19460 8766
rect 19628 9772 19740 9828
rect 19404 8206 19406 8258
rect 19458 8206 19460 8258
rect 18508 7534 18510 7586
rect 18562 7534 18564 7586
rect 18508 7522 18564 7534
rect 18844 8146 18900 8158
rect 18844 8094 18846 8146
rect 18898 8094 18900 8146
rect 18844 7588 18900 8094
rect 18844 7522 18900 7532
rect 19404 7252 19460 8206
rect 19516 8370 19572 8382
rect 19516 8318 19518 8370
rect 19570 8318 19572 8370
rect 19516 8148 19572 8318
rect 19516 8082 19572 8092
rect 19516 7476 19572 7486
rect 19628 7476 19684 9772
rect 19740 9762 19796 9772
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19740 8930 19796 8942
rect 19740 8878 19742 8930
rect 19794 8878 19796 8930
rect 19740 8818 19796 8878
rect 19740 8766 19742 8818
rect 19794 8766 19796 8818
rect 19740 8754 19796 8766
rect 20524 8820 20580 8830
rect 20524 8818 20692 8820
rect 20524 8766 20526 8818
rect 20578 8766 20692 8818
rect 20524 8764 20692 8766
rect 20524 8754 20580 8764
rect 20076 8148 20132 8158
rect 20076 8054 20132 8092
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19516 7474 19684 7476
rect 19516 7422 19518 7474
rect 19570 7422 19684 7474
rect 19516 7420 19684 7422
rect 19516 7410 19572 7420
rect 20188 7364 20244 7374
rect 20188 7362 20468 7364
rect 20188 7310 20190 7362
rect 20242 7310 20468 7362
rect 20188 7308 20468 7310
rect 20188 7298 20244 7308
rect 19404 7196 19908 7252
rect 19852 6802 19908 7196
rect 19852 6750 19854 6802
rect 19906 6750 19908 6802
rect 19852 6738 19908 6750
rect 17948 6638 17950 6690
rect 18002 6638 18004 6690
rect 17948 6626 18004 6638
rect 15820 6514 15876 6524
rect 17724 6580 17780 6590
rect 17724 6486 17780 6524
rect 18508 6580 18564 6590
rect 16268 6466 16324 6478
rect 16268 6414 16270 6466
rect 16322 6414 16324 6466
rect 16268 6356 16324 6414
rect 15708 6300 16324 6356
rect 16828 6466 16884 6478
rect 16828 6414 16830 6466
rect 16882 6414 16884 6466
rect 16380 6018 16436 6030
rect 16380 5966 16382 6018
rect 16434 5966 16436 6018
rect 15372 5236 15428 5246
rect 15260 5234 15652 5236
rect 15260 5182 15374 5234
rect 15426 5182 15652 5234
rect 15260 5180 15652 5182
rect 15372 5170 15428 5180
rect 15596 5122 15652 5180
rect 16380 5234 16436 5966
rect 16716 6020 16772 6030
rect 16828 6020 16884 6414
rect 16716 6018 16884 6020
rect 16716 5966 16718 6018
rect 16770 5966 16884 6018
rect 16716 5964 16884 5966
rect 16716 5954 16772 5964
rect 16380 5182 16382 5234
rect 16434 5182 16436 5234
rect 16380 5170 16436 5182
rect 18508 5234 18564 6524
rect 20412 6578 20468 7308
rect 20636 6690 20692 8764
rect 20748 8370 20804 11454
rect 21420 11508 21476 11518
rect 21420 11414 21476 11452
rect 20860 10500 20916 10510
rect 21532 10500 21588 12124
rect 21644 11620 21700 12910
rect 21868 12852 21924 12862
rect 21868 12758 21924 12796
rect 21644 11554 21700 11564
rect 20860 10498 21588 10500
rect 20860 10446 20862 10498
rect 20914 10446 21588 10498
rect 20860 10444 21588 10446
rect 20860 10434 20916 10444
rect 21532 9828 21588 10444
rect 22092 10052 22148 15092
rect 22204 14756 22260 14766
rect 22204 14530 22260 14700
rect 22204 14478 22206 14530
rect 22258 14478 22260 14530
rect 22204 14466 22260 14478
rect 22204 13748 22260 13758
rect 22316 13748 22372 16828
rect 22764 17444 22820 17454
rect 22652 15876 22708 15886
rect 22652 15782 22708 15820
rect 22204 13746 22372 13748
rect 22204 13694 22206 13746
rect 22258 13694 22372 13746
rect 22204 13692 22372 13694
rect 22428 15428 22484 15438
rect 22204 13682 22260 13692
rect 22316 13522 22372 13534
rect 22316 13470 22318 13522
rect 22370 13470 22372 13522
rect 22204 13412 22260 13422
rect 22204 13186 22260 13356
rect 22204 13134 22206 13186
rect 22258 13134 22260 13186
rect 22204 13122 22260 13134
rect 22316 13074 22372 13470
rect 22316 13022 22318 13074
rect 22370 13022 22372 13074
rect 22316 13010 22372 13022
rect 22428 12964 22484 15372
rect 22540 14532 22596 14542
rect 22540 14530 22708 14532
rect 22540 14478 22542 14530
rect 22594 14478 22708 14530
rect 22540 14476 22708 14478
rect 22540 14466 22596 14476
rect 22652 13970 22708 14476
rect 22764 14530 22820 17388
rect 22876 17106 22932 18956
rect 22988 17556 23044 17566
rect 22988 17462 23044 17500
rect 22876 17054 22878 17106
rect 22930 17054 22932 17106
rect 22876 16098 22932 17054
rect 23100 16884 23156 19516
rect 23324 19348 23380 19740
rect 23772 19684 23828 21868
rect 23884 21700 23940 22094
rect 23884 20468 23940 21644
rect 24332 21586 24388 23436
rect 24444 22932 24500 24332
rect 24556 23604 24612 24782
rect 24780 24724 24836 24734
rect 24780 24722 24948 24724
rect 24780 24670 24782 24722
rect 24834 24670 24948 24722
rect 24780 24668 24948 24670
rect 24780 24658 24836 24668
rect 24892 23940 24948 24668
rect 24892 23846 24948 23884
rect 24556 23538 24612 23548
rect 25004 23716 25060 23726
rect 24444 22838 24500 22876
rect 25004 22484 25060 23660
rect 24668 22428 25060 22484
rect 24556 21812 24612 21822
rect 24556 21698 24612 21756
rect 24556 21646 24558 21698
rect 24610 21646 24612 21698
rect 24556 21634 24612 21646
rect 24332 21534 24334 21586
rect 24386 21534 24388 21586
rect 24332 21522 24388 21534
rect 23884 20402 23940 20412
rect 23996 21362 24052 21374
rect 23996 21310 23998 21362
rect 24050 21310 24052 21362
rect 23548 19628 23828 19684
rect 23548 19458 23604 19628
rect 23548 19406 23550 19458
rect 23602 19406 23604 19458
rect 23548 19394 23604 19406
rect 23324 19254 23380 19292
rect 23212 19124 23268 19134
rect 23212 18674 23268 19068
rect 23884 19012 23940 19022
rect 23884 18918 23940 18956
rect 23996 18676 24052 21310
rect 24108 20804 24164 20814
rect 24108 20802 24276 20804
rect 24108 20750 24110 20802
rect 24162 20750 24276 20802
rect 24108 20748 24276 20750
rect 24108 20738 24164 20748
rect 24108 20580 24164 20590
rect 24108 20130 24164 20524
rect 24220 20244 24276 20748
rect 24556 20578 24612 20590
rect 24556 20526 24558 20578
rect 24610 20526 24612 20578
rect 24556 20468 24612 20526
rect 24556 20402 24612 20412
rect 24668 20244 24724 22428
rect 24892 22258 24948 22270
rect 24892 22206 24894 22258
rect 24946 22206 24948 22258
rect 24892 21924 24948 22206
rect 24892 21858 24948 21868
rect 25004 22146 25060 22158
rect 25004 22094 25006 22146
rect 25058 22094 25060 22146
rect 25004 21700 25060 22094
rect 25116 22036 25172 25004
rect 25676 24722 25732 25340
rect 26236 25396 26292 26236
rect 26236 25330 26292 25340
rect 26236 24948 26292 24958
rect 26236 24854 26292 24892
rect 25676 24670 25678 24722
rect 25730 24670 25732 24722
rect 25676 24658 25732 24670
rect 25228 24610 25284 24622
rect 25228 24558 25230 24610
rect 25282 24558 25284 24610
rect 25228 24052 25284 24558
rect 26460 24500 26516 26350
rect 27916 25508 27972 25518
rect 28252 25508 28308 28140
rect 28588 26292 28644 28702
rect 28588 26226 28644 26236
rect 27916 25506 28308 25508
rect 27916 25454 27918 25506
rect 27970 25454 28254 25506
rect 28306 25454 28308 25506
rect 27916 25452 28308 25454
rect 27916 25442 27972 25452
rect 28252 25442 28308 25452
rect 28588 26068 28644 26078
rect 27580 25282 27636 25294
rect 27580 25230 27582 25282
rect 27634 25230 27636 25282
rect 26572 24612 26628 24622
rect 26572 24610 26740 24612
rect 26572 24558 26574 24610
rect 26626 24558 26740 24610
rect 26572 24556 26740 24558
rect 26572 24546 26628 24556
rect 25228 23986 25284 23996
rect 25452 24444 26516 24500
rect 25340 23940 25396 23950
rect 25452 23940 25508 24444
rect 25340 23938 25508 23940
rect 25340 23886 25342 23938
rect 25394 23886 25508 23938
rect 25340 23884 25508 23886
rect 25564 24162 25620 24174
rect 25564 24110 25566 24162
rect 25618 24110 25620 24162
rect 25340 23874 25396 23884
rect 25228 23042 25284 23054
rect 25228 22990 25230 23042
rect 25282 22990 25284 23042
rect 25228 22596 25284 22990
rect 25228 22530 25284 22540
rect 25564 22820 25620 24110
rect 26124 23940 26180 23950
rect 26124 23938 26628 23940
rect 26124 23886 26126 23938
rect 26178 23886 26628 23938
rect 26124 23884 26628 23886
rect 26124 23874 26180 23884
rect 26348 23714 26404 23726
rect 26348 23662 26350 23714
rect 26402 23662 26404 23714
rect 26348 23268 26404 23662
rect 26348 23202 26404 23212
rect 25228 22260 25284 22270
rect 25228 22166 25284 22204
rect 25116 21980 25284 22036
rect 25228 21924 25284 21980
rect 25228 21868 25396 21924
rect 25004 21634 25060 21644
rect 25116 21812 25172 21822
rect 25116 21588 25172 21756
rect 25228 21588 25284 21598
rect 25116 21586 25284 21588
rect 25116 21534 25230 21586
rect 25282 21534 25284 21586
rect 25116 21532 25284 21534
rect 25228 21522 25284 21532
rect 25116 20802 25172 20814
rect 25116 20750 25118 20802
rect 25170 20750 25172 20802
rect 24220 20188 24388 20244
rect 24108 20078 24110 20130
rect 24162 20078 24164 20130
rect 24108 20066 24164 20078
rect 24220 20018 24276 20030
rect 24220 19966 24222 20018
rect 24274 19966 24276 20018
rect 24220 19796 24276 19966
rect 24220 19730 24276 19740
rect 24332 19572 24388 20188
rect 24556 20188 24948 20244
rect 24556 20130 24612 20188
rect 24556 20078 24558 20130
rect 24610 20078 24612 20130
rect 24556 20066 24612 20078
rect 24668 20020 24724 20030
rect 24668 19926 24724 19964
rect 24892 19572 24948 20188
rect 25116 19796 25172 20750
rect 25340 20132 25396 21868
rect 25564 21812 25620 22764
rect 25676 22596 25732 22606
rect 25676 22482 25732 22540
rect 26572 22594 26628 23884
rect 26572 22542 26574 22594
rect 26626 22542 26628 22594
rect 26572 22530 26628 22542
rect 25676 22430 25678 22482
rect 25730 22430 25732 22482
rect 25676 22418 25732 22430
rect 26684 22484 26740 24556
rect 27356 23268 27412 23278
rect 27356 23174 27412 23212
rect 27580 23156 27636 25230
rect 28588 25282 28644 26012
rect 28588 25230 28590 25282
rect 28642 25230 28644 25282
rect 27916 24948 27972 24958
rect 27916 23714 27972 24892
rect 27916 23662 27918 23714
rect 27970 23662 27972 23714
rect 27916 23156 27972 23662
rect 28364 23714 28420 23726
rect 28364 23662 28366 23714
rect 28418 23662 28420 23714
rect 28140 23156 28196 23166
rect 28364 23156 28420 23662
rect 28588 23548 28644 25230
rect 28700 24834 28756 29148
rect 29148 28754 29204 29148
rect 29148 28702 29150 28754
rect 29202 28702 29204 28754
rect 29148 28690 29204 28702
rect 29708 28756 29764 29262
rect 29932 29204 29988 29374
rect 30268 29204 30324 29214
rect 29932 29202 30324 29204
rect 29932 29150 30270 29202
rect 30322 29150 30324 29202
rect 29932 29148 30324 29150
rect 30268 29138 30324 29148
rect 30380 29204 30436 29484
rect 30828 29446 30884 29484
rect 31948 29426 32004 29438
rect 31948 29374 31950 29426
rect 32002 29374 32004 29426
rect 30716 29204 30772 29214
rect 30380 29202 30772 29204
rect 30380 29150 30718 29202
rect 30770 29150 30772 29202
rect 30380 29148 30772 29150
rect 29708 28690 29764 28700
rect 30268 28644 30324 28654
rect 30380 28644 30436 29148
rect 30716 29138 30772 29148
rect 31276 28756 31332 28766
rect 31276 28662 31332 28700
rect 30324 28588 30436 28644
rect 30268 28578 30324 28588
rect 30156 28420 30212 28430
rect 30156 27970 30212 28364
rect 31948 28084 32004 29374
rect 32060 28642 32116 30940
rect 32172 29428 32228 29438
rect 32172 29334 32228 29372
rect 32284 29204 32340 31724
rect 32396 31668 32452 31678
rect 32396 29650 32452 31612
rect 32508 30996 32564 31006
rect 32508 30902 32564 30940
rect 33180 30996 33236 31006
rect 32396 29598 32398 29650
rect 32450 29598 32452 29650
rect 32396 29586 32452 29598
rect 33180 29650 33236 30940
rect 33180 29598 33182 29650
rect 33234 29598 33236 29650
rect 33180 29586 33236 29598
rect 32620 29426 32676 29438
rect 32620 29374 32622 29426
rect 32674 29374 32676 29426
rect 32620 29316 32676 29374
rect 32620 29250 32676 29260
rect 32060 28590 32062 28642
rect 32114 28590 32116 28642
rect 32060 28578 32116 28590
rect 32172 29148 32340 29204
rect 31948 28018 32004 28028
rect 30156 27918 30158 27970
rect 30210 27918 30212 27970
rect 30156 27906 30212 27918
rect 28812 27858 28868 27870
rect 28812 27806 28814 27858
rect 28866 27806 28868 27858
rect 28812 27076 28868 27806
rect 29372 27858 29428 27870
rect 29372 27806 29374 27858
rect 29426 27806 29428 27858
rect 28812 27010 28868 27020
rect 29260 27076 29316 27086
rect 29260 26908 29316 27020
rect 29372 26908 29428 27806
rect 29708 26962 29764 26974
rect 29708 26910 29710 26962
rect 29762 26910 29764 26962
rect 29708 26908 29764 26910
rect 29260 26852 29764 26908
rect 28700 24782 28702 24834
rect 28754 24782 28756 24834
rect 28700 24770 28756 24782
rect 29148 26178 29204 26190
rect 29148 26126 29150 26178
rect 29202 26126 29204 26178
rect 29148 24500 29204 26126
rect 29372 24948 29428 24958
rect 29484 24948 29540 26852
rect 29596 26292 29652 26302
rect 29596 25956 29652 26236
rect 30716 26180 30772 26190
rect 29596 25900 30100 25956
rect 29932 25506 29988 25518
rect 29932 25454 29934 25506
rect 29986 25454 29988 25506
rect 29596 25284 29652 25294
rect 29932 25284 29988 25454
rect 29596 25282 29988 25284
rect 29596 25230 29598 25282
rect 29650 25230 29988 25282
rect 29596 25228 29988 25230
rect 29596 24948 29652 25228
rect 29428 24892 29652 24948
rect 29372 24722 29428 24892
rect 29372 24670 29374 24722
rect 29426 24670 29428 24722
rect 29372 24658 29428 24670
rect 29932 24724 29988 24734
rect 30044 24724 30100 25900
rect 30716 25618 30772 26124
rect 30716 25566 30718 25618
rect 30770 25566 30772 25618
rect 30716 25554 30772 25566
rect 29932 24722 30100 24724
rect 29932 24670 29934 24722
rect 29986 24670 30100 24722
rect 29932 24668 30100 24670
rect 30156 24834 30212 24846
rect 30156 24782 30158 24834
rect 30210 24782 30212 24834
rect 29932 24658 29988 24668
rect 28588 23492 28868 23548
rect 27916 23154 28420 23156
rect 27916 23102 28142 23154
rect 28194 23102 28420 23154
rect 27916 23100 28420 23102
rect 26908 22596 26964 22606
rect 26908 22502 26964 22540
rect 26684 22418 26740 22428
rect 27468 22258 27524 22270
rect 27468 22206 27470 22258
rect 27522 22206 27524 22258
rect 25788 22146 25844 22158
rect 25788 22094 25790 22146
rect 25842 22094 25844 22146
rect 25788 21812 25844 22094
rect 25564 21698 25620 21756
rect 25564 21646 25566 21698
rect 25618 21646 25620 21698
rect 25564 21634 25620 21646
rect 25676 21756 25844 21812
rect 26348 22148 26404 22158
rect 25676 20244 25732 21756
rect 26236 21700 26292 21710
rect 25788 21698 26292 21700
rect 25788 21646 26238 21698
rect 26290 21646 26292 21698
rect 25788 21644 26292 21646
rect 25788 20914 25844 21644
rect 26236 21634 26292 21644
rect 25900 21476 25956 21486
rect 25900 21382 25956 21420
rect 25788 20862 25790 20914
rect 25842 20862 25844 20914
rect 25788 20850 25844 20862
rect 25676 20188 26068 20244
rect 25564 20132 25620 20142
rect 25340 20130 25732 20132
rect 25340 20078 25566 20130
rect 25618 20078 25732 20130
rect 25340 20076 25732 20078
rect 25564 20066 25620 20076
rect 25228 20020 25284 20030
rect 25228 19926 25284 19964
rect 25564 19908 25620 19918
rect 25340 19796 25396 19806
rect 25116 19740 25284 19796
rect 25228 19572 25284 19740
rect 25396 19740 25508 19796
rect 25340 19730 25396 19740
rect 24332 19516 24500 19572
rect 24892 19516 25172 19572
rect 25228 19516 25396 19572
rect 24332 19348 24388 19358
rect 24332 19254 24388 19292
rect 24444 18900 24500 19516
rect 24892 19010 24948 19022
rect 24892 18958 24894 19010
rect 24946 18958 24948 19010
rect 24892 18900 24948 18958
rect 24444 18844 24836 18900
rect 23212 18622 23214 18674
rect 23266 18622 23268 18674
rect 23212 18340 23268 18622
rect 23660 18620 24052 18676
rect 24108 18676 24164 18686
rect 23212 18274 23268 18284
rect 23324 18564 23380 18574
rect 23324 17554 23380 18508
rect 23324 17502 23326 17554
rect 23378 17502 23380 17554
rect 23212 17444 23268 17454
rect 23212 17106 23268 17388
rect 23212 17054 23214 17106
rect 23266 17054 23268 17106
rect 23212 17042 23268 17054
rect 23324 16996 23380 17502
rect 23548 18562 23604 18574
rect 23548 18510 23550 18562
rect 23602 18510 23604 18562
rect 23548 17332 23604 18510
rect 23548 17266 23604 17276
rect 23660 17220 23716 18620
rect 23996 18450 24052 18462
rect 23996 18398 23998 18450
rect 24050 18398 24052 18450
rect 23996 18340 24052 18398
rect 23996 18274 24052 18284
rect 24108 18116 24164 18620
rect 24444 18676 24500 18686
rect 24220 18562 24276 18574
rect 24220 18510 24222 18562
rect 24274 18510 24276 18562
rect 24220 18340 24276 18510
rect 24220 18274 24276 18284
rect 24108 18060 24276 18116
rect 24108 17668 24164 17678
rect 24108 17574 24164 17612
rect 24108 17442 24164 17454
rect 24108 17390 24110 17442
rect 24162 17390 24164 17442
rect 24108 17220 24164 17390
rect 23660 17154 23716 17164
rect 23772 17164 24164 17220
rect 23772 17106 23828 17164
rect 23772 17054 23774 17106
rect 23826 17054 23828 17106
rect 23772 17042 23828 17054
rect 23996 16996 24052 17006
rect 24220 16996 24276 18060
rect 24444 17890 24500 18620
rect 24444 17838 24446 17890
rect 24498 17838 24500 17890
rect 24444 17826 24500 17838
rect 24444 17668 24500 17678
rect 24444 17220 24500 17612
rect 24668 17554 24724 17566
rect 24668 17502 24670 17554
rect 24722 17502 24724 17554
rect 24668 17444 24724 17502
rect 24668 17378 24724 17388
rect 24444 17154 24500 17164
rect 24668 17108 24724 17118
rect 23324 16940 23492 16996
rect 23100 16828 23380 16884
rect 22876 16046 22878 16098
rect 22930 16046 22932 16098
rect 22876 16034 22932 16046
rect 23212 15874 23268 15886
rect 23212 15822 23214 15874
rect 23266 15822 23268 15874
rect 22876 15652 22932 15662
rect 22876 14642 22932 15596
rect 22988 15204 23044 15242
rect 22988 15138 23044 15148
rect 23212 14756 23268 15822
rect 23212 14690 23268 14700
rect 22876 14590 22878 14642
rect 22930 14590 22932 14642
rect 22876 14578 22932 14590
rect 22764 14478 22766 14530
rect 22818 14478 22820 14530
rect 22764 14466 22820 14478
rect 22988 14420 23044 14430
rect 22652 13918 22654 13970
rect 22706 13918 22708 13970
rect 22652 13906 22708 13918
rect 22876 14418 23044 14420
rect 22876 14366 22990 14418
rect 23042 14366 23044 14418
rect 22876 14364 23044 14366
rect 22652 13748 22708 13758
rect 22652 13654 22708 13692
rect 22540 12964 22596 12974
rect 22428 12962 22596 12964
rect 22428 12910 22542 12962
rect 22594 12910 22596 12962
rect 22428 12908 22596 12910
rect 22540 12740 22596 12908
rect 22540 12674 22596 12684
rect 22764 12850 22820 12862
rect 22764 12798 22766 12850
rect 22818 12798 22820 12850
rect 22316 12068 22372 12078
rect 22316 12066 22596 12068
rect 22316 12014 22318 12066
rect 22370 12014 22596 12066
rect 22316 12012 22596 12014
rect 22316 12002 22372 12012
rect 22204 11396 22260 11406
rect 22204 11302 22260 11340
rect 22540 11282 22596 12012
rect 22540 11230 22542 11282
rect 22594 11230 22596 11282
rect 22540 11218 22596 11230
rect 22764 11060 22820 12798
rect 22876 11508 22932 14364
rect 22988 14354 23044 14364
rect 22988 12852 23044 12862
rect 23212 12852 23268 12862
rect 22988 12850 23268 12852
rect 22988 12798 22990 12850
rect 23042 12798 23214 12850
rect 23266 12798 23268 12850
rect 22988 12796 23268 12798
rect 22988 12786 23044 12796
rect 23212 12786 23268 12796
rect 23324 12852 23380 16828
rect 23436 12962 23492 16940
rect 23884 16994 24276 16996
rect 23884 16942 23998 16994
rect 24050 16942 24276 16994
rect 23884 16940 24276 16942
rect 24556 16996 24612 17006
rect 23548 16882 23604 16894
rect 23548 16830 23550 16882
rect 23602 16830 23604 16882
rect 23548 15652 23604 16830
rect 23660 16772 23716 16782
rect 23660 16678 23716 16716
rect 23884 16548 23940 16940
rect 23996 16930 24052 16940
rect 24556 16902 24612 16940
rect 24444 16882 24500 16894
rect 24444 16830 24446 16882
rect 24498 16830 24500 16882
rect 24444 16772 24500 16830
rect 24444 16706 24500 16716
rect 23660 16492 23940 16548
rect 24220 16548 24276 16558
rect 23660 15986 23716 16492
rect 23660 15934 23662 15986
rect 23714 15934 23716 15986
rect 23660 15922 23716 15934
rect 23772 16212 23828 16222
rect 23548 15586 23604 15596
rect 23772 15538 23828 16156
rect 23996 16212 24052 16222
rect 23996 16118 24052 16156
rect 23772 15486 23774 15538
rect 23826 15486 23828 15538
rect 23772 15428 23828 15486
rect 23772 15362 23828 15372
rect 23884 15874 23940 15886
rect 23884 15822 23886 15874
rect 23938 15822 23940 15874
rect 23884 14980 23940 15822
rect 24108 15874 24164 15886
rect 24108 15822 24110 15874
rect 24162 15822 24164 15874
rect 24108 15540 24164 15822
rect 23884 14914 23940 14924
rect 23996 15484 24164 15540
rect 23884 14756 23940 14766
rect 23548 14532 23604 14542
rect 23548 14438 23604 14476
rect 23548 13746 23604 13758
rect 23548 13694 23550 13746
rect 23602 13694 23604 13746
rect 23548 13076 23604 13694
rect 23884 13746 23940 14700
rect 23996 13970 24052 15484
rect 24220 15314 24276 16492
rect 24556 16100 24612 16110
rect 24668 16100 24724 17052
rect 24780 17106 24836 18844
rect 24892 18116 24948 18844
rect 24892 18050 24948 18060
rect 24892 17556 24948 17566
rect 24892 17462 24948 17500
rect 24780 17054 24782 17106
rect 24834 17054 24836 17106
rect 24780 17042 24836 17054
rect 24892 16436 24948 16446
rect 24892 16210 24948 16380
rect 24892 16158 24894 16210
rect 24946 16158 24948 16210
rect 24892 16146 24948 16158
rect 24612 16044 24724 16100
rect 24556 15986 24612 16044
rect 24556 15934 24558 15986
rect 24610 15934 24612 15986
rect 24556 15922 24612 15934
rect 24220 15262 24222 15314
rect 24274 15262 24276 15314
rect 24220 15250 24276 15262
rect 24444 15876 24500 15886
rect 23996 13918 23998 13970
rect 24050 13918 24052 13970
rect 23996 13906 24052 13918
rect 24108 14644 24164 14654
rect 23884 13694 23886 13746
rect 23938 13694 23940 13746
rect 23884 13682 23940 13694
rect 24108 13746 24164 14588
rect 24108 13694 24110 13746
rect 24162 13694 24164 13746
rect 24108 13682 24164 13694
rect 24444 14642 24500 15820
rect 24780 15874 24836 15886
rect 24780 15822 24782 15874
rect 24834 15822 24836 15874
rect 24780 15540 24836 15822
rect 24780 15474 24836 15484
rect 25004 15874 25060 15886
rect 25004 15822 25006 15874
rect 25058 15822 25060 15874
rect 24444 14590 24446 14642
rect 24498 14590 24500 14642
rect 23996 13524 24052 13534
rect 23996 13430 24052 13468
rect 24332 13188 24388 13198
rect 24332 13094 24388 13132
rect 23548 13010 23604 13020
rect 23884 13076 23940 13086
rect 23436 12910 23438 12962
rect 23490 12910 23492 12962
rect 23436 12898 23492 12910
rect 23660 12962 23716 12974
rect 23660 12910 23662 12962
rect 23714 12910 23716 12962
rect 23324 12786 23380 12796
rect 23660 12516 23716 12910
rect 23660 12450 23716 12460
rect 23772 12964 23828 12974
rect 23548 12404 23604 12414
rect 23100 12348 23548 12404
rect 23100 12180 23156 12348
rect 23548 12310 23604 12348
rect 23100 12086 23156 12124
rect 23772 12180 23828 12908
rect 23772 12114 23828 12124
rect 23884 11618 23940 13020
rect 23996 12964 24052 12974
rect 24444 12964 24500 14590
rect 24556 15316 24612 15326
rect 24556 15202 24612 15260
rect 24556 15150 24558 15202
rect 24610 15150 24612 15202
rect 24556 13188 24612 15150
rect 25004 13972 25060 15822
rect 25004 13906 25060 13916
rect 25116 13748 25172 19516
rect 25340 19012 25396 19516
rect 25228 18676 25284 18714
rect 25228 18610 25284 18620
rect 25228 18450 25284 18462
rect 25228 18398 25230 18450
rect 25282 18398 25284 18450
rect 25228 18340 25284 18398
rect 25340 18452 25396 18956
rect 25340 18386 25396 18396
rect 25228 17668 25284 18284
rect 25340 17892 25396 17902
rect 25452 17892 25508 19740
rect 25564 18450 25620 19852
rect 25676 18900 25732 20076
rect 25900 20020 25956 20030
rect 25900 19906 25956 19964
rect 25900 19854 25902 19906
rect 25954 19854 25956 19906
rect 25900 19842 25956 19854
rect 25676 18834 25732 18844
rect 26012 18562 26068 20188
rect 26348 19460 26404 22092
rect 27020 21812 27076 21822
rect 27020 21718 27076 21756
rect 27468 21700 27524 22206
rect 27580 21924 27636 23100
rect 27692 22370 27748 22382
rect 27692 22318 27694 22370
rect 27746 22318 27748 22370
rect 27692 22260 27748 22318
rect 27692 22194 27748 22204
rect 27580 21812 27636 21868
rect 27692 21812 27748 21822
rect 27580 21810 27748 21812
rect 27580 21758 27694 21810
rect 27746 21758 27748 21810
rect 27580 21756 27748 21758
rect 27692 21746 27748 21756
rect 27468 21634 27524 21644
rect 28028 21700 28084 21710
rect 26572 21588 26628 21598
rect 26572 21586 26852 21588
rect 26572 21534 26574 21586
rect 26626 21534 26852 21586
rect 26572 21532 26852 21534
rect 26572 21522 26628 21532
rect 26796 20242 26852 21532
rect 27916 20916 27972 20926
rect 26796 20190 26798 20242
rect 26850 20190 26852 20242
rect 26796 20178 26852 20190
rect 27132 20914 27972 20916
rect 27132 20862 27918 20914
rect 27970 20862 27972 20914
rect 27132 20860 27972 20862
rect 27132 20020 27188 20860
rect 27916 20850 27972 20860
rect 28028 20692 28084 21644
rect 27692 20636 28084 20692
rect 27692 20130 27748 20636
rect 28140 20580 28196 23100
rect 28588 23042 28644 23054
rect 28588 22990 28590 23042
rect 28642 22990 28644 23042
rect 28476 22484 28532 22494
rect 28588 22484 28644 22990
rect 28532 22428 28644 22484
rect 28476 22390 28532 22428
rect 28588 22146 28644 22158
rect 28588 22094 28590 22146
rect 28642 22094 28644 22146
rect 28476 21924 28532 21934
rect 28476 21810 28532 21868
rect 28476 21758 28478 21810
rect 28530 21758 28532 21810
rect 28476 21746 28532 21758
rect 28364 20580 28420 20590
rect 28140 20578 28420 20580
rect 28140 20526 28366 20578
rect 28418 20526 28420 20578
rect 28140 20524 28420 20526
rect 27692 20078 27694 20130
rect 27746 20078 27748 20130
rect 27692 20066 27748 20078
rect 27916 20132 27972 20142
rect 26012 18510 26014 18562
rect 26066 18510 26068 18562
rect 26012 18498 26068 18510
rect 26236 19404 26404 19460
rect 27020 20018 27188 20020
rect 27020 19966 27134 20018
rect 27186 19966 27188 20018
rect 27020 19964 27188 19966
rect 27020 19458 27076 19964
rect 27132 19954 27188 19964
rect 27804 20020 27860 20030
rect 27020 19406 27022 19458
rect 27074 19406 27076 19458
rect 25564 18398 25566 18450
rect 25618 18398 25620 18450
rect 25564 18386 25620 18398
rect 25676 18450 25732 18462
rect 25676 18398 25678 18450
rect 25730 18398 25732 18450
rect 25340 17890 25508 17892
rect 25340 17838 25342 17890
rect 25394 17838 25508 17890
rect 25340 17836 25508 17838
rect 25340 17826 25396 17836
rect 25340 17668 25396 17678
rect 25228 17612 25340 17668
rect 25340 17602 25396 17612
rect 25452 17554 25508 17566
rect 25452 17502 25454 17554
rect 25506 17502 25508 17554
rect 25340 17442 25396 17454
rect 25340 17390 25342 17442
rect 25394 17390 25396 17442
rect 25340 16436 25396 17390
rect 25340 16370 25396 16380
rect 25452 16212 25508 17502
rect 25676 16996 25732 18398
rect 25900 18452 25956 18462
rect 25564 16940 25732 16996
rect 25788 16996 25844 17006
rect 25900 16996 25956 18396
rect 26124 17668 26180 17678
rect 26012 16996 26068 17006
rect 25900 16994 26068 16996
rect 25900 16942 26014 16994
rect 26066 16942 26068 16994
rect 25900 16940 26068 16942
rect 25564 16884 25620 16940
rect 25564 16818 25620 16828
rect 25452 16146 25508 16156
rect 25676 16772 25732 16782
rect 25228 16100 25284 16110
rect 25228 16006 25284 16044
rect 25676 16098 25732 16716
rect 25788 16210 25844 16940
rect 26012 16930 26068 16940
rect 25900 16660 25956 16670
rect 25956 16604 26068 16660
rect 25900 16594 25956 16604
rect 25788 16158 25790 16210
rect 25842 16158 25844 16210
rect 25788 16146 25844 16158
rect 25676 16046 25678 16098
rect 25730 16046 25732 16098
rect 25676 16034 25732 16046
rect 25788 15988 25844 15998
rect 25676 15428 25732 15438
rect 25676 15314 25732 15372
rect 25676 15262 25678 15314
rect 25730 15262 25732 15314
rect 25564 15092 25620 15102
rect 25564 14532 25620 15036
rect 25564 13970 25620 14476
rect 25564 13918 25566 13970
rect 25618 13918 25620 13970
rect 25564 13906 25620 13918
rect 25116 13692 25508 13748
rect 25340 13524 25396 13534
rect 24556 13132 24948 13188
rect 24444 12908 24724 12964
rect 23996 12738 24052 12908
rect 23996 12686 23998 12738
rect 24050 12686 24052 12738
rect 23996 12674 24052 12686
rect 24444 12738 24500 12750
rect 24444 12686 24446 12738
rect 24498 12686 24500 12738
rect 24444 12516 24500 12686
rect 24556 12738 24612 12750
rect 24556 12686 24558 12738
rect 24610 12686 24612 12738
rect 24556 12628 24612 12686
rect 24556 12562 24612 12572
rect 24444 12450 24500 12460
rect 24668 12404 24724 12908
rect 24108 11844 24164 11854
rect 23884 11566 23886 11618
rect 23938 11566 23940 11618
rect 23884 11554 23940 11566
rect 23996 11788 24108 11844
rect 22876 11452 23156 11508
rect 22876 11284 22932 11294
rect 22876 11190 22932 11228
rect 22988 11170 23044 11182
rect 22988 11118 22990 11170
rect 23042 11118 23044 11170
rect 22988 11060 23044 11118
rect 22764 11004 23044 11060
rect 22764 10724 22820 10734
rect 22092 9986 22148 9996
rect 22204 10722 22820 10724
rect 22204 10670 22766 10722
rect 22818 10670 22820 10722
rect 22204 10668 22820 10670
rect 22204 9938 22260 10668
rect 22764 10658 22820 10668
rect 22988 10612 23044 10622
rect 22204 9886 22206 9938
rect 22258 9886 22260 9938
rect 22204 9874 22260 9886
rect 22876 10610 23044 10612
rect 22876 10558 22990 10610
rect 23042 10558 23044 10610
rect 22876 10556 23044 10558
rect 21532 9734 21588 9772
rect 22876 9716 22932 10556
rect 22988 10546 23044 10556
rect 22204 9660 22932 9716
rect 22204 9266 22260 9660
rect 23100 9604 23156 11452
rect 23996 9940 24052 11788
rect 24108 11778 24164 11788
rect 24108 11508 24164 11518
rect 24108 10836 24164 11452
rect 24220 11396 24276 11406
rect 24220 11394 24388 11396
rect 24220 11342 24222 11394
rect 24274 11342 24388 11394
rect 24220 11340 24388 11342
rect 24220 11330 24276 11340
rect 24220 10836 24276 10846
rect 24108 10834 24276 10836
rect 24108 10782 24222 10834
rect 24274 10782 24276 10834
rect 24108 10780 24276 10782
rect 24220 10770 24276 10780
rect 22204 9214 22206 9266
rect 22258 9214 22260 9266
rect 22204 9202 22260 9214
rect 22764 9548 23156 9604
rect 23884 9884 24052 9940
rect 24108 10052 24164 10062
rect 21532 9154 21588 9166
rect 21532 9102 21534 9154
rect 21586 9102 21588 9154
rect 20748 8318 20750 8370
rect 20802 8318 20804 8370
rect 20748 8260 20804 8318
rect 20748 8194 20804 8204
rect 20860 8818 20916 8830
rect 20860 8766 20862 8818
rect 20914 8766 20916 8818
rect 20860 8596 20916 8766
rect 20636 6638 20638 6690
rect 20690 6638 20692 6690
rect 20636 6626 20692 6638
rect 20412 6526 20414 6578
rect 20466 6526 20468 6578
rect 20412 6514 20468 6526
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20860 5908 20916 8540
rect 21532 8372 21588 9102
rect 21644 9044 21700 9054
rect 21644 8950 21700 8988
rect 22540 8818 22596 8830
rect 22540 8766 22542 8818
rect 22594 8766 22596 8818
rect 22540 8708 22596 8766
rect 22540 8642 22596 8652
rect 22204 8482 22260 8494
rect 22204 8430 22206 8482
rect 22258 8430 22260 8482
rect 21532 8306 21588 8316
rect 21644 8370 21700 8382
rect 21644 8318 21646 8370
rect 21698 8318 21700 8370
rect 21644 8260 21700 8318
rect 21644 8194 21700 8204
rect 21980 8258 22036 8270
rect 21980 8206 21982 8258
rect 22034 8206 22036 8258
rect 21980 8148 22036 8206
rect 21980 7700 22036 8092
rect 21980 7634 22036 7644
rect 22092 6916 22148 6926
rect 21980 6860 22092 6916
rect 21980 6018 22036 6860
rect 22092 6850 22148 6860
rect 21980 5966 21982 6018
rect 22034 5966 22036 6018
rect 21980 5954 22036 5966
rect 22092 6692 22148 6702
rect 21420 5908 21476 5918
rect 20860 5906 21476 5908
rect 20860 5854 21422 5906
rect 21474 5854 21476 5906
rect 20860 5852 21476 5854
rect 21420 5842 21476 5852
rect 21084 5684 21140 5694
rect 18508 5182 18510 5234
rect 18562 5182 18564 5234
rect 18508 5170 18564 5182
rect 20412 5682 21140 5684
rect 20412 5630 21086 5682
rect 21138 5630 21140 5682
rect 20412 5628 21140 5630
rect 15596 5070 15598 5122
rect 15650 5070 15652 5122
rect 15596 5058 15652 5070
rect 20412 5122 20468 5628
rect 21084 5618 21140 5628
rect 21308 5684 21364 5694
rect 20412 5070 20414 5122
rect 20466 5070 20468 5122
rect 20412 5058 20468 5070
rect 21308 5122 21364 5628
rect 21308 5070 21310 5122
rect 21362 5070 21364 5122
rect 21308 5058 21364 5070
rect 21644 5124 21700 5134
rect 20524 5012 20580 5022
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20524 4338 20580 4956
rect 21644 5010 21700 5068
rect 21644 4958 21646 5010
rect 21698 4958 21700 5010
rect 21644 4946 21700 4958
rect 22092 5122 22148 6636
rect 22204 6020 22260 8430
rect 22316 8372 22372 8382
rect 22316 7362 22372 8316
rect 22764 8370 22820 9548
rect 23212 9156 23268 9166
rect 23212 9062 23268 9100
rect 23324 9044 23380 9054
rect 23772 9044 23828 9054
rect 23380 9042 23828 9044
rect 23380 8990 23774 9042
rect 23826 8990 23828 9042
rect 23380 8988 23828 8990
rect 23324 8950 23380 8988
rect 23772 8978 23828 8988
rect 23100 8708 23156 8718
rect 22764 8318 22766 8370
rect 22818 8318 22820 8370
rect 22764 8306 22820 8318
rect 22988 8652 23100 8708
rect 22876 7700 22932 7710
rect 22876 7606 22932 7644
rect 22316 7310 22318 7362
rect 22370 7310 22372 7362
rect 22316 7298 22372 7310
rect 22540 6692 22596 6702
rect 22540 6598 22596 6636
rect 22204 5906 22260 5964
rect 22204 5854 22206 5906
rect 22258 5854 22260 5906
rect 22204 5842 22260 5854
rect 22988 5908 23044 8652
rect 23100 8642 23156 8652
rect 23100 8372 23156 8382
rect 23100 8278 23156 8316
rect 23324 8260 23380 8270
rect 23324 7698 23380 8204
rect 23884 8258 23940 9884
rect 24108 9044 24164 9996
rect 24332 9938 24388 11340
rect 24668 10724 24724 12348
rect 24892 11394 24948 13132
rect 25228 12962 25284 12974
rect 25228 12910 25230 12962
rect 25282 12910 25284 12962
rect 25228 12852 25284 12910
rect 25228 12786 25284 12796
rect 25340 11620 25396 13468
rect 25452 13076 25508 13692
rect 25452 12982 25508 13020
rect 25676 12404 25732 15262
rect 25788 15202 25844 15932
rect 25788 15150 25790 15202
rect 25842 15150 25844 15202
rect 25788 13076 25844 15150
rect 25900 15874 25956 15886
rect 25900 15822 25902 15874
rect 25954 15822 25956 15874
rect 25900 14308 25956 15822
rect 25900 14242 25956 14252
rect 26012 13860 26068 16604
rect 26124 14420 26180 17612
rect 26236 15988 26292 19404
rect 27020 19394 27076 19406
rect 26684 19348 26740 19358
rect 26348 19346 26740 19348
rect 26348 19294 26686 19346
rect 26738 19294 26740 19346
rect 26348 19292 26740 19294
rect 26348 17890 26404 19292
rect 26684 19282 26740 19292
rect 26796 19236 26852 19246
rect 26796 19122 26852 19180
rect 26796 19070 26798 19122
rect 26850 19070 26852 19122
rect 26796 19058 26852 19070
rect 26348 17838 26350 17890
rect 26402 17838 26404 17890
rect 26348 17826 26404 17838
rect 27692 18452 27748 18462
rect 27692 17780 27748 18396
rect 27356 17778 27748 17780
rect 27356 17726 27694 17778
rect 27746 17726 27748 17778
rect 27356 17724 27748 17726
rect 26460 17666 26516 17678
rect 26460 17614 26462 17666
rect 26514 17614 26516 17666
rect 26348 16996 26404 17006
rect 26348 16322 26404 16940
rect 26460 16884 26516 17614
rect 26796 17554 26852 17566
rect 26796 17502 26798 17554
rect 26850 17502 26852 17554
rect 26684 17442 26740 17454
rect 26684 17390 26686 17442
rect 26738 17390 26740 17442
rect 26460 16818 26516 16828
rect 26572 17220 26628 17230
rect 26348 16270 26350 16322
rect 26402 16270 26404 16322
rect 26348 16258 26404 16270
rect 26572 16212 26628 17164
rect 26684 16884 26740 17390
rect 26684 16818 26740 16828
rect 26684 16324 26740 16334
rect 26684 16230 26740 16268
rect 26572 16146 26628 16156
rect 26796 15988 26852 17502
rect 26236 15922 26292 15932
rect 26348 15932 26852 15988
rect 26908 17444 26964 17454
rect 26236 15652 26292 15662
rect 26236 15426 26292 15596
rect 26236 15374 26238 15426
rect 26290 15374 26292 15426
rect 26236 15362 26292 15374
rect 26236 14868 26292 14878
rect 26236 14644 26292 14812
rect 26236 14530 26292 14588
rect 26236 14478 26238 14530
rect 26290 14478 26292 14530
rect 26236 14466 26292 14478
rect 26124 14354 26180 14364
rect 26236 14308 26292 14318
rect 26236 14214 26292 14252
rect 26124 13860 26180 13870
rect 26012 13858 26180 13860
rect 26012 13806 26126 13858
rect 26178 13806 26180 13858
rect 26012 13804 26180 13806
rect 26124 13794 26180 13804
rect 25900 13748 25956 13758
rect 25900 13746 26068 13748
rect 25900 13694 25902 13746
rect 25954 13694 26068 13746
rect 25900 13692 26068 13694
rect 25900 13682 25956 13692
rect 25788 13020 25956 13076
rect 25788 12850 25844 12862
rect 25788 12798 25790 12850
rect 25842 12798 25844 12850
rect 25788 12740 25844 12798
rect 25788 12674 25844 12684
rect 25788 12404 25844 12414
rect 25676 12348 25788 12404
rect 25340 11564 25732 11620
rect 25676 11508 25732 11564
rect 25676 11414 25732 11452
rect 24892 11342 24894 11394
rect 24946 11342 24948 11394
rect 24892 11330 24948 11342
rect 25004 11282 25060 11294
rect 25004 11230 25006 11282
rect 25058 11230 25060 11282
rect 24668 10668 24836 10724
rect 24668 10498 24724 10510
rect 24668 10446 24670 10498
rect 24722 10446 24724 10498
rect 24668 10276 24724 10446
rect 24668 10210 24724 10220
rect 24332 9886 24334 9938
rect 24386 9886 24388 9938
rect 24332 9156 24388 9886
rect 24780 9826 24836 10668
rect 24780 9774 24782 9826
rect 24834 9774 24836 9826
rect 24780 9268 24836 9774
rect 24332 9090 24388 9100
rect 24668 9212 24780 9268
rect 24108 9042 24276 9044
rect 24108 8990 24110 9042
rect 24162 8990 24276 9042
rect 24108 8988 24276 8990
rect 24108 8978 24164 8988
rect 23884 8206 23886 8258
rect 23938 8206 23940 8258
rect 23884 8194 23940 8206
rect 23996 8930 24052 8942
rect 23996 8878 23998 8930
rect 24050 8878 24052 8930
rect 23996 8260 24052 8878
rect 24220 8932 24276 8988
rect 24220 8876 24500 8932
rect 24444 8370 24500 8876
rect 24444 8318 24446 8370
rect 24498 8318 24500 8370
rect 24444 8306 24500 8318
rect 23996 8194 24052 8204
rect 23324 7646 23326 7698
rect 23378 7646 23380 7698
rect 23324 7634 23380 7646
rect 23660 8146 23716 8158
rect 23660 8094 23662 8146
rect 23714 8094 23716 8146
rect 23660 6916 23716 8094
rect 23436 6860 23660 6916
rect 23324 6020 23380 6030
rect 23324 5926 23380 5964
rect 23100 5908 23156 5918
rect 22988 5906 23156 5908
rect 22988 5854 23102 5906
rect 23154 5854 23156 5906
rect 22988 5852 23156 5854
rect 23100 5842 23156 5852
rect 22764 5684 22820 5694
rect 22764 5590 22820 5628
rect 22092 5070 22094 5122
rect 22146 5070 22148 5122
rect 22092 5012 22148 5070
rect 22764 5124 22820 5134
rect 22764 5030 22820 5068
rect 22092 4946 22148 4956
rect 20748 4900 20804 4910
rect 20748 4898 21252 4900
rect 20748 4846 20750 4898
rect 20802 4846 21252 4898
rect 20748 4844 21252 4846
rect 20748 4834 20804 4844
rect 21196 4450 21252 4844
rect 21196 4398 21198 4450
rect 21250 4398 21252 4450
rect 21196 4386 21252 4398
rect 20524 4286 20526 4338
rect 20578 4286 20580 4338
rect 20524 4274 20580 4286
rect 23324 4228 23380 4238
rect 23436 4228 23492 6860
rect 23660 6850 23716 6860
rect 24668 6692 24724 9212
rect 24780 9202 24836 9212
rect 24668 6598 24724 6636
rect 23884 6020 23940 6030
rect 25004 6020 25060 11230
rect 25564 11284 25620 11294
rect 25340 10722 25396 10734
rect 25340 10670 25342 10722
rect 25394 10670 25396 10722
rect 25340 9940 25396 10670
rect 25564 10610 25620 11228
rect 25564 10558 25566 10610
rect 25618 10558 25620 10610
rect 25564 10276 25620 10558
rect 25564 10210 25620 10220
rect 25340 9884 25620 9940
rect 25452 9714 25508 9726
rect 25452 9662 25454 9714
rect 25506 9662 25508 9714
rect 25340 9268 25396 9278
rect 25340 8484 25396 9212
rect 25340 8418 25396 8428
rect 25452 8146 25508 9662
rect 25564 8596 25620 9884
rect 25788 9044 25844 12348
rect 25900 10612 25956 13020
rect 26012 10836 26068 13692
rect 26124 13076 26180 13086
rect 26124 12178 26180 13020
rect 26236 13074 26292 13086
rect 26236 13022 26238 13074
rect 26290 13022 26292 13074
rect 26236 12628 26292 13022
rect 26348 12964 26404 15932
rect 26572 15764 26628 15774
rect 26908 15764 26964 17388
rect 27132 17442 27188 17454
rect 27132 17390 27134 17442
rect 27186 17390 27188 17442
rect 27132 16548 27188 17390
rect 26572 15314 26628 15708
rect 26572 15262 26574 15314
rect 26626 15262 26628 15314
rect 26572 15250 26628 15262
rect 26684 15708 26964 15764
rect 27020 15764 27076 15774
rect 26684 14756 26740 15708
rect 27020 15652 27076 15708
rect 26796 15596 27076 15652
rect 26796 15090 26852 15596
rect 27132 15540 27188 16492
rect 27356 16098 27412 17724
rect 27692 17714 27748 17724
rect 27356 16046 27358 16098
rect 27410 16046 27412 16098
rect 27356 16034 27412 16046
rect 27804 16882 27860 19964
rect 27916 20018 27972 20076
rect 27916 19966 27918 20018
rect 27970 19966 27972 20018
rect 27916 19124 27972 19966
rect 27916 19058 27972 19068
rect 28364 20132 28420 20524
rect 28364 20018 28420 20076
rect 28364 19966 28366 20018
rect 28418 19966 28420 20018
rect 28028 19012 28084 19022
rect 28364 19012 28420 19966
rect 28084 18956 28420 19012
rect 28028 18918 28084 18956
rect 28364 18452 28420 18490
rect 28364 18386 28420 18396
rect 28028 18228 28084 18238
rect 28028 18134 28084 18172
rect 28364 18226 28420 18238
rect 28364 18174 28366 18226
rect 28418 18174 28420 18226
rect 28364 17892 28420 18174
rect 28364 17826 28420 17836
rect 28588 17668 28644 22094
rect 28588 17602 28644 17612
rect 28364 17444 28420 17454
rect 28140 16996 28196 17006
rect 28140 16902 28196 16940
rect 28364 16994 28420 17388
rect 28364 16942 28366 16994
rect 28418 16942 28420 16994
rect 28364 16930 28420 16942
rect 28700 17220 28756 17230
rect 27804 16830 27806 16882
rect 27858 16830 27860 16882
rect 27468 15988 27524 15998
rect 27468 15894 27524 15932
rect 27804 15876 27860 16830
rect 28588 16884 28644 16894
rect 28588 16790 28644 16828
rect 28700 16882 28756 17164
rect 28700 16830 28702 16882
rect 28754 16830 28756 16882
rect 28700 16818 28756 16830
rect 28252 16772 28308 16782
rect 28252 16678 28308 16716
rect 28140 16324 28196 16334
rect 28028 15876 28084 15886
rect 27804 15874 28084 15876
rect 27804 15822 28030 15874
rect 28082 15822 28084 15874
rect 27804 15820 28084 15822
rect 26796 15038 26798 15090
rect 26850 15038 26852 15090
rect 26796 15026 26852 15038
rect 26908 15484 27188 15540
rect 27244 15540 27300 15550
rect 26684 14700 26852 14756
rect 26572 14532 26628 14542
rect 26572 14530 26740 14532
rect 26572 14478 26574 14530
rect 26626 14478 26740 14530
rect 26572 14476 26740 14478
rect 26572 14466 26628 14476
rect 26460 14420 26516 14430
rect 26460 13748 26516 14364
rect 26684 13970 26740 14476
rect 26796 14530 26852 14700
rect 26796 14478 26798 14530
rect 26850 14478 26852 14530
rect 26796 14466 26852 14478
rect 26908 14308 26964 15484
rect 27244 15446 27300 15484
rect 27020 15314 27076 15326
rect 27020 15262 27022 15314
rect 27074 15262 27076 15314
rect 27020 14756 27076 15262
rect 27356 15316 27412 15326
rect 27916 15316 27972 15326
rect 27356 15314 27972 15316
rect 27356 15262 27358 15314
rect 27410 15262 27918 15314
rect 27970 15262 27972 15314
rect 27356 15260 27972 15262
rect 27356 15250 27412 15260
rect 27916 15250 27972 15260
rect 27132 15204 27188 15214
rect 27468 15148 27636 15204
rect 27132 15092 27300 15148
rect 27468 15092 27524 15148
rect 27580 15092 27748 15148
rect 27244 15036 27524 15092
rect 27580 14980 27636 14990
rect 27020 14690 27076 14700
rect 27244 14868 27300 14878
rect 27020 14420 27076 14430
rect 27020 14326 27076 14364
rect 26684 13918 26686 13970
rect 26738 13918 26740 13970
rect 26684 13906 26740 13918
rect 26796 14252 26964 14308
rect 26460 13682 26516 13692
rect 26460 13524 26516 13534
rect 26460 13430 26516 13468
rect 26684 12964 26740 12974
rect 26796 12964 26852 14252
rect 27020 13972 27076 13982
rect 27020 13878 27076 13916
rect 27244 13746 27300 14812
rect 27244 13694 27246 13746
rect 27298 13694 27300 13746
rect 27244 13682 27300 13694
rect 27468 14756 27524 14766
rect 27468 13746 27524 14700
rect 27580 14308 27636 14924
rect 27692 14530 27748 15092
rect 28028 15092 28084 15820
rect 28028 15026 28084 15036
rect 28028 14756 28084 14766
rect 28140 14756 28196 16268
rect 28588 15428 28644 15438
rect 28588 15334 28644 15372
rect 28252 15316 28308 15326
rect 28252 15222 28308 15260
rect 28476 15092 28532 15102
rect 28028 14754 28196 14756
rect 28028 14702 28030 14754
rect 28082 14702 28196 14754
rect 28028 14700 28196 14702
rect 28252 14756 28308 14766
rect 28028 14690 28084 14700
rect 27692 14478 27694 14530
rect 27746 14478 27748 14530
rect 27692 14466 27748 14478
rect 28252 14530 28308 14700
rect 28252 14478 28254 14530
rect 28306 14478 28308 14530
rect 28252 14466 28308 14478
rect 28476 14530 28532 15036
rect 28476 14478 28478 14530
rect 28530 14478 28532 14530
rect 28476 14466 28532 14478
rect 27692 14308 27748 14318
rect 27580 14306 27748 14308
rect 27580 14254 27694 14306
rect 27746 14254 27748 14306
rect 27580 14252 27748 14254
rect 27692 14242 27748 14252
rect 28812 13972 28868 23492
rect 29148 21924 29204 24444
rect 29260 23938 29316 23950
rect 29260 23886 29262 23938
rect 29314 23886 29316 23938
rect 29260 22594 29316 23886
rect 29484 23714 29540 23726
rect 29484 23662 29486 23714
rect 29538 23662 29540 23714
rect 29484 23268 29540 23662
rect 29484 23202 29540 23212
rect 29260 22542 29262 22594
rect 29314 22542 29316 22594
rect 29260 22530 29316 22542
rect 29596 22484 29652 22494
rect 30156 22484 30212 24782
rect 30716 23268 30772 23278
rect 30716 23174 30772 23212
rect 29596 22390 29652 22428
rect 30044 22428 30212 22484
rect 31388 23154 31444 23166
rect 31388 23102 31390 23154
rect 31442 23102 31444 23154
rect 30044 22372 30100 22428
rect 29820 22260 29876 22270
rect 29820 22166 29876 22204
rect 30044 21924 30100 22316
rect 31164 22372 31220 22382
rect 31388 22372 31444 23102
rect 32172 22932 32228 29148
rect 33404 28866 33460 31836
rect 33516 31780 33572 31836
rect 33516 31714 33572 31724
rect 33628 30212 33684 37772
rect 33964 37826 34020 37838
rect 33964 37774 33966 37826
rect 34018 37774 34020 37826
rect 33964 37716 34020 37774
rect 34188 37828 34244 37838
rect 34636 37828 34692 37838
rect 34188 37734 34244 37772
rect 34300 37826 34692 37828
rect 34300 37774 34638 37826
rect 34690 37774 34692 37826
rect 34300 37772 34692 37774
rect 33964 37650 34020 37660
rect 34300 37492 34356 37772
rect 34636 37762 34692 37772
rect 34748 37826 34804 37838
rect 34748 37774 34750 37826
rect 34802 37774 34804 37826
rect 33852 37436 34356 37492
rect 34412 37604 34468 37614
rect 33852 37378 33908 37436
rect 33852 37326 33854 37378
rect 33906 37326 33908 37378
rect 33852 37314 33908 37326
rect 33740 36484 33796 36494
rect 33740 36390 33796 36428
rect 34412 35810 34468 37548
rect 34748 37492 34804 37774
rect 34748 37426 34804 37436
rect 34860 36484 34916 38612
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35532 37828 35588 41134
rect 35756 41076 35812 41086
rect 35756 40982 35812 41020
rect 35644 40962 35700 40974
rect 35644 40910 35646 40962
rect 35698 40910 35700 40962
rect 35644 40514 35700 40910
rect 35644 40462 35646 40514
rect 35698 40462 35700 40514
rect 35644 40450 35700 40462
rect 36092 39732 36148 41916
rect 36540 41906 36596 41918
rect 36428 41076 36484 41086
rect 36428 40982 36484 41020
rect 36204 40964 36260 40974
rect 36204 40870 36260 40908
rect 36316 40962 36372 40974
rect 36316 40910 36318 40962
rect 36370 40910 36372 40962
rect 36316 40068 36372 40910
rect 36316 40002 36372 40012
rect 36428 39732 36484 39742
rect 36092 39730 36484 39732
rect 36092 39678 36430 39730
rect 36482 39678 36484 39730
rect 36092 39676 36484 39678
rect 36092 38164 36148 39676
rect 36428 39620 36484 39676
rect 36428 39554 36484 39564
rect 36652 38724 36708 46510
rect 37324 45444 37380 45454
rect 37324 44994 37380 45388
rect 37324 44942 37326 44994
rect 37378 44942 37380 44994
rect 37324 44930 37380 44942
rect 37548 44098 37604 44110
rect 37548 44046 37550 44098
rect 37602 44046 37604 44098
rect 37548 43764 37604 44046
rect 37548 43698 37604 43708
rect 36988 42644 37044 42654
rect 36988 42550 37044 42588
rect 37100 42530 37156 42542
rect 37100 42478 37102 42530
rect 37154 42478 37156 42530
rect 37100 42308 37156 42478
rect 37212 42532 37268 42542
rect 37212 42438 37268 42476
rect 37100 42242 37156 42252
rect 37212 42196 37268 42206
rect 37212 41972 37268 42140
rect 36988 41916 37268 41972
rect 36988 41186 37044 41916
rect 36988 41134 36990 41186
rect 37042 41134 37044 41186
rect 36988 41122 37044 41134
rect 37100 41076 37156 41086
rect 37100 40982 37156 41020
rect 37212 40964 37268 40974
rect 37212 40870 37268 40908
rect 37436 40962 37492 40974
rect 37436 40910 37438 40962
rect 37490 40910 37492 40962
rect 37436 40852 37492 40910
rect 37436 40786 37492 40796
rect 37100 39620 37156 39630
rect 37100 39526 37156 39564
rect 37660 39508 37716 47068
rect 40348 46676 40404 47180
rect 41132 46788 41188 46798
rect 41020 46786 41188 46788
rect 41020 46734 41134 46786
rect 41186 46734 41188 46786
rect 41020 46732 41188 46734
rect 41020 46676 41076 46732
rect 41132 46722 41188 46732
rect 40348 46674 41076 46676
rect 40348 46622 40350 46674
rect 40402 46622 41076 46674
rect 40348 46620 41076 46622
rect 40348 46610 40404 46620
rect 38780 46564 38836 46574
rect 38780 46470 38836 46508
rect 40908 46452 40964 46462
rect 40460 46450 40964 46452
rect 40460 46398 40910 46450
rect 40962 46398 40964 46450
rect 40460 46396 40964 46398
rect 38892 46004 38948 46014
rect 39676 46004 39732 46014
rect 38892 46002 39732 46004
rect 38892 45950 38894 46002
rect 38946 45950 39678 46002
rect 39730 45950 39732 46002
rect 38892 45948 39732 45950
rect 38668 45892 38724 45902
rect 38332 45890 38724 45892
rect 38332 45838 38670 45890
rect 38722 45838 38724 45890
rect 38332 45836 38724 45838
rect 38332 45444 38388 45836
rect 38668 45826 38724 45836
rect 38332 45330 38388 45388
rect 38332 45278 38334 45330
rect 38386 45278 38388 45330
rect 38332 45266 38388 45278
rect 37996 45218 38052 45230
rect 37996 45166 37998 45218
rect 38050 45166 38052 45218
rect 37772 44100 37828 44110
rect 37772 43426 37828 44044
rect 37996 43540 38052 45166
rect 38780 45108 38836 45118
rect 38556 44322 38612 44334
rect 38556 44270 38558 44322
rect 38610 44270 38612 44322
rect 38332 44212 38388 44222
rect 38332 44118 38388 44156
rect 38556 44100 38612 44270
rect 38556 44034 38612 44044
rect 37996 43474 38052 43484
rect 37772 43374 37774 43426
rect 37826 43374 37828 43426
rect 37772 43362 37828 43374
rect 38780 43092 38836 45052
rect 38892 43538 38948 45948
rect 39676 45938 39732 45948
rect 39340 45778 39396 45790
rect 39340 45726 39342 45778
rect 39394 45726 39396 45778
rect 39340 45332 39396 45726
rect 40460 45444 40516 46396
rect 40908 46386 40964 46396
rect 40348 45388 40516 45444
rect 39340 45276 39844 45332
rect 39676 45108 39732 45118
rect 39676 45014 39732 45052
rect 39788 44996 39844 45276
rect 40348 45218 40404 45388
rect 40348 45166 40350 45218
rect 40402 45166 40404 45218
rect 40348 45154 40404 45166
rect 40796 45108 40852 45118
rect 40012 44996 40068 45006
rect 39788 44994 40068 44996
rect 39788 44942 40014 44994
rect 40066 44942 40068 44994
rect 39788 44940 40068 44942
rect 39452 44322 39508 44334
rect 39452 44270 39454 44322
rect 39506 44270 39508 44322
rect 39452 44100 39508 44270
rect 39452 44034 39508 44044
rect 39900 44322 39956 44334
rect 39900 44270 39902 44322
rect 39954 44270 39956 44322
rect 39900 43876 39956 44270
rect 39900 43810 39956 43820
rect 39676 43764 39732 43774
rect 38892 43486 38894 43538
rect 38946 43486 38948 43538
rect 38892 43316 38948 43486
rect 38892 43250 38948 43260
rect 39004 43650 39060 43662
rect 39004 43598 39006 43650
rect 39058 43598 39060 43650
rect 39004 43540 39060 43598
rect 39228 43652 39284 43662
rect 39228 43558 39284 43596
rect 39676 43650 39732 43708
rect 39676 43598 39678 43650
rect 39730 43598 39732 43650
rect 39676 43586 39732 43598
rect 39004 43428 39060 43484
rect 39452 43538 39508 43550
rect 39452 43486 39454 43538
rect 39506 43486 39508 43538
rect 39452 43428 39508 43486
rect 39004 43372 39508 43428
rect 39564 43540 39620 43550
rect 38780 43036 38948 43092
rect 38668 42308 38724 42318
rect 38444 41972 38500 41982
rect 38108 41524 38164 41534
rect 38108 40962 38164 41468
rect 38444 41074 38500 41916
rect 38668 41858 38724 42252
rect 38668 41806 38670 41858
rect 38722 41806 38724 41858
rect 38668 41794 38724 41806
rect 38444 41022 38446 41074
rect 38498 41022 38500 41074
rect 38444 41010 38500 41022
rect 38108 40910 38110 40962
rect 38162 40910 38164 40962
rect 38108 40852 38164 40910
rect 38108 40786 38164 40796
rect 38780 40962 38836 40974
rect 38780 40910 38782 40962
rect 38834 40910 38836 40962
rect 37772 40404 37828 40414
rect 37772 40290 37828 40348
rect 38780 40404 38836 40910
rect 38780 40338 38836 40348
rect 37772 40238 37774 40290
rect 37826 40238 37828 40290
rect 37772 40226 37828 40238
rect 37772 40068 37828 40078
rect 37772 39730 37828 40012
rect 37772 39678 37774 39730
rect 37826 39678 37828 39730
rect 37772 39666 37828 39678
rect 37660 39442 37716 39452
rect 36652 38658 36708 38668
rect 36988 38948 37044 38958
rect 36540 38612 36596 38622
rect 36204 38164 36260 38174
rect 36092 38162 36260 38164
rect 36092 38110 36206 38162
rect 36258 38110 36260 38162
rect 36092 38108 36260 38110
rect 36204 38098 36260 38108
rect 35532 37762 35588 37772
rect 36428 37716 36484 37726
rect 36428 37492 36484 37660
rect 35868 37490 36484 37492
rect 35868 37438 36430 37490
rect 36482 37438 36484 37490
rect 35868 37436 36484 37438
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 34412 35758 34414 35810
rect 34466 35758 34468 35810
rect 34412 35746 34468 35758
rect 34636 36428 34916 36484
rect 34636 35812 34692 36428
rect 35868 36370 35924 37436
rect 36428 37426 36484 37436
rect 36204 37268 36260 37278
rect 36204 37174 36260 37212
rect 36540 37266 36596 38556
rect 36540 37214 36542 37266
rect 36594 37214 36596 37266
rect 35980 37154 36036 37166
rect 35980 37102 35982 37154
rect 36034 37102 36036 37154
rect 35980 36484 36036 37102
rect 36540 37044 36596 37214
rect 36876 38500 36932 38510
rect 36876 37268 36932 38444
rect 36988 37492 37044 38892
rect 37100 38946 37156 38958
rect 37100 38894 37102 38946
rect 37154 38894 37156 38946
rect 37100 37716 37156 38894
rect 37884 38948 37940 38958
rect 38444 38948 38500 38958
rect 37884 38946 38164 38948
rect 37884 38894 37886 38946
rect 37938 38894 38164 38946
rect 37884 38892 38164 38894
rect 37884 38882 37940 38892
rect 37772 38834 37828 38846
rect 37772 38782 37774 38834
rect 37826 38782 37828 38834
rect 37212 38722 37268 38734
rect 37212 38670 37214 38722
rect 37266 38670 37268 38722
rect 37212 38276 37268 38670
rect 37324 38722 37380 38734
rect 37324 38670 37326 38722
rect 37378 38670 37380 38722
rect 37324 38612 37380 38670
rect 37324 38546 37380 38556
rect 37772 38500 37828 38782
rect 37884 38612 37940 38622
rect 37884 38518 37940 38556
rect 37772 38434 37828 38444
rect 37212 38220 37940 38276
rect 37100 37650 37156 37660
rect 37660 37938 37716 37950
rect 37660 37886 37662 37938
rect 37714 37886 37716 37938
rect 37212 37604 37268 37614
rect 36988 37436 37156 37492
rect 37100 37378 37156 37436
rect 37100 37326 37102 37378
rect 37154 37326 37156 37378
rect 36876 37266 37044 37268
rect 36876 37214 36878 37266
rect 36930 37214 37044 37266
rect 36876 37212 37044 37214
rect 36876 37202 36932 37212
rect 36652 37044 36708 37054
rect 36540 36988 36652 37044
rect 36652 36978 36708 36988
rect 36988 36708 37044 37212
rect 37100 37044 37156 37326
rect 37212 37378 37268 37548
rect 37660 37490 37716 37886
rect 37660 37438 37662 37490
rect 37714 37438 37716 37490
rect 37660 37426 37716 37438
rect 37212 37326 37214 37378
rect 37266 37326 37268 37378
rect 37212 37268 37268 37326
rect 37212 37202 37268 37212
rect 37100 36988 37604 37044
rect 36988 36652 37492 36708
rect 36092 36484 36148 36494
rect 35980 36428 36092 36484
rect 36092 36390 36148 36428
rect 36988 36484 37044 36494
rect 36988 36390 37044 36428
rect 37212 36484 37268 36494
rect 37212 36390 37268 36428
rect 35868 36318 35870 36370
rect 35922 36318 35924 36370
rect 35868 36306 35924 36318
rect 34076 35700 34132 35710
rect 34076 34914 34132 35644
rect 34636 35698 34692 35756
rect 36988 35812 37044 35822
rect 37436 35812 37492 36652
rect 37548 36706 37604 36988
rect 37548 36654 37550 36706
rect 37602 36654 37604 36706
rect 37548 36642 37604 36654
rect 37884 36482 37940 38220
rect 37996 38052 38052 38062
rect 38108 38052 38164 38892
rect 38444 38854 38500 38892
rect 38332 38836 38388 38846
rect 38332 38742 38388 38780
rect 38668 38834 38724 38846
rect 38668 38782 38670 38834
rect 38722 38782 38724 38834
rect 38332 38052 38388 38062
rect 38108 38050 38388 38052
rect 38108 37998 38334 38050
rect 38386 37998 38388 38050
rect 38108 37996 38388 37998
rect 37996 36594 38052 37996
rect 37996 36542 37998 36594
rect 38050 36542 38052 36594
rect 37996 36530 38052 36542
rect 38108 36820 38164 36830
rect 37884 36430 37886 36482
rect 37938 36430 37940 36482
rect 37884 36418 37940 36430
rect 38108 36482 38164 36764
rect 38332 36596 38388 37996
rect 38444 37268 38500 37278
rect 38668 37268 38724 38782
rect 38444 37266 38724 37268
rect 38444 37214 38446 37266
rect 38498 37214 38724 37266
rect 38444 37212 38724 37214
rect 38780 38836 38836 38846
rect 38780 37604 38836 38780
rect 38892 38162 38948 43036
rect 39004 41970 39060 43372
rect 39564 43316 39620 43484
rect 39004 41918 39006 41970
rect 39058 41918 39060 41970
rect 39004 41906 39060 41918
rect 39228 43260 39620 43316
rect 39788 43316 39844 43326
rect 39228 41970 39284 43260
rect 39788 43222 39844 43260
rect 40012 42644 40068 44940
rect 40124 44324 40180 44334
rect 40124 44230 40180 44268
rect 40460 44322 40516 44334
rect 40460 44270 40462 44322
rect 40514 44270 40516 44322
rect 40236 44212 40292 44222
rect 40236 43650 40292 44156
rect 40236 43598 40238 43650
rect 40290 43598 40292 43650
rect 40236 43540 40292 43598
rect 40236 43474 40292 43484
rect 40348 43876 40404 43886
rect 40348 43538 40404 43820
rect 40348 43486 40350 43538
rect 40402 43486 40404 43538
rect 40348 43428 40404 43486
rect 40348 43362 40404 43372
rect 40460 43652 40516 44270
rect 40796 44322 40852 45052
rect 41020 44772 41076 46620
rect 41244 46452 41300 46462
rect 41244 46358 41300 46396
rect 41580 45892 41636 47404
rect 42140 47346 42196 47358
rect 42140 47294 42142 47346
rect 42194 47294 42196 47346
rect 42140 46900 42196 47294
rect 42140 46834 42196 46844
rect 44604 46676 44660 49644
rect 44940 49028 44996 49038
rect 45052 49028 45108 50652
rect 45500 50642 45556 50652
rect 45948 50428 46004 52668
rect 46620 52500 46676 52894
rect 46620 52434 46676 52444
rect 47404 52500 47460 52510
rect 46620 52276 46676 52286
rect 46620 52182 46676 52220
rect 46508 52164 46564 52174
rect 46508 52070 46564 52108
rect 46732 52162 46788 52174
rect 46732 52110 46734 52162
rect 46786 52110 46788 52162
rect 46172 51940 46228 51950
rect 46172 51938 46452 51940
rect 46172 51886 46174 51938
rect 46226 51886 46452 51938
rect 46172 51884 46452 51886
rect 46172 51874 46228 51884
rect 46060 51490 46116 51502
rect 46060 51438 46062 51490
rect 46114 51438 46116 51490
rect 46060 51380 46116 51438
rect 46396 51380 46452 51884
rect 46620 51604 46676 51614
rect 46620 51510 46676 51548
rect 46508 51380 46564 51390
rect 46396 51378 46564 51380
rect 46396 51326 46510 51378
rect 46562 51326 46564 51378
rect 46396 51324 46564 51326
rect 46060 51314 46116 51324
rect 46508 51314 46564 51324
rect 46732 50428 46788 52110
rect 46956 52164 47012 52174
rect 46956 51828 47012 52108
rect 47068 52052 47124 52062
rect 47068 51958 47124 51996
rect 47404 51938 47460 52444
rect 47740 52164 47796 53790
rect 47964 53172 48020 53182
rect 48076 53172 48132 54348
rect 48412 53732 48468 54348
rect 50092 53844 50148 53854
rect 48412 53730 48580 53732
rect 48412 53678 48414 53730
rect 48466 53678 48580 53730
rect 48412 53676 48580 53678
rect 48412 53666 48468 53676
rect 47964 53170 48132 53172
rect 47964 53118 47966 53170
rect 48018 53118 48132 53170
rect 47964 53116 48132 53118
rect 47964 53106 48020 53116
rect 48076 52164 48132 52174
rect 47740 52162 48132 52164
rect 47740 52110 47742 52162
rect 47794 52110 48078 52162
rect 48130 52110 48132 52162
rect 47740 52108 48132 52110
rect 47740 52098 47796 52108
rect 48076 52098 48132 52108
rect 48188 52164 48244 52174
rect 47404 51886 47406 51938
rect 47458 51886 47460 51938
rect 46956 51772 47124 51828
rect 47068 51378 47124 51772
rect 47404 51604 47460 51886
rect 47404 51548 48020 51604
rect 47068 51326 47070 51378
rect 47122 51326 47124 51378
rect 47068 51314 47124 51326
rect 47180 51490 47236 51502
rect 47180 51438 47182 51490
rect 47234 51438 47236 51490
rect 47180 51380 47236 51438
rect 47180 51314 47236 51324
rect 47740 51380 47796 51390
rect 45948 50372 46116 50428
rect 44940 49026 45108 49028
rect 44940 48974 44942 49026
rect 44994 48974 45108 49026
rect 44940 48972 45108 48974
rect 45388 49698 45444 49710
rect 45388 49646 45390 49698
rect 45442 49646 45444 49698
rect 44940 48962 44996 48972
rect 45388 48356 45444 49646
rect 46060 49140 46116 50372
rect 45612 48914 45668 48926
rect 45612 48862 45614 48914
rect 45666 48862 45668 48914
rect 45612 48468 45668 48862
rect 45836 48468 45892 48478
rect 45612 48466 45892 48468
rect 45612 48414 45838 48466
rect 45890 48414 45892 48466
rect 45612 48412 45892 48414
rect 45836 48402 45892 48412
rect 45388 48290 45444 48300
rect 46060 48242 46116 49084
rect 46060 48190 46062 48242
rect 46114 48190 46116 48242
rect 46060 48178 46116 48190
rect 46284 50372 46788 50428
rect 47292 50594 47348 50606
rect 47292 50542 47294 50594
rect 47346 50542 47348 50594
rect 46172 48132 46228 48142
rect 46172 48038 46228 48076
rect 44828 47572 44884 47582
rect 44604 46610 44660 46620
rect 44716 47516 44828 47572
rect 44380 46564 44436 46574
rect 44380 46470 44436 46508
rect 41804 46452 41860 46462
rect 41804 46002 41860 46396
rect 44604 46452 44660 46462
rect 44716 46452 44772 47516
rect 44828 47478 44884 47516
rect 45164 47572 45220 47582
rect 45500 47572 45556 47582
rect 45164 47570 45332 47572
rect 45164 47518 45166 47570
rect 45218 47518 45332 47570
rect 45164 47516 45332 47518
rect 45164 47506 45220 47516
rect 45052 47236 45108 47246
rect 44940 46676 44996 46686
rect 44940 46582 44996 46620
rect 45052 46564 45108 47180
rect 45164 46900 45220 46910
rect 45164 46564 45220 46844
rect 45276 46788 45332 47516
rect 45500 47458 45556 47516
rect 46284 47572 46340 50372
rect 47068 49812 47124 49822
rect 47292 49812 47348 50542
rect 47124 49756 47348 49812
rect 47068 49718 47124 49756
rect 47740 49140 47796 51324
rect 47964 51378 48020 51548
rect 47964 51326 47966 51378
rect 48018 51326 48020 51378
rect 47964 49700 48020 51326
rect 48076 51490 48132 51502
rect 48076 51438 48078 51490
rect 48130 51438 48132 51490
rect 48076 51380 48132 51438
rect 48076 51314 48132 51324
rect 48076 51154 48132 51166
rect 48076 51102 48078 51154
rect 48130 51102 48132 51154
rect 48076 49924 48132 51102
rect 48188 50594 48244 52108
rect 48300 52052 48356 52062
rect 48300 50706 48356 51996
rect 48300 50654 48302 50706
rect 48354 50654 48356 50706
rect 48300 50642 48356 50654
rect 48524 50708 48580 53676
rect 49196 53620 49252 53630
rect 48972 53618 49252 53620
rect 48972 53566 49198 53618
rect 49250 53566 49252 53618
rect 48972 53564 49252 53566
rect 48972 53170 49028 53564
rect 49196 53554 49252 53564
rect 48972 53118 48974 53170
rect 49026 53118 49028 53170
rect 48972 53106 49028 53118
rect 48748 52946 48804 52958
rect 50092 52948 50148 53788
rect 51324 53844 51380 53854
rect 51324 53750 51380 53788
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 48748 52894 48750 52946
rect 48802 52894 48804 52946
rect 48748 52724 48804 52894
rect 49644 52946 50148 52948
rect 49644 52894 50094 52946
rect 50146 52894 50148 52946
rect 49644 52892 50148 52894
rect 49084 52836 49140 52846
rect 49420 52836 49476 52846
rect 49084 52834 49476 52836
rect 49084 52782 49086 52834
rect 49138 52782 49422 52834
rect 49474 52782 49476 52834
rect 49084 52780 49476 52782
rect 49084 52770 49140 52780
rect 49420 52770 49476 52780
rect 48748 52658 48804 52668
rect 49644 52612 49700 52892
rect 50092 52882 50148 52892
rect 50316 52836 50372 52846
rect 50316 52834 50932 52836
rect 50316 52782 50318 52834
rect 50370 52782 50932 52834
rect 50316 52780 50932 52782
rect 50316 52770 50372 52780
rect 48860 52556 49700 52612
rect 48860 51490 48916 52556
rect 48860 51438 48862 51490
rect 48914 51438 48916 51490
rect 48860 51426 48916 51438
rect 49420 52388 49476 52398
rect 49420 51938 49476 52332
rect 49420 51886 49422 51938
rect 49474 51886 49476 51938
rect 49196 51380 49252 51390
rect 49252 51324 49364 51380
rect 49196 51286 49252 51324
rect 48188 50542 48190 50594
rect 48242 50542 48244 50594
rect 48188 50530 48244 50542
rect 48412 50596 48468 50606
rect 48412 50502 48468 50540
rect 48524 50428 48580 50652
rect 48748 51154 48804 51166
rect 48748 51102 48750 51154
rect 48802 51102 48804 51154
rect 48748 50596 48804 51102
rect 48748 50530 48804 50540
rect 48860 50594 48916 50606
rect 48860 50542 48862 50594
rect 48914 50542 48916 50594
rect 48076 49858 48132 49868
rect 48300 50372 48580 50428
rect 48860 50428 48916 50542
rect 48860 50372 49028 50428
rect 47964 49634 48020 49644
rect 47516 49138 48132 49140
rect 47516 49086 47742 49138
rect 47794 49086 48132 49138
rect 47516 49084 48132 49086
rect 45500 47406 45502 47458
rect 45554 47406 45556 47458
rect 45500 47394 45556 47406
rect 45836 47460 45892 47470
rect 45836 47366 45892 47404
rect 46172 47460 46228 47470
rect 46284 47460 46340 47516
rect 46172 47458 46340 47460
rect 46172 47406 46174 47458
rect 46226 47406 46340 47458
rect 46172 47404 46340 47406
rect 46172 47394 46228 47404
rect 45724 47348 45780 47358
rect 45612 47236 45668 47246
rect 45612 47142 45668 47180
rect 45276 46732 45668 46788
rect 45612 46674 45668 46732
rect 45612 46622 45614 46674
rect 45666 46622 45668 46674
rect 45612 46610 45668 46622
rect 45276 46564 45332 46574
rect 45164 46562 45332 46564
rect 45164 46510 45278 46562
rect 45330 46510 45332 46562
rect 45164 46508 45332 46510
rect 45052 46498 45108 46508
rect 45276 46498 45332 46508
rect 45500 46564 45556 46574
rect 44604 46450 44772 46452
rect 44604 46398 44606 46450
rect 44658 46398 44772 46450
rect 44604 46396 44772 46398
rect 45388 46452 45444 46462
rect 44604 46386 44660 46396
rect 45388 46358 45444 46396
rect 41804 45950 41806 46002
rect 41858 45950 41860 46002
rect 41804 45938 41860 45950
rect 41468 45108 41524 45118
rect 41580 45108 41636 45836
rect 42588 45892 42644 45902
rect 42588 45798 42644 45836
rect 43036 45892 43092 45902
rect 43036 45798 43092 45836
rect 44940 45892 44996 45902
rect 44940 45668 44996 45836
rect 45500 45890 45556 46508
rect 45500 45838 45502 45890
rect 45554 45838 45556 45890
rect 45500 45826 45556 45838
rect 45724 46450 45780 47292
rect 46284 46564 46340 47404
rect 46396 48356 46452 48366
rect 46396 47572 46452 48300
rect 47068 48356 47124 48366
rect 46620 48242 46676 48254
rect 46620 48190 46622 48242
rect 46674 48190 46676 48242
rect 46620 47684 46676 48190
rect 47068 48242 47124 48300
rect 47068 48190 47070 48242
rect 47122 48190 47124 48242
rect 47068 48178 47124 48190
rect 47180 48242 47236 48254
rect 47180 48190 47182 48242
rect 47234 48190 47236 48242
rect 47180 47684 47236 48190
rect 47404 48132 47460 48142
rect 47404 48038 47460 48076
rect 46620 47628 47236 47684
rect 46396 47516 46788 47572
rect 46396 47458 46452 47516
rect 46396 47406 46398 47458
rect 46450 47406 46452 47458
rect 46396 47394 46452 47406
rect 46620 47348 46676 47358
rect 46620 47254 46676 47292
rect 46508 47234 46564 47246
rect 46508 47182 46510 47234
rect 46562 47182 46564 47234
rect 46508 46788 46564 47182
rect 46508 46722 46564 46732
rect 46732 46786 46788 47516
rect 46844 47348 46900 47628
rect 47292 47460 47348 47470
rect 47292 47366 47348 47404
rect 47516 47458 47572 49084
rect 47740 49074 47796 49084
rect 47852 48356 47908 48366
rect 47852 48262 47908 48300
rect 47628 48242 47684 48254
rect 47628 48190 47630 48242
rect 47682 48190 47684 48242
rect 47628 47572 47684 48190
rect 48076 48242 48132 49084
rect 48300 49138 48356 50372
rect 48748 49924 48804 49934
rect 48748 49830 48804 49868
rect 48972 49810 49028 50372
rect 48972 49758 48974 49810
rect 49026 49758 49028 49810
rect 48972 49476 49028 49758
rect 49084 50036 49140 50046
rect 49084 49698 49140 49980
rect 49084 49646 49086 49698
rect 49138 49646 49140 49698
rect 49084 49634 49140 49646
rect 48972 49410 49028 49420
rect 48300 49086 48302 49138
rect 48354 49086 48356 49138
rect 48300 49074 48356 49086
rect 48748 49252 48804 49262
rect 48076 48190 48078 48242
rect 48130 48190 48132 48242
rect 48076 48178 48132 48190
rect 47964 47572 48020 47582
rect 48524 47572 48580 47582
rect 47628 47570 48580 47572
rect 47628 47518 47966 47570
rect 48018 47518 48526 47570
rect 48578 47518 48580 47570
rect 47628 47516 48580 47518
rect 47964 47506 48020 47516
rect 48524 47506 48580 47516
rect 47516 47406 47518 47458
rect 47570 47406 47572 47458
rect 47516 47394 47572 47406
rect 46844 47282 46900 47292
rect 48300 47348 48356 47358
rect 48300 47254 48356 47292
rect 46732 46734 46734 46786
rect 46786 46734 46788 46786
rect 46732 46722 46788 46734
rect 47740 47012 47796 47022
rect 46620 46674 46676 46686
rect 46620 46622 46622 46674
rect 46674 46622 46676 46674
rect 46620 46564 46676 46622
rect 46844 46676 46900 46686
rect 46844 46582 46900 46620
rect 47292 46676 47348 46686
rect 47292 46582 47348 46620
rect 45724 46398 45726 46450
rect 45778 46398 45780 46450
rect 45724 45778 45780 46398
rect 46172 46508 46676 46564
rect 46172 46002 46228 46508
rect 47740 46452 47796 46956
rect 48748 47012 48804 49196
rect 49308 49028 49364 51324
rect 49420 51378 49476 51886
rect 49644 51602 49700 52556
rect 49980 52724 50036 52734
rect 49644 51550 49646 51602
rect 49698 51550 49700 51602
rect 49644 51538 49700 51550
rect 49756 52164 49812 52174
rect 49756 51938 49812 52108
rect 49756 51886 49758 51938
rect 49810 51886 49812 51938
rect 49756 51380 49812 51886
rect 49420 51326 49422 51378
rect 49474 51326 49476 51378
rect 49420 51268 49476 51326
rect 49420 51202 49476 51212
rect 49644 51324 49812 51380
rect 49980 51378 50036 52668
rect 50316 52164 50372 52174
rect 50204 52162 50372 52164
rect 50204 52110 50318 52162
rect 50370 52110 50372 52162
rect 50204 52108 50372 52110
rect 49980 51326 49982 51378
rect 50034 51326 50036 51378
rect 49644 50482 49700 51324
rect 49980 51314 50036 51326
rect 50092 52050 50148 52062
rect 50092 51998 50094 52050
rect 50146 51998 50148 52050
rect 49756 51154 49812 51166
rect 49756 51102 49758 51154
rect 49810 51102 49812 51154
rect 49756 50932 49812 51102
rect 49756 50866 49812 50876
rect 49644 50430 49646 50482
rect 49698 50430 49700 50482
rect 49644 50418 49700 50430
rect 49868 50484 49924 50494
rect 50092 50484 50148 51998
rect 50204 51380 50260 52108
rect 50316 52098 50372 52108
rect 50428 52164 50484 52174
rect 50540 52164 50596 52174
rect 50484 52162 50596 52164
rect 50484 52110 50542 52162
rect 50594 52110 50596 52162
rect 50484 52108 50596 52110
rect 50204 51314 50260 51324
rect 50316 51938 50372 51950
rect 50316 51886 50318 51938
rect 50370 51886 50372 51938
rect 50316 51378 50372 51886
rect 50316 51326 50318 51378
rect 50370 51326 50372 51378
rect 50316 51314 50372 51326
rect 50428 51378 50484 52108
rect 50540 52098 50596 52108
rect 50876 52162 50932 52780
rect 50876 52110 50878 52162
rect 50930 52110 50932 52162
rect 50876 52098 50932 52110
rect 51100 52164 51156 52174
rect 51100 52050 51156 52108
rect 51100 51998 51102 52050
rect 51154 51998 51156 52050
rect 51100 51986 51156 51998
rect 51212 52050 51268 52062
rect 51212 51998 51214 52050
rect 51266 51998 51268 52050
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 51212 51604 51268 51998
rect 51212 51538 51268 51548
rect 50652 51492 50708 51502
rect 50652 51398 50708 51436
rect 53228 51492 53284 51502
rect 50428 51326 50430 51378
rect 50482 51326 50484 51378
rect 50428 51314 50484 51326
rect 50764 51380 50820 51418
rect 53228 51398 53284 51436
rect 50820 51324 50932 51380
rect 50764 51314 50820 51324
rect 50764 51156 50820 51166
rect 50316 50932 50372 50942
rect 50316 50706 50372 50876
rect 50316 50654 50318 50706
rect 50370 50654 50372 50706
rect 50316 50642 50372 50654
rect 50764 50820 50820 51100
rect 50764 50594 50820 50764
rect 50764 50542 50766 50594
rect 50818 50542 50820 50594
rect 50764 50530 50820 50542
rect 49868 50482 50148 50484
rect 49868 50430 49870 50482
rect 49922 50430 50148 50482
rect 49868 50428 50148 50430
rect 49756 50370 49812 50382
rect 49756 50318 49758 50370
rect 49810 50318 49812 50370
rect 49756 49924 49812 50318
rect 49868 50036 49924 50428
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 49868 49970 49924 49980
rect 49756 49858 49812 49868
rect 50764 49924 50820 49934
rect 50764 49830 50820 49868
rect 49868 49810 49924 49822
rect 49868 49758 49870 49810
rect 49922 49758 49924 49810
rect 49308 49026 49588 49028
rect 49308 48974 49310 49026
rect 49362 48974 49588 49026
rect 49308 48972 49588 48974
rect 49308 48962 49364 48972
rect 49084 48804 49140 48814
rect 48972 48802 49140 48804
rect 48972 48750 49086 48802
rect 49138 48750 49140 48802
rect 48972 48748 49140 48750
rect 48972 48692 49028 48748
rect 49084 48738 49140 48748
rect 48860 47572 48916 47582
rect 48860 47478 48916 47516
rect 48972 47124 49028 48636
rect 49196 48468 49252 48478
rect 49196 48130 49252 48412
rect 49532 48466 49588 48972
rect 49644 48804 49700 48814
rect 49644 48710 49700 48748
rect 49532 48414 49534 48466
rect 49586 48414 49588 48466
rect 49532 48402 49588 48414
rect 49868 48244 49924 49758
rect 50876 49812 50932 51324
rect 53900 51378 53956 51390
rect 53900 51326 53902 51378
rect 53954 51326 53956 51378
rect 51100 51268 51156 51278
rect 51100 51174 51156 51212
rect 51996 51268 52052 51278
rect 51996 50820 52052 51212
rect 51660 50708 51716 50718
rect 51660 50614 51716 50652
rect 51884 50596 51940 50606
rect 51212 50484 51268 50494
rect 51100 50482 51268 50484
rect 51100 50430 51214 50482
rect 51266 50430 51268 50482
rect 51100 50428 51268 50430
rect 50988 49812 51044 49822
rect 50876 49810 51044 49812
rect 50876 49758 50990 49810
rect 51042 49758 51044 49810
rect 50876 49756 51044 49758
rect 51100 49812 51156 50428
rect 51212 50418 51268 50428
rect 51548 50484 51604 50494
rect 51548 50034 51604 50428
rect 51548 49982 51550 50034
rect 51602 49982 51604 50034
rect 51548 49970 51604 49982
rect 51884 49922 51940 50540
rect 51996 50034 52052 50764
rect 52108 50708 52164 50718
rect 52108 50614 52164 50652
rect 52668 50708 52724 50718
rect 52668 50594 52724 50652
rect 53900 50708 53956 51326
rect 53900 50642 53956 50652
rect 55580 51268 55636 51278
rect 55580 50706 55636 51212
rect 55580 50654 55582 50706
rect 55634 50654 55636 50706
rect 55580 50642 55636 50654
rect 52668 50542 52670 50594
rect 52722 50542 52724 50594
rect 52668 50530 52724 50542
rect 53452 50484 53508 50494
rect 53452 50390 53508 50428
rect 51996 49982 51998 50034
rect 52050 49982 52052 50034
rect 51996 49970 52052 49982
rect 52220 50036 52276 50046
rect 52220 49942 52276 49980
rect 51884 49870 51886 49922
rect 51938 49870 51940 49922
rect 51884 49858 51940 49870
rect 51212 49812 51268 49822
rect 51100 49810 51268 49812
rect 51100 49758 51214 49810
rect 51266 49758 51268 49810
rect 51100 49756 51268 49758
rect 49980 49700 50036 49710
rect 50988 49700 51044 49756
rect 51212 49746 51268 49756
rect 51324 49810 51380 49822
rect 51324 49758 51326 49810
rect 51378 49758 51380 49810
rect 50988 49644 51156 49700
rect 49980 49606 50036 49644
rect 50316 49140 50372 49150
rect 50092 49028 50148 49038
rect 49980 48802 50036 48814
rect 49980 48750 49982 48802
rect 50034 48750 50036 48802
rect 49980 48692 50036 48750
rect 49980 48626 50036 48636
rect 49196 48078 49198 48130
rect 49250 48078 49252 48130
rect 48972 47058 49028 47068
rect 49084 48018 49140 48030
rect 49084 47966 49086 48018
rect 49138 47966 49140 48018
rect 49084 47570 49140 47966
rect 49084 47518 49086 47570
rect 49138 47518 49140 47570
rect 48748 46946 48804 46956
rect 48076 46900 48132 46910
rect 48076 46898 48356 46900
rect 48076 46846 48078 46898
rect 48130 46846 48356 46898
rect 48076 46844 48356 46846
rect 48076 46834 48132 46844
rect 47964 46788 48020 46798
rect 47964 46674 48020 46732
rect 47964 46622 47966 46674
rect 48018 46622 48020 46674
rect 47964 46610 48020 46622
rect 48076 46676 48132 46686
rect 48076 46582 48132 46620
rect 47740 46358 47796 46396
rect 46172 45950 46174 46002
rect 46226 45950 46228 46002
rect 46172 45938 46228 45950
rect 48300 46002 48356 46844
rect 48860 46676 48916 46686
rect 48860 46582 48916 46620
rect 49084 46676 49140 47518
rect 49084 46582 49140 46620
rect 48300 45950 48302 46002
rect 48354 45950 48356 46002
rect 48300 45938 48356 45950
rect 45724 45726 45726 45778
rect 45778 45726 45780 45778
rect 45724 45714 45780 45726
rect 49084 45892 49140 45902
rect 49196 45892 49252 48078
rect 49308 48188 49924 48244
rect 50092 48242 50148 48972
rect 50092 48190 50094 48242
rect 50146 48190 50148 48242
rect 49308 48018 49364 48188
rect 50092 48178 50148 48190
rect 50204 48916 50260 48926
rect 49308 47966 49310 48018
rect 49362 47966 49364 48018
rect 49308 47954 49364 47966
rect 49868 48020 49924 48030
rect 50204 48020 50260 48860
rect 50316 48914 50372 49084
rect 50988 49138 51044 49150
rect 50988 49086 50990 49138
rect 51042 49086 51044 49138
rect 50652 49028 50708 49038
rect 50316 48862 50318 48914
rect 50370 48862 50372 48914
rect 50316 48850 50372 48862
rect 50540 49026 50708 49028
rect 50540 48974 50654 49026
rect 50706 48974 50708 49026
rect 50540 48972 50708 48974
rect 50540 48916 50596 48972
rect 50652 48962 50708 48972
rect 50876 49028 50932 49038
rect 50540 48850 50596 48860
rect 50876 48914 50932 48972
rect 50876 48862 50878 48914
rect 50930 48862 50932 48914
rect 49868 48018 50260 48020
rect 49868 47966 49870 48018
rect 49922 47966 50260 48018
rect 49868 47964 50260 47966
rect 50428 48804 50484 48814
rect 49868 47348 49924 47964
rect 50428 47682 50484 48748
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50540 48468 50596 48478
rect 50540 48242 50596 48412
rect 50876 48468 50932 48862
rect 50876 48402 50932 48412
rect 50540 48190 50542 48242
rect 50594 48190 50596 48242
rect 50540 48178 50596 48190
rect 50988 48020 51044 49086
rect 51100 48804 51156 49644
rect 51324 49252 51380 49758
rect 51324 49186 51380 49196
rect 51100 48738 51156 48748
rect 53452 48468 53508 48478
rect 51324 48132 51380 48142
rect 50428 47630 50430 47682
rect 50482 47630 50484 47682
rect 50428 47618 50484 47630
rect 50540 47964 51044 48020
rect 51100 48130 51380 48132
rect 51100 48078 51326 48130
rect 51378 48078 51380 48130
rect 51100 48076 51380 48078
rect 50540 47682 50596 47964
rect 50540 47630 50542 47682
rect 50594 47630 50596 47682
rect 50540 47618 50596 47630
rect 50876 47684 50932 47694
rect 51100 47684 51156 48076
rect 51324 48066 51380 48076
rect 53452 48130 53508 48412
rect 53452 48078 53454 48130
rect 53506 48078 53508 48130
rect 53452 48066 53508 48078
rect 50876 47682 51156 47684
rect 50876 47630 50878 47682
rect 50930 47630 51156 47682
rect 50876 47628 51156 47630
rect 50876 47618 50932 47628
rect 50764 47458 50820 47470
rect 50764 47406 50766 47458
rect 50818 47406 50820 47458
rect 49868 47282 49924 47292
rect 50428 47348 50484 47358
rect 49644 47234 49700 47246
rect 49644 47182 49646 47234
rect 49698 47182 49700 47234
rect 49644 47124 49700 47182
rect 49644 47058 49700 47068
rect 49980 47234 50036 47246
rect 49980 47182 49982 47234
rect 50034 47182 50036 47234
rect 49980 47012 50036 47182
rect 49980 46946 50036 46956
rect 50204 46898 50260 46910
rect 50204 46846 50206 46898
rect 50258 46846 50260 46898
rect 49756 46676 49812 46686
rect 50092 46676 50148 46686
rect 49756 46674 50148 46676
rect 49756 46622 49758 46674
rect 49810 46622 50094 46674
rect 50146 46622 50148 46674
rect 49756 46620 50148 46622
rect 49756 46610 49812 46620
rect 50092 46610 50148 46620
rect 49084 45890 49252 45892
rect 49084 45838 49086 45890
rect 49138 45838 49252 45890
rect 49084 45836 49252 45838
rect 45052 45668 45108 45678
rect 44940 45666 45108 45668
rect 44940 45614 45054 45666
rect 45106 45614 45108 45666
rect 44940 45612 45108 45614
rect 44940 45444 44996 45612
rect 45052 45602 45108 45612
rect 44940 45330 44996 45388
rect 44940 45278 44942 45330
rect 44994 45278 44996 45330
rect 44940 45266 44996 45278
rect 47628 45332 47684 45342
rect 41468 45106 41636 45108
rect 41468 45054 41470 45106
rect 41522 45054 41636 45106
rect 41468 45052 41636 45054
rect 41468 45042 41524 45052
rect 41132 44994 41188 45006
rect 41132 44942 41134 44994
rect 41186 44942 41188 44994
rect 41132 44884 41188 44942
rect 42140 44996 42196 45006
rect 42140 44994 42420 44996
rect 42140 44942 42142 44994
rect 42194 44942 42420 44994
rect 42140 44940 42420 44942
rect 42140 44930 42196 44940
rect 41132 44828 41412 44884
rect 41020 44716 41300 44772
rect 40796 44270 40798 44322
rect 40850 44270 40852 44322
rect 40796 43876 40852 44270
rect 41020 44324 41076 44334
rect 41076 44268 41188 44324
rect 41020 44258 41076 44268
rect 40908 44100 40964 44110
rect 40908 44006 40964 44044
rect 41020 44098 41076 44110
rect 41020 44046 41022 44098
rect 41074 44046 41076 44098
rect 40796 43810 40852 43820
rect 41020 43764 41076 44046
rect 41020 43698 41076 43708
rect 40236 43314 40292 43326
rect 40236 43262 40238 43314
rect 40290 43262 40292 43314
rect 40236 42754 40292 43262
rect 40236 42702 40238 42754
rect 40290 42702 40292 42754
rect 40236 42690 40292 42702
rect 40124 42644 40180 42654
rect 40012 42588 40124 42644
rect 40124 42578 40180 42588
rect 40348 42644 40404 42654
rect 40460 42644 40516 43596
rect 40796 43540 40852 43550
rect 40572 43538 40852 43540
rect 40572 43486 40798 43538
rect 40850 43486 40852 43538
rect 40572 43484 40852 43486
rect 40572 42754 40628 43484
rect 40796 43474 40852 43484
rect 41132 43316 41188 44268
rect 40572 42702 40574 42754
rect 40626 42702 40628 42754
rect 40572 42690 40628 42702
rect 40796 43260 41188 43316
rect 40796 42754 40852 43260
rect 41244 43204 41300 44716
rect 40796 42702 40798 42754
rect 40850 42702 40852 42754
rect 40796 42690 40852 42702
rect 41020 43148 41300 43204
rect 41356 44322 41412 44828
rect 42364 44434 42420 44940
rect 42364 44382 42366 44434
rect 42418 44382 42420 44434
rect 42364 44370 42420 44382
rect 44380 44994 44436 45006
rect 44380 44942 44382 44994
rect 44434 44942 44436 44994
rect 41356 44270 41358 44322
rect 41410 44270 41412 44322
rect 40348 42642 40516 42644
rect 40348 42590 40350 42642
rect 40402 42590 40516 42642
rect 40348 42588 40516 42590
rect 40908 42644 40964 42654
rect 40348 42578 40404 42588
rect 40908 42550 40964 42588
rect 39788 42084 39844 42094
rect 40124 42084 40180 42094
rect 39788 42082 40180 42084
rect 39788 42030 39790 42082
rect 39842 42030 40126 42082
rect 40178 42030 40180 42082
rect 39788 42028 40180 42030
rect 39788 42018 39844 42028
rect 40124 42018 40180 42028
rect 40236 42082 40292 42094
rect 40236 42030 40238 42082
rect 40290 42030 40292 42082
rect 39228 41918 39230 41970
rect 39282 41918 39284 41970
rect 39228 41906 39284 41918
rect 39676 41972 39732 41982
rect 39452 41746 39508 41758
rect 39452 41694 39454 41746
rect 39506 41694 39508 41746
rect 39228 41300 39284 41310
rect 39228 41206 39284 41244
rect 39452 40964 39508 41694
rect 39564 41748 39620 41758
rect 39564 41410 39620 41692
rect 39564 41358 39566 41410
rect 39618 41358 39620 41410
rect 39564 41346 39620 41358
rect 39452 40516 39508 40908
rect 39676 40964 39732 41916
rect 40236 41860 40292 42030
rect 40460 41972 40516 41982
rect 39900 41804 40292 41860
rect 40348 41970 40516 41972
rect 40348 41918 40462 41970
rect 40514 41918 40516 41970
rect 40348 41916 40516 41918
rect 39900 41410 39956 41804
rect 40348 41748 40404 41916
rect 40460 41906 40516 41916
rect 39900 41358 39902 41410
rect 39954 41358 39956 41410
rect 39900 41346 39956 41358
rect 40124 41692 40404 41748
rect 39788 41300 39844 41310
rect 39788 41074 39844 41244
rect 39788 41022 39790 41074
rect 39842 41022 39844 41074
rect 39788 41010 39844 41022
rect 39676 40898 39732 40908
rect 40012 40516 40068 40526
rect 39452 40514 40068 40516
rect 39452 40462 40014 40514
rect 40066 40462 40068 40514
rect 39452 40460 40068 40462
rect 40012 40180 40068 40460
rect 40012 40114 40068 40124
rect 39900 39730 39956 39742
rect 39900 39678 39902 39730
rect 39954 39678 39956 39730
rect 39900 39620 39956 39678
rect 39900 39554 39956 39564
rect 40124 38668 40180 41692
rect 40348 40402 40404 40414
rect 40348 40350 40350 40402
rect 40402 40350 40404 40402
rect 40348 39620 40404 40350
rect 40348 39554 40404 39564
rect 41020 38668 41076 43148
rect 41132 42532 41188 42542
rect 41132 42438 41188 42476
rect 41356 42308 41412 44270
rect 41692 44324 41748 44334
rect 41692 44230 41748 44268
rect 42140 44322 42196 44334
rect 42140 44270 42142 44322
rect 42194 44270 42196 44322
rect 41804 44212 41860 44222
rect 41804 44118 41860 44156
rect 41916 44100 41972 44110
rect 42140 44100 42196 44270
rect 42476 44324 42532 44334
rect 42476 44230 42532 44268
rect 42700 44322 42756 44334
rect 42700 44270 42702 44322
rect 42754 44270 42756 44322
rect 42700 44212 42756 44270
rect 42700 44146 42756 44156
rect 41972 44044 42196 44100
rect 41916 44006 41972 44044
rect 42252 43876 42308 43886
rect 41580 43540 41636 43550
rect 41580 43446 41636 43484
rect 41804 43428 41860 43438
rect 41804 43334 41860 43372
rect 41244 42252 41412 42308
rect 41916 43314 41972 43326
rect 41916 43262 41918 43314
rect 41970 43262 41972 43314
rect 41916 42754 41972 43262
rect 41916 42702 41918 42754
rect 41970 42702 41972 42754
rect 41244 39284 41300 42252
rect 41804 42196 41860 42206
rect 41356 42194 41860 42196
rect 41356 42142 41806 42194
rect 41858 42142 41860 42194
rect 41356 42140 41860 42142
rect 41356 39844 41412 42140
rect 41804 42130 41860 42140
rect 41692 41970 41748 41982
rect 41692 41918 41694 41970
rect 41746 41918 41748 41970
rect 41692 41188 41748 41918
rect 41916 41972 41972 42702
rect 42252 42756 42308 43820
rect 44380 43428 44436 44942
rect 44828 44436 44884 44446
rect 47628 44436 47684 45276
rect 49084 45332 49140 45836
rect 49196 45332 49252 45342
rect 49140 45330 49588 45332
rect 49140 45278 49198 45330
rect 49250 45278 49588 45330
rect 49140 45276 49588 45278
rect 49084 45266 49140 45276
rect 49196 45266 49252 45276
rect 49532 45106 49588 45276
rect 50204 45220 50260 46846
rect 50316 46452 50372 46462
rect 50428 46452 50484 47292
rect 50764 47236 50820 47406
rect 50764 47170 50820 47180
rect 51324 47236 51380 47246
rect 51324 47142 51380 47180
rect 51772 47236 51828 47246
rect 51772 47142 51828 47180
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50540 46900 50596 46910
rect 50540 46674 50596 46844
rect 50540 46622 50542 46674
rect 50594 46622 50596 46674
rect 50540 46610 50596 46622
rect 51772 46676 51828 46686
rect 51772 46582 51828 46620
rect 51884 46676 51940 46686
rect 51884 46674 52052 46676
rect 51884 46622 51886 46674
rect 51938 46622 52052 46674
rect 51884 46620 52052 46622
rect 51884 46610 51940 46620
rect 50316 46450 50484 46452
rect 50316 46398 50318 46450
rect 50370 46398 50484 46450
rect 50316 46396 50484 46398
rect 50316 46386 50372 46396
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 51996 45332 52052 46620
rect 51996 45276 52500 45332
rect 50316 45220 50372 45230
rect 50204 45218 50372 45220
rect 50204 45166 50318 45218
rect 50370 45166 50372 45218
rect 50204 45164 50372 45166
rect 50316 45154 50372 45164
rect 49532 45054 49534 45106
rect 49586 45054 49588 45106
rect 49532 45042 49588 45054
rect 52444 44994 52500 45276
rect 52444 44942 52446 44994
rect 52498 44942 52500 44994
rect 52444 44930 52500 44942
rect 48188 44436 48244 44446
rect 44884 44380 44996 44436
rect 44828 44342 44884 44380
rect 44940 43652 44996 44380
rect 47628 44434 48244 44436
rect 47628 44382 48190 44434
rect 48242 44382 48244 44434
rect 47628 44380 48244 44382
rect 47628 44322 47684 44380
rect 47628 44270 47630 44322
rect 47682 44270 47684 44322
rect 47628 44258 47684 44270
rect 46956 44212 47012 44222
rect 44940 43538 44996 43596
rect 46508 44210 47012 44212
rect 46508 44158 46958 44210
rect 47010 44158 47012 44210
rect 46508 44156 47012 44158
rect 46508 43650 46564 44156
rect 46956 44146 47012 44156
rect 48188 43762 48244 44380
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 48188 43710 48190 43762
rect 48242 43710 48244 43762
rect 46508 43598 46510 43650
rect 46562 43598 46564 43650
rect 46508 43586 46564 43598
rect 47068 43652 47124 43662
rect 47068 43558 47124 43596
rect 44940 43486 44942 43538
rect 44994 43486 44996 43538
rect 44940 43474 44996 43486
rect 45612 43540 45668 43550
rect 45948 43540 46004 43550
rect 45612 43538 46004 43540
rect 45612 43486 45614 43538
rect 45666 43486 45950 43538
rect 46002 43486 46004 43538
rect 45612 43484 46004 43486
rect 45612 43474 45668 43484
rect 45948 43474 46004 43484
rect 48188 43540 48244 43710
rect 49980 43652 50036 43662
rect 48860 43540 48916 43550
rect 48188 43474 48244 43484
rect 48636 43484 48860 43540
rect 44716 43428 44772 43438
rect 43484 43316 43540 43326
rect 42252 42662 42308 42700
rect 43036 42754 43092 42766
rect 43036 42702 43038 42754
rect 43090 42702 43092 42754
rect 42812 42642 42868 42654
rect 42812 42590 42814 42642
rect 42866 42590 42868 42642
rect 42364 42530 42420 42542
rect 42364 42478 42366 42530
rect 42418 42478 42420 42530
rect 42252 41972 42308 41982
rect 41916 41970 42308 41972
rect 41916 41918 42254 41970
rect 42306 41918 42308 41970
rect 41916 41916 42308 41918
rect 42252 41906 42308 41916
rect 41804 41748 41860 41758
rect 41804 41654 41860 41692
rect 42364 41412 42420 42478
rect 42476 42532 42532 42542
rect 42812 42532 42868 42590
rect 42532 42476 42868 42532
rect 42476 42438 42532 42476
rect 43036 41972 43092 42702
rect 43372 42532 43428 42542
rect 43372 42438 43428 42476
rect 43372 41972 43428 41982
rect 43036 41970 43428 41972
rect 43036 41918 43374 41970
rect 43426 41918 43428 41970
rect 43036 41916 43428 41918
rect 43372 41748 43428 41916
rect 43372 41682 43428 41692
rect 43484 41524 43540 43260
rect 43372 41468 43540 41524
rect 44156 41970 44212 41982
rect 44156 41918 44158 41970
rect 44210 41918 44212 41970
rect 42364 41356 42868 41412
rect 41692 41132 42196 41188
rect 41580 41076 41636 41086
rect 41580 40982 41636 41020
rect 41468 40962 41524 40974
rect 41468 40910 41470 40962
rect 41522 40910 41524 40962
rect 41468 40628 41524 40910
rect 41692 40964 41748 40974
rect 41692 40870 41748 40908
rect 41916 40964 41972 40974
rect 41916 40962 42084 40964
rect 41916 40910 41918 40962
rect 41970 40910 42084 40962
rect 41916 40908 42084 40910
rect 41916 40898 41972 40908
rect 41916 40628 41972 40638
rect 41468 40572 41916 40628
rect 41468 40404 41524 40414
rect 41468 40310 41524 40348
rect 41916 40402 41972 40572
rect 41916 40350 41918 40402
rect 41970 40350 41972 40402
rect 41916 40338 41972 40350
rect 42028 39844 42084 40908
rect 42140 40514 42196 41132
rect 42588 41074 42644 41086
rect 42588 41022 42590 41074
rect 42642 41022 42644 41074
rect 42588 40964 42644 41022
rect 42588 40898 42644 40908
rect 42140 40462 42142 40514
rect 42194 40462 42196 40514
rect 42140 40404 42196 40462
rect 42812 40516 42868 41356
rect 42140 40338 42196 40348
rect 42700 40404 42756 40414
rect 42700 40310 42756 40348
rect 41356 39788 41524 39844
rect 42028 39788 42756 39844
rect 41356 39620 41412 39630
rect 41356 39526 41412 39564
rect 41468 39508 41524 39788
rect 41468 39442 41524 39452
rect 41692 39730 41748 39742
rect 41692 39678 41694 39730
rect 41746 39678 41748 39730
rect 41244 39228 41524 39284
rect 38892 38110 38894 38162
rect 38946 38110 38948 38162
rect 38892 38098 38948 38110
rect 40012 38612 40180 38668
rect 40348 38612 40404 38622
rect 39228 38052 39284 38090
rect 39228 37986 39284 37996
rect 38444 37202 38500 37212
rect 38332 36540 38500 36596
rect 38108 36430 38110 36482
rect 38162 36430 38164 36482
rect 38108 36418 38164 36430
rect 37548 35812 37604 35822
rect 37436 35810 38164 35812
rect 37436 35758 37550 35810
rect 37602 35758 38164 35810
rect 37436 35756 38164 35758
rect 34636 35646 34638 35698
rect 34690 35646 34692 35698
rect 34636 35634 34692 35646
rect 34972 35700 35028 35710
rect 34860 35588 34916 35598
rect 34860 35474 34916 35532
rect 34860 35422 34862 35474
rect 34914 35422 34916 35474
rect 34860 35364 34916 35422
rect 34860 35298 34916 35308
rect 34972 35476 35028 35644
rect 36764 35700 36820 35710
rect 36652 35588 36708 35598
rect 35084 35476 35140 35486
rect 34972 35474 35140 35476
rect 34972 35422 35086 35474
rect 35138 35422 35140 35474
rect 34972 35420 35140 35422
rect 34076 34862 34078 34914
rect 34130 34862 34132 34914
rect 34076 34850 34132 34862
rect 34412 34916 34468 34926
rect 34860 34916 34916 34926
rect 34412 34914 34916 34916
rect 34412 34862 34414 34914
rect 34466 34862 34862 34914
rect 34914 34862 34916 34914
rect 34412 34860 34916 34862
rect 34412 34850 34468 34860
rect 34860 34850 34916 34860
rect 34972 34914 35028 35420
rect 35084 35410 35140 35420
rect 35532 35476 35588 35486
rect 35532 35382 35588 35420
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34972 34862 34974 34914
rect 35026 34862 35028 34914
rect 33852 34802 33908 34814
rect 33852 34750 33854 34802
rect 33906 34750 33908 34802
rect 33852 34692 33908 34750
rect 33852 34626 33908 34636
rect 33964 34690 34020 34702
rect 33964 34638 33966 34690
rect 34018 34638 34020 34690
rect 33852 34244 33908 34254
rect 33964 34244 34020 34638
rect 33852 34242 34020 34244
rect 33852 34190 33854 34242
rect 33906 34190 34020 34242
rect 33852 34188 34020 34190
rect 34748 34692 34804 34702
rect 33852 34178 33908 34188
rect 34748 34020 34804 34636
rect 34748 33954 34804 33964
rect 33852 33460 33908 33470
rect 33852 33366 33908 33404
rect 34300 33124 34356 33134
rect 34300 33122 34468 33124
rect 34300 33070 34302 33122
rect 34354 33070 34468 33122
rect 34300 33068 34468 33070
rect 34300 33058 34356 33068
rect 34188 32788 34244 32798
rect 34188 32694 34244 32732
rect 33740 31892 33796 31902
rect 33740 30996 33796 31836
rect 34412 31892 34468 33068
rect 34972 32788 35028 34862
rect 35308 34916 35364 34926
rect 35308 34822 35364 34860
rect 36652 34916 36708 35532
rect 36764 35586 36820 35644
rect 36988 35698 37044 35756
rect 37548 35746 37604 35756
rect 36988 35646 36990 35698
rect 37042 35646 37044 35698
rect 36988 35634 37044 35646
rect 36764 35534 36766 35586
rect 36818 35534 36820 35586
rect 36764 35522 36820 35534
rect 38108 35586 38164 35756
rect 38444 35700 38500 36540
rect 38556 36484 38612 36494
rect 38780 36484 38836 37548
rect 39676 37492 39732 37502
rect 40012 37492 40068 38612
rect 40124 38162 40180 38174
rect 40124 38110 40126 38162
rect 40178 38110 40180 38162
rect 40124 38052 40180 38110
rect 40124 37986 40180 37996
rect 39732 37436 39956 37492
rect 40012 37436 40180 37492
rect 39676 37398 39732 37436
rect 38892 37268 38948 37278
rect 38892 37174 38948 37212
rect 39004 37156 39060 37166
rect 39452 37156 39508 37166
rect 39004 37154 39508 37156
rect 39004 37102 39006 37154
rect 39058 37102 39454 37154
rect 39506 37102 39508 37154
rect 39004 37100 39508 37102
rect 39004 37090 39060 37100
rect 39452 37090 39508 37100
rect 39788 37042 39844 37054
rect 39788 36990 39790 37042
rect 39842 36990 39844 37042
rect 38892 36820 38948 36830
rect 38892 36706 38948 36764
rect 38892 36654 38894 36706
rect 38946 36654 38948 36706
rect 38892 36642 38948 36654
rect 39788 36708 39844 36990
rect 39788 36642 39844 36652
rect 38556 36482 38836 36484
rect 38556 36430 38558 36482
rect 38610 36430 38836 36482
rect 38556 36428 38836 36430
rect 39676 36482 39732 36494
rect 39676 36430 39678 36482
rect 39730 36430 39732 36482
rect 38556 36418 38612 36428
rect 39004 36370 39060 36382
rect 39004 36318 39006 36370
rect 39058 36318 39060 36370
rect 38892 36260 38948 36270
rect 38892 36166 38948 36204
rect 39004 35924 39060 36318
rect 39676 35924 39732 36430
rect 38892 35868 39060 35924
rect 39564 35868 39732 35924
rect 39900 35924 39956 37436
rect 40012 37268 40068 37278
rect 40012 37174 40068 37212
rect 40124 36148 40180 37436
rect 40236 37378 40292 37390
rect 40236 37326 40238 37378
rect 40290 37326 40292 37378
rect 40236 36820 40292 37326
rect 40348 37378 40404 38556
rect 40348 37326 40350 37378
rect 40402 37326 40404 37378
rect 40348 37314 40404 37326
rect 40908 38612 41076 38668
rect 41468 39060 41524 39228
rect 40236 36754 40292 36764
rect 40460 36708 40516 36718
rect 40460 36594 40516 36652
rect 40460 36542 40462 36594
rect 40514 36542 40516 36594
rect 40460 36530 40516 36542
rect 40124 36092 40292 36148
rect 40124 35924 40180 35934
rect 39900 35922 40180 35924
rect 39900 35870 40126 35922
rect 40178 35870 40180 35922
rect 39900 35868 40180 35870
rect 38556 35700 38612 35710
rect 38444 35698 38612 35700
rect 38444 35646 38558 35698
rect 38610 35646 38612 35698
rect 38444 35644 38612 35646
rect 38108 35534 38110 35586
rect 38162 35534 38164 35586
rect 38108 35522 38164 35534
rect 37548 35026 37604 35038
rect 37548 34974 37550 35026
rect 37602 34974 37604 35026
rect 36652 34354 36708 34860
rect 37212 34916 37268 34926
rect 37212 34822 37268 34860
rect 36652 34302 36654 34354
rect 36706 34302 36708 34354
rect 36652 34290 36708 34302
rect 36988 34804 37044 34814
rect 36764 34132 36820 34142
rect 36764 34038 36820 34076
rect 35980 34020 36036 34030
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35084 33460 35140 33470
rect 35084 33236 35140 33404
rect 35532 33348 35588 33358
rect 35532 33254 35588 33292
rect 35980 33348 36036 33964
rect 36652 34020 36708 34030
rect 36652 33906 36708 33964
rect 36652 33854 36654 33906
rect 36706 33854 36708 33906
rect 36652 33842 36708 33854
rect 35980 33282 36036 33292
rect 35084 33234 35364 33236
rect 35084 33182 35086 33234
rect 35138 33182 35364 33234
rect 35084 33180 35364 33182
rect 35084 33170 35140 33180
rect 35084 32788 35140 32798
rect 34972 32786 35140 32788
rect 34972 32734 35086 32786
rect 35138 32734 35140 32786
rect 34972 32732 35140 32734
rect 35084 32722 35140 32732
rect 35308 32562 35364 33180
rect 35644 33234 35700 33246
rect 35644 33182 35646 33234
rect 35698 33182 35700 33234
rect 35420 32900 35476 32910
rect 35476 32844 35588 32900
rect 35420 32834 35476 32844
rect 35308 32510 35310 32562
rect 35362 32510 35364 32562
rect 35308 32498 35364 32510
rect 34748 32450 34804 32462
rect 34748 32398 34750 32450
rect 34802 32398 34804 32450
rect 34748 32004 34804 32398
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34748 31938 34804 31948
rect 34412 31826 34468 31836
rect 34188 31778 34244 31790
rect 34188 31726 34190 31778
rect 34242 31726 34244 31778
rect 33852 31668 33908 31678
rect 33852 31574 33908 31612
rect 33740 30902 33796 30940
rect 34188 30436 34244 31726
rect 34300 31780 34356 31818
rect 34300 31714 34356 31724
rect 34524 31778 34580 31790
rect 34524 31726 34526 31778
rect 34578 31726 34580 31778
rect 34300 31554 34356 31566
rect 34300 31502 34302 31554
rect 34354 31502 34356 31554
rect 34300 31108 34356 31502
rect 34524 31556 34580 31726
rect 34524 31490 34580 31500
rect 34748 31666 34804 31678
rect 34748 31614 34750 31666
rect 34802 31614 34804 31666
rect 34412 31108 34468 31118
rect 34300 31106 34468 31108
rect 34300 31054 34414 31106
rect 34466 31054 34468 31106
rect 34300 31052 34468 31054
rect 34412 31042 34468 31052
rect 34748 30548 34804 31614
rect 35532 31668 35588 32844
rect 35644 32676 35700 33182
rect 35644 32610 35700 32620
rect 36204 33122 36260 33134
rect 36204 33070 36206 33122
rect 36258 33070 36260 33122
rect 35196 31556 35252 31566
rect 35196 30884 35252 31500
rect 35196 30818 35252 30828
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 34748 30492 35140 30548
rect 35196 30538 35460 30548
rect 34188 30380 34916 30436
rect 33628 30210 33908 30212
rect 33628 30158 33630 30210
rect 33682 30158 33908 30210
rect 33628 30156 33908 30158
rect 33628 30146 33684 30156
rect 33852 30100 33908 30156
rect 33628 29988 33684 29998
rect 33628 29428 33684 29932
rect 33516 29316 33572 29326
rect 33516 29222 33572 29260
rect 33404 28814 33406 28866
rect 33458 28814 33460 28866
rect 33404 28756 33460 28814
rect 32620 28644 32676 28654
rect 32956 28644 33012 28654
rect 33180 28644 33236 28654
rect 32620 28642 33012 28644
rect 32620 28590 32622 28642
rect 32674 28590 32958 28642
rect 33010 28590 33012 28642
rect 32620 28588 33012 28590
rect 32620 28578 32676 28588
rect 32508 28530 32564 28542
rect 32508 28478 32510 28530
rect 32562 28478 32564 28530
rect 32396 27748 32452 27758
rect 32508 27748 32564 28478
rect 32844 28420 32900 28430
rect 32844 28326 32900 28364
rect 32956 27860 33012 28588
rect 32956 27794 33012 27804
rect 33068 28642 33236 28644
rect 33068 28590 33182 28642
rect 33234 28590 33236 28642
rect 33068 28588 33236 28590
rect 32396 27746 32564 27748
rect 32396 27694 32398 27746
rect 32450 27694 32564 27746
rect 32396 27692 32564 27694
rect 32396 27076 32452 27692
rect 32396 27010 32452 27020
rect 33068 27188 33124 28588
rect 33180 28578 33236 28588
rect 33404 28084 33460 28700
rect 32844 26852 32900 26862
rect 32508 26796 32844 26852
rect 32508 26514 32564 26796
rect 32844 26786 32900 26796
rect 32508 26462 32510 26514
rect 32562 26462 32564 26514
rect 32508 26450 32564 26462
rect 32956 26740 33012 26750
rect 32844 25620 32900 25630
rect 32956 25620 33012 26684
rect 33068 26516 33124 27132
rect 33180 28028 33460 28084
rect 33516 28868 33572 28878
rect 33180 26908 33236 28028
rect 33404 27860 33460 27870
rect 33404 27766 33460 27804
rect 33292 27746 33348 27758
rect 33292 27694 33294 27746
rect 33346 27694 33348 27746
rect 33292 27636 33348 27694
rect 33516 27636 33572 28812
rect 33292 27580 33572 27636
rect 33516 27186 33572 27580
rect 33516 27134 33518 27186
rect 33570 27134 33572 27186
rect 33516 27122 33572 27134
rect 33628 28642 33684 29372
rect 33628 28590 33630 28642
rect 33682 28590 33684 28642
rect 33404 27076 33460 27086
rect 33404 26982 33460 27020
rect 33180 26852 33572 26908
rect 33180 26786 33236 26796
rect 33068 26460 33348 26516
rect 33068 26292 33124 26302
rect 33068 26198 33124 26236
rect 33292 26290 33348 26460
rect 33292 26238 33294 26290
rect 33346 26238 33348 26290
rect 33292 26226 33348 26238
rect 33516 26290 33572 26852
rect 33516 26238 33518 26290
rect 33570 26238 33572 26290
rect 33516 26226 33572 26238
rect 33180 26180 33236 26190
rect 33180 26086 33236 26124
rect 32844 25618 33012 25620
rect 32844 25566 32846 25618
rect 32898 25566 33012 25618
rect 32844 25564 33012 25566
rect 33516 25956 33572 25966
rect 32844 25554 32900 25564
rect 33180 24052 33236 24062
rect 33180 23958 33236 23996
rect 33516 23380 33572 25900
rect 33628 25618 33684 28590
rect 33852 27748 33908 30044
rect 34860 29650 34916 30380
rect 34860 29598 34862 29650
rect 34914 29598 34916 29650
rect 34860 29586 34916 29598
rect 34972 30324 35028 30334
rect 34188 29428 34244 29438
rect 34188 29334 34244 29372
rect 34636 29428 34692 29438
rect 34412 29316 34468 29326
rect 34412 29314 34580 29316
rect 34412 29262 34414 29314
rect 34466 29262 34580 29314
rect 34412 29260 34580 29262
rect 34412 29250 34468 29260
rect 33964 28644 34020 28654
rect 33964 28642 34468 28644
rect 33964 28590 33966 28642
rect 34018 28590 34468 28642
rect 33964 28588 34468 28590
rect 33964 28578 34020 28588
rect 34412 28084 34468 28588
rect 34524 28642 34580 29260
rect 34524 28590 34526 28642
rect 34578 28590 34580 28642
rect 34524 28196 34580 28590
rect 34636 28418 34692 29372
rect 34860 28644 34916 28654
rect 34972 28644 35028 30268
rect 35084 29428 35140 30492
rect 35420 29988 35476 29998
rect 35420 29538 35476 29932
rect 35420 29486 35422 29538
rect 35474 29486 35476 29538
rect 35420 29474 35476 29486
rect 35084 29362 35140 29372
rect 35196 29316 35252 29326
rect 35196 29222 35252 29260
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 28868 35252 28878
rect 35196 28774 35252 28812
rect 34860 28642 35028 28644
rect 34860 28590 34862 28642
rect 34914 28590 35028 28642
rect 34860 28588 35028 28590
rect 34860 28578 34916 28588
rect 35308 28530 35364 28542
rect 35308 28478 35310 28530
rect 35362 28478 35364 28530
rect 34636 28366 34638 28418
rect 34690 28366 34692 28418
rect 34636 28354 34692 28366
rect 35196 28418 35252 28430
rect 35196 28366 35198 28418
rect 35250 28366 35252 28418
rect 34524 28140 34692 28196
rect 34412 28028 34580 28084
rect 34524 27970 34580 28028
rect 34524 27918 34526 27970
rect 34578 27918 34580 27970
rect 34524 27906 34580 27918
rect 34076 27860 34132 27870
rect 34300 27860 34356 27870
rect 34076 27858 34356 27860
rect 34076 27806 34078 27858
rect 34130 27806 34302 27858
rect 34354 27806 34356 27858
rect 34076 27804 34356 27806
rect 34076 27794 34132 27804
rect 34300 27794 34356 27804
rect 34412 27860 34468 27870
rect 33740 27692 33908 27748
rect 33740 26516 33796 27692
rect 34412 27636 34468 27804
rect 34188 27580 34468 27636
rect 34188 27076 34244 27580
rect 34524 27300 34580 27310
rect 34636 27300 34692 28140
rect 34860 28084 34916 28094
rect 34524 27298 34692 27300
rect 34524 27246 34526 27298
rect 34578 27246 34692 27298
rect 34524 27244 34692 27246
rect 34748 27858 34804 27870
rect 34748 27806 34750 27858
rect 34802 27806 34804 27858
rect 34524 27234 34580 27244
rect 34412 27076 34468 27086
rect 33852 26962 33908 26974
rect 33852 26910 33854 26962
rect 33906 26910 33908 26962
rect 33852 26908 33908 26910
rect 34188 26962 34244 27020
rect 34188 26910 34190 26962
rect 34242 26910 34244 26962
rect 33852 26852 34132 26908
rect 34188 26898 34244 26910
rect 34300 27074 34468 27076
rect 34300 27022 34414 27074
rect 34466 27022 34468 27074
rect 34300 27020 34468 27022
rect 34300 26964 34356 27020
rect 34412 27010 34468 27020
rect 34636 27076 34692 27086
rect 34636 26908 34692 27020
rect 34300 26898 34356 26908
rect 33740 26460 33908 26516
rect 33740 26292 33796 26302
rect 33740 26198 33796 26236
rect 33628 25566 33630 25618
rect 33682 25566 33684 25618
rect 33628 25554 33684 25566
rect 33852 24612 33908 26460
rect 33964 26290 34020 26302
rect 33964 26238 33966 26290
rect 34018 26238 34020 26290
rect 33964 26180 34020 26238
rect 33964 26114 34020 26124
rect 33964 25396 34020 25406
rect 34076 25396 34132 26852
rect 34412 26852 34692 26908
rect 34748 26908 34804 27806
rect 34860 27858 34916 28028
rect 34860 27806 34862 27858
rect 34914 27806 34916 27858
rect 34860 27794 34916 27806
rect 35196 27860 35252 28366
rect 35196 27794 35252 27804
rect 35308 27636 35364 28478
rect 35532 27858 35588 31612
rect 36204 31892 36260 33070
rect 36988 32900 37044 34748
rect 37100 34130 37156 34142
rect 37100 34078 37102 34130
rect 37154 34078 37156 34130
rect 37100 34020 37156 34078
rect 37548 34132 37604 34974
rect 38444 34692 38500 34702
rect 37548 34066 37604 34076
rect 38220 34690 38500 34692
rect 38220 34638 38446 34690
rect 38498 34638 38500 34690
rect 38220 34636 38500 34638
rect 38220 34132 38276 34636
rect 38444 34626 38500 34636
rect 38220 34130 38388 34132
rect 38220 34078 38222 34130
rect 38274 34078 38388 34130
rect 38220 34076 38388 34078
rect 38220 34066 38276 34076
rect 37100 33954 37156 33964
rect 37436 33346 37492 33358
rect 37436 33294 37438 33346
rect 37490 33294 37492 33346
rect 36988 32786 37044 32844
rect 36988 32734 36990 32786
rect 37042 32734 37044 32786
rect 36988 32722 37044 32734
rect 37100 33124 37156 33134
rect 37436 33124 37492 33294
rect 38220 33236 38276 33246
rect 37100 33122 37492 33124
rect 37100 33070 37102 33122
rect 37154 33070 37492 33122
rect 37100 33068 37492 33070
rect 37660 33234 38276 33236
rect 37660 33182 38222 33234
rect 38274 33182 38276 33234
rect 37660 33180 38276 33182
rect 37100 31892 37156 33068
rect 37660 32786 37716 33180
rect 38220 33170 38276 33180
rect 38108 32788 38164 32798
rect 38332 32788 38388 34076
rect 38556 33906 38612 35644
rect 38892 35700 38948 35868
rect 38892 35634 38948 35644
rect 39004 35700 39060 35710
rect 39340 35700 39396 35710
rect 39004 35698 39396 35700
rect 39004 35646 39006 35698
rect 39058 35646 39342 35698
rect 39394 35646 39396 35698
rect 39004 35644 39396 35646
rect 39004 35634 39060 35644
rect 39340 35634 39396 35644
rect 39340 34916 39396 34926
rect 39564 34916 39620 35868
rect 39676 35700 39732 35710
rect 39900 35700 39956 35868
rect 40124 35858 40180 35868
rect 40236 35700 40292 36092
rect 39676 35698 39956 35700
rect 39676 35646 39678 35698
rect 39730 35646 39956 35698
rect 39676 35644 39956 35646
rect 40124 35644 40292 35700
rect 39676 35634 39732 35644
rect 39676 35476 39732 35486
rect 39676 35474 40068 35476
rect 39676 35422 39678 35474
rect 39730 35422 40068 35474
rect 39676 35420 40068 35422
rect 39676 35410 39732 35420
rect 40012 35026 40068 35420
rect 40012 34974 40014 35026
rect 40066 34974 40068 35026
rect 40012 34962 40068 34974
rect 39340 34914 39620 34916
rect 39340 34862 39342 34914
rect 39394 34862 39620 34914
rect 39340 34860 39620 34862
rect 39340 34850 39396 34860
rect 39564 34692 39620 34860
rect 39564 34626 39620 34636
rect 38556 33854 38558 33906
rect 38610 33854 38612 33906
rect 38556 33842 38612 33854
rect 39340 34130 39396 34142
rect 39340 34078 39342 34130
rect 39394 34078 39396 34130
rect 37660 32734 37662 32786
rect 37714 32734 37716 32786
rect 37660 32722 37716 32734
rect 37884 32786 38388 32788
rect 37884 32734 38110 32786
rect 38162 32734 38388 32786
rect 37884 32732 38388 32734
rect 38556 33572 38612 33582
rect 38556 32900 38612 33516
rect 38556 32786 38612 32844
rect 38556 32734 38558 32786
rect 38610 32734 38612 32786
rect 37436 32676 37492 32686
rect 37436 32582 37492 32620
rect 37324 32562 37380 32574
rect 37324 32510 37326 32562
rect 37378 32510 37380 32562
rect 37324 32340 37380 32510
rect 37884 32562 37940 32732
rect 38108 32722 38164 32732
rect 38556 32722 38612 32734
rect 38444 32676 38500 32686
rect 37884 32510 37886 32562
rect 37938 32510 37940 32562
rect 37884 32498 37940 32510
rect 38332 32564 38388 32574
rect 38444 32564 38500 32620
rect 38332 32562 38500 32564
rect 38332 32510 38334 32562
rect 38386 32510 38500 32562
rect 38332 32508 38500 32510
rect 39340 32564 39396 34078
rect 38332 32498 38388 32508
rect 39340 32498 39396 32508
rect 38220 32450 38276 32462
rect 38220 32398 38222 32450
rect 38274 32398 38276 32450
rect 38220 32340 38276 32398
rect 37324 32284 38276 32340
rect 35980 31556 36036 31566
rect 36204 31556 36260 31836
rect 36988 31836 37156 31892
rect 37548 32002 37604 32014
rect 37548 31950 37550 32002
rect 37602 31950 37604 32002
rect 37548 31892 37604 31950
rect 36036 31500 36260 31556
rect 36428 31556 36484 31566
rect 35980 31462 36036 31500
rect 36428 31444 36484 31500
rect 36428 31388 36708 31444
rect 36652 30996 36708 31388
rect 36876 30996 36932 31006
rect 36988 30996 37044 31836
rect 37548 31826 37604 31836
rect 38108 31892 38164 31902
rect 37436 31778 37492 31790
rect 37436 31726 37438 31778
rect 37490 31726 37492 31778
rect 36652 30994 37044 30996
rect 36652 30942 36878 30994
rect 36930 30942 37044 30994
rect 36652 30940 37044 30942
rect 37100 31666 37156 31678
rect 37100 31614 37102 31666
rect 37154 31614 37156 31666
rect 36540 30882 36596 30894
rect 36540 30830 36542 30882
rect 36594 30830 36596 30882
rect 36092 30436 36148 30446
rect 36092 30342 36148 30380
rect 35756 30324 35812 30334
rect 35756 30230 35812 30268
rect 36540 30212 36596 30830
rect 36540 30146 36596 30156
rect 35980 29988 36036 29998
rect 35980 29894 36036 29932
rect 36092 28756 36148 28766
rect 36316 28756 36372 28766
rect 36148 28700 36260 28756
rect 36092 28690 36148 28700
rect 35980 28644 36036 28654
rect 35756 28420 35812 28430
rect 35756 28418 35924 28420
rect 35756 28366 35758 28418
rect 35810 28366 35924 28418
rect 35756 28364 35924 28366
rect 35756 28354 35812 28364
rect 35532 27806 35534 27858
rect 35586 27806 35588 27858
rect 35532 27794 35588 27806
rect 35644 28084 35700 28094
rect 35084 27580 35364 27636
rect 34860 27188 34916 27198
rect 34916 27132 35028 27188
rect 34860 27122 34916 27132
rect 34972 26908 35028 27132
rect 35084 27076 35140 27580
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35084 27010 35140 27020
rect 35196 27300 35252 27310
rect 35196 26964 35252 27244
rect 35644 27076 35700 28028
rect 35644 27010 35700 27020
rect 35756 27634 35812 27646
rect 35756 27582 35758 27634
rect 35810 27582 35812 27634
rect 34748 26852 34916 26908
rect 34972 26852 35140 26908
rect 34300 26404 34356 26414
rect 33964 25394 34132 25396
rect 33964 25342 33966 25394
rect 34018 25342 34132 25394
rect 33964 25340 34132 25342
rect 34188 26290 34244 26302
rect 34188 26238 34190 26290
rect 34242 26238 34244 26290
rect 34188 25506 34244 26238
rect 34188 25454 34190 25506
rect 34242 25454 34244 25506
rect 33964 25330 34020 25340
rect 34076 25172 34132 25182
rect 33964 24612 34020 24622
rect 33852 24556 33964 24612
rect 33964 24518 34020 24556
rect 33852 24052 33908 24062
rect 33628 23380 33684 23390
rect 33516 23324 33628 23380
rect 33628 23286 33684 23324
rect 33852 23266 33908 23996
rect 34076 23380 34132 25116
rect 34188 24052 34244 25454
rect 34188 23986 34244 23996
rect 34300 23938 34356 26348
rect 34300 23886 34302 23938
rect 34354 23886 34356 23938
rect 34300 23874 34356 23886
rect 34412 23940 34468 26852
rect 34860 26514 34916 26852
rect 35084 26850 35140 26852
rect 35084 26798 35086 26850
rect 35138 26798 35140 26850
rect 35084 26786 35140 26798
rect 34860 26462 34862 26514
rect 34914 26462 34916 26514
rect 34748 26402 34804 26414
rect 34748 26350 34750 26402
rect 34802 26350 34804 26402
rect 34524 26290 34580 26302
rect 34524 26238 34526 26290
rect 34578 26238 34580 26290
rect 34524 25620 34580 26238
rect 34524 24164 34580 25564
rect 34748 25396 34804 26350
rect 34860 26292 34916 26462
rect 35084 26404 35140 26414
rect 35084 26310 35140 26348
rect 35196 26402 35252 26908
rect 35196 26350 35198 26402
rect 35250 26350 35252 26402
rect 35196 26338 35252 26350
rect 35532 26852 35588 26862
rect 35532 26292 35588 26796
rect 35756 26740 35812 27582
rect 35756 26674 35812 26684
rect 35868 27188 35924 28364
rect 35868 26962 35924 27132
rect 35868 26910 35870 26962
rect 35922 26910 35924 26962
rect 35756 26292 35812 26302
rect 35532 26290 35812 26292
rect 35532 26238 35758 26290
rect 35810 26238 35812 26290
rect 35532 26236 35812 26238
rect 34860 26226 34916 26236
rect 34972 26180 35028 26190
rect 35028 26124 35140 26180
rect 34972 26114 35028 26124
rect 34860 25396 34916 25406
rect 34748 25394 34916 25396
rect 34748 25342 34862 25394
rect 34914 25342 34916 25394
rect 34748 25340 34916 25342
rect 34860 25284 34916 25340
rect 34860 25218 34916 25228
rect 34860 24612 34916 24622
rect 34524 24108 34804 24164
rect 34636 23940 34692 23950
rect 34412 23938 34692 23940
rect 34412 23886 34638 23938
rect 34690 23886 34692 23938
rect 34412 23884 34692 23886
rect 34636 23716 34692 23884
rect 34636 23650 34692 23660
rect 34748 23492 34804 24108
rect 34524 23436 34804 23492
rect 34076 23324 34244 23380
rect 33852 23214 33854 23266
rect 33906 23214 33908 23266
rect 33852 23202 33908 23214
rect 34076 23156 34132 23166
rect 32172 22866 32228 22876
rect 33964 23154 34132 23156
rect 33964 23102 34078 23154
rect 34130 23102 34132 23154
rect 33964 23100 34132 23102
rect 31164 22370 31444 22372
rect 31164 22318 31166 22370
rect 31218 22318 31444 22370
rect 31164 22316 31444 22318
rect 29148 21868 29540 21924
rect 29372 20804 29428 20814
rect 29260 20802 29428 20804
rect 29260 20750 29374 20802
rect 29426 20750 29428 20802
rect 29260 20748 29428 20750
rect 29148 20578 29204 20590
rect 29148 20526 29150 20578
rect 29202 20526 29204 20578
rect 29148 20130 29204 20526
rect 29148 20078 29150 20130
rect 29202 20078 29204 20130
rect 29148 20066 29204 20078
rect 29260 19458 29316 20748
rect 29372 20738 29428 20748
rect 29260 19406 29262 19458
rect 29314 19406 29316 19458
rect 29260 19394 29316 19406
rect 29484 18900 29540 21868
rect 29596 21868 30100 21924
rect 29596 21586 29652 21868
rect 30044 21812 30100 21868
rect 30380 22258 30436 22270
rect 30380 22206 30382 22258
rect 30434 22206 30436 22258
rect 30268 21812 30324 21822
rect 30044 21810 30324 21812
rect 30044 21758 30270 21810
rect 30322 21758 30324 21810
rect 30044 21756 30324 21758
rect 30268 21746 30324 21756
rect 29596 21534 29598 21586
rect 29650 21534 29652 21586
rect 29596 21522 29652 21534
rect 29820 21698 29876 21710
rect 29820 21646 29822 21698
rect 29874 21646 29876 21698
rect 29820 21588 29876 21646
rect 30380 21588 30436 22206
rect 29820 21532 30436 21588
rect 29596 19908 29652 19918
rect 29596 19460 29652 19852
rect 29596 19458 29988 19460
rect 29596 19406 29598 19458
rect 29650 19406 29988 19458
rect 29596 19404 29988 19406
rect 29596 19394 29652 19404
rect 29820 19124 29876 19134
rect 29820 19030 29876 19068
rect 29484 18844 29876 18900
rect 29372 18564 29428 18574
rect 29148 17668 29204 17678
rect 29148 17574 29204 17612
rect 29372 17666 29428 18508
rect 29708 18562 29764 18574
rect 29708 18510 29710 18562
rect 29762 18510 29764 18562
rect 29708 18452 29764 18510
rect 29708 18386 29764 18396
rect 29596 18228 29652 18238
rect 29372 17614 29374 17666
rect 29426 17614 29428 17666
rect 29260 17442 29316 17454
rect 29260 17390 29262 17442
rect 29314 17390 29316 17442
rect 29260 16324 29316 17390
rect 29260 16258 29316 16268
rect 29148 16100 29204 16138
rect 29148 16034 29204 16044
rect 29148 15874 29204 15886
rect 29148 15822 29150 15874
rect 29202 15822 29204 15874
rect 29148 15764 29204 15822
rect 29148 15698 29204 15708
rect 29372 15764 29428 17614
rect 29484 18226 29652 18228
rect 29484 18174 29598 18226
rect 29650 18174 29652 18226
rect 29484 18172 29652 18174
rect 29484 16322 29540 18172
rect 29596 18162 29652 18172
rect 29596 17892 29652 17902
rect 29596 17798 29652 17836
rect 29708 17666 29764 17678
rect 29708 17614 29710 17666
rect 29762 17614 29764 17666
rect 29484 16270 29486 16322
rect 29538 16270 29540 16322
rect 29484 16258 29540 16270
rect 29596 16770 29652 16782
rect 29596 16718 29598 16770
rect 29650 16718 29652 16770
rect 29596 15988 29652 16718
rect 29708 16212 29764 17614
rect 29708 16146 29764 16156
rect 29596 15922 29652 15932
rect 29708 15986 29764 15998
rect 29708 15934 29710 15986
rect 29762 15934 29764 15986
rect 29708 15764 29764 15934
rect 29372 15708 29764 15764
rect 29036 15428 29092 15438
rect 29036 15334 29092 15372
rect 29372 15148 29428 15708
rect 29260 15092 29428 15148
rect 29484 15204 29540 15214
rect 29148 13972 29204 13982
rect 28700 13970 29204 13972
rect 28700 13918 28814 13970
rect 28866 13918 29150 13970
rect 29202 13918 29204 13970
rect 28700 13916 29204 13918
rect 27468 13694 27470 13746
rect 27522 13694 27524 13746
rect 27468 13682 27524 13694
rect 27804 13748 27860 13758
rect 27804 13654 27860 13692
rect 27020 13524 27076 13534
rect 27020 13186 27076 13468
rect 27356 13524 27412 13534
rect 27356 13522 27524 13524
rect 27356 13470 27358 13522
rect 27410 13470 27524 13522
rect 27356 13468 27524 13470
rect 27356 13458 27412 13468
rect 27020 13134 27022 13186
rect 27074 13134 27076 13186
rect 27020 13122 27076 13134
rect 26348 12908 26628 12964
rect 26236 12562 26292 12572
rect 26124 12126 26126 12178
rect 26178 12126 26180 12178
rect 26124 11506 26180 12126
rect 26236 12404 26292 12414
rect 26236 12180 26292 12348
rect 26348 12180 26404 12190
rect 26236 12178 26404 12180
rect 26236 12126 26350 12178
rect 26402 12126 26404 12178
rect 26236 12124 26404 12126
rect 26348 12114 26404 12124
rect 26124 11454 26126 11506
rect 26178 11454 26180 11506
rect 26124 11442 26180 11454
rect 26236 11508 26292 11518
rect 26236 11396 26292 11452
rect 26236 11394 26516 11396
rect 26236 11342 26238 11394
rect 26290 11342 26516 11394
rect 26236 11340 26516 11342
rect 26236 11330 26292 11340
rect 26012 10780 26404 10836
rect 26012 10612 26068 10622
rect 25900 10610 26068 10612
rect 25900 10558 26014 10610
rect 26066 10558 26068 10610
rect 25900 10556 26068 10558
rect 26012 10546 26068 10556
rect 25564 8530 25620 8540
rect 25676 8988 25844 9044
rect 25452 8094 25454 8146
rect 25506 8094 25508 8146
rect 25452 8082 25508 8094
rect 25676 7700 25732 8988
rect 25788 8818 25844 8830
rect 25788 8766 25790 8818
rect 25842 8766 25844 8818
rect 25788 8258 25844 8766
rect 26124 8818 26180 8830
rect 26124 8766 26126 8818
rect 26178 8766 26180 8818
rect 25788 8206 25790 8258
rect 25842 8206 25844 8258
rect 25788 8194 25844 8206
rect 26012 8596 26068 8606
rect 26124 8596 26180 8766
rect 26068 8540 26180 8596
rect 25676 7634 25732 7644
rect 25340 7586 25396 7598
rect 25340 7534 25342 7586
rect 25394 7534 25396 7586
rect 25340 6802 25396 7534
rect 25340 6750 25342 6802
rect 25394 6750 25396 6802
rect 25340 6738 25396 6750
rect 25676 7474 25732 7486
rect 25676 7422 25678 7474
rect 25730 7422 25732 7474
rect 25676 6130 25732 7422
rect 25676 6078 25678 6130
rect 25730 6078 25732 6130
rect 25676 6066 25732 6078
rect 23884 6018 25060 6020
rect 23884 5966 23886 6018
rect 23938 5966 25060 6018
rect 23884 5964 25060 5966
rect 23884 5954 23940 5964
rect 23772 5236 23828 5246
rect 23772 4562 23828 5180
rect 24892 5236 24948 5246
rect 25004 5236 25060 5964
rect 26012 5906 26068 8540
rect 26348 7698 26404 10780
rect 26460 10610 26516 11340
rect 26572 10836 26628 12908
rect 26684 12962 26852 12964
rect 26684 12910 26686 12962
rect 26738 12910 26852 12962
rect 26684 12908 26852 12910
rect 27356 12964 27412 12974
rect 26684 12898 26740 12908
rect 27356 12870 27412 12908
rect 27132 12852 27188 12862
rect 27132 12758 27188 12796
rect 27468 12404 27524 13468
rect 28364 12962 28420 12974
rect 28364 12910 28366 12962
rect 28418 12910 28420 12962
rect 28364 12516 28420 12910
rect 28588 12852 28644 12862
rect 28588 12758 28644 12796
rect 28364 12450 28420 12460
rect 27468 12338 27524 12348
rect 28252 12404 28308 12442
rect 28252 12338 28308 12348
rect 28252 12180 28308 12190
rect 28252 12086 28308 12124
rect 26908 12066 26964 12078
rect 26908 12014 26910 12066
rect 26962 12014 26964 12066
rect 26908 11396 26964 12014
rect 28476 11954 28532 11966
rect 28476 11902 28478 11954
rect 28530 11902 28532 11954
rect 28476 11732 28532 11902
rect 28476 11666 28532 11676
rect 26908 11330 26964 11340
rect 26796 11284 26852 11294
rect 26572 10770 26628 10780
rect 26684 11282 26852 11284
rect 26684 11230 26798 11282
rect 26850 11230 26852 11282
rect 26684 11228 26852 11230
rect 26460 10558 26462 10610
rect 26514 10558 26516 10610
rect 26460 10546 26516 10558
rect 26348 7646 26350 7698
rect 26402 7646 26404 7698
rect 26348 7634 26404 7646
rect 26684 7588 26740 11228
rect 26796 11218 26852 11228
rect 28700 11284 28756 13916
rect 28812 13906 28868 13916
rect 29148 13906 29204 13916
rect 29260 13748 29316 15092
rect 29484 13970 29540 15148
rect 29484 13918 29486 13970
rect 29538 13918 29540 13970
rect 29484 13906 29540 13918
rect 28812 13692 29316 13748
rect 28812 12290 28868 13692
rect 28812 12238 28814 12290
rect 28866 12238 28868 12290
rect 28812 12226 28868 12238
rect 29148 13074 29204 13086
rect 29148 13022 29150 13074
rect 29202 13022 29204 13074
rect 29148 12964 29204 13022
rect 29148 12292 29204 12908
rect 29596 12516 29652 12526
rect 29596 12402 29652 12460
rect 29596 12350 29598 12402
rect 29650 12350 29652 12402
rect 29596 12338 29652 12350
rect 29148 12226 29204 12236
rect 28700 11218 28756 11228
rect 29036 12178 29092 12190
rect 29036 12126 29038 12178
rect 29090 12126 29092 12178
rect 27132 10836 27188 10846
rect 27132 10742 27188 10780
rect 26796 10724 26852 10734
rect 26796 9042 26852 10668
rect 28588 10724 28644 10734
rect 28588 10630 28644 10668
rect 28924 10722 28980 10734
rect 28924 10670 28926 10722
rect 28978 10670 28980 10722
rect 27244 10498 27300 10510
rect 27244 10446 27246 10498
rect 27298 10446 27300 10498
rect 26908 9940 26964 9950
rect 26908 9154 26964 9884
rect 27244 9940 27300 10446
rect 27916 10388 27972 10398
rect 27916 10386 28084 10388
rect 27916 10334 27918 10386
rect 27970 10334 28084 10386
rect 27916 10332 28084 10334
rect 27916 10322 27972 10332
rect 27244 9874 27300 9884
rect 27580 9940 27636 9950
rect 27580 9846 27636 9884
rect 28028 9826 28084 10332
rect 28028 9774 28030 9826
rect 28082 9774 28084 9826
rect 28028 9762 28084 9774
rect 28252 10386 28308 10398
rect 28252 10334 28254 10386
rect 28306 10334 28308 10386
rect 26908 9102 26910 9154
rect 26962 9102 26964 9154
rect 26908 9090 26964 9102
rect 28252 9604 28308 10334
rect 28924 9940 28980 10670
rect 28924 9874 28980 9884
rect 26796 8990 26798 9042
rect 26850 8990 26852 9042
rect 26796 8978 26852 8990
rect 27804 9042 27860 9054
rect 27804 8990 27806 9042
rect 27858 8990 27860 9042
rect 27356 8260 27412 8270
rect 27356 8036 27412 8204
rect 27804 8036 27860 8990
rect 26460 7364 26516 7374
rect 26460 7362 26628 7364
rect 26460 7310 26462 7362
rect 26514 7310 26628 7362
rect 26460 7308 26628 7310
rect 26460 7298 26516 7308
rect 26572 6916 26628 7308
rect 26572 6018 26628 6860
rect 26572 5966 26574 6018
rect 26626 5966 26628 6018
rect 26572 5954 26628 5966
rect 26012 5854 26014 5906
rect 26066 5854 26068 5906
rect 26012 5842 26068 5854
rect 26684 5906 26740 7532
rect 26684 5854 26686 5906
rect 26738 5854 26740 5906
rect 26684 5842 26740 5854
rect 27244 8034 27860 8036
rect 27244 7982 27358 8034
rect 27410 7982 27806 8034
rect 27858 7982 27860 8034
rect 27244 7980 27860 7982
rect 27244 6804 27300 7980
rect 27356 7970 27412 7980
rect 27804 7970 27860 7980
rect 27916 8708 27972 8718
rect 28252 8708 28308 9548
rect 28364 9604 28420 9614
rect 28364 9602 28532 9604
rect 28364 9550 28366 9602
rect 28418 9550 28532 9602
rect 28364 9548 28532 9550
rect 28364 9538 28420 9548
rect 28476 9154 28532 9548
rect 28476 9102 28478 9154
rect 28530 9102 28532 9154
rect 28476 9090 28532 9102
rect 27972 8652 28308 8708
rect 27916 7474 27972 8652
rect 29036 8428 29092 12126
rect 29260 11508 29316 11518
rect 29708 11508 29764 11518
rect 29820 11508 29876 18844
rect 29932 18562 29988 19404
rect 30380 19124 30436 21532
rect 30380 19030 30436 19068
rect 30828 21476 30884 21486
rect 31164 21476 31220 22316
rect 31948 22258 32004 22270
rect 31948 22206 31950 22258
rect 32002 22206 32004 22258
rect 31948 21812 32004 22206
rect 33964 22148 34020 23100
rect 34076 23090 34132 23100
rect 33964 22082 34020 22092
rect 34076 22482 34132 22494
rect 34076 22430 34078 22482
rect 34130 22430 34132 22482
rect 34076 21924 34132 22430
rect 34188 22372 34244 23324
rect 34524 23154 34580 23436
rect 34524 23102 34526 23154
rect 34578 23102 34580 23154
rect 34524 23090 34580 23102
rect 34300 23042 34356 23054
rect 34300 22990 34302 23042
rect 34354 22990 34356 23042
rect 34300 22932 34356 22990
rect 34748 22932 34804 22942
rect 34300 22930 34804 22932
rect 34300 22878 34750 22930
rect 34802 22878 34804 22930
rect 34300 22876 34804 22878
rect 34748 22866 34804 22876
rect 34636 22372 34692 22382
rect 34188 22370 34692 22372
rect 34188 22318 34638 22370
rect 34690 22318 34692 22370
rect 34188 22316 34692 22318
rect 33516 21868 34132 21924
rect 34412 22148 34468 22158
rect 34412 21924 34468 22092
rect 32060 21812 32116 21822
rect 31948 21810 32116 21812
rect 31948 21758 32062 21810
rect 32114 21758 32116 21810
rect 31948 21756 32116 21758
rect 32060 21746 32116 21756
rect 32396 21588 32452 21598
rect 33180 21588 33236 21598
rect 32396 21586 33236 21588
rect 32396 21534 32398 21586
rect 32450 21534 33182 21586
rect 33234 21534 33236 21586
rect 32396 21532 33236 21534
rect 32396 21522 32452 21532
rect 33180 21522 33236 21532
rect 30828 21474 31220 21476
rect 30828 21422 30830 21474
rect 30882 21422 31220 21474
rect 30828 21420 31220 21422
rect 30828 20132 30884 21420
rect 33516 21362 33572 21868
rect 34412 21858 34468 21868
rect 34636 21812 34692 22316
rect 34748 22372 34804 22382
rect 34748 21812 34804 22316
rect 34860 22148 34916 24556
rect 34972 23380 35028 23390
rect 34972 23286 35028 23324
rect 35084 23042 35140 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35532 24948 35588 24958
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 23938 35252 23950
rect 35196 23886 35198 23938
rect 35250 23886 35252 23938
rect 35196 23716 35252 23886
rect 35196 23650 35252 23660
rect 35084 22990 35086 23042
rect 35138 22990 35140 23042
rect 35084 22978 35140 22990
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35532 22370 35588 24892
rect 35644 24836 35700 24846
rect 35644 23940 35700 24780
rect 35756 24610 35812 26236
rect 35868 24948 35924 26910
rect 35980 27970 36036 28588
rect 36204 28642 36260 28700
rect 36204 28590 36206 28642
rect 36258 28590 36260 28642
rect 36204 28578 36260 28590
rect 35980 27918 35982 27970
rect 36034 27918 36036 27970
rect 35980 25172 36036 27918
rect 36204 27972 36260 27982
rect 36316 27972 36372 28700
rect 36204 27970 36372 27972
rect 36204 27918 36206 27970
rect 36258 27918 36372 27970
rect 36204 27916 36372 27918
rect 36652 27972 36708 27982
rect 36204 27906 36260 27916
rect 36652 27878 36708 27916
rect 36540 27860 36596 27870
rect 36540 27766 36596 27804
rect 36092 27746 36148 27758
rect 36092 27694 36094 27746
rect 36146 27694 36148 27746
rect 36092 27524 36148 27694
rect 36092 27468 36372 27524
rect 36092 27076 36148 27086
rect 36092 26982 36148 27020
rect 36316 26908 36372 27468
rect 36316 26852 36484 26908
rect 36428 26402 36484 26852
rect 36876 26852 36932 30940
rect 37100 30436 37156 31614
rect 37436 31556 37492 31726
rect 37660 31778 37716 31790
rect 37660 31726 37662 31778
rect 37714 31726 37716 31778
rect 37660 31668 37716 31726
rect 37660 31602 37716 31612
rect 37436 31490 37492 31500
rect 37548 31554 37604 31566
rect 37548 31502 37550 31554
rect 37602 31502 37604 31554
rect 37548 31108 37604 31502
rect 37660 31108 37716 31118
rect 37548 31106 37716 31108
rect 37548 31054 37662 31106
rect 37714 31054 37716 31106
rect 37548 31052 37716 31054
rect 37660 31042 37716 31052
rect 37100 30370 37156 30380
rect 36988 30212 37044 30222
rect 36988 30118 37044 30156
rect 37324 30212 37380 30222
rect 37324 29428 37380 30156
rect 38108 30210 38164 31836
rect 38780 31892 38836 31902
rect 38780 31798 38836 31836
rect 40124 31780 40180 35644
rect 40236 35476 40292 35486
rect 40236 31892 40292 35420
rect 40908 35140 40964 38612
rect 41020 37492 41076 37502
rect 41020 37398 41076 37436
rect 40908 35074 40964 35084
rect 41020 35700 41076 35710
rect 41020 35028 41076 35644
rect 40348 34132 40404 34142
rect 40348 33460 40404 34076
rect 40348 33458 40964 33460
rect 40348 33406 40350 33458
rect 40402 33406 40964 33458
rect 40348 33404 40964 33406
rect 40348 33394 40404 33404
rect 40908 33346 40964 33404
rect 40908 33294 40910 33346
rect 40962 33294 40964 33346
rect 40908 33282 40964 33294
rect 41020 33234 41076 34972
rect 41020 33182 41022 33234
rect 41074 33182 41076 33234
rect 41020 33170 41076 33182
rect 41244 35140 41300 35150
rect 41244 32788 41300 35084
rect 41468 33572 41524 39004
rect 41692 38052 41748 39678
rect 42588 39618 42644 39630
rect 42588 39566 42590 39618
rect 42642 39566 42644 39618
rect 42028 39508 42084 39518
rect 42028 39414 42084 39452
rect 42588 39508 42644 39566
rect 42588 39442 42644 39452
rect 42140 39060 42196 39070
rect 42140 38966 42196 39004
rect 42476 38836 42532 38846
rect 42476 38742 42532 38780
rect 42700 38834 42756 39788
rect 42812 39730 42868 40460
rect 42924 41186 42980 41198
rect 42924 41134 42926 41186
rect 42978 41134 42980 41186
rect 42924 40068 42980 41134
rect 43260 41186 43316 41198
rect 43260 41134 43262 41186
rect 43314 41134 43316 41186
rect 42924 40002 42980 40012
rect 43036 40404 43092 40414
rect 42812 39678 42814 39730
rect 42866 39678 42868 39730
rect 42812 39666 42868 39678
rect 43036 39058 43092 40348
rect 43148 40292 43204 40302
rect 43148 40198 43204 40236
rect 43036 39006 43038 39058
rect 43090 39006 43092 39058
rect 43036 38994 43092 39006
rect 43260 40180 43316 41134
rect 42700 38782 42702 38834
rect 42754 38782 42756 38834
rect 42700 38164 42756 38782
rect 43260 38836 43316 40124
rect 43260 38770 43316 38780
rect 43372 38668 43428 41468
rect 43484 41300 43540 41310
rect 43484 40962 43540 41244
rect 44156 41300 44212 41918
rect 44156 41234 44212 41244
rect 44268 41076 44324 41086
rect 44268 40982 44324 41020
rect 43484 40910 43486 40962
rect 43538 40910 43540 40962
rect 43484 40898 43540 40910
rect 43708 40964 43764 40974
rect 44156 40964 44212 40974
rect 43708 40962 44212 40964
rect 43708 40910 43710 40962
rect 43762 40910 44158 40962
rect 44210 40910 44212 40962
rect 43708 40908 44212 40910
rect 43708 40898 43764 40908
rect 44156 40898 44212 40908
rect 44268 40516 44324 40526
rect 44268 40402 44324 40460
rect 44268 40350 44270 40402
rect 44322 40350 44324 40402
rect 44268 40338 44324 40350
rect 43932 40180 43988 40190
rect 43932 40086 43988 40124
rect 44380 40068 44436 43372
rect 44604 43426 44772 43428
rect 44604 43374 44718 43426
rect 44770 43374 44772 43426
rect 44604 43372 44772 43374
rect 44604 42644 44660 43372
rect 44716 43362 44772 43372
rect 47516 43426 47572 43438
rect 47516 43374 47518 43426
rect 47570 43374 47572 43426
rect 46172 43316 46228 43326
rect 46284 43316 46340 43326
rect 46172 43314 46284 43316
rect 46172 43262 46174 43314
rect 46226 43262 46284 43314
rect 46172 43260 46284 43262
rect 46172 43250 46228 43260
rect 45612 43092 45668 43102
rect 44492 40292 44548 40302
rect 44492 40198 44548 40236
rect 44604 40180 44660 42588
rect 45500 42756 45556 42766
rect 45052 42532 45108 42542
rect 45052 41970 45108 42476
rect 45052 41918 45054 41970
rect 45106 41918 45108 41970
rect 45052 41906 45108 41918
rect 45276 42420 45332 42430
rect 45164 41298 45220 41310
rect 45164 41246 45166 41298
rect 45218 41246 45220 41298
rect 45164 40628 45220 41246
rect 45164 40562 45220 40572
rect 45276 40740 45332 42364
rect 45500 41970 45556 42700
rect 45500 41918 45502 41970
rect 45554 41918 45556 41970
rect 45500 41906 45556 41918
rect 45612 42530 45668 43036
rect 46284 42868 46340 43260
rect 46396 43314 46452 43326
rect 46396 43262 46398 43314
rect 46450 43262 46452 43314
rect 46396 43092 46452 43262
rect 47516 43316 47572 43374
rect 47516 43250 47572 43260
rect 46396 43026 46452 43036
rect 47740 42980 47796 42990
rect 46284 42812 46452 42868
rect 46060 42644 46116 42654
rect 46060 42550 46116 42588
rect 45612 42478 45614 42530
rect 45666 42478 45668 42530
rect 45276 40626 45332 40684
rect 45276 40574 45278 40626
rect 45330 40574 45332 40626
rect 45276 40562 45332 40574
rect 44940 40516 44996 40526
rect 44940 40422 44996 40460
rect 44716 40402 44772 40414
rect 45612 40404 45668 42478
rect 45724 41524 45780 41534
rect 45780 41468 45892 41524
rect 45724 41458 45780 41468
rect 44716 40350 44718 40402
rect 44770 40350 44772 40402
rect 44716 40292 44772 40350
rect 45500 40348 45668 40404
rect 45836 40402 45892 41468
rect 45836 40350 45838 40402
rect 45890 40350 45892 40402
rect 44716 40236 44884 40292
rect 44604 40124 44772 40180
rect 44380 40012 44548 40068
rect 43484 39508 43540 39518
rect 43484 39506 43764 39508
rect 43484 39454 43486 39506
rect 43538 39454 43764 39506
rect 43484 39452 43764 39454
rect 43484 39442 43540 39452
rect 43708 38948 43764 39452
rect 44268 39394 44324 39406
rect 44268 39342 44270 39394
rect 44322 39342 44324 39394
rect 43820 39172 43876 39182
rect 43820 39058 43876 39116
rect 44268 39172 44324 39342
rect 44268 39106 44324 39116
rect 43820 39006 43822 39058
rect 43874 39006 43876 39058
rect 43820 38994 43876 39006
rect 44044 39060 44100 39070
rect 44044 38966 44100 39004
rect 43708 38854 43764 38892
rect 44268 38948 44324 38958
rect 44268 38854 44324 38892
rect 44492 38668 44548 40012
rect 42700 38098 42756 38108
rect 43148 38612 43428 38668
rect 44044 38612 44548 38668
rect 44604 38724 44660 38762
rect 44604 38658 44660 38668
rect 42924 38052 42980 38062
rect 41692 37986 41748 37996
rect 42812 38050 42980 38052
rect 42812 37998 42926 38050
rect 42978 37998 42980 38050
rect 42812 37996 42980 37998
rect 42252 37940 42308 37950
rect 42252 37846 42308 37884
rect 42812 37154 42868 37996
rect 42924 37986 42980 37996
rect 43148 37266 43204 38612
rect 43372 38052 43428 38062
rect 43372 37958 43428 37996
rect 43708 38052 43764 38062
rect 43708 37938 43764 37996
rect 43708 37886 43710 37938
rect 43762 37886 43764 37938
rect 43708 37874 43764 37886
rect 44044 37716 44100 38612
rect 44268 38164 44324 38174
rect 44268 38070 44324 38108
rect 44156 38052 44212 38062
rect 44156 37958 44212 37996
rect 44044 37660 44212 37716
rect 43148 37214 43150 37266
rect 43202 37214 43204 37266
rect 43148 37202 43204 37214
rect 43260 37378 43316 37390
rect 43260 37326 43262 37378
rect 43314 37326 43316 37378
rect 42812 37102 42814 37154
rect 42866 37102 42868 37154
rect 42588 36932 42644 36942
rect 42588 36594 42644 36876
rect 42588 36542 42590 36594
rect 42642 36542 42644 36594
rect 42588 36530 42644 36542
rect 42588 36372 42644 36382
rect 42140 35028 42196 35038
rect 42140 34934 42196 34972
rect 42588 34690 42644 36316
rect 42812 36260 42868 37102
rect 43148 36932 43204 36942
rect 43260 36932 43316 37326
rect 44156 37268 44212 37660
rect 44604 37490 44660 37502
rect 44604 37438 44606 37490
rect 44658 37438 44660 37490
rect 44268 37268 44324 37278
rect 44156 37266 44324 37268
rect 44156 37214 44270 37266
rect 44322 37214 44324 37266
rect 44156 37212 44324 37214
rect 44268 37202 44324 37212
rect 43204 36876 43316 36932
rect 43148 36866 43204 36876
rect 44492 36484 44548 36494
rect 43036 36260 43092 36270
rect 42812 36258 43092 36260
rect 42812 36206 43038 36258
rect 43090 36206 43092 36258
rect 42812 36204 43092 36206
rect 42588 34638 42590 34690
rect 42642 34638 42644 34690
rect 42588 34356 42644 34638
rect 41468 33506 41524 33516
rect 42364 34300 42644 34356
rect 42700 34692 42756 34702
rect 42028 33348 42084 33358
rect 42028 33254 42084 33292
rect 41916 33236 41972 33246
rect 41916 33122 41972 33180
rect 41916 33070 41918 33122
rect 41970 33070 41972 33122
rect 41916 33058 41972 33070
rect 41244 32786 41636 32788
rect 41244 32734 41246 32786
rect 41298 32734 41636 32786
rect 41244 32732 41636 32734
rect 41244 32722 41300 32732
rect 40684 31892 40740 31902
rect 40236 31836 40628 31892
rect 40124 31724 40404 31780
rect 38892 31668 38948 31678
rect 38892 31666 39844 31668
rect 38892 31614 38894 31666
rect 38946 31614 39844 31666
rect 38892 31612 39844 31614
rect 38892 31602 38948 31612
rect 38332 31556 38388 31566
rect 38332 31462 38388 31500
rect 38892 30884 38948 30894
rect 38892 30324 38948 30828
rect 39788 30882 39844 31612
rect 40348 31666 40404 31724
rect 40348 31614 40350 31666
rect 40402 31614 40404 31666
rect 40348 30996 40404 31614
rect 40572 31668 40628 31836
rect 40684 31890 41188 31892
rect 40684 31838 40686 31890
rect 40738 31838 41188 31890
rect 40684 31836 41188 31838
rect 40684 31826 40740 31836
rect 40572 31574 40628 31612
rect 40348 30930 40404 30940
rect 40460 31220 40516 31230
rect 39788 30830 39790 30882
rect 39842 30830 39844 30882
rect 39788 30818 39844 30830
rect 39564 30436 39620 30446
rect 39564 30342 39620 30380
rect 38108 30158 38110 30210
rect 38162 30158 38164 30210
rect 38108 30146 38164 30158
rect 38780 30212 38836 30222
rect 38780 30118 38836 30156
rect 37324 29362 37380 29372
rect 37996 29428 38052 29438
rect 37548 29092 37604 29102
rect 37100 28756 37156 28766
rect 37100 28662 37156 28700
rect 37548 28644 37604 29036
rect 37996 28756 38052 29372
rect 37996 28662 38052 28700
rect 37436 28642 37604 28644
rect 37436 28590 37550 28642
rect 37602 28590 37604 28642
rect 37436 28588 37604 28590
rect 37436 27298 37492 28588
rect 37548 28578 37604 28588
rect 38332 28644 38388 28654
rect 38332 28550 38388 28588
rect 38668 28532 38724 28542
rect 38668 28530 38836 28532
rect 38668 28478 38670 28530
rect 38722 28478 38836 28530
rect 38668 28476 38836 28478
rect 38668 28466 38724 28476
rect 38668 27860 38724 27870
rect 38780 27860 38836 28476
rect 37436 27246 37438 27298
rect 37490 27246 37492 27298
rect 37436 27234 37492 27246
rect 38556 27858 38836 27860
rect 38556 27806 38670 27858
rect 38722 27806 38836 27858
rect 38556 27804 38836 27806
rect 37212 27074 37268 27086
rect 37212 27022 37214 27074
rect 37266 27022 37268 27074
rect 36876 26786 36932 26796
rect 36988 26962 37044 26974
rect 36988 26910 36990 26962
rect 37042 26910 37044 26962
rect 36428 26350 36430 26402
rect 36482 26350 36484 26402
rect 36428 26338 36484 26350
rect 36988 25844 37044 26910
rect 37212 26908 37268 27022
rect 37548 27074 37604 27086
rect 37548 27022 37550 27074
rect 37602 27022 37604 27074
rect 37100 26850 37156 26862
rect 37212 26852 37492 26908
rect 37100 26798 37102 26850
rect 37154 26798 37156 26850
rect 37100 26740 37156 26798
rect 37100 26674 37156 26684
rect 36876 25788 37044 25844
rect 37324 26628 37380 26638
rect 36428 25620 36484 25630
rect 36428 25506 36484 25564
rect 36428 25454 36430 25506
rect 36482 25454 36484 25506
rect 36428 25442 36484 25454
rect 36876 25284 36932 25788
rect 37324 25732 37380 26572
rect 36988 25676 37380 25732
rect 36988 25506 37044 25676
rect 37436 25620 37492 26852
rect 36988 25454 36990 25506
rect 37042 25454 37044 25506
rect 36988 25442 37044 25454
rect 37100 25564 37492 25620
rect 37548 25620 37604 27022
rect 37996 27074 38052 27086
rect 37996 27022 37998 27074
rect 38050 27022 38052 27074
rect 36876 25228 37044 25284
rect 35980 25116 36484 25172
rect 35868 24892 36036 24948
rect 35756 24558 35758 24610
rect 35810 24558 35812 24610
rect 35756 24546 35812 24558
rect 35644 23938 35924 23940
rect 35644 23886 35646 23938
rect 35698 23886 35924 23938
rect 35644 23884 35924 23886
rect 35644 23874 35700 23884
rect 35756 22932 35812 22942
rect 35532 22318 35534 22370
rect 35586 22318 35588 22370
rect 35532 22306 35588 22318
rect 35644 22876 35756 22932
rect 35196 22148 35252 22158
rect 34860 22146 35252 22148
rect 34860 22094 35198 22146
rect 35250 22094 35252 22146
rect 34860 22092 35252 22094
rect 34972 21812 35028 21822
rect 34748 21810 35028 21812
rect 34748 21758 34974 21810
rect 35026 21758 35028 21810
rect 34748 21756 35028 21758
rect 34636 21746 34692 21756
rect 34972 21746 35028 21756
rect 33740 21698 33796 21710
rect 33740 21646 33742 21698
rect 33794 21646 33796 21698
rect 33740 21476 33796 21646
rect 33740 21410 33796 21420
rect 33852 21700 33908 21710
rect 34076 21700 34132 21710
rect 33908 21698 34132 21700
rect 33908 21646 34078 21698
rect 34130 21646 34132 21698
rect 33908 21644 34132 21646
rect 33516 21310 33518 21362
rect 33570 21310 33572 21362
rect 33516 21028 33572 21310
rect 32732 20972 33572 21028
rect 32508 20580 32564 20590
rect 32396 20578 32564 20580
rect 32396 20526 32510 20578
rect 32562 20526 32564 20578
rect 32396 20524 32564 20526
rect 30828 19236 30884 20076
rect 32060 20130 32116 20142
rect 32060 20078 32062 20130
rect 32114 20078 32116 20130
rect 31276 19908 31332 19918
rect 31276 19814 31332 19852
rect 31948 19348 32004 19358
rect 32060 19348 32116 20078
rect 32396 20130 32452 20524
rect 32508 20514 32564 20524
rect 32396 20078 32398 20130
rect 32450 20078 32452 20130
rect 32396 20066 32452 20078
rect 31948 19346 32116 19348
rect 31948 19294 31950 19346
rect 32002 19294 32116 19346
rect 31948 19292 32116 19294
rect 31948 19282 32004 19292
rect 31164 19236 31220 19246
rect 30828 19234 31220 19236
rect 30828 19182 31166 19234
rect 31218 19182 31220 19234
rect 30828 19180 31220 19182
rect 29932 18510 29934 18562
rect 29986 18510 29988 18562
rect 29932 18498 29988 18510
rect 30604 18788 30660 18798
rect 30380 17554 30436 17566
rect 30380 17502 30382 17554
rect 30434 17502 30436 17554
rect 30380 16322 30436 17502
rect 30604 17108 30660 18732
rect 30828 18674 30884 19180
rect 31164 19170 31220 19180
rect 30828 18622 30830 18674
rect 30882 18622 30884 18674
rect 30828 18610 30884 18622
rect 32396 18452 32452 18462
rect 32172 17668 32228 17678
rect 32172 17574 32228 17612
rect 31836 17556 31892 17566
rect 31836 17462 31892 17500
rect 32396 17554 32452 18396
rect 32396 17502 32398 17554
rect 32450 17502 32452 17554
rect 32396 17490 32452 17502
rect 32732 17554 32788 20972
rect 32844 20802 32900 20814
rect 32844 20750 32846 20802
rect 32898 20750 32900 20802
rect 32844 18788 32900 20750
rect 33068 20690 33124 20702
rect 33068 20638 33070 20690
rect 33122 20638 33124 20690
rect 33068 19796 33124 20638
rect 33628 20692 33684 20702
rect 33852 20692 33908 21644
rect 34076 21634 34132 21644
rect 35084 21588 35140 22092
rect 35196 22082 35252 22092
rect 35196 21812 35252 21822
rect 35532 21812 35588 21822
rect 35644 21812 35700 22876
rect 35756 22866 35812 22876
rect 35756 22372 35812 22382
rect 35756 22278 35812 22316
rect 35196 21718 35252 21756
rect 35308 21810 35700 21812
rect 35308 21758 35534 21810
rect 35586 21758 35700 21810
rect 35308 21756 35700 21758
rect 35756 22036 35812 22046
rect 35756 21810 35812 21980
rect 35756 21758 35758 21810
rect 35810 21758 35812 21810
rect 35308 21698 35364 21756
rect 35532 21746 35588 21756
rect 35756 21746 35812 21758
rect 35308 21646 35310 21698
rect 35362 21646 35364 21698
rect 35308 21634 35364 21646
rect 35868 21698 35924 23884
rect 35980 22820 36036 24892
rect 36316 24722 36372 24734
rect 36316 24670 36318 24722
rect 36370 24670 36372 24722
rect 36316 24612 36372 24670
rect 36316 24546 36372 24556
rect 36092 24052 36148 24062
rect 36092 23958 36148 23996
rect 36204 23828 36260 23838
rect 36204 23734 36260 23772
rect 36428 23828 36484 25116
rect 36428 23762 36484 23772
rect 36652 24276 36708 24286
rect 36316 23042 36372 23054
rect 36316 22990 36318 23042
rect 36370 22990 36372 23042
rect 35980 22764 36260 22820
rect 36204 22708 36260 22764
rect 35868 21646 35870 21698
rect 35922 21646 35924 21698
rect 35868 21634 35924 21646
rect 35980 22596 36036 22606
rect 35980 22370 36036 22540
rect 36204 22482 36260 22652
rect 36204 22430 36206 22482
rect 36258 22430 36260 22482
rect 36204 22418 36260 22430
rect 35980 22318 35982 22370
rect 36034 22318 36036 22370
rect 34860 21532 35140 21588
rect 34524 20804 34580 20814
rect 34524 20710 34580 20748
rect 33628 20690 33908 20692
rect 33628 20638 33630 20690
rect 33682 20638 33908 20690
rect 33628 20636 33908 20638
rect 33628 20626 33684 20636
rect 34748 20578 34804 20590
rect 34748 20526 34750 20578
rect 34802 20526 34804 20578
rect 34748 20132 34804 20526
rect 34748 20066 34804 20076
rect 34636 20018 34692 20030
rect 34636 19966 34638 20018
rect 34690 19966 34692 20018
rect 34300 19908 34356 19918
rect 34300 19814 34356 19852
rect 33068 19730 33124 19740
rect 34076 19346 34132 19358
rect 34076 19294 34078 19346
rect 34130 19294 34132 19346
rect 34076 18788 34132 19294
rect 32844 18732 34132 18788
rect 32732 17502 32734 17554
rect 32786 17502 32788 17554
rect 32732 17490 32788 17502
rect 33404 17778 33460 17790
rect 33404 17726 33406 17778
rect 33458 17726 33460 17778
rect 33404 17668 33460 17726
rect 30716 17444 30772 17454
rect 30716 17442 31780 17444
rect 30716 17390 30718 17442
rect 30770 17390 31780 17442
rect 30716 17388 31780 17390
rect 30716 17378 30772 17388
rect 30604 17042 30660 17052
rect 31724 16994 31780 17388
rect 31724 16942 31726 16994
rect 31778 16942 31780 16994
rect 31724 16930 31780 16942
rect 33404 16996 33460 17612
rect 33404 16930 33460 16940
rect 32508 16884 32564 16894
rect 32508 16790 32564 16828
rect 33180 16884 33236 16894
rect 33180 16790 33236 16828
rect 30380 16270 30382 16322
rect 30434 16270 30436 16322
rect 30380 16258 30436 16270
rect 30716 16660 30772 16670
rect 30716 16322 30772 16604
rect 30716 16270 30718 16322
rect 30770 16270 30772 16322
rect 29932 15988 29988 15998
rect 29932 15986 30100 15988
rect 29932 15934 29934 15986
rect 29986 15934 30100 15986
rect 29932 15932 30100 15934
rect 29932 15922 29988 15932
rect 29932 15764 29988 15774
rect 29932 15204 29988 15708
rect 29932 12178 29988 15148
rect 29932 12126 29934 12178
rect 29986 12126 29988 12178
rect 29932 11620 29988 12126
rect 29932 11554 29988 11564
rect 29260 11506 29876 11508
rect 29260 11454 29262 11506
rect 29314 11454 29710 11506
rect 29762 11454 29876 11506
rect 29260 11452 29876 11454
rect 29260 11442 29316 11452
rect 29484 10834 29540 11452
rect 29708 11442 29764 11452
rect 29484 10782 29486 10834
rect 29538 10782 29540 10834
rect 29484 9826 29540 10782
rect 29820 10722 29876 10734
rect 29820 10670 29822 10722
rect 29874 10670 29876 10722
rect 29820 10388 29876 10670
rect 29820 10322 29876 10332
rect 29932 10052 29988 10062
rect 30044 10052 30100 15932
rect 30716 15764 30772 16270
rect 30716 15698 30772 15708
rect 30940 15986 30996 15998
rect 30940 15934 30942 15986
rect 30994 15934 30996 15986
rect 30940 15652 30996 15934
rect 31276 15988 31332 15998
rect 31276 15894 31332 15932
rect 30940 15586 30996 15596
rect 31388 15652 31444 15662
rect 30940 15428 30996 15438
rect 30828 15092 30884 15102
rect 30604 15090 30884 15092
rect 30604 15038 30830 15090
rect 30882 15038 30884 15090
rect 30604 15036 30884 15038
rect 30604 14530 30660 15036
rect 30828 15026 30884 15036
rect 30940 14644 30996 15372
rect 31388 15426 31444 15596
rect 31388 15374 31390 15426
rect 31442 15374 31444 15426
rect 31388 15362 31444 15374
rect 31724 15428 31780 15438
rect 31724 15334 31780 15372
rect 31164 15092 31220 15102
rect 31164 15090 31444 15092
rect 31164 15038 31166 15090
rect 31218 15038 31444 15090
rect 31164 15036 31444 15038
rect 31164 15026 31220 15036
rect 31164 14644 31220 14654
rect 30940 14642 31220 14644
rect 30940 14590 31166 14642
rect 31218 14590 31220 14642
rect 30940 14588 31220 14590
rect 31164 14578 31220 14588
rect 30604 14478 30606 14530
rect 30658 14478 30660 14530
rect 30604 14466 30660 14478
rect 30828 14420 30884 14430
rect 30828 14326 30884 14364
rect 31276 12852 31332 12862
rect 31276 12758 31332 12796
rect 30268 12740 30324 12750
rect 30268 12290 30324 12684
rect 30268 12238 30270 12290
rect 30322 12238 30324 12290
rect 30268 12226 30324 12238
rect 30492 12292 30548 12302
rect 30492 12198 30548 12236
rect 30492 10724 30548 10734
rect 30492 10722 31108 10724
rect 30492 10670 30494 10722
rect 30546 10670 31108 10722
rect 30492 10668 31108 10670
rect 30492 10658 30548 10668
rect 30268 10610 30324 10622
rect 30268 10558 30270 10610
rect 30322 10558 30324 10610
rect 30268 10500 30324 10558
rect 30940 10500 30996 10510
rect 30268 10498 30996 10500
rect 30268 10446 30942 10498
rect 30994 10446 30996 10498
rect 30268 10444 30996 10446
rect 30940 10434 30996 10444
rect 29932 10050 30100 10052
rect 29932 9998 29934 10050
rect 29986 9998 30100 10050
rect 29932 9996 30100 9998
rect 29932 9986 29988 9996
rect 29820 9940 29876 9950
rect 29820 9846 29876 9884
rect 30604 9940 30660 9950
rect 29484 9774 29486 9826
rect 29538 9774 29540 9826
rect 29484 9762 29540 9774
rect 30268 9826 30324 9838
rect 30268 9774 30270 9826
rect 30322 9774 30324 9826
rect 29148 9604 29204 9614
rect 29148 9510 29204 9548
rect 30268 8428 30324 9774
rect 30604 8930 30660 9884
rect 31052 9938 31108 10668
rect 31276 10612 31332 10622
rect 31388 10612 31444 15036
rect 33292 14420 33348 14430
rect 33292 14326 33348 14364
rect 33180 14196 33236 14206
rect 33180 13970 33236 14140
rect 33180 13918 33182 13970
rect 33234 13918 33236 13970
rect 33180 13906 33236 13918
rect 33516 13746 33572 18732
rect 34076 18562 34132 18574
rect 34076 18510 34078 18562
rect 34130 18510 34132 18562
rect 33740 18452 33796 18462
rect 33628 18450 33796 18452
rect 33628 18398 33742 18450
rect 33794 18398 33796 18450
rect 33628 18396 33796 18398
rect 33628 17106 33684 18396
rect 33740 18386 33796 18396
rect 34076 17780 34132 18510
rect 34076 17714 34132 17724
rect 33628 17054 33630 17106
rect 33682 17054 33684 17106
rect 33628 17042 33684 17054
rect 34188 17108 34244 17118
rect 34188 16994 34244 17052
rect 34188 16942 34190 16994
rect 34242 16942 34244 16994
rect 34188 16930 34244 16942
rect 34524 16996 34580 17006
rect 34524 16902 34580 16940
rect 33852 16884 33908 16894
rect 33852 14532 33908 16828
rect 34636 16884 34692 19966
rect 34860 20020 34916 21532
rect 35756 21476 35812 21486
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 20804 35252 20814
rect 35196 20710 35252 20748
rect 35532 20804 35588 20814
rect 35532 20802 35700 20804
rect 35532 20750 35534 20802
rect 35586 20750 35700 20802
rect 35532 20748 35700 20750
rect 35532 20738 35588 20748
rect 35308 20132 35364 20142
rect 35308 20038 35364 20076
rect 34860 19954 34916 19964
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35532 19234 35588 19246
rect 35532 19182 35534 19234
rect 35586 19182 35588 19234
rect 35196 19012 35252 19022
rect 34972 19010 35252 19012
rect 34972 18958 35198 19010
rect 35250 18958 35252 19010
rect 34972 18956 35252 18958
rect 34972 18450 35028 18956
rect 35196 18946 35252 18956
rect 34972 18398 34974 18450
rect 35026 18398 35028 18450
rect 34972 18386 35028 18398
rect 35196 18562 35252 18574
rect 35196 18510 35198 18562
rect 35250 18510 35252 18562
rect 35196 18452 35252 18510
rect 35196 18386 35252 18396
rect 35532 18340 35588 19182
rect 35644 18900 35700 20748
rect 35756 20690 35812 21420
rect 35756 20638 35758 20690
rect 35810 20638 35812 20690
rect 35756 20626 35812 20638
rect 35980 19908 36036 22318
rect 36316 21586 36372 22990
rect 36652 22596 36708 24220
rect 36988 24164 37044 25228
rect 37100 24724 37156 25564
rect 37548 25554 37604 25564
rect 37660 26852 37716 26862
rect 37660 25506 37716 26796
rect 37660 25454 37662 25506
rect 37714 25454 37716 25506
rect 37660 25442 37716 25454
rect 37884 25620 37940 25630
rect 37324 25396 37380 25406
rect 37324 25302 37380 25340
rect 37212 25282 37268 25294
rect 37212 25230 37214 25282
rect 37266 25230 37268 25282
rect 37212 24948 37268 25230
rect 37212 24882 37268 24892
rect 37884 24834 37940 25564
rect 37884 24782 37886 24834
rect 37938 24782 37940 24834
rect 37884 24770 37940 24782
rect 37212 24724 37268 24734
rect 37100 24722 37268 24724
rect 37100 24670 37214 24722
rect 37266 24670 37268 24722
rect 37100 24668 37268 24670
rect 36652 22530 36708 22540
rect 36876 24108 37044 24164
rect 36876 22372 36932 24108
rect 37212 24052 37268 24668
rect 37212 23986 37268 23996
rect 37436 24612 37492 24622
rect 36876 22306 36932 22316
rect 36988 23938 37044 23950
rect 36988 23886 36990 23938
rect 37042 23886 37044 23938
rect 36428 22260 36484 22270
rect 36428 22166 36484 22204
rect 36988 22260 37044 23886
rect 37100 23828 37156 23838
rect 37100 23734 37156 23772
rect 37212 23716 37268 23726
rect 37212 23622 37268 23660
rect 36988 22194 37044 22204
rect 37100 23492 37156 23502
rect 37100 22482 37156 23436
rect 37436 23154 37492 24556
rect 37996 24164 38052 27022
rect 38332 26852 38388 26862
rect 38332 26758 38388 26796
rect 38556 26178 38612 27804
rect 38668 27794 38724 27804
rect 38780 27188 38836 27198
rect 38780 27094 38836 27132
rect 38892 26628 38948 30268
rect 40460 30324 40516 31164
rect 41020 30882 41076 30894
rect 41020 30830 41022 30882
rect 41074 30830 41076 30882
rect 41020 30772 41076 30830
rect 39452 30210 39508 30222
rect 39452 30158 39454 30210
rect 39506 30158 39508 30210
rect 39228 30098 39284 30110
rect 39228 30046 39230 30098
rect 39282 30046 39284 30098
rect 39228 28532 39284 30046
rect 38892 26562 38948 26572
rect 39116 28476 39284 28532
rect 38892 26292 38948 26302
rect 38892 26290 39060 26292
rect 38892 26238 38894 26290
rect 38946 26238 39060 26290
rect 38892 26236 39060 26238
rect 38892 26226 38948 26236
rect 38556 26126 38558 26178
rect 38610 26126 38612 26178
rect 38556 26114 38612 26126
rect 38892 26068 38948 26078
rect 38668 26066 38948 26068
rect 38668 26014 38894 26066
rect 38946 26014 38948 26066
rect 38668 26012 38948 26014
rect 38668 25732 38724 26012
rect 38892 26002 38948 26012
rect 38444 25676 38724 25732
rect 38444 25618 38500 25676
rect 38444 25566 38446 25618
rect 38498 25566 38500 25618
rect 38444 25554 38500 25566
rect 38108 25396 38164 25406
rect 38164 25340 38500 25396
rect 38108 25330 38164 25340
rect 37996 24108 38388 24164
rect 37436 23102 37438 23154
rect 37490 23102 37492 23154
rect 37436 23090 37492 23102
rect 37996 23940 38052 23950
rect 37100 22430 37102 22482
rect 37154 22430 37156 22482
rect 36540 22148 36596 22158
rect 36540 22146 36932 22148
rect 36540 22094 36542 22146
rect 36594 22094 36932 22146
rect 36540 22092 36932 22094
rect 36540 22082 36596 22092
rect 36876 21700 36932 22092
rect 37100 22036 37156 22430
rect 37100 21970 37156 21980
rect 37212 22708 37268 22718
rect 36988 21700 37044 21710
rect 36876 21698 37044 21700
rect 36876 21646 36990 21698
rect 37042 21646 37044 21698
rect 36876 21644 37044 21646
rect 36988 21634 37044 21644
rect 36316 21534 36318 21586
rect 36370 21534 36372 21586
rect 35980 19842 36036 19852
rect 36092 20690 36148 20702
rect 36092 20638 36094 20690
rect 36146 20638 36148 20690
rect 35756 19796 35812 19806
rect 35756 19122 35812 19740
rect 35756 19070 35758 19122
rect 35810 19070 35812 19122
rect 35756 19058 35812 19070
rect 36092 19124 36148 20638
rect 36316 19908 36372 21534
rect 36316 19842 36372 19852
rect 37212 19346 37268 22652
rect 37324 22370 37380 22382
rect 37324 22318 37326 22370
rect 37378 22318 37380 22370
rect 37324 22260 37380 22318
rect 37996 22370 38052 23884
rect 38220 23380 38276 23390
rect 37996 22318 37998 22370
rect 38050 22318 38052 22370
rect 37996 22306 38052 22318
rect 38108 23324 38220 23380
rect 37324 20914 37380 22204
rect 37324 20862 37326 20914
rect 37378 20862 37380 20914
rect 37324 20850 37380 20862
rect 37660 21476 37716 21486
rect 37660 20914 37716 21420
rect 38108 21028 38164 23324
rect 38220 23314 38276 23324
rect 38332 23156 38388 24108
rect 38444 23378 38500 25340
rect 39004 25172 39060 26236
rect 38668 25116 39060 25172
rect 38556 24722 38612 24734
rect 38556 24670 38558 24722
rect 38610 24670 38612 24722
rect 38556 23492 38612 24670
rect 38556 23426 38612 23436
rect 38444 23326 38446 23378
rect 38498 23326 38500 23378
rect 38444 23314 38500 23326
rect 38556 23266 38612 23278
rect 38556 23214 38558 23266
rect 38610 23214 38612 23266
rect 38556 23156 38612 23214
rect 38332 23100 38612 23156
rect 38332 22932 38388 22942
rect 38332 22838 38388 22876
rect 38220 22484 38276 22494
rect 38220 22370 38276 22428
rect 38220 22318 38222 22370
rect 38274 22318 38276 22370
rect 38220 22306 38276 22318
rect 38332 21924 38388 21934
rect 38444 21924 38500 23100
rect 38668 23044 38724 25116
rect 39116 25060 39172 28476
rect 39340 28084 39396 28094
rect 39452 28084 39508 30158
rect 40124 30212 40180 30222
rect 40124 30118 40180 30156
rect 40460 30098 40516 30268
rect 40908 30716 41020 30772
rect 40796 30212 40852 30222
rect 40796 30118 40852 30156
rect 40460 30046 40462 30098
rect 40514 30046 40516 30098
rect 40460 30034 40516 30046
rect 39788 29986 39844 29998
rect 39788 29934 39790 29986
rect 39842 29934 39844 29986
rect 39676 28756 39732 28766
rect 39676 28662 39732 28700
rect 39788 28644 39844 29934
rect 40908 29092 40964 30716
rect 41020 30706 41076 30716
rect 41132 30212 41188 31836
rect 41244 31778 41300 31790
rect 41244 31726 41246 31778
rect 41298 31726 41300 31778
rect 41244 31108 41300 31726
rect 41244 31042 41300 31052
rect 41020 30210 41188 30212
rect 41020 30158 41134 30210
rect 41186 30158 41188 30210
rect 41020 30156 41188 30158
rect 41020 29426 41076 30156
rect 41132 30146 41188 30156
rect 41020 29374 41022 29426
rect 41074 29374 41076 29426
rect 41020 29362 41076 29374
rect 41244 29538 41300 29550
rect 41244 29486 41246 29538
rect 41298 29486 41300 29538
rect 40796 29036 40964 29092
rect 41244 29092 41300 29486
rect 40684 28756 40740 28766
rect 40012 28644 40068 28654
rect 39788 28642 40068 28644
rect 39788 28590 40014 28642
rect 40066 28590 40068 28642
rect 39788 28588 40068 28590
rect 39340 28082 39508 28084
rect 39340 28030 39342 28082
rect 39394 28030 39508 28082
rect 39340 28028 39508 28030
rect 39340 28018 39396 28028
rect 39228 27970 39284 27982
rect 39228 27918 39230 27970
rect 39282 27918 39284 27970
rect 39228 26908 39284 27918
rect 40012 27748 40068 28588
rect 40684 28642 40740 28700
rect 40684 28590 40686 28642
rect 40738 28590 40740 28642
rect 40684 28578 40740 28590
rect 40012 27682 40068 27692
rect 40348 28418 40404 28430
rect 40348 28366 40350 28418
rect 40402 28366 40404 28418
rect 39564 27188 39620 27198
rect 39228 26852 39396 26908
rect 39004 25004 39172 25060
rect 39228 26066 39284 26078
rect 39228 26014 39230 26066
rect 39282 26014 39284 26066
rect 39004 23378 39060 25004
rect 39228 24948 39284 26014
rect 39228 24882 39284 24892
rect 39116 24836 39172 24846
rect 39116 24742 39172 24780
rect 39004 23326 39006 23378
rect 39058 23326 39060 23378
rect 39004 23314 39060 23326
rect 38388 21868 38500 21924
rect 38556 22988 38724 23044
rect 38220 21028 38276 21038
rect 38108 21026 38276 21028
rect 38108 20974 38222 21026
rect 38274 20974 38276 21026
rect 38108 20972 38276 20974
rect 38220 20962 38276 20972
rect 37660 20862 37662 20914
rect 37714 20862 37716 20914
rect 37660 20850 37716 20862
rect 38108 20804 38164 20814
rect 38332 20804 38388 21868
rect 38444 21700 38500 21710
rect 38444 21026 38500 21644
rect 38444 20974 38446 21026
rect 38498 20974 38500 21026
rect 38444 20962 38500 20974
rect 38556 21026 38612 22988
rect 39228 21812 39284 21822
rect 39340 21812 39396 26852
rect 39564 23042 39620 27132
rect 40348 26908 40404 28366
rect 40348 26852 40516 26908
rect 40012 26628 40068 26638
rect 40236 26628 40292 26638
rect 39788 26292 39844 26302
rect 39788 26198 39844 26236
rect 39900 26178 39956 26190
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39788 25060 39844 25070
rect 39788 23154 39844 25004
rect 39900 23380 39956 26126
rect 39900 23314 39956 23324
rect 40012 24610 40068 26572
rect 40124 26572 40236 26628
rect 40124 26402 40180 26572
rect 40236 26562 40292 26572
rect 40124 26350 40126 26402
rect 40178 26350 40180 26402
rect 40124 26338 40180 26350
rect 40348 26290 40404 26302
rect 40348 26238 40350 26290
rect 40402 26238 40404 26290
rect 40348 25172 40404 26238
rect 40348 25106 40404 25116
rect 40012 24558 40014 24610
rect 40066 24558 40068 24610
rect 39788 23102 39790 23154
rect 39842 23102 39844 23154
rect 39788 23090 39844 23102
rect 39900 23154 39956 23166
rect 39900 23102 39902 23154
rect 39954 23102 39956 23154
rect 39564 22990 39566 23042
rect 39618 22990 39620 23042
rect 39564 22978 39620 22990
rect 39228 21810 39340 21812
rect 39228 21758 39230 21810
rect 39282 21758 39340 21810
rect 39228 21756 39340 21758
rect 38556 20974 38558 21026
rect 38610 20974 38612 21026
rect 38556 20962 38612 20974
rect 39116 21700 39172 21710
rect 38108 20802 38388 20804
rect 38108 20750 38110 20802
rect 38162 20750 38388 20802
rect 38108 20748 38388 20750
rect 39004 20802 39060 20814
rect 39004 20750 39006 20802
rect 39058 20750 39060 20802
rect 38108 20738 38164 20748
rect 37212 19294 37214 19346
rect 37266 19294 37268 19346
rect 37212 19282 37268 19294
rect 37436 19906 37492 19918
rect 37436 19854 37438 19906
rect 37490 19854 37492 19906
rect 36092 19030 36148 19068
rect 35644 18834 35700 18844
rect 36316 18900 36372 18910
rect 35532 18338 35700 18340
rect 35532 18286 35534 18338
rect 35586 18286 35700 18338
rect 35532 18284 35700 18286
rect 35532 18274 35588 18284
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35532 17780 35588 17790
rect 35644 17780 35700 18284
rect 35644 17724 36036 17780
rect 35532 17686 35588 17724
rect 34636 16818 34692 16828
rect 35532 17108 35588 17118
rect 33964 16660 34020 16670
rect 33964 16566 34020 16604
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35532 16324 35588 17052
rect 35308 16268 35588 16324
rect 35196 15874 35252 15886
rect 35196 15822 35198 15874
rect 35250 15822 35252 15874
rect 35084 15314 35140 15326
rect 35084 15262 35086 15314
rect 35138 15262 35140 15314
rect 35084 14756 35140 15262
rect 35196 15092 35252 15822
rect 35308 15092 35364 16268
rect 35532 16098 35588 16110
rect 35532 16046 35534 16098
rect 35586 16046 35588 16098
rect 35420 15428 35476 15438
rect 35420 15334 35476 15372
rect 35532 15204 35588 16046
rect 35756 15986 35812 15998
rect 35756 15934 35758 15986
rect 35810 15934 35812 15986
rect 35756 15540 35812 15934
rect 35756 15474 35812 15484
rect 35756 15204 35812 15214
rect 35532 15202 35812 15204
rect 35532 15150 35758 15202
rect 35810 15150 35812 15202
rect 35532 15148 35812 15150
rect 35980 15148 36036 17724
rect 36204 17668 36260 17678
rect 36204 16884 36260 17612
rect 36204 16818 36260 16828
rect 36316 15986 36372 18844
rect 37436 18900 37492 19854
rect 37884 19908 37940 19918
rect 37884 19814 37940 19852
rect 38556 19908 38612 19918
rect 37436 18834 37492 18844
rect 37660 18452 37716 18462
rect 37660 18358 37716 18396
rect 38444 18452 38500 18462
rect 38556 18452 38612 19852
rect 39004 19908 39060 20750
rect 39116 20242 39172 21644
rect 39228 21476 39284 21756
rect 39340 21718 39396 21756
rect 39900 22372 39956 23102
rect 39788 21588 39844 21598
rect 39900 21588 39956 22316
rect 40012 21700 40068 24558
rect 40348 24836 40404 24846
rect 40012 21634 40068 21644
rect 40236 23828 40292 23838
rect 40236 22484 40292 23772
rect 39788 21586 39956 21588
rect 39788 21534 39790 21586
rect 39842 21534 39956 21586
rect 39788 21532 39956 21534
rect 39228 21410 39284 21420
rect 39676 21476 39732 21486
rect 39676 20914 39732 21420
rect 39676 20862 39678 20914
rect 39730 20862 39732 20914
rect 39676 20850 39732 20862
rect 39116 20190 39118 20242
rect 39170 20190 39172 20242
rect 39116 20178 39172 20190
rect 39788 20018 39844 21532
rect 40236 21474 40292 22428
rect 40348 22482 40404 24780
rect 40460 23716 40516 26852
rect 40796 26068 40852 29036
rect 41244 29026 41300 29036
rect 41356 28756 41412 32732
rect 41580 32562 41636 32732
rect 41580 32510 41582 32562
rect 41634 32510 41636 32562
rect 41580 32498 41636 32510
rect 41804 32450 41860 32462
rect 41804 32398 41806 32450
rect 41858 32398 41860 32450
rect 41804 31892 41860 32398
rect 41916 32452 41972 32462
rect 41916 32358 41972 32396
rect 41916 31892 41972 31902
rect 41804 31890 41972 31892
rect 41804 31838 41918 31890
rect 41970 31838 41972 31890
rect 41804 31836 41972 31838
rect 41916 31826 41972 31836
rect 41916 31668 41972 31678
rect 41916 31106 41972 31612
rect 41916 31054 41918 31106
rect 41970 31054 41972 31106
rect 41916 31042 41972 31054
rect 41468 30994 41524 31006
rect 41468 30942 41470 30994
rect 41522 30942 41524 30994
rect 41468 30212 41524 30942
rect 42140 30996 42196 31006
rect 42140 30902 42196 30940
rect 41804 30212 41860 30222
rect 41524 30210 41860 30212
rect 41524 30158 41806 30210
rect 41858 30158 41860 30210
rect 41524 30156 41860 30158
rect 41468 30098 41524 30156
rect 41804 30146 41860 30156
rect 41468 30046 41470 30098
rect 41522 30046 41524 30098
rect 41468 30034 41524 30046
rect 42140 29986 42196 29998
rect 42140 29934 42142 29986
rect 42194 29934 42196 29986
rect 42140 29876 42196 29934
rect 42140 29810 42196 29820
rect 41356 28690 41412 28700
rect 41916 28644 41972 28654
rect 41020 28532 41076 28542
rect 41020 28530 41636 28532
rect 41020 28478 41022 28530
rect 41074 28478 41636 28530
rect 41020 28476 41636 28478
rect 41020 28466 41076 28476
rect 40908 28418 40964 28430
rect 40908 28366 40910 28418
rect 40962 28366 40964 28418
rect 40908 27186 40964 28366
rect 41580 27860 41636 28476
rect 41692 28084 41748 28094
rect 41916 28084 41972 28588
rect 42364 28644 42420 34300
rect 42588 34132 42644 34142
rect 42588 33234 42644 34076
rect 42700 34130 42756 34636
rect 42700 34078 42702 34130
rect 42754 34078 42756 34130
rect 42700 34066 42756 34078
rect 42924 34690 42980 34702
rect 42924 34638 42926 34690
rect 42978 34638 42980 34690
rect 42924 34468 42980 34638
rect 43036 34692 43092 36204
rect 44268 36260 44324 36270
rect 44380 36260 44436 36270
rect 44268 36258 44380 36260
rect 44268 36206 44270 36258
rect 44322 36206 44380 36258
rect 44268 36204 44380 36206
rect 44268 36194 44324 36204
rect 44044 35924 44100 35934
rect 43036 34626 43092 34636
rect 43148 35586 43204 35598
rect 43148 35534 43150 35586
rect 43202 35534 43204 35586
rect 43148 34468 43204 35534
rect 44044 35138 44100 35868
rect 44268 35588 44324 35598
rect 44268 35494 44324 35532
rect 44044 35086 44046 35138
rect 44098 35086 44100 35138
rect 44044 35074 44100 35086
rect 44156 35476 44212 35486
rect 44156 35138 44212 35420
rect 44156 35086 44158 35138
rect 44210 35086 44212 35138
rect 44156 35074 44212 35086
rect 43820 34914 43876 34926
rect 43820 34862 43822 34914
rect 43874 34862 43876 34914
rect 43596 34804 43652 34814
rect 43372 34692 43428 34702
rect 43372 34598 43428 34636
rect 42924 34412 43204 34468
rect 42588 33182 42590 33234
rect 42642 33182 42644 33234
rect 42588 33170 42644 33182
rect 42924 32900 42980 34412
rect 43372 34244 43428 34254
rect 43372 34150 43428 34188
rect 43596 33458 43652 34748
rect 43708 34802 43764 34814
rect 43708 34750 43710 34802
rect 43762 34750 43764 34802
rect 43708 33572 43764 34750
rect 43820 34580 43876 34862
rect 43820 34514 43876 34524
rect 43820 33572 43876 33582
rect 43708 33570 43876 33572
rect 43708 33518 43822 33570
rect 43874 33518 43876 33570
rect 43708 33516 43876 33518
rect 43820 33506 43876 33516
rect 43596 33406 43598 33458
rect 43650 33406 43652 33458
rect 43596 33394 43652 33406
rect 43484 33348 43540 33358
rect 43372 33346 43540 33348
rect 43372 33294 43486 33346
rect 43538 33294 43540 33346
rect 43372 33292 43540 33294
rect 43260 33124 43316 33134
rect 43372 33124 43428 33292
rect 43484 33282 43540 33292
rect 43260 33122 43428 33124
rect 43260 33070 43262 33122
rect 43314 33070 43428 33122
rect 43260 33068 43428 33070
rect 43260 33058 43316 33068
rect 42924 32834 42980 32844
rect 43260 32676 43316 32686
rect 43260 32582 43316 32620
rect 43036 32564 43092 32574
rect 42700 32562 43092 32564
rect 42700 32510 43038 32562
rect 43090 32510 43092 32562
rect 42700 32508 43092 32510
rect 42700 32450 42756 32508
rect 43036 32498 43092 32508
rect 42700 32398 42702 32450
rect 42754 32398 42756 32450
rect 42700 31556 42756 32398
rect 43148 32452 43204 32462
rect 43148 32358 43204 32396
rect 42476 30770 42532 30782
rect 42476 30718 42478 30770
rect 42530 30718 42532 30770
rect 42476 30212 42532 30718
rect 42700 30436 42756 31500
rect 43260 31668 43316 31678
rect 43260 30994 43316 31612
rect 43372 31220 43428 33068
rect 43372 31154 43428 31164
rect 43484 32674 43540 32686
rect 43484 32622 43486 32674
rect 43538 32622 43540 32674
rect 43484 31106 43540 32622
rect 44044 31892 44100 31902
rect 44044 31798 44100 31836
rect 44380 31668 44436 36204
rect 44044 31612 44436 31668
rect 44492 31668 44548 36428
rect 44604 34244 44660 37438
rect 44716 36260 44772 40124
rect 44828 39508 44884 40236
rect 45388 39620 45444 39630
rect 45388 39526 45444 39564
rect 44828 39442 44884 39452
rect 45164 38836 45220 38846
rect 45164 38742 45220 38780
rect 45500 38388 45556 40348
rect 45612 40180 45668 40190
rect 45612 39730 45668 40124
rect 45612 39678 45614 39730
rect 45666 39678 45668 39730
rect 45612 39666 45668 39678
rect 45724 40068 45780 40078
rect 45724 39508 45780 40012
rect 45612 39452 45780 39508
rect 45612 39058 45668 39452
rect 45612 39006 45614 39058
rect 45666 39006 45668 39058
rect 45612 38836 45668 39006
rect 45724 39284 45780 39294
rect 45724 39058 45780 39228
rect 45836 39172 45892 40350
rect 46172 40514 46228 40526
rect 46172 40462 46174 40514
rect 46226 40462 46228 40514
rect 46172 40068 46228 40462
rect 46172 40002 46228 40012
rect 46060 39620 46116 39630
rect 46284 39620 46340 39630
rect 46060 39618 46340 39620
rect 46060 39566 46062 39618
rect 46114 39566 46286 39618
rect 46338 39566 46340 39618
rect 46060 39564 46340 39566
rect 46060 39554 46116 39564
rect 46284 39554 46340 39564
rect 46284 39172 46340 39182
rect 45836 39116 46228 39172
rect 45724 39006 45726 39058
rect 45778 39006 45780 39058
rect 45724 38994 45780 39006
rect 45612 38770 45668 38780
rect 45836 38948 45892 38958
rect 45836 38834 45892 38892
rect 45836 38782 45838 38834
rect 45890 38782 45892 38834
rect 45836 38770 45892 38782
rect 45948 38836 46004 38846
rect 45724 38724 45780 38734
rect 45500 38322 45556 38332
rect 45612 38612 45780 38668
rect 44828 38164 44884 38174
rect 44828 38050 44884 38108
rect 45052 38164 45108 38174
rect 45052 38070 45108 38108
rect 44828 37998 44830 38050
rect 44882 37998 44884 38050
rect 44828 37378 44884 37998
rect 45276 38050 45332 38062
rect 45276 37998 45278 38050
rect 45330 37998 45332 38050
rect 44940 37940 44996 37950
rect 45276 37940 45332 37998
rect 44940 37846 44996 37884
rect 45052 37884 45332 37940
rect 45388 38050 45444 38062
rect 45388 37998 45390 38050
rect 45442 37998 45444 38050
rect 45388 37940 45444 37998
rect 44828 37326 44830 37378
rect 44882 37326 44884 37378
rect 44828 37314 44884 37326
rect 45052 37156 45108 37884
rect 45388 37874 45444 37884
rect 45500 38052 45556 38062
rect 45052 37090 45108 37100
rect 45164 37266 45220 37278
rect 45388 37268 45444 37278
rect 45164 37214 45166 37266
rect 45218 37214 45220 37266
rect 45164 36484 45220 37214
rect 45164 36418 45220 36428
rect 45276 37266 45444 37268
rect 45276 37214 45390 37266
rect 45442 37214 45444 37266
rect 45276 37212 45444 37214
rect 44828 36370 44884 36382
rect 44828 36318 44830 36370
rect 44882 36318 44884 36370
rect 44828 36260 44884 36318
rect 45164 36260 45220 36270
rect 45276 36260 45332 37212
rect 45388 37202 45444 37212
rect 45500 36706 45556 37996
rect 45612 37380 45668 38612
rect 45836 38050 45892 38062
rect 45836 37998 45838 38050
rect 45890 37998 45892 38050
rect 45724 37380 45780 37390
rect 45612 37378 45780 37380
rect 45612 37326 45726 37378
rect 45778 37326 45780 37378
rect 45612 37324 45780 37326
rect 45724 37314 45780 37324
rect 45612 37156 45668 37166
rect 45836 37156 45892 37998
rect 45612 37154 45892 37156
rect 45612 37102 45614 37154
rect 45666 37102 45892 37154
rect 45612 37100 45892 37102
rect 45612 37090 45668 37100
rect 45500 36654 45502 36706
rect 45554 36654 45556 36706
rect 45500 36642 45556 36654
rect 45836 36484 45892 36494
rect 45948 36484 46004 38780
rect 46172 38668 46228 39116
rect 46284 39058 46340 39116
rect 46284 39006 46286 39058
rect 46338 39006 46340 39058
rect 46284 38994 46340 39006
rect 46396 38668 46452 42812
rect 47404 42530 47460 42542
rect 47404 42478 47406 42530
rect 47458 42478 47460 42530
rect 47404 42308 47460 42478
rect 47404 42242 47460 42252
rect 47740 42530 47796 42924
rect 47740 42478 47742 42530
rect 47794 42478 47796 42530
rect 46732 41860 46788 41870
rect 46732 41766 46788 41804
rect 47180 41860 47236 41870
rect 47180 41858 47460 41860
rect 47180 41806 47182 41858
rect 47234 41806 47460 41858
rect 47180 41804 47460 41806
rect 47180 41794 47236 41804
rect 47292 41076 47348 41086
rect 46620 41074 47348 41076
rect 46620 41022 47294 41074
rect 47346 41022 47348 41074
rect 46620 41020 47348 41022
rect 46508 40628 46564 40638
rect 46508 40534 46564 40572
rect 46508 39396 46564 39406
rect 46508 38946 46564 39340
rect 46620 39394 46676 41020
rect 47292 41010 47348 41020
rect 46844 40740 46900 40750
rect 46844 40626 46900 40684
rect 47404 40740 47460 41804
rect 47740 41636 47796 42478
rect 47740 41570 47796 41580
rect 48636 41300 48692 43484
rect 48860 43446 48916 43484
rect 49532 43428 49588 43438
rect 49196 43426 49588 43428
rect 49196 43374 49534 43426
rect 49586 43374 49588 43426
rect 49196 43372 49588 43374
rect 48860 42754 48916 42766
rect 48860 42702 48862 42754
rect 48914 42702 48916 42754
rect 48748 42308 48804 42318
rect 48860 42308 48916 42702
rect 49084 42756 49140 42766
rect 49084 42662 49140 42700
rect 48804 42252 48916 42308
rect 48748 42242 48804 42252
rect 48076 41298 48692 41300
rect 48076 41246 48638 41298
rect 48690 41246 48692 41298
rect 48076 41244 48692 41246
rect 48076 41186 48132 41244
rect 48636 41234 48692 41244
rect 48748 41858 48804 41870
rect 48748 41806 48750 41858
rect 48802 41806 48804 41858
rect 48076 41134 48078 41186
rect 48130 41134 48132 41186
rect 48076 41122 48132 41134
rect 47460 40684 47684 40740
rect 47404 40674 47460 40684
rect 46844 40574 46846 40626
rect 46898 40574 46900 40626
rect 46844 40562 46900 40574
rect 47628 40626 47684 40684
rect 47628 40574 47630 40626
rect 47682 40574 47684 40626
rect 47628 40562 47684 40574
rect 47180 40514 47236 40526
rect 47180 40462 47182 40514
rect 47234 40462 47236 40514
rect 46732 39620 46788 39630
rect 46732 39526 46788 39564
rect 46844 39618 46900 39630
rect 46844 39566 46846 39618
rect 46898 39566 46900 39618
rect 46620 39342 46622 39394
rect 46674 39342 46676 39394
rect 46620 39330 46676 39342
rect 46844 39284 46900 39566
rect 46844 39218 46900 39228
rect 46956 39508 47012 39518
rect 46956 39060 47012 39452
rect 47180 39284 47236 40462
rect 48076 40404 48132 40414
rect 47180 39218 47236 39228
rect 47404 40180 47460 40190
rect 46508 38894 46510 38946
rect 46562 38894 46564 38946
rect 46508 38882 46564 38894
rect 46620 39004 47012 39060
rect 46172 38612 46340 38668
rect 46396 38612 46564 38668
rect 45836 36482 46004 36484
rect 45836 36430 45838 36482
rect 45890 36430 46004 36482
rect 45836 36428 46004 36430
rect 46060 38164 46116 38174
rect 46060 37828 46116 38108
rect 46172 37828 46228 37838
rect 46060 37826 46228 37828
rect 46060 37774 46174 37826
rect 46226 37774 46228 37826
rect 46060 37772 46228 37774
rect 44772 36204 44884 36260
rect 44940 36258 45332 36260
rect 44940 36206 45166 36258
rect 45218 36206 45332 36258
rect 44940 36204 45332 36206
rect 45612 36260 45668 36270
rect 44716 36194 44772 36204
rect 44716 35810 44772 35822
rect 44716 35758 44718 35810
rect 44770 35758 44772 35810
rect 44716 35476 44772 35758
rect 44716 35410 44772 35420
rect 44940 35698 44996 36204
rect 45164 36194 45220 36204
rect 45612 36166 45668 36204
rect 45164 35924 45220 35934
rect 45164 35830 45220 35868
rect 44940 35646 44942 35698
rect 44994 35646 44996 35698
rect 44828 34804 44884 34814
rect 44828 34710 44884 34748
rect 44940 34580 44996 35646
rect 45724 35700 45780 35710
rect 45052 35586 45108 35598
rect 45052 35534 45054 35586
rect 45106 35534 45108 35586
rect 45052 34914 45108 35534
rect 45500 35588 45556 35598
rect 45276 35026 45332 35038
rect 45276 34974 45278 35026
rect 45330 34974 45332 35026
rect 45052 34862 45054 34914
rect 45106 34862 45108 34914
rect 45052 34850 45108 34862
rect 45164 34916 45220 34926
rect 45276 34916 45332 34974
rect 45220 34860 45332 34916
rect 45388 34916 45444 34926
rect 45164 34850 45220 34860
rect 44940 34514 44996 34524
rect 44604 34188 45108 34244
rect 45052 32786 45108 34188
rect 45388 34020 45444 34860
rect 45500 34914 45556 35532
rect 45612 35586 45668 35598
rect 45612 35534 45614 35586
rect 45666 35534 45668 35586
rect 45612 35476 45668 35534
rect 45612 35410 45668 35420
rect 45500 34862 45502 34914
rect 45554 34862 45556 34914
rect 45500 34356 45556 34862
rect 45724 34914 45780 35644
rect 45724 34862 45726 34914
rect 45778 34862 45780 34914
rect 45724 34850 45780 34862
rect 45500 34290 45556 34300
rect 45612 34690 45668 34702
rect 45612 34638 45614 34690
rect 45666 34638 45668 34690
rect 45612 34244 45668 34638
rect 45612 34178 45668 34188
rect 45500 34020 45556 34030
rect 45836 34020 45892 36428
rect 45948 35588 46004 35598
rect 46060 35588 46116 37772
rect 46172 37762 46228 37772
rect 46172 36484 46228 36494
rect 46172 36390 46228 36428
rect 46004 35532 46116 35588
rect 46172 35700 46228 35710
rect 45948 35522 46004 35532
rect 46172 35138 46228 35644
rect 46172 35086 46174 35138
rect 46226 35086 46228 35138
rect 46172 35074 46228 35086
rect 46060 34916 46116 34926
rect 46060 34822 46116 34860
rect 45388 34018 45556 34020
rect 45388 33966 45502 34018
rect 45554 33966 45556 34018
rect 45388 33964 45556 33966
rect 45052 32734 45054 32786
rect 45106 32734 45108 32786
rect 45052 32722 45108 32734
rect 45388 33124 45444 33134
rect 45388 32786 45444 33068
rect 45388 32734 45390 32786
rect 45442 32734 45444 32786
rect 45388 32722 45444 32734
rect 45276 32674 45332 32686
rect 45276 32622 45278 32674
rect 45330 32622 45332 32674
rect 44828 32564 44884 32574
rect 44828 32470 44884 32508
rect 43484 31054 43486 31106
rect 43538 31054 43540 31106
rect 43484 31042 43540 31054
rect 43596 31106 43652 31118
rect 43596 31054 43598 31106
rect 43650 31054 43652 31106
rect 43260 30942 43262 30994
rect 43314 30942 43316 30994
rect 43260 30930 43316 30942
rect 43596 30996 43652 31054
rect 43596 30930 43652 30940
rect 43932 31106 43988 31118
rect 43932 31054 43934 31106
rect 43986 31054 43988 31106
rect 43932 30660 43988 31054
rect 43932 30594 43988 30604
rect 42644 30380 42756 30436
rect 42644 30212 42700 30380
rect 43148 30212 43204 30222
rect 42644 30156 42756 30212
rect 42476 28644 42532 30156
rect 42700 29988 42756 30156
rect 43148 30118 43204 30156
rect 42812 29988 42868 29998
rect 42700 29986 42868 29988
rect 42700 29934 42814 29986
rect 42866 29934 42868 29986
rect 42700 29932 42868 29934
rect 42588 28644 42644 28654
rect 42476 28642 42644 28644
rect 42476 28590 42590 28642
rect 42642 28590 42644 28642
rect 42476 28588 42644 28590
rect 42364 28578 42420 28588
rect 42588 28578 42644 28588
rect 41692 28082 41972 28084
rect 41692 28030 41694 28082
rect 41746 28030 41972 28082
rect 41692 28028 41972 28030
rect 41692 28018 41748 28028
rect 41804 27860 41860 27870
rect 41580 27858 41860 27860
rect 41580 27806 41806 27858
rect 41858 27806 41860 27858
rect 41580 27804 41860 27806
rect 41804 27794 41860 27804
rect 41916 27858 41972 27870
rect 41916 27806 41918 27858
rect 41970 27806 41972 27858
rect 40908 27134 40910 27186
rect 40962 27134 40964 27186
rect 40908 27122 40964 27134
rect 41916 27188 41972 27806
rect 41916 27122 41972 27132
rect 42028 27748 42084 27758
rect 41692 27074 41748 27086
rect 41692 27022 41694 27074
rect 41746 27022 41748 27074
rect 41692 26908 41748 27022
rect 42028 26908 42084 27692
rect 41692 26852 42084 26908
rect 42140 27746 42196 27758
rect 42140 27694 42142 27746
rect 42194 27694 42196 27746
rect 41916 26514 41972 26852
rect 42140 26628 42196 27694
rect 42364 27634 42420 27646
rect 42364 27582 42366 27634
rect 42418 27582 42420 27634
rect 42364 27186 42420 27582
rect 42364 27134 42366 27186
rect 42418 27134 42420 27186
rect 42364 27122 42420 27134
rect 42252 27074 42308 27086
rect 42252 27022 42254 27074
rect 42306 27022 42308 27074
rect 42252 26964 42308 27022
rect 42476 27076 42532 27086
rect 42364 26964 42420 26974
rect 42252 26908 42364 26964
rect 42364 26898 42420 26908
rect 42476 26962 42532 27020
rect 42476 26910 42478 26962
rect 42530 26910 42532 26962
rect 42140 26562 42196 26572
rect 41916 26462 41918 26514
rect 41970 26462 41972 26514
rect 41916 26450 41972 26462
rect 40796 26002 40852 26012
rect 40908 26290 40964 26302
rect 40908 26238 40910 26290
rect 40962 26238 40964 26290
rect 40572 25620 40628 25630
rect 40908 25620 40964 26238
rect 40572 25618 40964 25620
rect 40572 25566 40574 25618
rect 40626 25566 40964 25618
rect 40572 25564 40964 25566
rect 41020 26292 41076 26302
rect 40572 25060 40628 25564
rect 41020 25396 41076 26236
rect 40572 24994 40628 25004
rect 40796 25394 41076 25396
rect 40796 25342 41022 25394
rect 41074 25342 41076 25394
rect 40796 25340 41076 25342
rect 40460 23650 40516 23660
rect 40572 24164 40628 24174
rect 40796 24164 40852 25340
rect 41020 25330 41076 25340
rect 41356 26178 41412 26190
rect 41356 26126 41358 26178
rect 41410 26126 41412 26178
rect 41020 24948 41076 24958
rect 41020 24854 41076 24892
rect 41132 24948 41188 24958
rect 41356 24948 41412 26126
rect 42476 25618 42532 26910
rect 42476 25566 42478 25618
rect 42530 25566 42532 25618
rect 41916 25508 41972 25518
rect 41804 25506 41972 25508
rect 41804 25454 41918 25506
rect 41970 25454 41972 25506
rect 41804 25452 41972 25454
rect 41692 25396 41748 25406
rect 41692 25302 41748 25340
rect 41132 24946 41412 24948
rect 41132 24894 41134 24946
rect 41186 24894 41412 24946
rect 41132 24892 41412 24894
rect 41132 24882 41188 24892
rect 40908 24724 40964 24734
rect 40908 24630 40964 24668
rect 41356 24164 41412 24892
rect 41804 25172 41860 25452
rect 41916 25442 41972 25452
rect 42364 25506 42420 25518
rect 42364 25454 42366 25506
rect 42418 25454 42420 25506
rect 40796 24108 40964 24164
rect 40348 22430 40350 22482
rect 40402 22430 40404 22482
rect 40348 22418 40404 22430
rect 40572 22372 40628 24108
rect 40796 23940 40852 23950
rect 40796 23846 40852 23884
rect 40684 23828 40740 23838
rect 40684 23734 40740 23772
rect 40460 22370 40628 22372
rect 40460 22318 40574 22370
rect 40626 22318 40628 22370
rect 40460 22316 40628 22318
rect 40348 22258 40404 22270
rect 40348 22206 40350 22258
rect 40402 22206 40404 22258
rect 40348 21924 40404 22206
rect 40348 21858 40404 21868
rect 40348 21700 40404 21710
rect 40460 21700 40516 22316
rect 40572 22306 40628 22316
rect 40796 22372 40852 22382
rect 40796 22278 40852 22316
rect 40348 21698 40516 21700
rect 40348 21646 40350 21698
rect 40402 21646 40516 21698
rect 40348 21644 40516 21646
rect 40908 21698 40964 24108
rect 41356 24098 41412 24108
rect 41468 24722 41524 24734
rect 41468 24670 41470 24722
rect 41522 24670 41524 24722
rect 41356 23938 41412 23950
rect 41356 23886 41358 23938
rect 41410 23886 41412 23938
rect 41356 23828 41412 23886
rect 41356 23762 41412 23772
rect 41356 23380 41412 23390
rect 41468 23380 41524 24670
rect 41804 24162 41860 25116
rect 41916 25282 41972 25294
rect 41916 25230 41918 25282
rect 41970 25230 41972 25282
rect 41916 25060 41972 25230
rect 41916 25004 42084 25060
rect 41804 24110 41806 24162
rect 41858 24110 41860 24162
rect 41804 24098 41860 24110
rect 41916 24724 41972 24734
rect 42028 24724 42084 25004
rect 42252 24724 42308 24734
rect 42028 24722 42308 24724
rect 42028 24670 42254 24722
rect 42306 24670 42308 24722
rect 42028 24668 42308 24670
rect 41916 24610 41972 24668
rect 42252 24658 42308 24668
rect 41916 24558 41918 24610
rect 41970 24558 41972 24610
rect 41804 23940 41860 23950
rect 41804 23846 41860 23884
rect 41916 23604 41972 24558
rect 42252 24164 42308 24174
rect 42252 23938 42308 24108
rect 42252 23886 42254 23938
rect 42306 23886 42308 23938
rect 42252 23874 42308 23886
rect 42364 23940 42420 25454
rect 42476 25396 42532 25566
rect 42476 25330 42532 25340
rect 42700 24724 42756 29932
rect 42812 29922 42868 29932
rect 43484 29988 43540 29998
rect 43372 28644 43428 28654
rect 43372 28550 43428 28588
rect 42924 28418 42980 28430
rect 43484 28420 43540 29932
rect 43708 29316 43764 29326
rect 43708 29222 43764 29260
rect 43932 28644 43988 28654
rect 44044 28644 44100 31612
rect 44492 31602 44548 31612
rect 44940 31554 44996 31566
rect 44940 31502 44942 31554
rect 44994 31502 44996 31554
rect 44268 31276 44884 31332
rect 44156 30996 44212 31006
rect 44156 30902 44212 30940
rect 44268 30994 44324 31276
rect 44268 30942 44270 30994
rect 44322 30942 44324 30994
rect 44268 30930 44324 30942
rect 44716 31106 44772 31118
rect 44716 31054 44718 31106
rect 44770 31054 44772 31106
rect 44716 30996 44772 31054
rect 44716 30930 44772 30940
rect 44828 30994 44884 31276
rect 44940 31108 44996 31502
rect 44940 31042 44996 31052
rect 44828 30942 44830 30994
rect 44882 30942 44884 30994
rect 44716 30770 44772 30782
rect 44716 30718 44718 30770
rect 44770 30718 44772 30770
rect 44716 30660 44772 30718
rect 44716 29988 44772 30604
rect 44716 29922 44772 29932
rect 44828 29652 44884 30942
rect 45276 30548 45332 32622
rect 45500 32340 45556 33964
rect 45612 33964 45892 34020
rect 45948 34692 46004 34702
rect 45948 34018 46004 34636
rect 45948 33966 45950 34018
rect 46002 33966 46004 34018
rect 45612 32562 45668 33964
rect 45948 33908 46004 33966
rect 45948 33852 46228 33908
rect 46172 33460 46228 33852
rect 46284 33796 46340 38612
rect 46508 36708 46564 38612
rect 46620 38610 46676 39004
rect 46732 38836 46788 38846
rect 46732 38668 46788 38780
rect 46844 38836 46900 38846
rect 47068 38836 47124 38846
rect 46844 38834 47068 38836
rect 46844 38782 46846 38834
rect 46898 38782 47068 38834
rect 46844 38780 47068 38782
rect 46844 38770 46900 38780
rect 47068 38722 47124 38780
rect 47068 38670 47070 38722
rect 47122 38670 47124 38722
rect 46732 38612 47012 38668
rect 47068 38658 47124 38670
rect 47404 38834 47460 40124
rect 48076 39620 48132 40348
rect 48076 39554 48132 39564
rect 48188 39730 48244 39742
rect 48748 39732 48804 41806
rect 48972 41188 49028 41198
rect 48972 41094 49028 41132
rect 49196 40626 49252 43372
rect 49532 43362 49588 43372
rect 49868 43428 49924 43438
rect 49868 42756 49924 43372
rect 49868 42662 49924 42700
rect 49308 42644 49364 42654
rect 49308 42550 49364 42588
rect 49756 42644 49812 42654
rect 49420 41970 49476 41982
rect 49420 41918 49422 41970
rect 49474 41918 49476 41970
rect 49420 41860 49476 41918
rect 49756 41970 49812 42588
rect 49756 41918 49758 41970
rect 49810 41918 49812 41970
rect 49756 41906 49812 41918
rect 49420 41794 49476 41804
rect 49756 41636 49812 41646
rect 49756 41076 49812 41580
rect 49868 41412 49924 41422
rect 49980 41412 50036 43596
rect 52108 43652 52164 43662
rect 52108 43558 52164 43596
rect 51996 43538 52052 43550
rect 51996 43486 51998 43538
rect 52050 43486 52052 43538
rect 51660 43428 51716 43438
rect 51660 43334 51716 43372
rect 50540 42980 50596 42990
rect 50540 42866 50596 42924
rect 50540 42814 50542 42866
rect 50594 42814 50596 42866
rect 50540 42802 50596 42814
rect 51996 42868 52052 43486
rect 51996 42802 52052 42812
rect 52108 43314 52164 43326
rect 52108 43262 52110 43314
rect 52162 43262 52164 43314
rect 50764 42754 50820 42766
rect 50764 42702 50766 42754
rect 50818 42702 50820 42754
rect 50204 42532 50260 42542
rect 50764 42532 50820 42702
rect 49868 41410 50036 41412
rect 49868 41358 49870 41410
rect 49922 41358 50036 41410
rect 49868 41356 50036 41358
rect 50092 42530 50820 42532
rect 50092 42478 50206 42530
rect 50258 42478 50820 42530
rect 50092 42476 50820 42478
rect 50988 42644 51044 42654
rect 49868 41346 49924 41356
rect 49868 41076 49924 41086
rect 49756 41074 49924 41076
rect 49756 41022 49870 41074
rect 49922 41022 49924 41074
rect 49756 41020 49924 41022
rect 49868 41010 49924 41020
rect 49980 41076 50036 41086
rect 50092 41076 50148 42476
rect 50204 42466 50260 42476
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50764 41858 50820 41870
rect 50764 41806 50766 41858
rect 50818 41806 50820 41858
rect 50316 41188 50372 41198
rect 50540 41188 50596 41198
rect 50316 41094 50372 41132
rect 50428 41186 50596 41188
rect 50428 41134 50542 41186
rect 50594 41134 50596 41186
rect 50428 41132 50596 41134
rect 49980 41074 50148 41076
rect 49980 41022 49982 41074
rect 50034 41022 50148 41074
rect 49980 41020 50148 41022
rect 49980 41010 50036 41020
rect 49532 40964 49588 40974
rect 49196 40574 49198 40626
rect 49250 40574 49252 40626
rect 49196 40562 49252 40574
rect 49420 40962 49588 40964
rect 49420 40910 49534 40962
rect 49586 40910 49588 40962
rect 49420 40908 49588 40910
rect 49420 40628 49476 40908
rect 49532 40898 49588 40908
rect 48188 39678 48190 39730
rect 48242 39678 48244 39730
rect 47516 39396 47572 39406
rect 47516 39394 47796 39396
rect 47516 39342 47518 39394
rect 47570 39342 47796 39394
rect 47516 39340 47796 39342
rect 47516 39330 47572 39340
rect 47404 38782 47406 38834
rect 47458 38782 47460 38834
rect 47404 38668 47460 38782
rect 47740 39172 47796 39340
rect 47628 38724 47684 38762
rect 47404 38612 47572 38668
rect 47628 38658 47684 38668
rect 46620 38558 46622 38610
rect 46674 38558 46676 38610
rect 46620 38546 46676 38558
rect 46956 38500 47012 38612
rect 46956 38444 47124 38500
rect 46620 38388 46676 38398
rect 46620 38050 46676 38332
rect 46620 37998 46622 38050
rect 46674 37998 46676 38050
rect 46620 37156 46676 37998
rect 47068 37826 47124 38444
rect 47516 38052 47572 38612
rect 47628 38052 47684 38062
rect 47516 38050 47684 38052
rect 47516 37998 47630 38050
rect 47682 37998 47684 38050
rect 47516 37996 47684 37998
rect 47628 37986 47684 37996
rect 47068 37774 47070 37826
rect 47122 37774 47124 37826
rect 47068 37380 47124 37774
rect 47628 37492 47684 37530
rect 47628 37426 47684 37436
rect 46620 37090 46676 37100
rect 46956 37324 47124 37380
rect 46508 36370 46564 36652
rect 46956 36484 47012 37324
rect 47628 37268 47684 37278
rect 47404 37212 47628 37268
rect 47068 37154 47124 37166
rect 47068 37102 47070 37154
rect 47122 37102 47124 37154
rect 47068 37042 47124 37102
rect 47068 36990 47070 37042
rect 47122 36990 47124 37042
rect 47068 36978 47124 36990
rect 46956 36418 47012 36428
rect 47068 36820 47124 36830
rect 46508 36318 46510 36370
rect 46562 36318 46564 36370
rect 46508 36306 46564 36318
rect 46732 36260 46788 36270
rect 46788 36204 47012 36260
rect 46732 36194 46788 36204
rect 46732 35700 46788 35710
rect 46732 35606 46788 35644
rect 46620 34804 46676 34814
rect 46620 34710 46676 34748
rect 46956 34354 47012 36204
rect 47068 35698 47124 36764
rect 47068 35646 47070 35698
rect 47122 35646 47124 35698
rect 47068 35588 47124 35646
rect 47292 36482 47348 36494
rect 47292 36430 47294 36482
rect 47346 36430 47348 36482
rect 47292 35700 47348 36430
rect 47292 35634 47348 35644
rect 47068 35522 47124 35532
rect 46956 34302 46958 34354
rect 47010 34302 47012 34354
rect 46956 34290 47012 34302
rect 46732 34132 46788 34142
rect 46732 34038 46788 34076
rect 47180 34130 47236 34142
rect 47180 34078 47182 34130
rect 47234 34078 47236 34130
rect 47068 34018 47124 34030
rect 47068 33966 47070 34018
rect 47122 33966 47124 34018
rect 46284 33740 46788 33796
rect 46172 33404 46452 33460
rect 46060 33348 46116 33358
rect 45836 33234 45892 33246
rect 45836 33182 45838 33234
rect 45890 33182 45892 33234
rect 45836 33124 45892 33182
rect 46060 33234 46116 33292
rect 46060 33182 46062 33234
rect 46114 33182 46116 33234
rect 46060 33170 46116 33182
rect 45836 33058 45892 33068
rect 45948 33122 46004 33134
rect 45948 33070 45950 33122
rect 46002 33070 46004 33122
rect 45612 32510 45614 32562
rect 45666 32510 45668 32562
rect 45612 32498 45668 32510
rect 45724 32786 45780 32798
rect 45724 32734 45726 32786
rect 45778 32734 45780 32786
rect 45724 32564 45780 32734
rect 45724 32498 45780 32508
rect 45836 32340 45892 32350
rect 45500 32338 45892 32340
rect 45500 32286 45838 32338
rect 45890 32286 45892 32338
rect 45500 32284 45892 32286
rect 45836 32274 45892 32284
rect 45948 32004 46004 33070
rect 46396 32900 46452 33404
rect 46508 33236 46564 33246
rect 46508 33142 46564 33180
rect 46620 33124 46676 33134
rect 46620 33030 46676 33068
rect 46396 32844 46676 32900
rect 46060 32340 46116 32350
rect 46060 32246 46116 32284
rect 46284 32340 46340 32350
rect 46284 32338 46564 32340
rect 46284 32286 46286 32338
rect 46338 32286 46564 32338
rect 46284 32284 46564 32286
rect 46284 32274 46340 32284
rect 45500 31948 46452 32004
rect 45500 30994 45556 31948
rect 45500 30942 45502 30994
rect 45554 30942 45556 30994
rect 45500 30930 45556 30942
rect 45612 31780 45668 31790
rect 45276 30482 45332 30492
rect 45388 30770 45444 30782
rect 45388 30718 45390 30770
rect 45442 30718 45444 30770
rect 45388 30436 45444 30718
rect 45388 30370 45444 30380
rect 45500 30324 45556 30334
rect 44828 29586 44884 29596
rect 45052 30210 45108 30222
rect 45052 30158 45054 30210
rect 45106 30158 45108 30210
rect 45052 29876 45108 30158
rect 45164 30098 45220 30110
rect 45164 30046 45166 30098
rect 45218 30046 45220 30098
rect 45164 29988 45220 30046
rect 45164 29922 45220 29932
rect 45276 29986 45332 29998
rect 45276 29934 45278 29986
rect 45330 29934 45332 29986
rect 44156 29428 44212 29438
rect 44156 29334 44212 29372
rect 42924 28366 42926 28418
rect 42978 28366 42980 28418
rect 42924 27300 42980 28366
rect 43372 28364 43540 28420
rect 43820 28588 43932 28644
rect 43988 28588 44100 28644
rect 44940 28980 44996 28990
rect 43036 27858 43092 27870
rect 43036 27806 43038 27858
rect 43090 27806 43092 27858
rect 43036 27748 43092 27806
rect 43036 27682 43092 27692
rect 42924 27074 42980 27244
rect 42924 27022 42926 27074
rect 42978 27022 42980 27074
rect 42924 27010 42980 27022
rect 43036 27188 43092 27198
rect 42700 24658 42756 24668
rect 42812 26290 42868 26302
rect 42812 26238 42814 26290
rect 42866 26238 42868 26290
rect 42812 25956 42868 26238
rect 42812 24722 42868 25900
rect 43036 25508 43092 27132
rect 43148 26962 43204 26974
rect 43148 26910 43150 26962
rect 43202 26910 43204 26962
rect 43148 26292 43204 26910
rect 43260 26964 43316 27002
rect 43260 26898 43316 26908
rect 43148 26226 43204 26236
rect 43260 25618 43316 25630
rect 43260 25566 43262 25618
rect 43314 25566 43316 25618
rect 43148 25508 43204 25518
rect 43036 25452 43148 25508
rect 43148 25414 43204 25452
rect 42812 24670 42814 24722
rect 42866 24670 42868 24722
rect 42812 24658 42868 24670
rect 43260 24162 43316 25566
rect 43260 24110 43262 24162
rect 43314 24110 43316 24162
rect 43260 24098 43316 24110
rect 42364 23874 42420 23884
rect 42588 24050 42644 24062
rect 42588 23998 42590 24050
rect 42642 23998 42644 24050
rect 41916 23538 41972 23548
rect 41356 23378 41468 23380
rect 41356 23326 41358 23378
rect 41410 23326 41468 23378
rect 41356 23324 41468 23326
rect 41356 23314 41412 23324
rect 41468 23286 41524 23324
rect 42588 23378 42644 23998
rect 42588 23326 42590 23378
rect 42642 23326 42644 23378
rect 42588 23314 42644 23326
rect 42924 23940 42980 23950
rect 42028 23268 42084 23278
rect 42028 23174 42084 23212
rect 42924 23266 42980 23884
rect 42924 23214 42926 23266
rect 42978 23214 42980 23266
rect 42924 23202 42980 23214
rect 43036 23716 43092 23726
rect 41692 23154 41748 23166
rect 41692 23102 41694 23154
rect 41746 23102 41748 23154
rect 41692 22372 41748 23102
rect 41804 23156 41860 23166
rect 41804 23062 41860 23100
rect 42364 23154 42420 23166
rect 42364 23102 42366 23154
rect 42418 23102 42420 23154
rect 41692 22306 41748 22316
rect 41580 22258 41636 22270
rect 41580 22206 41582 22258
rect 41634 22206 41636 22258
rect 41580 21924 41636 22206
rect 42364 22148 42420 23102
rect 42588 22820 42644 22830
rect 42588 22482 42644 22764
rect 42588 22430 42590 22482
rect 42642 22430 42644 22482
rect 42588 22418 42644 22430
rect 42924 22148 42980 22158
rect 42364 22082 42420 22092
rect 42700 22146 42980 22148
rect 42700 22094 42926 22146
rect 42978 22094 42980 22146
rect 42700 22092 42980 22094
rect 41580 21858 41636 21868
rect 42476 21924 42532 21934
rect 42700 21924 42756 22092
rect 42924 22082 42980 22092
rect 43036 21924 43092 23660
rect 43372 22484 43428 28364
rect 43708 27746 43764 27758
rect 43708 27694 43710 27746
rect 43762 27694 43764 27746
rect 43708 27300 43764 27694
rect 43596 27244 43764 27300
rect 43484 26962 43540 26974
rect 43484 26910 43486 26962
rect 43538 26910 43540 26962
rect 43484 26404 43540 26910
rect 43596 26908 43652 27244
rect 43708 27076 43764 27086
rect 43820 27076 43876 28588
rect 43932 28550 43988 28588
rect 44828 27300 44884 27310
rect 44716 27244 44828 27300
rect 43708 27074 43876 27076
rect 43708 27022 43710 27074
rect 43762 27022 43876 27074
rect 43708 27020 43876 27022
rect 44156 27076 44212 27086
rect 43708 27010 43764 27020
rect 44156 26982 44212 27020
rect 44044 26962 44100 26974
rect 44044 26910 44046 26962
rect 44098 26910 44100 26962
rect 43596 26852 43876 26908
rect 43820 26516 43876 26852
rect 43820 26450 43876 26460
rect 43484 26338 43540 26348
rect 43932 26404 43988 26414
rect 43820 24052 43876 24062
rect 43820 23938 43876 23996
rect 43820 23886 43822 23938
rect 43874 23886 43876 23938
rect 43708 23826 43764 23838
rect 43708 23774 43710 23826
rect 43762 23774 43764 23826
rect 43708 23380 43764 23774
rect 42532 21868 42756 21924
rect 42924 21868 43092 21924
rect 43260 22428 43428 22484
rect 43484 23324 43764 23380
rect 43484 23268 43540 23324
rect 43260 21924 43316 22428
rect 43484 22372 43540 23212
rect 43708 23156 43764 23166
rect 43820 23156 43876 23886
rect 43932 23938 43988 26348
rect 44044 26290 44100 26910
rect 44716 26908 44772 27244
rect 44828 27234 44884 27244
rect 44828 27076 44884 27086
rect 44940 27076 44996 28924
rect 44828 27074 44996 27076
rect 44828 27022 44830 27074
rect 44882 27022 44996 27074
rect 44828 27020 44996 27022
rect 44828 27010 44884 27020
rect 44716 26852 44884 26908
rect 44044 26238 44046 26290
rect 44098 26238 44100 26290
rect 44044 26226 44100 26238
rect 44268 26628 44324 26638
rect 44268 24276 44324 26572
rect 44716 26628 44772 26638
rect 44716 26514 44772 26572
rect 44716 26462 44718 26514
rect 44770 26462 44772 26514
rect 44716 26450 44772 26462
rect 44380 26292 44436 26302
rect 44380 26198 44436 26236
rect 44828 25506 44884 26852
rect 44828 25454 44830 25506
rect 44882 25454 44884 25506
rect 44828 25442 44884 25454
rect 44716 25284 44772 25294
rect 44716 24946 44772 25228
rect 44716 24894 44718 24946
rect 44770 24894 44772 24946
rect 44716 24882 44772 24894
rect 44940 25172 44996 25182
rect 44940 24722 44996 25116
rect 45052 24836 45108 29820
rect 45164 29428 45220 29438
rect 45276 29428 45332 29934
rect 45164 29426 45332 29428
rect 45164 29374 45166 29426
rect 45218 29374 45332 29426
rect 45164 29372 45332 29374
rect 45164 29362 45220 29372
rect 45276 29204 45332 29214
rect 45500 29204 45556 30268
rect 45612 30210 45668 31724
rect 46284 31778 46340 31790
rect 46284 31726 46286 31778
rect 46338 31726 46340 31778
rect 45836 31666 45892 31678
rect 45836 31614 45838 31666
rect 45890 31614 45892 31666
rect 45836 31444 45892 31614
rect 45836 31378 45892 31388
rect 45836 31220 45892 31230
rect 45836 31106 45892 31164
rect 46284 31220 46340 31726
rect 46284 31154 46340 31164
rect 45836 31054 45838 31106
rect 45890 31054 45892 31106
rect 45836 31042 45892 31054
rect 46396 30994 46452 31948
rect 46396 30942 46398 30994
rect 46450 30942 46452 30994
rect 46396 30930 46452 30942
rect 45612 30158 45614 30210
rect 45666 30158 45668 30210
rect 45612 29764 45668 30158
rect 45724 30770 45780 30782
rect 45724 30718 45726 30770
rect 45778 30718 45780 30770
rect 45724 30548 45780 30718
rect 46284 30770 46340 30782
rect 46284 30718 46286 30770
rect 46338 30718 46340 30770
rect 46284 30548 46340 30718
rect 45724 30492 46340 30548
rect 46396 30548 46452 30558
rect 45724 29986 45780 30492
rect 45724 29934 45726 29986
rect 45778 29934 45780 29986
rect 45724 29922 45780 29934
rect 46284 30210 46340 30222
rect 46284 30158 46286 30210
rect 46338 30158 46340 30210
rect 45612 29708 46004 29764
rect 45836 29538 45892 29550
rect 45836 29486 45838 29538
rect 45890 29486 45892 29538
rect 45836 29316 45892 29486
rect 45836 29250 45892 29260
rect 45164 28642 45220 28654
rect 45164 28590 45166 28642
rect 45218 28590 45220 28642
rect 45164 27748 45220 28590
rect 45164 27682 45220 27692
rect 45276 25506 45332 29148
rect 45388 29148 45556 29204
rect 45388 26908 45444 29148
rect 45500 28980 45556 28990
rect 45948 28980 46004 29708
rect 46060 29426 46116 29438
rect 46060 29374 46062 29426
rect 46114 29374 46116 29426
rect 46060 29204 46116 29374
rect 46060 29138 46116 29148
rect 46284 28980 46340 30158
rect 46396 29764 46452 30492
rect 46508 30212 46564 32284
rect 46620 31108 46676 32844
rect 46620 31042 46676 31052
rect 46620 30770 46676 30782
rect 46620 30718 46622 30770
rect 46674 30718 46676 30770
rect 46620 30436 46676 30718
rect 46620 30370 46676 30380
rect 46732 30324 46788 33740
rect 46844 33348 46900 33358
rect 46844 33254 46900 33292
rect 47068 32562 47124 33966
rect 47180 33124 47236 34078
rect 47180 33058 47236 33068
rect 47404 32900 47460 37212
rect 47628 37202 47684 37212
rect 47516 37044 47572 37054
rect 47740 37044 47796 39116
rect 48188 39060 48244 39678
rect 48524 39676 48804 39732
rect 48524 39618 48580 39676
rect 48524 39566 48526 39618
rect 48578 39566 48580 39618
rect 48524 39554 48580 39566
rect 48748 39396 48804 39676
rect 48972 40402 49028 40414
rect 48972 40350 48974 40402
rect 49026 40350 49028 40402
rect 48972 39730 49028 40350
rect 49196 40404 49252 40414
rect 49420 40404 49476 40572
rect 49252 40348 49476 40404
rect 49532 40404 49588 40414
rect 49532 40402 49812 40404
rect 49532 40350 49534 40402
rect 49586 40350 49812 40402
rect 49532 40348 49812 40350
rect 49196 40310 49252 40348
rect 49532 40338 49588 40348
rect 48972 39678 48974 39730
rect 49026 39678 49028 39730
rect 48972 39666 49028 39678
rect 49756 39396 49812 40348
rect 49980 40290 50036 40302
rect 49980 40238 49982 40290
rect 50034 40238 50036 40290
rect 49980 40180 50036 40238
rect 49980 40114 50036 40124
rect 49868 39620 49924 39630
rect 49868 39526 49924 39564
rect 50092 39620 50148 41020
rect 49756 39340 50036 39396
rect 48524 39284 48580 39294
rect 48300 39060 48356 39070
rect 48188 39058 48356 39060
rect 48188 39006 48302 39058
rect 48354 39006 48356 39058
rect 48188 39004 48356 39006
rect 48300 38994 48356 39004
rect 48076 38948 48132 38958
rect 48076 38854 48132 38892
rect 47964 38836 48020 38846
rect 47964 38742 48020 38780
rect 48524 38724 48580 39228
rect 48748 38948 48804 39340
rect 49868 39060 49924 39070
rect 48748 38882 48804 38892
rect 49196 39004 49700 39060
rect 49196 38946 49252 39004
rect 49196 38894 49198 38946
rect 49250 38894 49252 38946
rect 49196 38882 49252 38894
rect 49308 38836 49364 38846
rect 49308 38742 49364 38780
rect 49532 38836 49588 38846
rect 48188 37268 48244 37278
rect 48524 37268 48580 38668
rect 48188 37266 48468 37268
rect 48188 37214 48190 37266
rect 48242 37214 48468 37266
rect 48188 37212 48468 37214
rect 48188 37202 48244 37212
rect 47516 37042 47796 37044
rect 47516 36990 47518 37042
rect 47570 36990 47796 37042
rect 47516 36988 47796 36990
rect 47852 37044 47908 37054
rect 48188 37044 48244 37054
rect 47852 37042 48020 37044
rect 47852 36990 47854 37042
rect 47906 36990 48020 37042
rect 47852 36988 48020 36990
rect 47516 36484 47572 36988
rect 47852 36978 47908 36988
rect 47628 36820 47684 36830
rect 47628 36594 47684 36764
rect 47628 36542 47630 36594
rect 47682 36542 47684 36594
rect 47628 36530 47684 36542
rect 47740 36706 47796 36718
rect 47740 36654 47742 36706
rect 47794 36654 47796 36706
rect 47516 34468 47572 36428
rect 47740 36036 47796 36654
rect 47516 34402 47572 34412
rect 47628 35980 47740 36036
rect 47628 34244 47684 35980
rect 47740 35970 47796 35980
rect 47852 36260 47908 36270
rect 47740 35812 47796 35822
rect 47740 35698 47796 35756
rect 47852 35810 47908 36204
rect 47852 35758 47854 35810
rect 47906 35758 47908 35810
rect 47852 35746 47908 35758
rect 47740 35646 47742 35698
rect 47794 35646 47796 35698
rect 47740 35634 47796 35646
rect 47852 35588 47908 35598
rect 47852 34914 47908 35532
rect 47852 34862 47854 34914
rect 47906 34862 47908 34914
rect 47852 34850 47908 34862
rect 47964 34354 48020 36988
rect 48188 36950 48244 36988
rect 48076 36484 48132 36494
rect 48076 36390 48132 36428
rect 48188 36372 48244 36382
rect 48076 36148 48132 36158
rect 48076 35922 48132 36092
rect 48076 35870 48078 35922
rect 48130 35870 48132 35922
rect 48076 35858 48132 35870
rect 48188 35810 48244 36316
rect 48188 35758 48190 35810
rect 48242 35758 48244 35810
rect 48188 35746 48244 35758
rect 48076 35700 48132 35710
rect 48076 35308 48132 35644
rect 48076 35252 48356 35308
rect 47964 34302 47966 34354
rect 48018 34302 48020 34354
rect 47964 34290 48020 34302
rect 47852 34244 47908 34254
rect 47628 34242 47908 34244
rect 47628 34190 47854 34242
rect 47906 34190 47908 34242
rect 47628 34188 47908 34190
rect 47852 34178 47908 34188
rect 48076 34244 48132 34254
rect 48076 34150 48132 34188
rect 47516 34132 47572 34142
rect 47516 34038 47572 34076
rect 47068 32510 47070 32562
rect 47122 32510 47124 32562
rect 47068 32498 47124 32510
rect 47292 32844 47460 32900
rect 46956 32452 47012 32462
rect 46732 30258 46788 30268
rect 46844 32396 46956 32452
rect 46508 30156 46676 30212
rect 46620 29988 46676 30156
rect 46844 30210 46900 32396
rect 46956 32386 47012 32396
rect 47180 32004 47236 32014
rect 47068 31948 47180 32004
rect 46956 31890 47012 31902
rect 46956 31838 46958 31890
rect 47010 31838 47012 31890
rect 46956 31780 47012 31838
rect 46956 31714 47012 31724
rect 46956 31554 47012 31566
rect 46956 31502 46958 31554
rect 47010 31502 47012 31554
rect 46956 30884 47012 31502
rect 47068 31218 47124 31948
rect 47180 31938 47236 31948
rect 47068 31166 47070 31218
rect 47122 31166 47124 31218
rect 47068 31154 47124 31166
rect 47180 31666 47236 31678
rect 47180 31614 47182 31666
rect 47234 31614 47236 31666
rect 46956 30818 47012 30828
rect 46844 30158 46846 30210
rect 46898 30158 46900 30210
rect 46844 30146 46900 30158
rect 46956 30098 47012 30110
rect 46956 30046 46958 30098
rect 47010 30046 47012 30098
rect 46956 29988 47012 30046
rect 46620 29932 47012 29988
rect 46396 29708 46788 29764
rect 46508 29538 46564 29550
rect 46508 29486 46510 29538
rect 46562 29486 46564 29538
rect 46508 29428 46564 29486
rect 46508 29362 46564 29372
rect 46620 29426 46676 29438
rect 46620 29374 46622 29426
rect 46674 29374 46676 29426
rect 45948 28924 46228 28980
rect 46284 28924 46452 28980
rect 45500 28754 45556 28924
rect 45724 28868 45780 28878
rect 45500 28702 45502 28754
rect 45554 28702 45556 28754
rect 45500 28690 45556 28702
rect 45612 28812 45724 28868
rect 45612 28754 45668 28812
rect 45724 28802 45780 28812
rect 46172 28866 46228 28924
rect 46172 28814 46174 28866
rect 46226 28814 46228 28866
rect 46172 28802 46228 28814
rect 45612 28702 45614 28754
rect 45666 28702 45668 28754
rect 45612 28690 45668 28702
rect 46284 28756 46340 28766
rect 45948 28644 46004 28654
rect 46284 28644 46340 28700
rect 45948 28642 46340 28644
rect 45948 28590 45950 28642
rect 46002 28590 46340 28642
rect 45948 28588 46340 28590
rect 45948 28578 46004 28588
rect 45948 28308 46004 28318
rect 45836 27746 45892 27758
rect 45836 27694 45838 27746
rect 45890 27694 45892 27746
rect 45836 27636 45892 27694
rect 45836 27570 45892 27580
rect 45948 26962 46004 28252
rect 46284 28084 46340 28094
rect 46396 28084 46452 28924
rect 46620 28868 46676 29374
rect 46620 28802 46676 28812
rect 46284 28082 46452 28084
rect 46284 28030 46286 28082
rect 46338 28030 46452 28082
rect 46284 28028 46452 28030
rect 46508 28420 46564 28430
rect 46284 28018 46340 28028
rect 46508 27076 46564 28364
rect 46508 27010 46564 27020
rect 46620 28084 46676 28094
rect 45948 26910 45950 26962
rect 46002 26910 46004 26962
rect 45388 26852 45556 26908
rect 45948 26898 46004 26910
rect 45500 26796 45780 26852
rect 45388 26404 45444 26414
rect 45388 26310 45444 26348
rect 45276 25454 45278 25506
rect 45330 25454 45332 25506
rect 45276 25442 45332 25454
rect 45500 26180 45556 26190
rect 45500 25620 45556 26124
rect 45724 25844 45780 26796
rect 46396 26516 46452 26526
rect 46396 26422 46452 26460
rect 45724 25778 45780 25788
rect 45836 26404 45892 26414
rect 45836 25620 45892 26348
rect 46620 26402 46676 28028
rect 46732 27970 46788 29708
rect 46844 28866 46900 29932
rect 47180 29428 47236 31614
rect 47180 29362 47236 29372
rect 46844 28814 46846 28866
rect 46898 28814 46900 28866
rect 46844 28084 46900 28814
rect 46956 29314 47012 29326
rect 46956 29262 46958 29314
rect 47010 29262 47012 29314
rect 46956 28756 47012 29262
rect 46956 28690 47012 28700
rect 46844 28018 46900 28028
rect 46956 28530 47012 28542
rect 46956 28478 46958 28530
rect 47010 28478 47012 28530
rect 46732 27918 46734 27970
rect 46786 27918 46788 27970
rect 46732 27186 46788 27918
rect 46844 27858 46900 27870
rect 46844 27806 46846 27858
rect 46898 27806 46900 27858
rect 46844 27412 46900 27806
rect 46844 27346 46900 27356
rect 46956 27858 47012 28478
rect 47292 28532 47348 32844
rect 47404 32676 47460 32686
rect 47404 32582 47460 32620
rect 47628 32562 47684 32574
rect 47628 32510 47630 32562
rect 47682 32510 47684 32562
rect 47516 32452 47572 32462
rect 47516 32358 47572 32396
rect 47628 32116 47684 32510
rect 47628 32050 47684 32060
rect 48076 32564 48132 32574
rect 48076 32004 48132 32508
rect 48188 32450 48244 32462
rect 48188 32398 48190 32450
rect 48242 32398 48244 32450
rect 48188 32228 48244 32398
rect 48188 32162 48244 32172
rect 48076 31778 48132 31948
rect 48076 31726 48078 31778
rect 48130 31726 48132 31778
rect 48076 31714 48132 31726
rect 48300 31666 48356 35252
rect 48412 35252 48468 37212
rect 48524 37202 48580 37212
rect 48748 38610 48804 38622
rect 48748 38558 48750 38610
rect 48802 38558 48804 38610
rect 48524 36484 48580 36494
rect 48748 36484 48804 38558
rect 48860 38612 48916 38622
rect 48860 38050 48916 38556
rect 48860 37998 48862 38050
rect 48914 37998 48916 38050
rect 48860 37986 48916 37998
rect 49532 38050 49588 38780
rect 49644 38668 49700 39004
rect 49868 38966 49924 39004
rect 49980 39058 50036 39340
rect 49980 39006 49982 39058
rect 50034 39006 50036 39058
rect 49980 38994 50036 39006
rect 50092 39058 50148 39564
rect 50092 39006 50094 39058
rect 50146 39006 50148 39058
rect 50092 38994 50148 39006
rect 50204 41076 50260 41086
rect 50204 39730 50260 41020
rect 50428 40292 50484 41132
rect 50540 41122 50596 41132
rect 50764 41076 50820 41806
rect 50988 41188 51044 42588
rect 51100 42644 51156 42654
rect 51436 42644 51492 42654
rect 51100 42642 51492 42644
rect 51100 42590 51102 42642
rect 51154 42590 51438 42642
rect 51490 42590 51492 42642
rect 51100 42588 51492 42590
rect 51100 42578 51156 42588
rect 51436 42578 51492 42588
rect 51660 42644 51716 42654
rect 51996 42644 52052 42654
rect 51660 42550 51716 42588
rect 51884 42642 52052 42644
rect 51884 42590 51998 42642
rect 52050 42590 52052 42642
rect 51884 42588 52052 42590
rect 51548 42532 51604 42542
rect 51548 41860 51604 42476
rect 51772 42530 51828 42542
rect 51772 42478 51774 42530
rect 51826 42478 51828 42530
rect 51772 41970 51828 42478
rect 51772 41918 51774 41970
rect 51826 41918 51828 41970
rect 51772 41906 51828 41918
rect 51436 41804 51604 41860
rect 51884 41860 51940 42588
rect 51996 42578 52052 42588
rect 51212 41188 51268 41198
rect 50988 41186 51268 41188
rect 50988 41134 51214 41186
rect 51266 41134 51268 41186
rect 50988 41132 51268 41134
rect 51212 41122 51268 41132
rect 51436 41186 51492 41804
rect 51884 41794 51940 41804
rect 51996 42084 52052 42094
rect 51436 41134 51438 41186
rect 51490 41134 51492 41186
rect 50764 41010 50820 41020
rect 50876 40964 50932 40974
rect 51436 40964 51492 41134
rect 51548 41412 51604 41422
rect 51548 41186 51604 41356
rect 51996 41410 52052 42028
rect 52108 41972 52164 43262
rect 52780 42980 52836 42990
rect 52332 42978 52836 42980
rect 52332 42926 52782 42978
rect 52834 42926 52836 42978
rect 52332 42924 52836 42926
rect 52220 41972 52276 41982
rect 52108 41916 52220 41972
rect 52220 41906 52276 41916
rect 52332 41970 52388 42924
rect 52780 42914 52836 42924
rect 52332 41918 52334 41970
rect 52386 41918 52388 41970
rect 52332 41906 52388 41918
rect 52668 42756 52724 42766
rect 51996 41358 51998 41410
rect 52050 41358 52052 41410
rect 51996 41346 52052 41358
rect 52668 41412 52724 42700
rect 52780 42532 52836 42542
rect 52780 42438 52836 42476
rect 53788 42532 53844 42542
rect 53116 42194 53172 42206
rect 53116 42142 53118 42194
rect 53170 42142 53172 42194
rect 53004 42084 53060 42094
rect 53004 41990 53060 42028
rect 52780 41970 52836 41982
rect 52780 41918 52782 41970
rect 52834 41918 52836 41970
rect 52780 41860 52836 41918
rect 52780 41794 52836 41804
rect 52780 41412 52836 41422
rect 52724 41410 52836 41412
rect 52724 41358 52782 41410
rect 52834 41358 52836 41410
rect 52724 41356 52836 41358
rect 52668 41318 52724 41356
rect 52780 41346 52836 41356
rect 51548 41134 51550 41186
rect 51602 41134 51604 41186
rect 51548 41122 51604 41134
rect 52892 41074 52948 41086
rect 52892 41022 52894 41074
rect 52946 41022 52948 41074
rect 50876 40962 51492 40964
rect 50876 40910 50878 40962
rect 50930 40910 51492 40962
rect 50876 40908 51492 40910
rect 52780 40964 52836 40974
rect 50876 40898 50932 40908
rect 52780 40870 52836 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 51436 40628 51492 40638
rect 52108 40628 52164 40638
rect 51436 40626 51940 40628
rect 51436 40574 51438 40626
rect 51490 40574 51940 40626
rect 51436 40572 51940 40574
rect 51436 40562 51492 40572
rect 50428 40226 50484 40236
rect 50540 40516 50596 40526
rect 50204 39678 50206 39730
rect 50258 39678 50260 39730
rect 50204 38668 50260 39678
rect 50316 40180 50372 40190
rect 50316 39060 50372 40124
rect 50540 39730 50596 40460
rect 51884 40514 51940 40572
rect 51884 40462 51886 40514
rect 51938 40462 51940 40514
rect 51884 40450 51940 40462
rect 50764 40404 50820 40414
rect 50764 40310 50820 40348
rect 50876 40402 50932 40414
rect 50876 40350 50878 40402
rect 50930 40350 50932 40402
rect 50876 39844 50932 40350
rect 51324 40402 51380 40414
rect 51548 40404 51604 40414
rect 52108 40404 52164 40572
rect 52444 40516 52500 40526
rect 52892 40516 52948 41022
rect 52444 40422 52500 40460
rect 52780 40460 52948 40516
rect 51324 40350 51326 40402
rect 51378 40350 51380 40402
rect 51324 40292 51380 40350
rect 51324 40226 51380 40236
rect 51436 40402 51604 40404
rect 51436 40350 51550 40402
rect 51602 40350 51604 40402
rect 51436 40348 51604 40350
rect 51436 40180 51492 40348
rect 51548 40338 51604 40348
rect 51996 40402 52164 40404
rect 51996 40350 52110 40402
rect 52162 40350 52164 40402
rect 51996 40348 52164 40350
rect 51436 40114 51492 40124
rect 51884 40292 51940 40302
rect 50540 39678 50542 39730
rect 50594 39678 50596 39730
rect 50540 39666 50596 39678
rect 50764 39788 50932 39844
rect 50764 39508 50820 39788
rect 51884 39732 51940 40236
rect 50876 39620 50932 39630
rect 50876 39526 50932 39564
rect 50316 38994 50372 39004
rect 50428 39452 50820 39508
rect 51100 39506 51156 39518
rect 51100 39454 51102 39506
rect 51154 39454 51156 39506
rect 49644 38612 50260 38668
rect 50428 38834 50484 39452
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50428 38782 50430 38834
rect 50482 38782 50484 38834
rect 50428 38724 50484 38782
rect 50428 38658 50484 38668
rect 50988 38724 51044 38734
rect 49532 37998 49534 38050
rect 49586 37998 49588 38050
rect 49532 37986 49588 37998
rect 49868 38276 49924 38286
rect 48524 36482 48804 36484
rect 48524 36430 48526 36482
rect 48578 36430 48804 36482
rect 48524 36428 48804 36430
rect 49644 37492 49700 37502
rect 49644 36482 49700 37436
rect 49644 36430 49646 36482
rect 49698 36430 49700 36482
rect 48524 35924 48580 36428
rect 49084 36372 49140 36382
rect 49084 36278 49140 36316
rect 48636 36260 48692 36270
rect 48636 36166 48692 36204
rect 48748 36260 48804 36270
rect 48748 36258 48916 36260
rect 48748 36206 48750 36258
rect 48802 36206 48916 36258
rect 48748 36204 48916 36206
rect 48748 36194 48804 36204
rect 48524 35858 48580 35868
rect 48748 36036 48804 36046
rect 48748 35698 48804 35980
rect 48748 35646 48750 35698
rect 48802 35646 48804 35698
rect 48748 35634 48804 35646
rect 48860 35476 48916 36204
rect 49196 36258 49252 36270
rect 49196 36206 49198 36258
rect 49250 36206 49252 36258
rect 49196 35812 49252 36206
rect 49308 36260 49364 36270
rect 49308 36166 49364 36204
rect 49196 35746 49252 35756
rect 48860 35410 48916 35420
rect 49420 35700 49476 35710
rect 49084 35252 49140 35262
rect 48412 35196 49028 35252
rect 48412 34916 48468 34926
rect 48412 34822 48468 34860
rect 48972 33570 49028 35196
rect 48972 33518 48974 33570
rect 49026 33518 49028 33570
rect 48972 33506 49028 33518
rect 49084 34132 49140 35196
rect 49420 35026 49476 35644
rect 49420 34974 49422 35026
rect 49474 34974 49476 35026
rect 49420 34962 49476 34974
rect 49532 35698 49588 35710
rect 49532 35646 49534 35698
rect 49586 35646 49588 35698
rect 49532 35588 49588 35646
rect 49420 34692 49476 34702
rect 48860 33460 48916 33470
rect 48860 32564 48916 33404
rect 49084 33234 49140 34076
rect 49084 33182 49086 33234
rect 49138 33182 49140 33234
rect 49084 33170 49140 33182
rect 49196 34468 49252 34478
rect 48860 32470 48916 32508
rect 49084 32788 49140 32798
rect 49196 32788 49252 34412
rect 49308 33572 49364 33582
rect 49420 33572 49476 34636
rect 49532 34244 49588 35532
rect 49532 33684 49588 34188
rect 49532 33618 49588 33628
rect 49308 33570 49476 33572
rect 49308 33518 49310 33570
rect 49362 33518 49476 33570
rect 49308 33516 49476 33518
rect 49308 33506 49364 33516
rect 49084 32786 49252 32788
rect 49084 32734 49086 32786
rect 49138 32734 49252 32786
rect 49084 32732 49252 32734
rect 48300 31614 48302 31666
rect 48354 31614 48356 31666
rect 48300 31556 48356 31614
rect 48300 31490 48356 31500
rect 48412 32340 48468 32350
rect 47516 31220 47572 31230
rect 47516 31126 47572 31164
rect 48076 30996 48132 31006
rect 48076 30994 48244 30996
rect 48076 30942 48078 30994
rect 48130 30942 48244 30994
rect 48076 30940 48244 30942
rect 48076 30930 48132 30940
rect 47628 30210 47684 30222
rect 47628 30158 47630 30210
rect 47682 30158 47684 30210
rect 47516 29652 47572 29662
rect 47516 29558 47572 29596
rect 47292 28466 47348 28476
rect 47628 28308 47684 30158
rect 47964 30098 48020 30110
rect 47964 30046 47966 30098
rect 48018 30046 48020 30098
rect 47852 29316 47908 29326
rect 47852 29222 47908 29260
rect 47628 28242 47684 28252
rect 47740 29092 47796 29102
rect 47628 28084 47684 28094
rect 47628 27990 47684 28028
rect 47404 27860 47460 27870
rect 46956 27806 46958 27858
rect 47010 27806 47012 27858
rect 46956 27636 47012 27806
rect 46732 27134 46734 27186
rect 46786 27134 46788 27186
rect 46732 27122 46788 27134
rect 46620 26350 46622 26402
rect 46674 26350 46676 26402
rect 46620 26338 46676 26350
rect 46844 26404 46900 26414
rect 46844 26310 46900 26348
rect 46284 26292 46340 26302
rect 46284 26198 46340 26236
rect 45500 25506 45556 25564
rect 45500 25454 45502 25506
rect 45554 25454 45556 25506
rect 45500 25442 45556 25454
rect 45724 25618 45892 25620
rect 45724 25566 45838 25618
rect 45890 25566 45892 25618
rect 45724 25564 45892 25566
rect 45388 25284 45444 25294
rect 45052 24770 45108 24780
rect 45276 25282 45444 25284
rect 45276 25230 45390 25282
rect 45442 25230 45444 25282
rect 45276 25228 45444 25230
rect 44940 24670 44942 24722
rect 44994 24670 44996 24722
rect 44940 24658 44996 24670
rect 44268 24220 44436 24276
rect 43932 23886 43934 23938
rect 43986 23886 43988 23938
rect 43932 23874 43988 23886
rect 43764 23100 43876 23156
rect 43708 23062 43764 23100
rect 43484 22278 43540 22316
rect 43596 22820 43652 22830
rect 43372 22258 43428 22270
rect 43372 22206 43374 22258
rect 43426 22206 43428 22258
rect 43372 22148 43428 22206
rect 43372 22082 43428 22092
rect 43596 22036 43652 22764
rect 44268 22708 44324 22718
rect 44268 22482 44324 22652
rect 44268 22430 44270 22482
rect 44322 22430 44324 22482
rect 44268 22418 44324 22430
rect 43708 22370 43764 22382
rect 43708 22318 43710 22370
rect 43762 22318 43764 22370
rect 43708 22260 43764 22318
rect 43708 22194 43764 22204
rect 43596 21980 43764 22036
rect 43260 21868 43652 21924
rect 40908 21646 40910 21698
rect 40962 21646 40964 21698
rect 40348 21634 40404 21644
rect 40236 21422 40238 21474
rect 40290 21422 40292 21474
rect 40236 21410 40292 21422
rect 40908 20804 40964 21646
rect 42364 21700 42420 21710
rect 40908 20738 40964 20748
rect 41244 21588 41300 21598
rect 41244 20242 41300 21532
rect 42140 21588 42196 21598
rect 42140 21494 42196 21532
rect 41244 20190 41246 20242
rect 41298 20190 41300 20242
rect 41244 20178 41300 20190
rect 41804 20914 41860 20926
rect 41804 20862 41806 20914
rect 41858 20862 41860 20914
rect 40348 20132 40404 20142
rect 40348 20038 40404 20076
rect 41132 20132 41188 20142
rect 41132 20038 41188 20076
rect 41804 20132 41860 20862
rect 42252 20916 42308 20926
rect 42252 20822 42308 20860
rect 42140 20804 42196 20814
rect 42140 20710 42196 20748
rect 42364 20802 42420 21644
rect 42476 21586 42532 21868
rect 42476 21534 42478 21586
rect 42530 21534 42532 21586
rect 42476 21522 42532 21534
rect 42924 21586 42980 21868
rect 42924 21534 42926 21586
rect 42978 21534 42980 21586
rect 42364 20750 42366 20802
rect 42418 20750 42420 20802
rect 42364 20738 42420 20750
rect 42812 20914 42868 20926
rect 42812 20862 42814 20914
rect 42866 20862 42868 20914
rect 42812 20802 42868 20862
rect 42812 20750 42814 20802
rect 42866 20750 42868 20802
rect 42812 20738 42868 20750
rect 42924 20580 42980 21534
rect 43148 21588 43204 21598
rect 43148 21494 43204 21532
rect 43036 21476 43092 21486
rect 43036 21382 43092 21420
rect 43372 21476 43428 21486
rect 43372 21382 43428 21420
rect 43596 21026 43652 21868
rect 43708 21586 43764 21980
rect 44380 21700 44436 24220
rect 44828 24052 44884 24062
rect 44716 23268 44772 23278
rect 44716 22148 44772 23212
rect 44828 22482 44884 23996
rect 44940 23940 44996 23950
rect 45164 23940 45220 23950
rect 44940 23846 44996 23884
rect 45052 23938 45220 23940
rect 45052 23886 45166 23938
rect 45218 23886 45220 23938
rect 45052 23884 45220 23886
rect 45276 23940 45332 25228
rect 45388 25218 45444 25228
rect 45724 24834 45780 25564
rect 45836 25554 45892 25564
rect 46060 25844 46116 25854
rect 45724 24782 45726 24834
rect 45778 24782 45780 24834
rect 45724 24770 45780 24782
rect 45948 24612 46004 24622
rect 45388 24276 45444 24286
rect 45388 24162 45444 24220
rect 45388 24110 45390 24162
rect 45442 24110 45444 24162
rect 45388 24098 45444 24110
rect 45500 23996 45780 24052
rect 45500 23940 45556 23996
rect 45276 23884 45556 23940
rect 44940 22708 44996 22718
rect 45052 22708 45108 23884
rect 45164 23874 45220 23884
rect 45612 23826 45668 23838
rect 45612 23774 45614 23826
rect 45666 23774 45668 23826
rect 45500 23714 45556 23726
rect 45500 23662 45502 23714
rect 45554 23662 45556 23714
rect 44996 22652 45108 22708
rect 45164 23154 45220 23166
rect 45164 23102 45166 23154
rect 45218 23102 45220 23154
rect 44940 22642 44996 22652
rect 44828 22430 44830 22482
rect 44882 22430 44884 22482
rect 44828 22418 44884 22430
rect 44716 22082 44772 22092
rect 45164 22372 45220 23102
rect 45164 21810 45220 22316
rect 45276 22708 45332 22718
rect 45276 22370 45332 22652
rect 45276 22318 45278 22370
rect 45330 22318 45332 22370
rect 45276 22260 45332 22318
rect 45276 22194 45332 22204
rect 45164 21758 45166 21810
rect 45218 21758 45220 21810
rect 45164 21746 45220 21758
rect 44380 21606 44436 21644
rect 43708 21534 43710 21586
rect 43762 21534 43764 21586
rect 43708 21522 43764 21534
rect 43932 21586 43988 21598
rect 43932 21534 43934 21586
rect 43986 21534 43988 21586
rect 43596 20974 43598 21026
rect 43650 20974 43652 21026
rect 43596 20914 43652 20974
rect 43596 20862 43598 20914
rect 43650 20862 43652 20914
rect 43596 20850 43652 20862
rect 43932 20804 43988 21534
rect 44492 21586 44548 21598
rect 44492 21534 44494 21586
rect 44546 21534 44548 21586
rect 44156 21476 44212 21486
rect 44156 21382 44212 21420
rect 44492 20916 44548 21534
rect 45276 21476 45332 21486
rect 45276 21382 45332 21420
rect 44492 20850 44548 20860
rect 43932 20738 43988 20748
rect 44940 20804 44996 20814
rect 43260 20580 43316 20590
rect 42924 20524 43260 20580
rect 43260 20486 43316 20524
rect 41804 20066 41860 20076
rect 39788 19966 39790 20018
rect 39842 19966 39844 20018
rect 39788 19954 39844 19966
rect 44940 20018 44996 20748
rect 45500 20132 45556 23662
rect 45612 23044 45668 23774
rect 45724 23266 45780 23996
rect 45948 23938 46004 24556
rect 45948 23886 45950 23938
rect 46002 23886 46004 23938
rect 45948 23874 46004 23886
rect 46060 23380 46116 25788
rect 46732 25620 46788 25630
rect 46732 25526 46788 25564
rect 46396 25396 46452 25406
rect 46620 25396 46676 25406
rect 46396 25394 46620 25396
rect 46396 25342 46398 25394
rect 46450 25342 46620 25394
rect 46396 25340 46620 25342
rect 46396 25330 46452 25340
rect 46620 25330 46676 25340
rect 46956 25396 47012 27580
rect 47180 27858 47460 27860
rect 47180 27806 47406 27858
rect 47458 27806 47460 27858
rect 47180 27804 47460 27806
rect 47180 26514 47236 27804
rect 47404 27794 47460 27804
rect 47180 26462 47182 26514
rect 47234 26462 47236 26514
rect 47180 26292 47236 26462
rect 47516 27746 47572 27758
rect 47516 27694 47518 27746
rect 47570 27694 47572 27746
rect 47516 26404 47572 27694
rect 47516 26338 47572 26348
rect 47740 27188 47796 29036
rect 47852 28532 47908 28542
rect 47852 28084 47908 28476
rect 47852 27990 47908 28028
rect 47964 27188 48020 30046
rect 48076 29540 48132 29550
rect 48076 29446 48132 29484
rect 48188 28644 48244 30940
rect 48188 28578 48244 28588
rect 48412 27972 48468 32284
rect 48972 32004 49028 32014
rect 48972 31910 49028 31948
rect 48860 31668 48916 31678
rect 48748 31612 48860 31668
rect 48636 31108 48692 31118
rect 48636 28754 48692 31052
rect 48748 31106 48804 31612
rect 48860 31574 48916 31612
rect 48748 31054 48750 31106
rect 48802 31054 48804 31106
rect 48748 31042 48804 31054
rect 48972 31556 49028 31566
rect 48860 30996 48916 31006
rect 48860 30902 48916 30940
rect 48972 30772 49028 31500
rect 49084 31220 49140 32732
rect 49420 32676 49476 32686
rect 49420 31780 49476 32620
rect 49532 32676 49588 32686
rect 49644 32676 49700 36430
rect 49756 35252 49812 35262
rect 49756 35026 49812 35196
rect 49756 34974 49758 35026
rect 49810 34974 49812 35026
rect 49756 34962 49812 34974
rect 49868 34018 49924 38220
rect 50204 38050 50260 38612
rect 50876 38276 50932 38286
rect 50876 38182 50932 38220
rect 50204 37998 50206 38050
rect 50258 37998 50260 38050
rect 50204 37986 50260 37998
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50092 37266 50148 37278
rect 50092 37214 50094 37266
rect 50146 37214 50148 37266
rect 49980 37154 50036 37166
rect 49980 37102 49982 37154
rect 50034 37102 50036 37154
rect 49980 36596 50036 37102
rect 49980 36148 50036 36540
rect 49980 36082 50036 36092
rect 49868 33966 49870 34018
rect 49922 33966 49924 34018
rect 49868 33954 49924 33966
rect 49980 35924 50036 35934
rect 49980 33458 50036 35868
rect 50092 35700 50148 37214
rect 50764 36708 50820 36718
rect 50652 36596 50708 36606
rect 50316 36482 50372 36494
rect 50316 36430 50318 36482
rect 50370 36430 50372 36482
rect 50092 35634 50148 35644
rect 50204 36372 50260 36382
rect 50204 34914 50260 36316
rect 50316 36260 50372 36430
rect 50540 36484 50596 36522
rect 50540 36418 50596 36428
rect 50652 36482 50708 36540
rect 50652 36430 50654 36482
rect 50706 36430 50708 36482
rect 50652 36418 50708 36430
rect 50764 36372 50820 36652
rect 50876 36596 50932 36606
rect 50988 36596 51044 38668
rect 51100 38722 51156 39454
rect 51884 39506 51940 39676
rect 51884 39454 51886 39506
rect 51938 39454 51940 39506
rect 51884 39442 51940 39454
rect 51436 39396 51492 39406
rect 51436 39302 51492 39340
rect 51996 39284 52052 40348
rect 52108 40338 52164 40348
rect 52332 40292 52388 40302
rect 52332 40198 52388 40236
rect 52668 39732 52724 39742
rect 52780 39732 52836 40460
rect 52892 40290 52948 40302
rect 52892 40238 52894 40290
rect 52946 40238 52948 40290
rect 52892 40180 52948 40238
rect 52892 40114 52948 40124
rect 52724 39676 52836 39732
rect 52668 39638 52724 39676
rect 51100 38670 51102 38722
rect 51154 38670 51156 38722
rect 51100 38276 51156 38670
rect 51884 39228 52052 39284
rect 51100 38220 51492 38276
rect 51324 38052 51380 38062
rect 50876 36594 51044 36596
rect 50876 36542 50878 36594
rect 50930 36542 51044 36594
rect 50876 36540 51044 36542
rect 51100 38050 51380 38052
rect 51100 37998 51326 38050
rect 51378 37998 51380 38050
rect 51100 37996 51380 37998
rect 51436 38052 51492 38220
rect 51772 38052 51828 38062
rect 51436 38050 51828 38052
rect 51436 37998 51774 38050
rect 51826 37998 51828 38050
rect 51436 37996 51828 37998
rect 50876 36530 50932 36540
rect 50988 36372 51044 36382
rect 50764 36370 51044 36372
rect 50764 36318 50990 36370
rect 51042 36318 51044 36370
rect 50764 36316 51044 36318
rect 50316 36194 50372 36204
rect 50556 36092 50820 36102
rect 50204 34862 50206 34914
rect 50258 34862 50260 34914
rect 50204 34850 50260 34862
rect 50316 36036 50372 36046
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50316 34692 50372 35980
rect 50876 35924 50932 36316
rect 50988 36306 51044 36316
rect 50876 35858 50932 35868
rect 50652 35700 50708 35710
rect 50652 35606 50708 35644
rect 51100 35588 51156 37996
rect 51324 37986 51380 37996
rect 50652 35476 50708 35486
rect 50652 34914 50708 35420
rect 50652 34862 50654 34914
rect 50706 34862 50708 34914
rect 50652 34850 50708 34862
rect 51100 34802 51156 35532
rect 51100 34750 51102 34802
rect 51154 34750 51156 34802
rect 51100 34738 51156 34750
rect 51212 37266 51268 37278
rect 51212 37214 51214 37266
rect 51266 37214 51268 37266
rect 50092 34636 50372 34692
rect 50988 34690 51044 34702
rect 50988 34638 50990 34690
rect 51042 34638 51044 34690
rect 50092 33572 50148 34636
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50316 34132 50372 34142
rect 50316 34038 50372 34076
rect 50988 34130 51044 34638
rect 50988 34078 50990 34130
rect 51042 34078 51044 34130
rect 50988 34066 51044 34078
rect 50204 33908 50260 33918
rect 50204 33906 50484 33908
rect 50204 33854 50206 33906
rect 50258 33854 50484 33906
rect 50204 33852 50484 33854
rect 50204 33842 50260 33852
rect 50316 33684 50372 33694
rect 50204 33572 50260 33582
rect 50092 33570 50260 33572
rect 50092 33518 50206 33570
rect 50258 33518 50260 33570
rect 50092 33516 50260 33518
rect 50204 33506 50260 33516
rect 49980 33406 49982 33458
rect 50034 33406 50036 33458
rect 49980 33394 50036 33406
rect 50316 33346 50372 33628
rect 50316 33294 50318 33346
rect 50370 33294 50372 33346
rect 50316 33282 50372 33294
rect 49868 32788 49924 32798
rect 49868 32786 50372 32788
rect 49868 32734 49870 32786
rect 49922 32734 50372 32786
rect 49868 32732 50372 32734
rect 49868 32722 49924 32732
rect 49532 32674 49700 32676
rect 49532 32622 49534 32674
rect 49586 32622 49700 32674
rect 49532 32620 49700 32622
rect 50316 32674 50372 32732
rect 50316 32622 50318 32674
rect 50370 32622 50372 32674
rect 49532 32228 49588 32620
rect 50316 32610 50372 32622
rect 49756 32564 49812 32574
rect 49868 32564 49924 32574
rect 49756 32562 49868 32564
rect 49756 32510 49758 32562
rect 49810 32510 49868 32562
rect 49756 32508 49868 32510
rect 49756 32498 49812 32508
rect 49532 32162 49588 32172
rect 49420 31686 49476 31724
rect 49644 32116 49700 32126
rect 49644 31778 49700 32060
rect 49644 31726 49646 31778
rect 49698 31726 49700 31778
rect 49084 31154 49140 31164
rect 49196 31444 49252 31454
rect 48636 28702 48638 28754
rect 48690 28702 48692 28754
rect 48636 28690 48692 28702
rect 48748 30716 49028 30772
rect 49084 30994 49140 31006
rect 49084 30942 49086 30994
rect 49138 30942 49140 30994
rect 48412 27906 48468 27916
rect 47964 27132 48468 27188
rect 47740 26402 47796 27132
rect 47740 26350 47742 26402
rect 47794 26350 47796 26402
rect 47740 26338 47796 26350
rect 47964 26964 48020 26974
rect 47180 26226 47236 26236
rect 47516 26068 47572 26078
rect 47516 26066 47796 26068
rect 47516 26014 47518 26066
rect 47570 26014 47796 26066
rect 47516 26012 47796 26014
rect 47516 26002 47572 26012
rect 47516 25620 47572 25630
rect 46956 25330 47012 25340
rect 47404 25508 47460 25518
rect 47292 25284 47348 25294
rect 47292 25190 47348 25228
rect 46620 24836 46676 24846
rect 46620 24742 46676 24780
rect 47292 24836 47348 24846
rect 46844 24722 46900 24734
rect 46844 24670 46846 24722
rect 46898 24670 46900 24722
rect 46284 24052 46340 24062
rect 46284 23958 46340 23996
rect 46508 23940 46564 23950
rect 46508 23846 46564 23884
rect 46060 23314 46116 23324
rect 45724 23214 45726 23266
rect 45778 23214 45780 23266
rect 45724 23202 45780 23214
rect 45948 23154 46004 23166
rect 45948 23102 45950 23154
rect 46002 23102 46004 23154
rect 45948 23044 46004 23102
rect 46396 23156 46452 23166
rect 46396 23062 46452 23100
rect 45612 22988 46004 23044
rect 45948 22932 46004 22988
rect 45948 22866 46004 22876
rect 46172 23042 46228 23054
rect 46172 22990 46174 23042
rect 46226 22990 46228 23042
rect 46172 22596 46228 22990
rect 46732 23042 46788 23054
rect 46732 22990 46734 23042
rect 46786 22990 46788 23042
rect 46508 22932 46564 22942
rect 46564 22876 46676 22932
rect 46508 22866 46564 22876
rect 45836 22540 46228 22596
rect 46620 22594 46676 22876
rect 46620 22542 46622 22594
rect 46674 22542 46676 22594
rect 45724 22482 45780 22494
rect 45724 22430 45726 22482
rect 45778 22430 45780 22482
rect 45612 20916 45668 20926
rect 45724 20916 45780 22430
rect 45836 22258 45892 22540
rect 46620 22530 46676 22542
rect 46732 22596 46788 22990
rect 46732 22530 46788 22540
rect 46844 22484 46900 24670
rect 47292 24722 47348 24780
rect 47292 24670 47294 24722
rect 47346 24670 47348 24722
rect 47068 24612 47124 24622
rect 47068 24518 47124 24556
rect 47180 24052 47236 24062
rect 47180 23958 47236 23996
rect 47292 23716 47348 24670
rect 47404 24724 47460 25452
rect 47516 25506 47572 25564
rect 47740 25618 47796 26012
rect 47740 25566 47742 25618
rect 47794 25566 47796 25618
rect 47740 25554 47796 25566
rect 47852 25844 47908 25854
rect 47516 25454 47518 25506
rect 47570 25454 47572 25506
rect 47516 25442 47572 25454
rect 47740 25396 47796 25406
rect 47516 24724 47572 24734
rect 47404 24722 47572 24724
rect 47404 24670 47518 24722
rect 47570 24670 47572 24722
rect 47404 24668 47572 24670
rect 47516 24658 47572 24668
rect 47740 24722 47796 25340
rect 47740 24670 47742 24722
rect 47794 24670 47796 24722
rect 47740 24658 47796 24670
rect 47852 24388 47908 25788
rect 47964 25506 48020 26908
rect 48188 26516 48244 26526
rect 48244 26460 48356 26516
rect 48188 26450 48244 26460
rect 48300 26402 48356 26460
rect 48300 26350 48302 26402
rect 48354 26350 48356 26402
rect 48300 26338 48356 26350
rect 47964 25454 47966 25506
rect 48018 25454 48020 25506
rect 47964 25442 48020 25454
rect 48076 25506 48132 25518
rect 48076 25454 48078 25506
rect 48130 25454 48132 25506
rect 48076 24724 48132 25454
rect 47628 24332 47908 24388
rect 47628 24050 47684 24332
rect 47628 23998 47630 24050
rect 47682 23998 47684 24050
rect 47628 23986 47684 23998
rect 47740 24164 47796 24174
rect 47516 23940 47572 23950
rect 47516 23846 47572 23884
rect 46956 23660 47348 23716
rect 47404 23828 47460 23838
rect 46956 22594 47012 23660
rect 46956 22542 46958 22594
rect 47010 22542 47012 22594
rect 46956 22530 47012 22542
rect 47068 23492 47124 23502
rect 47068 23156 47124 23436
rect 47404 23378 47460 23772
rect 47740 23492 47796 24108
rect 47404 23326 47406 23378
rect 47458 23326 47460 23378
rect 47404 23314 47460 23326
rect 47628 23436 47796 23492
rect 47180 23156 47236 23166
rect 47068 23154 47236 23156
rect 47068 23102 47182 23154
rect 47234 23102 47236 23154
rect 47068 23100 47236 23102
rect 46844 22418 46900 22428
rect 46060 22372 46116 22382
rect 47068 22372 47124 23100
rect 47180 23090 47236 23100
rect 47516 23156 47572 23166
rect 47292 23042 47348 23054
rect 47292 22990 47294 23042
rect 47346 22990 47348 23042
rect 47180 22484 47236 22494
rect 47180 22390 47236 22428
rect 46060 22278 46116 22316
rect 46956 22316 47124 22372
rect 47292 22372 47348 22990
rect 47516 22594 47572 23100
rect 47516 22542 47518 22594
rect 47570 22542 47572 22594
rect 47516 22530 47572 22542
rect 45836 22206 45838 22258
rect 45890 22206 45892 22258
rect 45836 22194 45892 22206
rect 46844 21812 46900 21822
rect 46956 21812 47012 22316
rect 47292 22306 47348 22316
rect 47628 22258 47684 23436
rect 47740 23156 47796 23166
rect 47740 23062 47796 23100
rect 47852 22932 47908 24332
rect 47964 24668 48076 24724
rect 47964 23044 48020 24668
rect 48076 24658 48132 24668
rect 48076 24498 48132 24510
rect 48076 24446 48078 24498
rect 48130 24446 48132 24498
rect 48076 23268 48132 24446
rect 48300 23940 48356 23950
rect 48076 23202 48132 23212
rect 48188 23380 48244 23390
rect 48188 23156 48244 23324
rect 48188 23090 48244 23100
rect 47964 22988 48132 23044
rect 47628 22206 47630 22258
rect 47682 22206 47684 22258
rect 47628 22194 47684 22206
rect 47740 22876 47908 22932
rect 47740 22260 47796 22876
rect 48076 22708 48132 22988
rect 47852 22652 48132 22708
rect 47852 22482 47908 22652
rect 47852 22430 47854 22482
rect 47906 22430 47908 22482
rect 47852 22418 47908 22430
rect 48188 22484 48244 22494
rect 47740 22204 48020 22260
rect 46844 21810 47012 21812
rect 46844 21758 46846 21810
rect 46898 21758 47012 21810
rect 46844 21756 47012 21758
rect 47404 22148 47460 22158
rect 47404 21810 47460 22092
rect 47740 21924 47796 22204
rect 47404 21758 47406 21810
rect 47458 21758 47460 21810
rect 46844 21746 46900 21756
rect 47404 21746 47460 21758
rect 47516 21868 47796 21924
rect 47852 22036 47908 22046
rect 47180 21588 47236 21598
rect 47516 21588 47572 21868
rect 47852 21812 47908 21980
rect 47740 21810 47908 21812
rect 47740 21758 47854 21810
rect 47906 21758 47908 21810
rect 47740 21756 47908 21758
rect 47180 21586 47572 21588
rect 47180 21534 47182 21586
rect 47234 21534 47572 21586
rect 47180 21532 47572 21534
rect 47180 21522 47236 21532
rect 45612 20914 45780 20916
rect 45612 20862 45614 20914
rect 45666 20862 45780 20914
rect 45612 20860 45780 20862
rect 45612 20850 45668 20860
rect 47516 20692 47572 21532
rect 47628 21586 47684 21598
rect 47628 21534 47630 21586
rect 47682 21534 47684 21586
rect 47628 21476 47684 21534
rect 47628 21410 47684 21420
rect 47740 20914 47796 21756
rect 47852 21746 47908 21756
rect 47964 21698 48020 22204
rect 47964 21646 47966 21698
rect 48018 21646 48020 21698
rect 47964 21634 48020 21646
rect 47740 20862 47742 20914
rect 47794 20862 47796 20914
rect 47740 20850 47796 20862
rect 48188 20914 48244 22428
rect 48300 22260 48356 23884
rect 48412 22482 48468 27132
rect 48524 27074 48580 27086
rect 48524 27022 48526 27074
rect 48578 27022 48580 27074
rect 48524 25844 48580 27022
rect 48748 27076 48804 30716
rect 49084 30436 49140 30942
rect 49196 30994 49252 31388
rect 49196 30942 49198 30994
rect 49250 30942 49252 30994
rect 49196 30930 49252 30942
rect 49532 31444 49588 31454
rect 49084 30370 49140 30380
rect 48972 30210 49028 30222
rect 48972 30158 48974 30210
rect 49026 30158 49028 30210
rect 48860 30100 48916 30110
rect 48860 29652 48916 30044
rect 48972 29764 49028 30158
rect 48972 29708 49364 29764
rect 49308 29652 49364 29708
rect 48860 29650 49252 29652
rect 48860 29598 48862 29650
rect 48914 29598 49252 29650
rect 48860 29596 49252 29598
rect 48860 29586 48916 29596
rect 49196 28644 49252 29596
rect 49308 29586 49364 29596
rect 49308 28644 49364 28654
rect 49196 28588 49308 28644
rect 49196 27858 49252 28588
rect 49308 28550 49364 28588
rect 49196 27806 49198 27858
rect 49250 27806 49252 27858
rect 49196 27794 49252 27806
rect 49420 27188 49476 27198
rect 49420 27094 49476 27132
rect 48860 27076 48916 27086
rect 48748 27074 48916 27076
rect 48748 27022 48862 27074
rect 48914 27022 48916 27074
rect 48748 27020 48916 27022
rect 48524 25778 48580 25788
rect 48636 26962 48692 26974
rect 48636 26910 48638 26962
rect 48690 26910 48692 26962
rect 48636 25620 48692 26910
rect 48748 26964 48804 27020
rect 48860 27010 48916 27020
rect 48748 26898 48804 26908
rect 49196 26964 49252 26974
rect 49196 26962 49364 26964
rect 49196 26910 49198 26962
rect 49250 26910 49364 26962
rect 49196 26908 49364 26910
rect 49196 26898 49252 26908
rect 48748 26404 48804 26414
rect 48860 26404 48916 26414
rect 48748 26402 48860 26404
rect 48748 26350 48750 26402
rect 48802 26350 48860 26402
rect 48748 26348 48860 26350
rect 48748 26338 48804 26348
rect 48524 25564 48692 25620
rect 48524 23268 48580 25564
rect 48860 25506 48916 26348
rect 49308 26404 49364 26908
rect 49308 26338 49364 26348
rect 49420 26516 49476 26526
rect 49084 26292 49140 26302
rect 49084 26198 49140 26236
rect 49420 26290 49476 26460
rect 49420 26238 49422 26290
rect 49474 26238 49476 26290
rect 49420 26226 49476 26238
rect 49532 25956 49588 31388
rect 49644 31220 49700 31726
rect 49644 31154 49700 31164
rect 49756 31554 49812 31566
rect 49756 31502 49758 31554
rect 49810 31502 49812 31554
rect 49644 29652 49700 29662
rect 49644 29538 49700 29596
rect 49644 29486 49646 29538
rect 49698 29486 49700 29538
rect 49644 29474 49700 29486
rect 49756 29540 49812 31502
rect 49868 30884 49924 32508
rect 49980 32562 50036 32574
rect 49980 32510 49982 32562
rect 50034 32510 50036 32562
rect 49980 32004 50036 32510
rect 49980 31938 50036 31948
rect 49980 31666 50036 31678
rect 49980 31614 49982 31666
rect 50034 31614 50036 31666
rect 49980 31332 50036 31614
rect 50428 31668 50484 33852
rect 51212 33460 51268 37214
rect 51324 36482 51380 36494
rect 51324 36430 51326 36482
rect 51378 36430 51380 36482
rect 51324 34916 51380 36430
rect 51660 36370 51716 37996
rect 51772 37986 51828 37996
rect 51660 36318 51662 36370
rect 51714 36318 51716 36370
rect 51660 36306 51716 36318
rect 51772 37266 51828 37278
rect 51772 37214 51774 37266
rect 51826 37214 51828 37266
rect 51772 35924 51828 37214
rect 51324 34850 51380 34860
rect 51436 35868 51828 35924
rect 51436 35586 51492 35868
rect 51436 35534 51438 35586
rect 51490 35534 51492 35586
rect 51436 34132 51492 35534
rect 51436 34066 51492 34076
rect 51884 33908 51940 39228
rect 52220 38276 52276 38286
rect 52220 37266 52276 38220
rect 52220 37214 52222 37266
rect 52274 37214 52276 37266
rect 52220 37202 52276 37214
rect 52668 38050 52724 38062
rect 52668 37998 52670 38050
rect 52722 37998 52724 38050
rect 52556 36708 52612 36718
rect 51996 36484 52052 36494
rect 51996 36370 52052 36428
rect 51996 36318 51998 36370
rect 52050 36318 52052 36370
rect 51996 36306 52052 36318
rect 52556 36258 52612 36652
rect 52556 36206 52558 36258
rect 52610 36206 52612 36258
rect 52556 36148 52612 36206
rect 51996 36092 52612 36148
rect 51996 34690 52052 36092
rect 52108 35700 52164 35710
rect 52668 35700 52724 37998
rect 53116 38050 53172 42142
rect 53788 42082 53844 42476
rect 53788 42030 53790 42082
rect 53842 42030 53844 42082
rect 53788 42018 53844 42030
rect 53676 41972 53732 41982
rect 53676 41878 53732 41916
rect 53340 40964 53396 40974
rect 53340 40870 53396 40908
rect 53788 40628 53844 40638
rect 53788 40534 53844 40572
rect 53452 40404 53508 40414
rect 53452 40310 53508 40348
rect 54012 40404 54068 40414
rect 54012 38836 54068 40348
rect 54796 40292 54852 40302
rect 54796 39730 54852 40236
rect 54796 39678 54798 39730
rect 54850 39678 54852 39730
rect 54796 39666 54852 39678
rect 54012 38742 54068 38780
rect 55468 39618 55524 39630
rect 55468 39566 55470 39618
rect 55522 39566 55524 39618
rect 55468 38836 55524 39566
rect 55468 38770 55524 38780
rect 55580 39396 55636 39406
rect 53228 38724 53284 38734
rect 53228 38630 53284 38668
rect 53116 37998 53118 38050
rect 53170 37998 53172 38050
rect 53116 37492 53172 37998
rect 52108 35698 52724 35700
rect 52108 35646 52110 35698
rect 52162 35646 52724 35698
rect 52108 35644 52724 35646
rect 52780 37436 53116 37492
rect 52108 35634 52164 35644
rect 52108 35140 52164 35150
rect 52108 34914 52164 35084
rect 52108 34862 52110 34914
rect 52162 34862 52164 34914
rect 52108 34850 52164 34862
rect 51996 34638 51998 34690
rect 52050 34638 52052 34690
rect 51996 34626 52052 34638
rect 52108 34692 52164 34702
rect 52220 34692 52276 35644
rect 52164 34636 52276 34692
rect 52108 34626 52164 34636
rect 51212 33394 51268 33404
rect 51324 33852 51940 33908
rect 51100 33122 51156 33134
rect 51100 33070 51102 33122
rect 51154 33070 51156 33122
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50540 32564 50596 32574
rect 50540 32470 50596 32508
rect 50876 32562 50932 32574
rect 50876 32510 50878 32562
rect 50930 32510 50932 32562
rect 50764 32450 50820 32462
rect 50764 32398 50766 32450
rect 50818 32398 50820 32450
rect 50764 32116 50820 32398
rect 50764 32050 50820 32060
rect 50876 32004 50932 32510
rect 51100 32340 51156 33070
rect 51100 32274 51156 32284
rect 51324 31948 51380 33852
rect 52108 33348 52164 33358
rect 52108 33122 52164 33292
rect 52780 33234 52836 37436
rect 53116 37426 53172 37436
rect 53788 37492 53844 37502
rect 53788 37398 53844 37436
rect 54908 37380 54964 37390
rect 53116 37268 53172 37278
rect 53004 36820 53060 36830
rect 53004 36706 53060 36764
rect 53004 36654 53006 36706
rect 53058 36654 53060 36706
rect 53004 36642 53060 36654
rect 53116 35140 53172 37212
rect 54684 37266 54740 37278
rect 54684 37214 54686 37266
rect 54738 37214 54740 37266
rect 53452 37156 53508 37166
rect 53452 37062 53508 37100
rect 54236 37154 54292 37166
rect 54236 37102 54238 37154
rect 54290 37102 54292 37154
rect 54236 36820 54292 37102
rect 54236 36754 54292 36764
rect 54684 37156 54740 37214
rect 54684 36594 54740 37100
rect 54908 37266 54964 37324
rect 54908 37214 54910 37266
rect 54962 37214 54964 37266
rect 54908 36708 54964 37214
rect 55356 37268 55412 37278
rect 55356 37174 55412 37212
rect 55132 37154 55188 37166
rect 55132 37102 55134 37154
rect 55186 37102 55188 37154
rect 54908 36642 54964 36652
rect 55020 37044 55076 37054
rect 54684 36542 54686 36594
rect 54738 36542 54740 36594
rect 54684 36530 54740 36542
rect 53228 36484 53284 36494
rect 53452 36484 53508 36494
rect 54908 36484 54964 36494
rect 53284 36428 53396 36484
rect 53228 36390 53284 36428
rect 53228 35698 53284 35710
rect 53228 35646 53230 35698
rect 53282 35646 53284 35698
rect 53228 35252 53284 35646
rect 53228 35186 53284 35196
rect 53116 35046 53172 35084
rect 52892 35028 52948 35038
rect 52892 34692 52948 34972
rect 52892 34626 52948 34636
rect 53340 34914 53396 36428
rect 53452 36482 53732 36484
rect 53452 36430 53454 36482
rect 53506 36430 53732 36482
rect 53452 36428 53732 36430
rect 53452 36418 53508 36428
rect 53340 34862 53342 34914
rect 53394 34862 53396 34914
rect 53228 34130 53284 34142
rect 53228 34078 53230 34130
rect 53282 34078 53284 34130
rect 53228 34020 53284 34078
rect 53228 33954 53284 33964
rect 53340 33346 53396 34862
rect 53676 34916 53732 36428
rect 53900 36260 53956 36270
rect 53900 36166 53956 36204
rect 54572 35924 54628 35934
rect 54628 35868 54740 35924
rect 54572 35858 54628 35868
rect 54012 35810 54068 35822
rect 54012 35758 54014 35810
rect 54066 35758 54068 35810
rect 53788 34916 53844 34926
rect 53676 34860 53788 34916
rect 53788 34822 53844 34860
rect 54012 34356 54068 35758
rect 54012 34262 54068 34300
rect 54348 35698 54404 35710
rect 54348 35646 54350 35698
rect 54402 35646 54404 35698
rect 54348 34692 54404 35646
rect 54572 35252 54628 35262
rect 54572 35138 54628 35196
rect 54572 35086 54574 35138
rect 54626 35086 54628 35138
rect 54572 35074 54628 35086
rect 54460 35028 54516 35038
rect 54460 34934 54516 34972
rect 54460 34692 54516 34702
rect 54348 34690 54516 34692
rect 54348 34638 54462 34690
rect 54514 34638 54516 34690
rect 54348 34636 54516 34638
rect 54236 34244 54292 34254
rect 54348 34244 54404 34636
rect 54460 34626 54516 34636
rect 54236 34242 54404 34244
rect 54236 34190 54238 34242
rect 54290 34190 54404 34242
rect 54236 34188 54404 34190
rect 54684 34244 54740 35868
rect 54908 35364 54964 36428
rect 55020 36482 55076 36988
rect 55020 36430 55022 36482
rect 55074 36430 55076 36482
rect 55020 36418 55076 36430
rect 55132 35698 55188 37102
rect 55468 36372 55524 36382
rect 55468 36278 55524 36316
rect 55132 35646 55134 35698
rect 55186 35646 55188 35698
rect 55132 35634 55188 35646
rect 55356 35588 55412 35598
rect 54908 35298 54964 35308
rect 55244 35532 55356 35588
rect 55244 35252 55300 35532
rect 55356 35522 55412 35532
rect 55356 35364 55412 35374
rect 55356 35252 55524 35308
rect 55132 35196 55300 35252
rect 54796 34916 54852 34926
rect 54852 34860 55076 34916
rect 54796 34822 54852 34860
rect 54796 34244 54852 34254
rect 54684 34242 54852 34244
rect 54684 34190 54798 34242
rect 54850 34190 54852 34242
rect 54684 34188 54852 34190
rect 54236 34178 54292 34188
rect 54796 34178 54852 34188
rect 55020 34244 55076 34860
rect 55020 34150 55076 34188
rect 53340 33294 53342 33346
rect 53394 33294 53396 33346
rect 53340 33282 53396 33294
rect 53452 34130 53508 34142
rect 53452 34078 53454 34130
rect 53506 34078 53508 34130
rect 52780 33182 52782 33234
rect 52834 33182 52836 33234
rect 52780 33170 52836 33182
rect 52108 33070 52110 33122
rect 52162 33070 52164 33122
rect 52108 32788 52164 33070
rect 52108 32722 52164 32732
rect 52220 33124 52276 33134
rect 53228 33124 53284 33134
rect 52220 32786 52276 33068
rect 52220 32734 52222 32786
rect 52274 32734 52276 32786
rect 52220 32722 52276 32734
rect 53116 33122 53284 33124
rect 53116 33070 53230 33122
rect 53282 33070 53284 33122
rect 53116 33068 53284 33070
rect 51660 32562 51716 32574
rect 51660 32510 51662 32562
rect 51714 32510 51716 32562
rect 50876 31938 50932 31948
rect 51212 31892 51380 31948
rect 51436 32450 51492 32462
rect 51436 32398 51438 32450
rect 51490 32398 51492 32450
rect 50316 31556 50372 31566
rect 49980 31266 50036 31276
rect 50092 31554 50372 31556
rect 50092 31502 50318 31554
rect 50370 31502 50372 31554
rect 50092 31500 50372 31502
rect 49868 30882 50036 30884
rect 49868 30830 49870 30882
rect 49922 30830 50036 30882
rect 49868 30828 50036 30830
rect 49868 30818 49924 30828
rect 49980 30100 50036 30828
rect 49980 30034 50036 30044
rect 49756 29426 49812 29484
rect 49756 29374 49758 29426
rect 49810 29374 49812 29426
rect 49756 29362 49812 29374
rect 49980 29316 50036 29326
rect 50092 29316 50148 31500
rect 50316 31490 50372 31500
rect 50204 31332 50260 31342
rect 50204 30996 50260 31276
rect 50204 30930 50260 30940
rect 50036 29260 50148 29316
rect 50204 30210 50260 30222
rect 50204 30158 50206 30210
rect 50258 30158 50260 30210
rect 49980 29222 50036 29260
rect 50204 27412 50260 30158
rect 50428 30212 50484 31612
rect 50652 31778 50708 31790
rect 50652 31726 50654 31778
rect 50706 31726 50708 31778
rect 50652 31556 50708 31726
rect 50876 31780 50932 31790
rect 50876 31778 51044 31780
rect 50876 31726 50878 31778
rect 50930 31726 51044 31778
rect 50876 31724 51044 31726
rect 50876 31714 50932 31724
rect 50652 31490 50708 31500
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50988 31332 51044 31724
rect 50988 30996 51044 31276
rect 50988 30930 51044 30940
rect 51100 31220 51156 31230
rect 51100 30994 51156 31164
rect 51100 30942 51102 30994
rect 51154 30942 51156 30994
rect 51100 30930 51156 30942
rect 50540 30884 50596 30894
rect 50596 30828 50708 30884
rect 50540 30818 50596 30828
rect 50652 30324 50708 30828
rect 50540 30212 50596 30222
rect 50428 30210 50596 30212
rect 50428 30158 50542 30210
rect 50594 30158 50596 30210
rect 50428 30156 50596 30158
rect 50540 30146 50596 30156
rect 50652 29988 50708 30268
rect 50428 29932 50708 29988
rect 50876 29986 50932 29998
rect 50876 29934 50878 29986
rect 50930 29934 50932 29986
rect 50428 29652 50484 29932
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50428 29596 50596 29652
rect 50428 29428 50484 29438
rect 50428 29334 50484 29372
rect 50540 29426 50596 29596
rect 50540 29374 50542 29426
rect 50594 29374 50596 29426
rect 50540 28980 50596 29374
rect 50428 28924 50596 28980
rect 50316 28644 50372 28654
rect 50316 28550 50372 28588
rect 50428 28084 50484 28924
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50428 28028 50596 28084
rect 50428 27748 50484 27758
rect 50428 27654 50484 27692
rect 49644 27356 50260 27412
rect 49644 27186 49700 27356
rect 49644 27134 49646 27186
rect 49698 27134 49700 27186
rect 49644 27122 49700 27134
rect 49980 27188 50036 27198
rect 49868 27076 49924 27086
rect 49868 26982 49924 27020
rect 49980 26850 50036 27132
rect 50204 27186 50260 27356
rect 50204 27134 50206 27186
rect 50258 27134 50260 27186
rect 50204 27122 50260 27134
rect 50540 27636 50596 28028
rect 50540 27186 50596 27580
rect 50540 27134 50542 27186
rect 50594 27134 50596 27186
rect 50540 27122 50596 27134
rect 50652 27972 50708 27982
rect 50652 27524 50708 27916
rect 50652 27074 50708 27468
rect 50652 27022 50654 27074
rect 50706 27022 50708 27074
rect 50652 27010 50708 27022
rect 50876 26964 50932 29934
rect 51100 29428 51156 29438
rect 50988 28980 51044 28990
rect 50988 28642 51044 28924
rect 50988 28590 50990 28642
rect 51042 28590 51044 28642
rect 50988 28578 51044 28590
rect 51100 28418 51156 29372
rect 51100 28366 51102 28418
rect 51154 28366 51156 28418
rect 51100 28354 51156 28366
rect 51212 28084 51268 31892
rect 51436 31780 51492 32398
rect 51660 32340 51716 32510
rect 51772 32564 51828 32574
rect 52108 32564 52164 32574
rect 51772 32562 52164 32564
rect 51772 32510 51774 32562
rect 51826 32510 52110 32562
rect 52162 32510 52164 32562
rect 51772 32508 52164 32510
rect 51772 32498 51828 32508
rect 51660 32284 51828 32340
rect 51548 32004 51604 32042
rect 51772 31948 51828 32284
rect 51548 31938 51604 31948
rect 51660 31892 51828 31948
rect 51548 31780 51604 31790
rect 51436 31778 51604 31780
rect 51436 31726 51550 31778
rect 51602 31726 51604 31778
rect 51436 31724 51604 31726
rect 51436 30994 51492 31006
rect 51436 30942 51438 30994
rect 51490 30942 51492 30994
rect 51436 30884 51492 30942
rect 51436 30818 51492 30828
rect 51548 30548 51604 31724
rect 51660 31220 51716 31892
rect 51884 31778 51940 32508
rect 52108 32498 52164 32508
rect 51884 31726 51886 31778
rect 51938 31726 51940 31778
rect 51884 31714 51940 31726
rect 52108 32340 52164 32350
rect 52108 32004 52164 32284
rect 52108 31778 52164 31948
rect 52108 31726 52110 31778
rect 52162 31726 52164 31778
rect 52108 31714 52164 31726
rect 52668 31892 52724 31902
rect 52668 31780 52724 31836
rect 52668 31778 52836 31780
rect 52668 31726 52670 31778
rect 52722 31726 52836 31778
rect 52668 31724 52836 31726
rect 52668 31714 52724 31724
rect 51996 31668 52052 31678
rect 51996 31574 52052 31612
rect 52108 31556 52164 31566
rect 51660 31154 51716 31164
rect 51996 31332 52052 31342
rect 51996 30882 52052 31276
rect 51996 30830 51998 30882
rect 52050 30830 52052 30882
rect 51548 30492 51940 30548
rect 51660 30324 51716 30334
rect 51548 30100 51604 30110
rect 51548 30006 51604 30044
rect 51660 29650 51716 30268
rect 51660 29598 51662 29650
rect 51714 29598 51716 29650
rect 51660 29586 51716 29598
rect 51884 28308 51940 30492
rect 51996 28530 52052 30830
rect 52108 30324 52164 31500
rect 52108 29538 52164 30268
rect 52444 30994 52500 31006
rect 52444 30942 52446 30994
rect 52498 30942 52500 30994
rect 52444 30884 52500 30942
rect 52780 30994 52836 31724
rect 52780 30942 52782 30994
rect 52834 30942 52836 30994
rect 52780 30930 52836 30942
rect 53004 30996 53060 31006
rect 53004 30902 53060 30940
rect 52444 29652 52500 30828
rect 53116 30212 53172 33068
rect 53228 33058 53284 33068
rect 53340 32674 53396 32686
rect 53340 32622 53342 32674
rect 53394 32622 53396 32674
rect 53340 32116 53396 32622
rect 53228 32060 53396 32116
rect 53228 31890 53284 32060
rect 53228 31838 53230 31890
rect 53282 31838 53284 31890
rect 53228 31780 53284 31838
rect 53228 31714 53284 31724
rect 53340 31948 53396 31958
rect 53340 30996 53396 31892
rect 53452 31332 53508 34078
rect 55132 34132 55188 35196
rect 55244 35026 55300 35038
rect 55244 34974 55246 35026
rect 55298 34974 55300 35026
rect 55244 34356 55300 34974
rect 55244 34290 55300 34300
rect 55244 34132 55300 34142
rect 55132 34130 55300 34132
rect 55132 34078 55246 34130
rect 55298 34078 55300 34130
rect 55132 34076 55300 34078
rect 55244 34066 55300 34076
rect 55468 34130 55524 35252
rect 55580 34580 55636 39340
rect 57372 38836 57428 38846
rect 55692 37380 55748 37390
rect 55692 37286 55748 37324
rect 55804 37268 55860 37278
rect 55804 37174 55860 37212
rect 55692 37044 55748 37054
rect 55692 36950 55748 36988
rect 56364 36708 56420 36718
rect 56364 36706 56532 36708
rect 56364 36654 56366 36706
rect 56418 36654 56532 36706
rect 56364 36652 56532 36654
rect 56364 36642 56420 36652
rect 56364 36484 56420 36494
rect 56364 36390 56420 36428
rect 55804 36370 55860 36382
rect 55804 36318 55806 36370
rect 55858 36318 55860 36370
rect 55804 36260 55860 36318
rect 55804 36194 55860 36204
rect 56028 36370 56084 36382
rect 56028 36318 56030 36370
rect 56082 36318 56084 36370
rect 55804 35586 55860 35598
rect 55804 35534 55806 35586
rect 55858 35534 55860 35586
rect 55804 34692 55860 35534
rect 55804 34626 55860 34636
rect 55580 34514 55636 34524
rect 55468 34078 55470 34130
rect 55522 34078 55524 34130
rect 53900 34020 53956 34030
rect 53900 33926 53956 33964
rect 54908 34018 54964 34030
rect 54908 33966 54910 34018
rect 54962 33966 54964 34018
rect 54236 33908 54292 33918
rect 54236 33234 54292 33852
rect 54796 33684 54852 33694
rect 54796 33572 54852 33628
rect 54348 33570 54852 33572
rect 54348 33518 54798 33570
rect 54850 33518 54852 33570
rect 54348 33516 54852 33518
rect 54348 33346 54404 33516
rect 54796 33506 54852 33516
rect 54908 33572 54964 33966
rect 55468 33684 55524 34078
rect 54908 33506 54964 33516
rect 55356 33628 55524 33684
rect 55916 34356 55972 34366
rect 55916 34242 55972 34300
rect 55916 34190 55918 34242
rect 55970 34190 55972 34242
rect 55244 33458 55300 33470
rect 55244 33406 55246 33458
rect 55298 33406 55300 33458
rect 55244 33348 55300 33406
rect 54348 33294 54350 33346
rect 54402 33294 54404 33346
rect 54348 33282 54404 33294
rect 54684 33292 55300 33348
rect 55356 33348 55412 33628
rect 54236 33182 54238 33234
rect 54290 33182 54292 33234
rect 54236 33170 54292 33182
rect 54684 33234 54740 33292
rect 55356 33282 55412 33292
rect 54684 33182 54686 33234
rect 54738 33182 54740 33234
rect 54684 32676 54740 33182
rect 54796 32676 54852 32686
rect 54684 32674 54852 32676
rect 54684 32622 54798 32674
rect 54850 32622 54852 32674
rect 54684 32620 54852 32622
rect 54796 32610 54852 32620
rect 55916 32562 55972 34190
rect 56028 34354 56084 36318
rect 56252 36258 56308 36270
rect 56252 36206 56254 36258
rect 56306 36206 56308 36258
rect 56252 35028 56308 36206
rect 56252 34962 56308 34972
rect 56028 34302 56030 34354
rect 56082 34302 56084 34354
rect 56028 33908 56084 34302
rect 56476 34356 56532 36652
rect 57036 36484 57092 36494
rect 57036 36390 57092 36428
rect 56588 36372 56644 36382
rect 56588 35810 56644 36316
rect 56588 35758 56590 35810
rect 56642 35758 56644 35810
rect 56588 35746 56644 35758
rect 57372 35922 57428 38780
rect 57372 35870 57374 35922
rect 57426 35870 57428 35922
rect 56924 35698 56980 35710
rect 56924 35646 56926 35698
rect 56978 35646 56980 35698
rect 56700 35588 56756 35598
rect 56700 35494 56756 35532
rect 56924 35308 56980 35646
rect 57372 35474 57428 35870
rect 57484 36260 57540 36270
rect 57484 35812 57540 36204
rect 57484 35756 57988 35812
rect 57372 35422 57374 35474
rect 57426 35422 57428 35474
rect 57372 35410 57428 35422
rect 57820 35586 57876 35598
rect 57820 35534 57822 35586
rect 57874 35534 57876 35586
rect 57820 35308 57876 35534
rect 56924 35252 57876 35308
rect 57372 35028 57428 35038
rect 57372 34934 57428 34972
rect 56476 34290 56532 34300
rect 57260 34692 57316 34702
rect 56588 34244 56644 34254
rect 56588 34150 56644 34188
rect 57260 34242 57316 34636
rect 57372 34356 57428 34366
rect 57372 34262 57428 34300
rect 57260 34190 57262 34242
rect 57314 34190 57316 34242
rect 57260 34178 57316 34190
rect 57484 34242 57540 35252
rect 57932 34356 57988 35756
rect 58044 35474 58100 35486
rect 58044 35422 58046 35474
rect 58098 35422 58100 35474
rect 58044 34916 58100 35422
rect 58044 34914 58212 34916
rect 58044 34862 58046 34914
rect 58098 34862 58212 34914
rect 58044 34860 58212 34862
rect 58044 34850 58100 34860
rect 58044 34356 58100 34366
rect 57932 34354 58100 34356
rect 57932 34302 58046 34354
rect 58098 34302 58100 34354
rect 57932 34300 58100 34302
rect 58044 34290 58100 34300
rect 57484 34190 57486 34242
rect 57538 34190 57540 34242
rect 56028 33842 56084 33852
rect 56812 34130 56868 34142
rect 56812 34078 56814 34130
rect 56866 34078 56868 34130
rect 56812 33684 56868 34078
rect 56812 33618 56868 33628
rect 57372 33572 57428 33582
rect 57372 33458 57428 33516
rect 57372 33406 57374 33458
rect 57426 33406 57428 33458
rect 57372 33394 57428 33406
rect 55916 32510 55918 32562
rect 55970 32510 55972 32562
rect 55916 32498 55972 32510
rect 56700 33348 56756 33358
rect 56700 32786 56756 33292
rect 56700 32734 56702 32786
rect 56754 32734 56756 32786
rect 53452 31266 53508 31276
rect 53900 31890 53956 31902
rect 53900 31838 53902 31890
rect 53954 31838 53956 31890
rect 53676 31220 53732 31230
rect 53676 31126 53732 31164
rect 53900 30996 53956 31838
rect 56700 31778 56756 32734
rect 56700 31726 56702 31778
rect 56754 31726 56756 31778
rect 56028 31668 56084 31678
rect 56028 31574 56084 31612
rect 54460 31108 54516 31118
rect 54460 31014 54516 31052
rect 56700 31108 56756 31726
rect 56700 31042 56756 31052
rect 57148 32452 57204 32462
rect 57484 32452 57540 34190
rect 58156 33348 58212 34860
rect 58156 33254 58212 33292
rect 57148 32450 57540 32452
rect 57148 32398 57150 32450
rect 57202 32398 57540 32450
rect 57148 32396 57540 32398
rect 53340 30940 53508 30996
rect 53340 30770 53396 30782
rect 53340 30718 53342 30770
rect 53394 30718 53396 30770
rect 53340 30212 53396 30718
rect 53116 30210 53284 30212
rect 53116 30158 53118 30210
rect 53170 30158 53284 30210
rect 53116 30156 53284 30158
rect 53116 30146 53172 30156
rect 52892 29986 52948 29998
rect 52892 29934 52894 29986
rect 52946 29934 52948 29986
rect 52892 29652 52948 29934
rect 52108 29486 52110 29538
rect 52162 29486 52164 29538
rect 52108 28644 52164 29486
rect 52220 29596 52948 29652
rect 52220 29538 52276 29596
rect 52220 29486 52222 29538
rect 52274 29486 52276 29538
rect 52220 29474 52276 29486
rect 52444 29428 52500 29438
rect 52444 29334 52500 29372
rect 52668 29204 52724 29214
rect 52668 29110 52724 29148
rect 52668 28644 52724 28654
rect 52108 28642 52724 28644
rect 52108 28590 52110 28642
rect 52162 28590 52670 28642
rect 52722 28590 52724 28642
rect 52108 28588 52724 28590
rect 52108 28578 52164 28588
rect 52668 28578 52724 28588
rect 51996 28478 51998 28530
rect 52050 28478 52052 28530
rect 51996 28466 52052 28478
rect 52892 28530 52948 29596
rect 52892 28478 52894 28530
rect 52946 28478 52948 28530
rect 52892 28466 52948 28478
rect 53116 29426 53172 29438
rect 53116 29374 53118 29426
rect 53170 29374 53172 29426
rect 52668 28420 52724 28430
rect 51884 28252 52500 28308
rect 52108 28084 52164 28094
rect 51212 28028 52052 28084
rect 51660 27858 51716 27870
rect 51660 27806 51662 27858
rect 51714 27806 51716 27858
rect 51548 27300 51604 27310
rect 51660 27300 51716 27806
rect 51884 27860 51940 27870
rect 51884 27766 51940 27804
rect 51604 27244 51716 27300
rect 51772 27746 51828 27758
rect 51772 27694 51774 27746
rect 51826 27694 51828 27746
rect 51548 27074 51604 27244
rect 51548 27022 51550 27074
rect 51602 27022 51604 27074
rect 51548 27010 51604 27022
rect 50876 26908 51044 26964
rect 49980 26798 49982 26850
rect 50034 26798 50036 26850
rect 49980 26786 50036 26798
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 49644 26404 49700 26414
rect 49700 26348 49812 26404
rect 49644 26338 49700 26348
rect 49756 26292 49812 26348
rect 49980 26292 50036 26302
rect 49756 26290 49924 26292
rect 49756 26238 49758 26290
rect 49810 26238 49924 26290
rect 49756 26236 49924 26238
rect 49756 26226 49812 26236
rect 49644 26180 49700 26190
rect 49644 26086 49700 26124
rect 49532 25844 49588 25900
rect 49532 25788 49812 25844
rect 49756 25730 49812 25788
rect 49756 25678 49758 25730
rect 49810 25678 49812 25730
rect 49756 25666 49812 25678
rect 48860 25454 48862 25506
rect 48914 25454 48916 25506
rect 48860 25442 48916 25454
rect 49868 25508 49924 26236
rect 49980 25732 50036 26236
rect 50764 26292 50820 26302
rect 50764 26198 50820 26236
rect 50092 26180 50148 26190
rect 50876 26180 50932 26190
rect 50092 26178 50484 26180
rect 50092 26126 50094 26178
rect 50146 26126 50484 26178
rect 50092 26124 50484 26126
rect 50092 26114 50148 26124
rect 50092 25732 50148 25742
rect 49980 25730 50148 25732
rect 49980 25678 50094 25730
rect 50146 25678 50148 25730
rect 49980 25676 50148 25678
rect 50092 25666 50148 25676
rect 49980 25508 50036 25518
rect 49868 25506 50036 25508
rect 49868 25454 49982 25506
rect 50034 25454 50036 25506
rect 49868 25452 50036 25454
rect 49980 25442 50036 25452
rect 50428 25506 50484 26124
rect 50876 26086 50932 26124
rect 50988 26068 51044 26908
rect 51772 26516 51828 27694
rect 50988 26002 51044 26012
rect 51100 26460 51828 26516
rect 51996 27186 52052 28028
rect 52108 27990 52164 28028
rect 51996 27134 51998 27186
rect 52050 27134 52052 27186
rect 50876 25956 50932 25966
rect 50428 25454 50430 25506
rect 50482 25454 50484 25506
rect 50428 25442 50484 25454
rect 50764 25620 50820 25630
rect 49420 25396 49476 25406
rect 48636 25284 48692 25294
rect 48636 25190 48692 25228
rect 48972 25282 49028 25294
rect 48972 25230 48974 25282
rect 49026 25230 49028 25282
rect 48860 25172 48916 25182
rect 48748 24722 48804 24734
rect 48748 24670 48750 24722
rect 48802 24670 48804 24722
rect 48748 24164 48804 24670
rect 48860 24610 48916 25116
rect 48972 24836 49028 25230
rect 49084 25284 49140 25294
rect 49084 25190 49140 25228
rect 48972 24770 49028 24780
rect 49084 24724 49140 24734
rect 49084 24630 49140 24668
rect 48860 24558 48862 24610
rect 48914 24558 48916 24610
rect 48860 24546 48916 24558
rect 48748 24050 48804 24108
rect 48748 23998 48750 24050
rect 48802 23998 48804 24050
rect 48748 23986 48804 23998
rect 49084 23938 49140 23950
rect 49084 23886 49086 23938
rect 49138 23886 49140 23938
rect 49084 23268 49140 23886
rect 48524 23212 48916 23268
rect 48748 23042 48804 23054
rect 48748 22990 48750 23042
rect 48802 22990 48804 23042
rect 48748 22596 48804 22990
rect 48748 22530 48804 22540
rect 48412 22430 48414 22482
rect 48466 22430 48468 22482
rect 48412 22418 48468 22430
rect 48860 22370 48916 23212
rect 49084 23202 49140 23212
rect 49196 23826 49252 23838
rect 49196 23774 49198 23826
rect 49250 23774 49252 23826
rect 49196 23492 49252 23774
rect 49196 23156 49252 23436
rect 49308 23156 49364 23166
rect 49196 23154 49364 23156
rect 49196 23102 49310 23154
rect 49362 23102 49364 23154
rect 49196 23100 49364 23102
rect 48860 22318 48862 22370
rect 48914 22318 48916 22370
rect 48300 22166 48356 22204
rect 48524 22258 48580 22270
rect 48524 22206 48526 22258
rect 48578 22206 48580 22258
rect 48524 22148 48580 22206
rect 48524 22082 48580 22092
rect 48860 22036 48916 22318
rect 49196 22260 49252 22270
rect 49196 22166 49252 22204
rect 49308 22148 49364 23100
rect 49420 22484 49476 25340
rect 50092 25282 50148 25294
rect 50092 25230 50094 25282
rect 50146 25230 50148 25282
rect 49532 23940 49588 23950
rect 49532 23846 49588 23884
rect 50092 23940 50148 25230
rect 50764 25282 50820 25564
rect 50876 25506 50932 25900
rect 50876 25454 50878 25506
rect 50930 25454 50932 25506
rect 50876 25442 50932 25454
rect 51100 25506 51156 26460
rect 51436 26292 51492 26302
rect 51436 26198 51492 26236
rect 51100 25454 51102 25506
rect 51154 25454 51156 25506
rect 51100 25442 51156 25454
rect 51548 26178 51604 26190
rect 51548 26126 51550 26178
rect 51602 26126 51604 26178
rect 51548 25508 51604 26126
rect 51996 25956 52052 27134
rect 52332 27748 52388 27758
rect 52332 27076 52388 27692
rect 52444 27076 52500 28252
rect 52668 27970 52724 28364
rect 52780 28418 52836 28430
rect 52780 28366 52782 28418
rect 52834 28366 52836 28418
rect 52780 28084 52836 28366
rect 53116 28084 53172 29374
rect 53228 29316 53284 30156
rect 53340 29538 53396 30156
rect 53452 29876 53508 30940
rect 53900 30902 53956 30940
rect 54348 30660 54404 30670
rect 57148 30660 57204 32396
rect 54404 30604 54516 30660
rect 54348 30594 54404 30604
rect 53564 30324 53620 30334
rect 53564 30098 53620 30268
rect 53788 30212 53844 30222
rect 53788 30118 53844 30156
rect 53564 30046 53566 30098
rect 53618 30046 53620 30098
rect 53564 30034 53620 30046
rect 53452 29820 53620 29876
rect 53340 29486 53342 29538
rect 53394 29486 53396 29538
rect 53340 29474 53396 29486
rect 53452 29426 53508 29438
rect 53452 29374 53454 29426
rect 53506 29374 53508 29426
rect 53452 29316 53508 29374
rect 53228 29260 53508 29316
rect 53564 29204 53620 29820
rect 53676 29428 53732 29438
rect 53676 29334 53732 29372
rect 53452 29148 53620 29204
rect 54012 29314 54068 29326
rect 54012 29262 54014 29314
rect 54066 29262 54068 29314
rect 53228 28980 53284 28990
rect 53228 28642 53284 28924
rect 53228 28590 53230 28642
rect 53282 28590 53284 28642
rect 53228 28578 53284 28590
rect 52780 28028 52948 28084
rect 52668 27918 52670 27970
rect 52722 27918 52724 27970
rect 52668 27748 52724 27918
rect 52780 27860 52836 27870
rect 52780 27766 52836 27804
rect 52668 27682 52724 27692
rect 52780 27076 52836 27086
rect 52444 27074 52836 27076
rect 52444 27022 52782 27074
rect 52834 27022 52836 27074
rect 52444 27020 52836 27022
rect 52332 26290 52388 27020
rect 52332 26238 52334 26290
rect 52386 26238 52388 26290
rect 51996 25890 52052 25900
rect 52220 26068 52276 26078
rect 52108 25732 52164 25742
rect 51548 25442 51604 25452
rect 51996 25676 52108 25732
rect 50764 25230 50766 25282
rect 50818 25230 50820 25282
rect 50764 25218 50820 25230
rect 51436 25394 51492 25406
rect 51436 25342 51438 25394
rect 51490 25342 51492 25394
rect 51436 25284 51492 25342
rect 51996 25394 52052 25676
rect 52108 25666 52164 25676
rect 52108 25508 52164 25518
rect 52108 25414 52164 25452
rect 51996 25342 51998 25394
rect 52050 25342 52052 25394
rect 51996 25330 52052 25342
rect 51436 25218 51492 25228
rect 52108 25284 52164 25294
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50316 24724 50372 24734
rect 50316 24162 50372 24668
rect 50316 24110 50318 24162
rect 50370 24110 50372 24162
rect 50316 24098 50372 24110
rect 50652 24722 50708 24734
rect 50652 24670 50654 24722
rect 50706 24670 50708 24722
rect 50652 24052 50708 24670
rect 52108 24722 52164 25228
rect 52108 24670 52110 24722
rect 52162 24670 52164 24722
rect 52108 24658 52164 24670
rect 52220 24610 52276 26012
rect 52220 24558 52222 24610
rect 52274 24558 52276 24610
rect 52220 24546 52276 24558
rect 50652 23986 50708 23996
rect 50092 23874 50148 23884
rect 51100 23940 51156 23950
rect 51100 23846 51156 23884
rect 51660 23940 51716 23950
rect 51660 23846 51716 23884
rect 49756 23826 49812 23838
rect 49756 23774 49758 23826
rect 49810 23774 49812 23826
rect 49756 23492 49812 23774
rect 49756 23426 49812 23436
rect 49868 23826 49924 23838
rect 49868 23774 49870 23826
rect 49922 23774 49924 23826
rect 49644 23268 49700 23278
rect 49868 23268 49924 23774
rect 51772 23828 51828 23838
rect 51772 23734 51828 23772
rect 51548 23716 51604 23726
rect 51436 23660 51548 23716
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50876 23380 50932 23390
rect 49700 23212 49924 23268
rect 50428 23268 50484 23278
rect 49644 23154 49700 23212
rect 50428 23174 50484 23212
rect 49644 23102 49646 23154
rect 49698 23102 49700 23154
rect 49644 23090 49700 23102
rect 50092 23156 50148 23166
rect 50876 23156 50932 23324
rect 50092 22708 50148 23100
rect 50092 22642 50148 22652
rect 50540 23154 50932 23156
rect 50540 23102 50878 23154
rect 50930 23102 50932 23154
rect 50540 23100 50932 23102
rect 49644 22484 49700 22494
rect 49420 22482 49700 22484
rect 49420 22430 49646 22482
rect 49698 22430 49700 22482
rect 49420 22428 49700 22430
rect 49644 22418 49700 22428
rect 50428 22484 50484 22494
rect 50540 22484 50596 23100
rect 50876 23090 50932 23100
rect 50484 22428 50596 22484
rect 50876 22820 50932 22830
rect 50876 22484 50932 22764
rect 51436 22594 51492 23660
rect 51548 23650 51604 23660
rect 52332 23380 52388 26238
rect 52668 25508 52724 25518
rect 52668 25414 52724 25452
rect 52556 25396 52612 25406
rect 52332 23314 52388 23324
rect 52444 25284 52500 25294
rect 51548 23044 51604 23054
rect 51548 23042 51716 23044
rect 51548 22990 51550 23042
rect 51602 22990 51716 23042
rect 51548 22988 51716 22990
rect 51548 22978 51604 22988
rect 51436 22542 51438 22594
rect 51490 22542 51492 22594
rect 51436 22530 51492 22542
rect 50876 22482 51268 22484
rect 50876 22430 50878 22482
rect 50930 22430 51268 22482
rect 50876 22428 51268 22430
rect 50428 22390 50484 22428
rect 50876 22418 50932 22428
rect 51212 22370 51268 22428
rect 51212 22318 51214 22370
rect 51266 22318 51268 22370
rect 51212 22306 51268 22318
rect 49308 22082 49364 22092
rect 50876 22260 50932 22270
rect 48860 21970 48916 21980
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 48188 20862 48190 20914
rect 48242 20862 48244 20914
rect 48188 20804 48244 20862
rect 47516 20636 47796 20692
rect 45612 20132 45668 20142
rect 45500 20130 45668 20132
rect 45500 20078 45614 20130
rect 45666 20078 45668 20130
rect 45500 20076 45668 20078
rect 45612 20066 45668 20076
rect 44940 19966 44942 20018
rect 44994 19966 44996 20018
rect 44940 19954 44996 19966
rect 39004 19842 39060 19852
rect 39452 19908 39508 19918
rect 39452 19814 39508 19852
rect 47740 19906 47796 20636
rect 48188 20242 48244 20748
rect 50876 21474 50932 22204
rect 51660 22146 51716 22988
rect 52444 22820 52500 25228
rect 52444 22754 52500 22764
rect 51772 22596 51828 22606
rect 51772 22370 51828 22540
rect 51772 22318 51774 22370
rect 51826 22318 51828 22370
rect 51772 22306 51828 22318
rect 51996 22260 52052 22270
rect 51996 22166 52052 22204
rect 52556 22260 52612 25340
rect 52780 25284 52836 27020
rect 52892 25618 52948 28028
rect 53116 28018 53172 28028
rect 53340 28196 53396 28206
rect 53004 27970 53060 27982
rect 53004 27918 53006 27970
rect 53058 27918 53060 27970
rect 53004 27412 53060 27918
rect 53228 27412 53284 27422
rect 53340 27412 53396 28140
rect 53004 27356 53172 27412
rect 53004 27188 53060 27198
rect 53004 27094 53060 27132
rect 52892 25566 52894 25618
rect 52946 25566 52948 25618
rect 52892 25554 52948 25566
rect 53004 26178 53060 26190
rect 53004 26126 53006 26178
rect 53058 26126 53060 26178
rect 53004 25620 53060 26126
rect 53116 25732 53172 27356
rect 53284 27356 53396 27412
rect 53228 27074 53284 27356
rect 53228 27022 53230 27074
rect 53282 27022 53284 27074
rect 53228 27010 53284 27022
rect 53340 26964 53396 26974
rect 53340 26870 53396 26908
rect 53452 26962 53508 29148
rect 54012 28980 54068 29262
rect 54012 28914 54068 28924
rect 53900 28644 53956 28654
rect 53788 28642 53956 28644
rect 53788 28590 53902 28642
rect 53954 28590 53956 28642
rect 53788 28588 53956 28590
rect 53452 26910 53454 26962
rect 53506 26910 53508 26962
rect 53452 26516 53508 26910
rect 53340 25732 53396 25742
rect 53172 25676 53284 25732
rect 53116 25666 53172 25676
rect 53004 25554 53060 25564
rect 52780 25218 52836 25228
rect 53004 23940 53060 23950
rect 52668 23826 52724 23838
rect 52892 23828 52948 23838
rect 52668 23774 52670 23826
rect 52722 23774 52724 23826
rect 52668 23268 52724 23774
rect 52668 23202 52724 23212
rect 52780 23826 52948 23828
rect 52780 23774 52894 23826
rect 52946 23774 52948 23826
rect 52780 23772 52948 23774
rect 52668 22596 52724 22606
rect 52780 22596 52836 23772
rect 52892 23762 52948 23772
rect 53004 23714 53060 23884
rect 53004 23662 53006 23714
rect 53058 23662 53060 23714
rect 53004 23650 53060 23662
rect 53228 23548 53284 25676
rect 53340 23938 53396 25676
rect 53452 25396 53508 26460
rect 53564 27972 53620 27982
rect 53564 25506 53620 27916
rect 53788 27746 53844 28588
rect 53900 28578 53956 28588
rect 54348 27860 54404 27870
rect 54348 27766 54404 27804
rect 53788 27694 53790 27746
rect 53842 27694 53844 27746
rect 53788 27524 53844 27694
rect 53788 27458 53844 27468
rect 53564 25454 53566 25506
rect 53618 25454 53620 25506
rect 53564 25442 53620 25454
rect 53676 27076 53732 27086
rect 53452 25330 53508 25340
rect 53676 24948 53732 27020
rect 54124 27076 54180 27086
rect 54124 26982 54180 27020
rect 54236 25284 54292 25294
rect 54236 25190 54292 25228
rect 54124 24948 54180 24958
rect 53676 24946 54180 24948
rect 53676 24894 53678 24946
rect 53730 24894 54126 24946
rect 54178 24894 54180 24946
rect 53676 24892 54180 24894
rect 53676 24882 53732 24892
rect 54124 24882 54180 24892
rect 54348 24052 54404 24062
rect 54460 24052 54516 30604
rect 57148 30594 57204 30604
rect 54572 29428 54628 29438
rect 54572 29334 54628 29372
rect 57372 29428 57428 29438
rect 55020 29314 55076 29326
rect 55020 29262 55022 29314
rect 55074 29262 55076 29314
rect 54572 28644 54628 28654
rect 55020 28644 55076 29262
rect 55804 29204 55860 29214
rect 55244 28756 55300 28766
rect 55244 28662 55300 28700
rect 54572 28642 55076 28644
rect 54572 28590 54574 28642
rect 54626 28590 55076 28642
rect 54572 28588 55076 28590
rect 54572 27076 54628 28588
rect 55692 28196 55748 28206
rect 55132 28082 55188 28094
rect 55132 28030 55134 28082
rect 55186 28030 55188 28082
rect 55020 27972 55076 27982
rect 55132 27972 55188 28030
rect 55580 28084 55636 28094
rect 55580 27990 55636 28028
rect 55692 28082 55748 28140
rect 55692 28030 55694 28082
rect 55746 28030 55748 28082
rect 55692 28018 55748 28030
rect 55076 27916 55188 27972
rect 55020 27906 55076 27916
rect 54684 27858 54740 27870
rect 54684 27806 54686 27858
rect 54738 27806 54740 27858
rect 54684 27636 54740 27806
rect 54908 27858 54964 27870
rect 54908 27806 54910 27858
rect 54962 27806 54964 27858
rect 54684 27570 54740 27580
rect 54796 27634 54852 27646
rect 54796 27582 54798 27634
rect 54850 27582 54852 27634
rect 54572 27010 54628 27020
rect 54684 25956 54740 25966
rect 54684 25618 54740 25900
rect 54796 25732 54852 27582
rect 54908 27524 54964 27806
rect 54908 27458 54964 27468
rect 54908 26964 54964 26974
rect 54908 26870 54964 26908
rect 55132 26178 55188 27916
rect 55468 27748 55524 27758
rect 55468 27654 55524 27692
rect 55580 26516 55636 26526
rect 55580 26422 55636 26460
rect 55132 26126 55134 26178
rect 55186 26126 55188 26178
rect 55132 26114 55188 26126
rect 54796 25666 54852 25676
rect 54684 25566 54686 25618
rect 54738 25566 54740 25618
rect 54684 25554 54740 25566
rect 53340 23886 53342 23938
rect 53394 23886 53396 23938
rect 53340 23874 53396 23886
rect 53900 24050 54516 24052
rect 53900 23998 54350 24050
rect 54402 23998 54516 24050
rect 53900 23996 54516 23998
rect 53900 23938 53956 23996
rect 54348 23986 54404 23996
rect 53900 23886 53902 23938
rect 53954 23886 53956 23938
rect 53900 23874 53956 23886
rect 53564 23828 53620 23838
rect 53564 23734 53620 23772
rect 53676 23716 53732 23726
rect 53676 23622 53732 23660
rect 52724 22540 52836 22596
rect 52892 23492 53732 23548
rect 52668 22502 52724 22540
rect 52780 22372 52836 22382
rect 52892 22372 52948 23492
rect 53676 23042 53732 23492
rect 55804 23156 55860 29148
rect 57372 28754 57428 29372
rect 57372 28702 57374 28754
rect 57426 28702 57428 28754
rect 57372 28690 57428 28702
rect 56588 28196 56644 28206
rect 56588 28082 56644 28140
rect 56588 28030 56590 28082
rect 56642 28030 56644 28082
rect 56588 28018 56644 28030
rect 56700 27860 56756 27870
rect 56756 27804 57092 27860
rect 56700 27766 56756 27804
rect 57036 27186 57092 27804
rect 57036 27134 57038 27186
rect 57090 27134 57092 27186
rect 57036 27122 57092 27134
rect 55804 23090 55860 23100
rect 53676 22990 53678 23042
rect 53730 22990 53732 23042
rect 53676 22978 53732 22990
rect 52780 22370 52948 22372
rect 52780 22318 52782 22370
rect 52834 22318 52948 22370
rect 52780 22316 52948 22318
rect 52780 22306 52836 22316
rect 52556 22194 52612 22204
rect 51660 22094 51662 22146
rect 51714 22094 51716 22146
rect 51660 22082 51716 22094
rect 50876 21422 50878 21474
rect 50930 21422 50932 21474
rect 50876 20580 50932 21422
rect 50876 20514 50932 20524
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 48188 20190 48190 20242
rect 48242 20190 48244 20242
rect 48188 20178 48244 20190
rect 47740 19854 47742 19906
rect 47794 19854 47796 19906
rect 47740 19842 47796 19854
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 38444 18450 38612 18452
rect 38444 18398 38446 18450
rect 38498 18398 38612 18450
rect 38444 18396 38612 18398
rect 37100 17668 37156 17678
rect 38444 17668 38500 18396
rect 38892 18340 38948 18350
rect 38668 18338 38948 18340
rect 38668 18286 38894 18338
rect 38946 18286 38948 18338
rect 38668 18284 38948 18286
rect 38556 17668 38612 17678
rect 38444 17612 38556 17668
rect 37100 17574 37156 17612
rect 38556 17444 38612 17612
rect 38668 17444 38724 18284
rect 38892 18274 38948 18284
rect 38556 17388 38724 17444
rect 36316 15934 36318 15986
rect 36370 15934 36372 15986
rect 36316 15922 36372 15934
rect 36316 15540 36372 15550
rect 35756 15092 35924 15148
rect 35980 15092 36260 15148
rect 35308 15036 35700 15092
rect 35196 15026 35252 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 14756 35252 14766
rect 35084 14754 35252 14756
rect 35084 14702 35198 14754
rect 35250 14702 35252 14754
rect 35084 14700 35252 14702
rect 35196 14690 35252 14700
rect 33964 14532 34020 14542
rect 34524 14532 34580 14542
rect 33852 14530 34580 14532
rect 33852 14478 33966 14530
rect 34018 14478 34526 14530
rect 34578 14478 34580 14530
rect 33852 14476 34580 14478
rect 33516 13694 33518 13746
rect 33570 13694 33572 13746
rect 33516 13682 33572 13694
rect 33740 13858 33796 13870
rect 33740 13806 33742 13858
rect 33794 13806 33796 13858
rect 32060 12964 32116 12974
rect 32508 12964 32564 12974
rect 33068 12964 33124 12974
rect 32060 12962 33068 12964
rect 32060 12910 32062 12962
rect 32114 12910 32510 12962
rect 32562 12910 33068 12962
rect 32060 12908 33068 12910
rect 32060 12898 32116 12908
rect 32508 12898 32564 12908
rect 31500 12740 31556 12750
rect 31500 10722 31556 12684
rect 32060 12628 32116 12638
rect 31724 11844 31780 11854
rect 31724 11284 31780 11788
rect 31948 11732 32004 11742
rect 31948 11618 32004 11676
rect 31948 11566 31950 11618
rect 32002 11566 32004 11618
rect 31948 11554 32004 11566
rect 31724 11218 31780 11228
rect 32060 11284 32116 12572
rect 32508 12292 32564 12302
rect 32508 12198 32564 12236
rect 32284 12180 32340 12190
rect 32284 12178 32452 12180
rect 32284 12126 32286 12178
rect 32338 12126 32452 12178
rect 32284 12124 32452 12126
rect 32284 12114 32340 12124
rect 32396 11732 32452 12124
rect 33068 12178 33124 12908
rect 33740 12628 33796 13806
rect 33852 12964 33908 14476
rect 33964 14466 34020 14476
rect 34524 14466 34580 14476
rect 35532 14530 35588 14542
rect 35532 14478 35534 14530
rect 35586 14478 35588 14530
rect 33852 12898 33908 12908
rect 34188 13858 34244 13870
rect 34188 13806 34190 13858
rect 34242 13806 34244 13858
rect 33740 12562 33796 12572
rect 33852 12292 33908 12302
rect 33852 12198 33908 12236
rect 33068 12126 33070 12178
rect 33122 12126 33124 12178
rect 33068 12114 33124 12126
rect 34188 12068 34244 13806
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35532 13076 35588 14478
rect 35644 14420 35700 15036
rect 35756 14420 35812 14430
rect 35644 14418 35812 14420
rect 35644 14366 35758 14418
rect 35810 14366 35812 14418
rect 35644 14364 35812 14366
rect 35868 14420 35924 15092
rect 36092 14420 36148 14430
rect 35868 14418 36148 14420
rect 35868 14366 36094 14418
rect 36146 14366 36148 14418
rect 35868 14364 36148 14366
rect 35756 14354 35812 14364
rect 36092 14354 36148 14364
rect 35644 13748 35700 13758
rect 35644 13654 35700 13692
rect 35980 13748 36036 13758
rect 36204 13748 36260 15092
rect 36316 13858 36372 15484
rect 37884 15428 37940 15438
rect 37884 15334 37940 15372
rect 38668 15316 38724 17388
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 39116 15316 39172 15326
rect 38668 15314 39172 15316
rect 38668 15262 38670 15314
rect 38722 15262 39118 15314
rect 39170 15262 39172 15314
rect 38668 15260 39172 15262
rect 38668 15250 38724 15260
rect 36316 13806 36318 13858
rect 36370 13806 36372 13858
rect 36316 13794 36372 13806
rect 36540 13858 36596 13870
rect 36540 13806 36542 13858
rect 36594 13806 36596 13858
rect 35980 13746 36260 13748
rect 35980 13694 35982 13746
rect 36034 13694 36260 13746
rect 35980 13692 36260 13694
rect 35980 13682 36036 13692
rect 35532 13020 35700 13076
rect 32396 11676 33236 11732
rect 33180 11618 33236 11676
rect 33180 11566 33182 11618
rect 33234 11566 33236 11618
rect 33180 11554 33236 11566
rect 33516 11620 33572 11630
rect 33516 11526 33572 11564
rect 32060 11190 32116 11228
rect 32284 11282 32340 11294
rect 32284 11230 32286 11282
rect 32338 11230 32340 11282
rect 31500 10670 31502 10722
rect 31554 10670 31556 10722
rect 31500 10658 31556 10670
rect 32060 10724 32116 10734
rect 32284 10724 32340 11230
rect 34188 11282 34244 12012
rect 35532 12850 35588 12862
rect 35532 12798 35534 12850
rect 35586 12798 35588 12850
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 11620 35252 11630
rect 35532 11620 35588 12798
rect 35196 11618 35588 11620
rect 35196 11566 35198 11618
rect 35250 11566 35588 11618
rect 35196 11564 35588 11566
rect 35196 11554 35252 11564
rect 34188 11230 34190 11282
rect 34242 11230 34244 11282
rect 34188 11218 34244 11230
rect 34300 11394 34356 11406
rect 34300 11342 34302 11394
rect 34354 11342 34356 11394
rect 34300 11284 34356 11342
rect 34300 11218 34356 11228
rect 35532 11396 35588 11406
rect 35644 11396 35700 13020
rect 36316 12964 36372 12974
rect 36316 12870 36372 12908
rect 35868 12740 35924 12750
rect 35868 12646 35924 12684
rect 36540 12404 36596 13806
rect 36316 12348 36596 12404
rect 38444 12740 38500 12750
rect 35980 12068 36036 12078
rect 35980 11974 36036 12012
rect 36316 12066 36372 12348
rect 38444 12290 38500 12684
rect 38444 12238 38446 12290
rect 38498 12238 38500 12290
rect 38444 12226 38500 12238
rect 39116 12404 39172 15260
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 39676 12404 39732 12414
rect 39116 12402 39732 12404
rect 39116 12350 39678 12402
rect 39730 12350 39732 12402
rect 39116 12348 39732 12350
rect 39116 12178 39172 12348
rect 39676 12338 39732 12348
rect 39116 12126 39118 12178
rect 39170 12126 39172 12178
rect 39116 12114 39172 12126
rect 36316 12014 36318 12066
rect 36370 12014 36372 12066
rect 35532 11394 35700 11396
rect 35532 11342 35534 11394
rect 35586 11342 35700 11394
rect 35532 11340 35700 11342
rect 32060 10722 32340 10724
rect 32060 10670 32062 10722
rect 32114 10670 32340 10722
rect 32060 10668 32340 10670
rect 31276 10610 31444 10612
rect 31276 10558 31278 10610
rect 31330 10558 31444 10610
rect 31276 10556 31444 10558
rect 31276 10546 31332 10556
rect 31388 10388 31444 10556
rect 31388 10322 31444 10332
rect 31052 9886 31054 9938
rect 31106 9886 31108 9938
rect 31052 9874 31108 9886
rect 32060 9940 32116 10668
rect 35532 10388 35588 11340
rect 35756 11284 35812 11294
rect 35756 11190 35812 11228
rect 36316 11282 36372 12014
rect 36316 11230 36318 11282
rect 36370 11230 36372 11282
rect 36316 11218 36372 11230
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 35532 10322 35588 10332
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 33180 9940 33236 9950
rect 32060 9938 33236 9940
rect 32060 9886 33182 9938
rect 33234 9886 33236 9938
rect 32060 9884 33236 9886
rect 33180 9874 33236 9884
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 30604 8878 30606 8930
rect 30658 8878 30660 8930
rect 30604 8866 30660 8878
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 29036 8372 29204 8428
rect 29148 7698 29204 8372
rect 30156 8372 30324 8428
rect 29932 8260 29988 8270
rect 30156 8260 30212 8372
rect 29988 8204 30212 8260
rect 29932 8166 29988 8204
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 29148 7646 29150 7698
rect 29202 7646 29204 7698
rect 29148 7634 29204 7646
rect 28252 7588 28308 7598
rect 28252 7494 28308 7532
rect 28700 7586 28756 7598
rect 28700 7534 28702 7586
rect 28754 7534 28756 7586
rect 27916 7422 27918 7474
rect 27970 7422 27972 7474
rect 27916 7410 27972 7422
rect 28700 7364 28756 7534
rect 29260 7364 29316 7374
rect 28700 7362 29316 7364
rect 28700 7310 29262 7362
rect 29314 7310 29316 7362
rect 28700 7308 29316 7310
rect 27580 7252 27636 7262
rect 27580 7250 27860 7252
rect 27580 7198 27582 7250
rect 27634 7198 27860 7250
rect 27580 7196 27860 7198
rect 27580 7186 27636 7196
rect 27244 5906 27300 6748
rect 27468 6916 27524 6926
rect 27468 6802 27524 6860
rect 27468 6750 27470 6802
rect 27522 6750 27524 6802
rect 27468 6738 27524 6750
rect 27804 6690 27860 7196
rect 28588 6804 28644 6814
rect 28588 6710 28644 6748
rect 27804 6638 27806 6690
rect 27858 6638 27860 6690
rect 27804 6626 27860 6638
rect 28140 6468 28196 6478
rect 28028 6466 28196 6468
rect 28028 6414 28142 6466
rect 28194 6414 28196 6466
rect 28028 6412 28196 6414
rect 28028 6018 28084 6412
rect 28140 6402 28196 6412
rect 28028 5966 28030 6018
rect 28082 5966 28084 6018
rect 28028 5954 28084 5966
rect 27244 5854 27246 5906
rect 27298 5854 27300 5906
rect 24892 5234 25060 5236
rect 24892 5182 24894 5234
rect 24946 5182 25060 5234
rect 24892 5180 25060 5182
rect 25340 5236 25396 5246
rect 24892 5170 24948 5180
rect 25340 5142 25396 5180
rect 26796 5236 26852 5246
rect 26908 5236 26964 5246
rect 27244 5236 27300 5854
rect 29260 5796 29316 7308
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 30156 5796 30212 5806
rect 29260 5794 30212 5796
rect 29260 5742 30158 5794
rect 30210 5742 30212 5794
rect 29260 5740 30212 5742
rect 30156 5730 30212 5740
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 26852 5234 27300 5236
rect 26852 5182 26910 5234
rect 26962 5182 27300 5234
rect 26852 5180 27300 5182
rect 26796 5170 26852 5180
rect 26908 5170 26964 5180
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 23772 4510 23774 4562
rect 23826 4510 23828 4562
rect 23772 4498 23828 4510
rect 23324 4226 23492 4228
rect 23324 4174 23326 4226
rect 23378 4174 23492 4226
rect 23324 4172 23492 4174
rect 23324 4162 23380 4172
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
<< via2 >>
rect 4620 56306 4676 56308
rect 4620 56254 4622 56306
rect 4622 56254 4674 56306
rect 4674 56254 4676 56306
rect 4620 56252 4676 56254
rect 5516 56252 5572 56308
rect 5852 56194 5908 56196
rect 5852 56142 5854 56194
rect 5854 56142 5906 56194
rect 5906 56142 5908 56194
rect 5852 56140 5908 56142
rect 8428 56140 8484 56196
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4060 54796 4116 54852
rect 2380 54626 2436 54628
rect 2380 54574 2382 54626
rect 2382 54574 2434 54626
rect 2434 54574 2436 54626
rect 2380 54572 2436 54574
rect 3612 53676 3668 53732
rect 2492 52050 2548 52052
rect 2492 51998 2494 52050
rect 2494 51998 2546 52050
rect 2546 51998 2548 52050
rect 2492 51996 2548 51998
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 6972 54572 7028 54628
rect 4956 53676 5012 53732
rect 3836 52946 3892 52948
rect 3836 52894 3838 52946
rect 3838 52894 3890 52946
rect 3890 52894 3892 52946
rect 3836 52892 3892 52894
rect 4620 52946 4676 52948
rect 4620 52894 4622 52946
rect 4622 52894 4674 52946
rect 4674 52894 4676 52946
rect 4620 52892 4676 52894
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4844 52220 4900 52276
rect 4620 52108 4676 52164
rect 3724 51884 3780 51940
rect 4508 51996 4564 52052
rect 5180 53676 5236 53732
rect 5068 52444 5124 52500
rect 4956 52108 5012 52164
rect 4844 51154 4900 51156
rect 4844 51102 4846 51154
rect 4846 51102 4898 51154
rect 4898 51102 4900 51154
rect 4844 51100 4900 51102
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 2492 50428 2548 50484
rect 4620 49698 4676 49700
rect 4620 49646 4622 49698
rect 4622 49646 4674 49698
rect 4674 49646 4676 49698
rect 4620 49644 4676 49646
rect 5628 52162 5684 52164
rect 5628 52110 5630 52162
rect 5630 52110 5682 52162
rect 5682 52110 5684 52162
rect 5628 52108 5684 52110
rect 5740 51884 5796 51940
rect 5740 51100 5796 51156
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 1820 48636 1876 48692
rect 4732 48748 4788 48804
rect 2828 48524 2884 48580
rect 2940 48130 2996 48132
rect 2940 48078 2942 48130
rect 2942 48078 2994 48130
rect 2994 48078 2996 48130
rect 2940 48076 2996 48078
rect 3836 48076 3892 48132
rect 1596 46620 1652 46676
rect 5068 48636 5124 48692
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 5628 50482 5684 50484
rect 5628 50430 5630 50482
rect 5630 50430 5682 50482
rect 5682 50430 5684 50482
rect 5628 50428 5684 50430
rect 5740 50316 5796 50372
rect 6524 52946 6580 52948
rect 6524 52894 6526 52946
rect 6526 52894 6578 52946
rect 6578 52894 6580 52946
rect 6524 52892 6580 52894
rect 6748 53730 6804 53732
rect 6748 53678 6750 53730
rect 6750 53678 6802 53730
rect 6802 53678 6804 53730
rect 6748 53676 6804 53678
rect 7644 54626 7700 54628
rect 7644 54574 7646 54626
rect 7646 54574 7698 54626
rect 7698 54574 7700 54626
rect 7644 54572 7700 54574
rect 6748 52780 6804 52836
rect 6412 52444 6468 52500
rect 6972 52444 7028 52500
rect 7532 53116 7588 53172
rect 6636 51100 6692 51156
rect 6076 50316 6132 50372
rect 6188 50204 6244 50260
rect 5740 49810 5796 49812
rect 5740 49758 5742 49810
rect 5742 49758 5794 49810
rect 5794 49758 5796 49810
rect 5740 49756 5796 49758
rect 5404 48300 5460 48356
rect 5516 49698 5572 49700
rect 5516 49646 5518 49698
rect 5518 49646 5570 49698
rect 5570 49646 5572 49698
rect 5516 49644 5572 49646
rect 6076 49026 6132 49028
rect 6076 48974 6078 49026
rect 6078 48974 6130 49026
rect 6130 48974 6132 49026
rect 6076 48972 6132 48974
rect 6076 48748 6132 48804
rect 6188 48860 6244 48916
rect 6300 48300 6356 48356
rect 6636 48972 6692 49028
rect 6860 50316 6916 50372
rect 7420 52780 7476 52836
rect 7532 52946 7588 52948
rect 7532 52894 7534 52946
rect 7534 52894 7586 52946
rect 7586 52894 7588 52946
rect 7532 52892 7588 52894
rect 8316 52780 8372 52836
rect 7756 52220 7812 52276
rect 8092 51212 8148 51268
rect 7196 50204 7252 50260
rect 7084 49810 7140 49812
rect 7084 49758 7086 49810
rect 7086 49758 7138 49810
rect 7138 49758 7140 49810
rect 7084 49756 7140 49758
rect 7308 49644 7364 49700
rect 6972 48524 7028 48580
rect 7084 48748 7140 48804
rect 6636 48300 6692 48356
rect 6524 48188 6580 48244
rect 6412 48076 6468 48132
rect 2268 46786 2324 46788
rect 2268 46734 2270 46786
rect 2270 46734 2322 46786
rect 2322 46734 2324 46786
rect 2268 46732 2324 46734
rect 3276 46732 3332 46788
rect 2156 46620 2212 46676
rect 1708 45500 1764 45556
rect 2604 45500 2660 45556
rect 2492 45388 2548 45444
rect 2044 45052 2100 45108
rect 2380 44492 2436 44548
rect 4508 46786 4564 46788
rect 4508 46734 4510 46786
rect 4510 46734 4562 46786
rect 4562 46734 4564 46786
rect 4508 46732 4564 46734
rect 4172 46674 4228 46676
rect 4172 46622 4174 46674
rect 4174 46622 4226 46674
rect 4226 46622 4228 46674
rect 4172 46620 4228 46622
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 3948 45388 4004 45444
rect 5068 45276 5124 45332
rect 5404 45836 5460 45892
rect 6972 47964 7028 48020
rect 6636 47852 6692 47908
rect 15708 56194 15764 56196
rect 15708 56142 15710 56194
rect 15710 56142 15762 56194
rect 15762 56142 15764 56194
rect 15708 56140 15764 56142
rect 9100 54796 9156 54852
rect 8764 51266 8820 51268
rect 8764 51214 8766 51266
rect 8766 51214 8818 51266
rect 8818 51214 8820 51266
rect 8764 51212 8820 51214
rect 8876 50482 8932 50484
rect 8876 50430 8878 50482
rect 8878 50430 8930 50482
rect 8930 50430 8932 50482
rect 8876 50428 8932 50430
rect 7420 48860 7476 48916
rect 8092 49084 8148 49140
rect 7756 48300 7812 48356
rect 7308 47852 7364 47908
rect 3724 45106 3780 45108
rect 3724 45054 3726 45106
rect 3726 45054 3778 45106
rect 3778 45054 3780 45106
rect 3724 45052 3780 45054
rect 3276 44546 3332 44548
rect 3276 44494 3278 44546
rect 3278 44494 3330 44546
rect 3330 44494 3332 44546
rect 3276 44492 3332 44494
rect 4172 44492 4228 44548
rect 3052 44156 3108 44212
rect 1932 43820 1988 43876
rect 3836 44322 3892 44324
rect 3836 44270 3838 44322
rect 3838 44270 3890 44322
rect 3890 44270 3892 44322
rect 3836 44268 3892 44270
rect 3724 43820 3780 43876
rect 4060 43932 4116 43988
rect 3612 43372 3668 43428
rect 1820 42476 1876 42532
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4620 44434 4676 44436
rect 4620 44382 4622 44434
rect 4622 44382 4674 44434
rect 4674 44382 4676 44434
rect 4620 44380 4676 44382
rect 4956 44268 5012 44324
rect 4732 43932 4788 43988
rect 4396 43596 4452 43652
rect 5068 43650 5124 43652
rect 5068 43598 5070 43650
rect 5070 43598 5122 43650
rect 5122 43598 5124 43650
rect 5068 43596 5124 43598
rect 4620 43538 4676 43540
rect 4620 43486 4622 43538
rect 4622 43486 4674 43538
rect 4674 43486 4676 43538
rect 4620 43484 4676 43486
rect 4956 43426 5012 43428
rect 4956 43374 4958 43426
rect 4958 43374 5010 43426
rect 5010 43374 5012 43426
rect 4956 43372 5012 43374
rect 4844 43260 4900 43316
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 3948 41804 4004 41860
rect 4172 41804 4228 41860
rect 3836 41692 3892 41748
rect 3612 40962 3668 40964
rect 3612 40910 3614 40962
rect 3614 40910 3666 40962
rect 3666 40910 3668 40962
rect 3612 40908 3668 40910
rect 4620 41692 4676 41748
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 6972 45890 7028 45892
rect 6972 45838 6974 45890
rect 6974 45838 7026 45890
rect 7026 45838 7028 45890
rect 6972 45836 7028 45838
rect 7196 45778 7252 45780
rect 7196 45726 7198 45778
rect 7198 45726 7250 45778
rect 7250 45726 7252 45778
rect 7196 45724 7252 45726
rect 6860 45612 6916 45668
rect 5516 43260 5572 43316
rect 5628 44268 5684 44324
rect 5740 44210 5796 44212
rect 5740 44158 5742 44210
rect 5742 44158 5794 44210
rect 5794 44158 5796 44210
rect 5740 44156 5796 44158
rect 5964 45276 6020 45332
rect 5964 43372 6020 43428
rect 8092 48130 8148 48132
rect 8092 48078 8094 48130
rect 8094 48078 8146 48130
rect 8146 48078 8148 48130
rect 8092 48076 8148 48078
rect 7980 48018 8036 48020
rect 7980 47966 7982 48018
rect 7982 47966 8034 48018
rect 8034 47966 8036 48018
rect 7980 47964 8036 47966
rect 7644 45666 7700 45668
rect 7644 45614 7646 45666
rect 7646 45614 7698 45666
rect 7698 45614 7700 45666
rect 7644 45612 7700 45614
rect 7532 44940 7588 44996
rect 6300 44322 6356 44324
rect 6300 44270 6302 44322
rect 6302 44270 6354 44322
rect 6354 44270 6356 44322
rect 6300 44268 6356 44270
rect 6076 43484 6132 43540
rect 4956 42530 5012 42532
rect 4956 42478 4958 42530
rect 4958 42478 5010 42530
rect 5010 42478 5012 42530
rect 4956 42476 5012 42478
rect 4956 42028 5012 42084
rect 4956 41858 5012 41860
rect 4956 41806 4958 41858
rect 4958 41806 5010 41858
rect 5010 41806 5012 41858
rect 4956 41804 5012 41806
rect 4844 41244 4900 41300
rect 4284 41186 4340 41188
rect 4284 41134 4286 41186
rect 4286 41134 4338 41186
rect 4338 41134 4340 41186
rect 4284 41132 4340 41134
rect 4732 41132 4788 41188
rect 4172 40908 4228 40964
rect 2492 40572 2548 40628
rect 4508 40626 4564 40628
rect 4508 40574 4510 40626
rect 4510 40574 4562 40626
rect 4562 40574 4564 40626
rect 4508 40572 4564 40574
rect 3948 39564 4004 39620
rect 2828 39004 2884 39060
rect 1820 38668 1876 38724
rect 2492 38780 2548 38836
rect 3052 38946 3108 38948
rect 3052 38894 3054 38946
rect 3054 38894 3106 38946
rect 3106 38894 3108 38946
rect 3052 38892 3108 38894
rect 3724 38946 3780 38948
rect 3724 38894 3726 38946
rect 3726 38894 3778 38946
rect 3778 38894 3780 38946
rect 3724 38892 3780 38894
rect 3500 38834 3556 38836
rect 3500 38782 3502 38834
rect 3502 38782 3554 38834
rect 3554 38782 3556 38834
rect 3500 38780 3556 38782
rect 4620 40178 4676 40180
rect 4620 40126 4622 40178
rect 4622 40126 4674 40178
rect 4674 40126 4676 40178
rect 4620 40124 4676 40126
rect 5292 41356 5348 41412
rect 5516 41244 5572 41300
rect 4844 40402 4900 40404
rect 4844 40350 4846 40402
rect 4846 40350 4898 40402
rect 4898 40350 4900 40402
rect 4844 40348 4900 40350
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4620 39730 4676 39732
rect 4620 39678 4622 39730
rect 4622 39678 4674 39730
rect 4674 39678 4676 39730
rect 4620 39676 4676 39678
rect 4508 38946 4564 38948
rect 4508 38894 4510 38946
rect 4510 38894 4562 38946
rect 4562 38894 4564 38946
rect 4508 38892 4564 38894
rect 6076 42028 6132 42084
rect 5964 41804 6020 41860
rect 6076 41356 6132 41412
rect 5852 40348 5908 40404
rect 6188 41186 6244 41188
rect 6188 41134 6190 41186
rect 6190 41134 6242 41186
rect 6242 41134 6244 41186
rect 6188 41132 6244 41134
rect 6524 40460 6580 40516
rect 6412 40348 6468 40404
rect 6076 40124 6132 40180
rect 4844 39116 4900 39172
rect 4956 39676 5012 39732
rect 5516 39676 5572 39732
rect 5068 39394 5124 39396
rect 5068 39342 5070 39394
rect 5070 39342 5122 39394
rect 5122 39342 5124 39394
rect 5068 39340 5124 39342
rect 5068 38668 5124 38724
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4620 38220 4676 38276
rect 4620 37378 4676 37380
rect 4620 37326 4622 37378
rect 4622 37326 4674 37378
rect 4674 37326 4676 37378
rect 4620 37324 4676 37326
rect 5180 38892 5236 38948
rect 5852 39004 5908 39060
rect 5516 38946 5572 38948
rect 5516 38894 5518 38946
rect 5518 38894 5570 38946
rect 5570 38894 5572 38946
rect 5516 38892 5572 38894
rect 6300 39452 6356 39508
rect 5852 38780 5908 38836
rect 6300 38892 6356 38948
rect 6076 38780 6132 38836
rect 6636 39564 6692 39620
rect 8428 48300 8484 48356
rect 8316 48242 8372 48244
rect 8316 48190 8318 48242
rect 8318 48190 8370 48242
rect 8370 48190 8372 48242
rect 8316 48188 8372 48190
rect 8204 45276 8260 45332
rect 6860 41916 6916 41972
rect 8428 41970 8484 41972
rect 8428 41918 8430 41970
rect 8430 41918 8482 41970
rect 8482 41918 8484 41970
rect 8428 41916 8484 41918
rect 6860 41410 6916 41412
rect 6860 41358 6862 41410
rect 6862 41358 6914 41410
rect 6914 41358 6916 41410
rect 6860 41356 6916 41358
rect 7084 41244 7140 41300
rect 6972 41186 7028 41188
rect 6972 41134 6974 41186
rect 6974 41134 7026 41186
rect 7026 41134 7028 41186
rect 6972 41132 7028 41134
rect 7644 40514 7700 40516
rect 7644 40462 7646 40514
rect 7646 40462 7698 40514
rect 7698 40462 7700 40514
rect 7644 40460 7700 40462
rect 16268 55132 16324 55188
rect 17052 56140 17108 56196
rect 16828 55468 16884 55524
rect 16940 55356 16996 55412
rect 16828 55186 16884 55188
rect 16828 55134 16830 55186
rect 16830 55134 16882 55186
rect 16882 55134 16884 55186
rect 16828 55132 16884 55134
rect 16604 54738 16660 54740
rect 16604 54686 16606 54738
rect 16606 54686 16658 54738
rect 16658 54686 16660 54738
rect 16604 54684 16660 54686
rect 9660 53842 9716 53844
rect 9660 53790 9662 53842
rect 9662 53790 9714 53842
rect 9714 53790 9716 53842
rect 9660 53788 9716 53790
rect 11452 53788 11508 53844
rect 10780 53618 10836 53620
rect 10780 53566 10782 53618
rect 10782 53566 10834 53618
rect 10834 53566 10836 53618
rect 10780 53564 10836 53566
rect 9996 53116 10052 53172
rect 10444 52444 10500 52500
rect 10892 52444 10948 52500
rect 10332 52162 10388 52164
rect 10332 52110 10334 52162
rect 10334 52110 10386 52162
rect 10386 52110 10388 52162
rect 10332 52108 10388 52110
rect 11564 53058 11620 53060
rect 11564 53006 11566 53058
rect 11566 53006 11618 53058
rect 11618 53006 11620 53058
rect 11564 53004 11620 53006
rect 11676 52722 11732 52724
rect 11676 52670 11678 52722
rect 11678 52670 11730 52722
rect 11730 52670 11732 52722
rect 11676 52668 11732 52670
rect 11564 52162 11620 52164
rect 11564 52110 11566 52162
rect 11566 52110 11618 52162
rect 11618 52110 11620 52162
rect 11564 52108 11620 52110
rect 11788 51884 11844 51940
rect 12908 53676 12964 53732
rect 12796 53004 12852 53060
rect 12460 52668 12516 52724
rect 12460 52220 12516 52276
rect 12572 52162 12628 52164
rect 12572 52110 12574 52162
rect 12574 52110 12626 52162
rect 12626 52110 12628 52162
rect 12572 52108 12628 52110
rect 13020 52834 13076 52836
rect 13020 52782 13022 52834
rect 13022 52782 13074 52834
rect 13074 52782 13076 52834
rect 13020 52780 13076 52782
rect 12908 52444 12964 52500
rect 12460 51884 12516 51940
rect 9660 51212 9716 51268
rect 12124 50540 12180 50596
rect 11004 50316 11060 50372
rect 11900 50482 11956 50484
rect 11900 50430 11902 50482
rect 11902 50430 11954 50482
rect 11954 50430 11956 50482
rect 11900 50428 11956 50430
rect 11788 50316 11844 50372
rect 11340 49138 11396 49140
rect 11340 49086 11342 49138
rect 11342 49086 11394 49138
rect 11394 49086 11396 49138
rect 11340 49084 11396 49086
rect 11340 48412 11396 48468
rect 8764 44994 8820 44996
rect 8764 44942 8766 44994
rect 8766 44942 8818 44994
rect 8818 44942 8820 44994
rect 8764 44940 8820 44942
rect 8876 43596 8932 43652
rect 8876 43260 8932 43316
rect 8988 42140 9044 42196
rect 8876 41970 8932 41972
rect 8876 41918 8878 41970
rect 8878 41918 8930 41970
rect 8930 41918 8932 41970
rect 8876 41916 8932 41918
rect 8540 40572 8596 40628
rect 7196 39564 7252 39620
rect 7532 39506 7588 39508
rect 7532 39454 7534 39506
rect 7534 39454 7586 39506
rect 7586 39454 7588 39506
rect 7532 39452 7588 39454
rect 8316 39394 8372 39396
rect 8316 39342 8318 39394
rect 8318 39342 8370 39394
rect 8370 39342 8372 39394
rect 8316 39340 8372 39342
rect 6860 39116 6916 39172
rect 6748 39004 6804 39060
rect 6860 38834 6916 38836
rect 6860 38782 6862 38834
rect 6862 38782 6914 38834
rect 6914 38782 6916 38834
rect 6860 38780 6916 38782
rect 7756 39058 7812 39060
rect 7756 39006 7758 39058
rect 7758 39006 7810 39058
rect 7810 39006 7812 39058
rect 7756 39004 7812 39006
rect 7532 38834 7588 38836
rect 7532 38782 7534 38834
rect 7534 38782 7586 38834
rect 7586 38782 7588 38834
rect 7532 38780 7588 38782
rect 9996 48018 10052 48020
rect 9996 47966 9998 48018
rect 9998 47966 10050 48018
rect 10050 47966 10052 48018
rect 9996 47964 10052 47966
rect 10108 46396 10164 46452
rect 10668 47964 10724 48020
rect 9772 45778 9828 45780
rect 9772 45726 9774 45778
rect 9774 45726 9826 45778
rect 9826 45726 9828 45778
rect 9772 45724 9828 45726
rect 9660 45330 9716 45332
rect 9660 45278 9662 45330
rect 9662 45278 9714 45330
rect 9714 45278 9716 45330
rect 9660 45276 9716 45278
rect 11228 46562 11284 46564
rect 11228 46510 11230 46562
rect 11230 46510 11282 46562
rect 11282 46510 11284 46562
rect 11228 46508 11284 46510
rect 10444 46284 10500 46340
rect 13468 53730 13524 53732
rect 13468 53678 13470 53730
rect 13470 53678 13522 53730
rect 13522 53678 13524 53730
rect 13468 53676 13524 53678
rect 14364 53564 14420 53620
rect 13356 52444 13412 52500
rect 13580 51884 13636 51940
rect 12908 51100 12964 51156
rect 12460 50652 12516 50708
rect 12796 50594 12852 50596
rect 12796 50542 12798 50594
rect 12798 50542 12850 50594
rect 12850 50542 12852 50594
rect 12796 50540 12852 50542
rect 13580 51100 13636 51156
rect 13468 50594 13524 50596
rect 13468 50542 13470 50594
rect 13470 50542 13522 50594
rect 13522 50542 13524 50594
rect 13468 50540 13524 50542
rect 13804 52444 13860 52500
rect 14252 52834 14308 52836
rect 14252 52782 14254 52834
rect 14254 52782 14306 52834
rect 14306 52782 14308 52834
rect 14252 52780 14308 52782
rect 13916 51884 13972 51940
rect 13804 51212 13860 51268
rect 14252 51212 14308 51268
rect 16940 54290 16996 54292
rect 16940 54238 16942 54290
rect 16942 54238 16994 54290
rect 16994 54238 16996 54290
rect 16940 54236 16996 54238
rect 17612 56194 17668 56196
rect 17612 56142 17614 56194
rect 17614 56142 17666 56194
rect 17666 56142 17668 56194
rect 17612 56140 17668 56142
rect 17948 56140 18004 56196
rect 17500 56028 17556 56084
rect 17500 55468 17556 55524
rect 18620 56194 18676 56196
rect 18620 56142 18622 56194
rect 18622 56142 18674 56194
rect 18674 56142 18676 56194
rect 18620 56140 18676 56142
rect 17276 54236 17332 54292
rect 17500 53954 17556 53956
rect 17500 53902 17502 53954
rect 17502 53902 17554 53954
rect 17554 53902 17556 53954
rect 17500 53900 17556 53902
rect 17276 53730 17332 53732
rect 17276 53678 17278 53730
rect 17278 53678 17330 53730
rect 17330 53678 17332 53730
rect 17276 53676 17332 53678
rect 14588 52162 14644 52164
rect 14588 52110 14590 52162
rect 14590 52110 14642 52162
rect 14642 52110 14644 52162
rect 14588 52108 14644 52110
rect 14812 51884 14868 51940
rect 14588 51100 14644 51156
rect 14476 50652 14532 50708
rect 12460 49756 12516 49812
rect 12348 49084 12404 49140
rect 12460 49420 12516 49476
rect 12124 48860 12180 48916
rect 11564 46732 11620 46788
rect 11676 48300 11732 48356
rect 12012 46674 12068 46676
rect 12012 46622 12014 46674
rect 12014 46622 12066 46674
rect 12066 46622 12068 46674
rect 12012 46620 12068 46622
rect 11900 46562 11956 46564
rect 11900 46510 11902 46562
rect 11902 46510 11954 46562
rect 11954 46510 11956 46562
rect 11900 46508 11956 46510
rect 11228 46284 11284 46340
rect 11004 45836 11060 45892
rect 10556 45724 10612 45780
rect 10444 45106 10500 45108
rect 10444 45054 10446 45106
rect 10446 45054 10498 45106
rect 10498 45054 10500 45106
rect 10444 45052 10500 45054
rect 10780 45612 10836 45668
rect 10892 45276 10948 45332
rect 10108 43650 10164 43652
rect 10108 43598 10110 43650
rect 10110 43598 10162 43650
rect 10162 43598 10164 43650
rect 10108 43596 10164 43598
rect 10220 43484 10276 43540
rect 10668 44044 10724 44100
rect 10220 42252 10276 42308
rect 9660 41970 9716 41972
rect 9660 41918 9662 41970
rect 9662 41918 9714 41970
rect 9714 41918 9716 41970
rect 9660 41916 9716 41918
rect 11228 45500 11284 45556
rect 12236 48188 12292 48244
rect 12796 49196 12852 49252
rect 12684 49026 12740 49028
rect 12684 48974 12686 49026
rect 12686 48974 12738 49026
rect 12738 48974 12740 49026
rect 12684 48972 12740 48974
rect 12908 49084 12964 49140
rect 12684 47852 12740 47908
rect 12348 46844 12404 46900
rect 12684 46956 12740 47012
rect 11564 45612 11620 45668
rect 12124 45836 12180 45892
rect 11452 45388 11508 45444
rect 11340 45164 11396 45220
rect 11228 45052 11284 45108
rect 11004 43708 11060 43764
rect 11228 43538 11284 43540
rect 11228 43486 11230 43538
rect 11230 43486 11282 43538
rect 11282 43486 11284 43538
rect 11228 43484 11284 43486
rect 11116 43372 11172 43428
rect 11004 42866 11060 42868
rect 11004 42814 11006 42866
rect 11006 42814 11058 42866
rect 11058 42814 11060 42866
rect 11004 42812 11060 42814
rect 11788 45666 11844 45668
rect 11788 45614 11790 45666
rect 11790 45614 11842 45666
rect 11842 45614 11844 45666
rect 11788 45612 11844 45614
rect 12012 45388 12068 45444
rect 11900 45276 11956 45332
rect 11788 45164 11844 45220
rect 12572 45890 12628 45892
rect 12572 45838 12574 45890
rect 12574 45838 12626 45890
rect 12626 45838 12628 45890
rect 12572 45836 12628 45838
rect 13132 47292 13188 47348
rect 13020 47234 13076 47236
rect 13020 47182 13022 47234
rect 13022 47182 13074 47234
rect 13074 47182 13076 47234
rect 13020 47180 13076 47182
rect 12796 45836 12852 45892
rect 12684 45388 12740 45444
rect 13020 45388 13076 45444
rect 12684 45052 12740 45108
rect 12460 44268 12516 44324
rect 11788 43708 11844 43764
rect 11340 42700 11396 42756
rect 11788 43484 11844 43540
rect 12124 43762 12180 43764
rect 12124 43710 12126 43762
rect 12126 43710 12178 43762
rect 12178 43710 12180 43762
rect 12124 43708 12180 43710
rect 12684 44434 12740 44436
rect 12684 44382 12686 44434
rect 12686 44382 12738 44434
rect 12738 44382 12740 44434
rect 12684 44380 12740 44382
rect 12012 43484 12068 43540
rect 11564 41804 11620 41860
rect 12236 41858 12292 41860
rect 12236 41806 12238 41858
rect 12238 41806 12290 41858
rect 12290 41806 12292 41858
rect 12236 41804 12292 41806
rect 12572 41804 12628 41860
rect 13356 49420 13412 49476
rect 13804 49756 13860 49812
rect 13916 48972 13972 49028
rect 14364 49810 14420 49812
rect 14364 49758 14366 49810
rect 14366 49758 14418 49810
rect 14418 49758 14420 49810
rect 14364 49756 14420 49758
rect 13692 48748 13748 48804
rect 14140 47852 14196 47908
rect 13692 46956 13748 47012
rect 13916 47346 13972 47348
rect 13916 47294 13918 47346
rect 13918 47294 13970 47346
rect 13970 47294 13972 47346
rect 13916 47292 13972 47294
rect 13468 46844 13524 46900
rect 13468 46396 13524 46452
rect 13468 45276 13524 45332
rect 13580 45836 13636 45892
rect 13916 46732 13972 46788
rect 14028 46674 14084 46676
rect 14028 46622 14030 46674
rect 14030 46622 14082 46674
rect 14082 46622 14084 46674
rect 14028 46620 14084 46622
rect 15372 52220 15428 52276
rect 15484 52162 15540 52164
rect 15484 52110 15486 52162
rect 15486 52110 15538 52162
rect 15538 52110 15540 52162
rect 15484 52108 15540 52110
rect 15372 51490 15428 51492
rect 15372 51438 15374 51490
rect 15374 51438 15426 51490
rect 15426 51438 15428 51490
rect 15372 51436 15428 51438
rect 15260 51378 15316 51380
rect 15260 51326 15262 51378
rect 15262 51326 15314 51378
rect 15314 51326 15316 51378
rect 15260 51324 15316 51326
rect 15596 51378 15652 51380
rect 15596 51326 15598 51378
rect 15598 51326 15650 51378
rect 15650 51326 15652 51378
rect 15596 51324 15652 51326
rect 16492 51378 16548 51380
rect 16492 51326 16494 51378
rect 16494 51326 16546 51378
rect 16546 51326 16548 51378
rect 16492 51324 16548 51326
rect 16044 51266 16100 51268
rect 16044 51214 16046 51266
rect 16046 51214 16098 51266
rect 16098 51214 16100 51266
rect 16044 51212 16100 51214
rect 15036 50876 15092 50932
rect 14924 50482 14980 50484
rect 14924 50430 14926 50482
rect 14926 50430 14978 50482
rect 14978 50430 14980 50482
rect 14924 50428 14980 50430
rect 14812 49586 14868 49588
rect 14812 49534 14814 49586
rect 14814 49534 14866 49586
rect 14866 49534 14868 49586
rect 14812 49532 14868 49534
rect 16044 50988 16100 51044
rect 16268 51154 16324 51156
rect 16268 51102 16270 51154
rect 16270 51102 16322 51154
rect 16322 51102 16324 51154
rect 16268 51100 16324 51102
rect 14812 49196 14868 49252
rect 15148 48412 15204 48468
rect 14700 48242 14756 48244
rect 14700 48190 14702 48242
rect 14702 48190 14754 48242
rect 14754 48190 14756 48242
rect 14700 48188 14756 48190
rect 14588 47852 14644 47908
rect 15036 47628 15092 47684
rect 14588 47292 14644 47348
rect 14252 46562 14308 46564
rect 14252 46510 14254 46562
rect 14254 46510 14306 46562
rect 14306 46510 14308 46562
rect 14252 46508 14308 46510
rect 13916 46396 13972 46452
rect 14476 45724 14532 45780
rect 14140 45106 14196 45108
rect 14140 45054 14142 45106
rect 14142 45054 14194 45106
rect 14194 45054 14196 45106
rect 14140 45052 14196 45054
rect 14812 45890 14868 45892
rect 14812 45838 14814 45890
rect 14814 45838 14866 45890
rect 14866 45838 14868 45890
rect 14812 45836 14868 45838
rect 14700 45500 14756 45556
rect 15036 45500 15092 45556
rect 15820 49586 15876 49588
rect 15820 49534 15822 49586
rect 15822 49534 15874 49586
rect 15874 49534 15876 49586
rect 15820 49532 15876 49534
rect 15596 48354 15652 48356
rect 15596 48302 15598 48354
rect 15598 48302 15650 48354
rect 15650 48302 15652 48354
rect 15596 48300 15652 48302
rect 16156 48748 16212 48804
rect 15372 46060 15428 46116
rect 15372 45612 15428 45668
rect 15260 45500 15316 45556
rect 14812 45388 14868 45444
rect 15260 45276 15316 45332
rect 13804 44380 13860 44436
rect 13692 44098 13748 44100
rect 13692 44046 13694 44098
rect 13694 44046 13746 44098
rect 13746 44046 13748 44098
rect 13692 44044 13748 44046
rect 12908 43426 12964 43428
rect 12908 43374 12910 43426
rect 12910 43374 12962 43426
rect 12962 43374 12964 43426
rect 12908 43372 12964 43374
rect 13580 43148 13636 43204
rect 13580 42924 13636 42980
rect 13020 42812 13076 42868
rect 14476 44322 14532 44324
rect 14476 44270 14478 44322
rect 14478 44270 14530 44322
rect 14530 44270 14532 44322
rect 14476 44268 14532 44270
rect 15708 47740 15764 47796
rect 16492 51100 16548 51156
rect 17724 54684 17780 54740
rect 18284 55858 18340 55860
rect 18284 55806 18286 55858
rect 18286 55806 18338 55858
rect 18338 55806 18340 55858
rect 18284 55804 18340 55806
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 18844 55804 18900 55860
rect 18396 55468 18452 55524
rect 17948 54460 18004 54516
rect 18284 54514 18340 54516
rect 18284 54462 18286 54514
rect 18286 54462 18338 54514
rect 18338 54462 18340 54514
rect 18284 54460 18340 54462
rect 18844 55410 18900 55412
rect 18844 55358 18846 55410
rect 18846 55358 18898 55410
rect 18898 55358 18900 55410
rect 18844 55356 18900 55358
rect 19404 56028 19460 56084
rect 20188 56194 20244 56196
rect 20188 56142 20190 56194
rect 20190 56142 20242 56194
rect 20242 56142 20244 56194
rect 20188 56140 20244 56142
rect 21308 56194 21364 56196
rect 21308 56142 21310 56194
rect 21310 56142 21362 56194
rect 21362 56142 21364 56194
rect 21308 56140 21364 56142
rect 19852 55356 19908 55412
rect 19180 55244 19236 55300
rect 19068 55186 19124 55188
rect 19068 55134 19070 55186
rect 19070 55134 19122 55186
rect 19122 55134 19124 55186
rect 19068 55132 19124 55134
rect 18172 53900 18228 53956
rect 18396 53842 18452 53844
rect 18396 53790 18398 53842
rect 18398 53790 18450 53842
rect 18450 53790 18452 53842
rect 18396 53788 18452 53790
rect 18620 53730 18676 53732
rect 18620 53678 18622 53730
rect 18622 53678 18674 53730
rect 18674 53678 18676 53730
rect 18620 53676 18676 53678
rect 16828 51378 16884 51380
rect 16828 51326 16830 51378
rect 16830 51326 16882 51378
rect 16882 51326 16884 51378
rect 16828 51324 16884 51326
rect 16604 50876 16660 50932
rect 16828 50316 16884 50372
rect 16380 48972 16436 49028
rect 16604 49026 16660 49028
rect 16604 48974 16606 49026
rect 16606 48974 16658 49026
rect 16658 48974 16660 49026
rect 16604 48972 16660 48974
rect 16828 48748 16884 48804
rect 16716 47404 16772 47460
rect 16380 47346 16436 47348
rect 16380 47294 16382 47346
rect 16382 47294 16434 47346
rect 16434 47294 16436 47346
rect 16380 47292 16436 47294
rect 16604 47292 16660 47348
rect 15708 46396 15764 46452
rect 15820 46674 15876 46676
rect 15820 46622 15822 46674
rect 15822 46622 15874 46674
rect 15874 46622 15876 46674
rect 15820 46620 15876 46622
rect 15708 45778 15764 45780
rect 15708 45726 15710 45778
rect 15710 45726 15762 45778
rect 15762 45726 15764 45778
rect 15708 45724 15764 45726
rect 15820 45666 15876 45668
rect 15820 45614 15822 45666
rect 15822 45614 15874 45666
rect 15874 45614 15876 45666
rect 15820 45612 15876 45614
rect 15596 45388 15652 45444
rect 16156 46620 16212 46676
rect 16380 46450 16436 46452
rect 16380 46398 16382 46450
rect 16382 46398 16434 46450
rect 16434 46398 16436 46450
rect 16380 46396 16436 46398
rect 16044 45666 16100 45668
rect 16044 45614 16046 45666
rect 16046 45614 16098 45666
rect 16098 45614 16100 45666
rect 16044 45612 16100 45614
rect 15932 44492 15988 44548
rect 15820 44268 15876 44324
rect 14028 43708 14084 43764
rect 13804 43372 13860 43428
rect 14924 44098 14980 44100
rect 14924 44046 14926 44098
rect 14926 44046 14978 44098
rect 14978 44046 14980 44098
rect 14924 44044 14980 44046
rect 15484 44098 15540 44100
rect 15484 44046 15486 44098
rect 15486 44046 15538 44098
rect 15538 44046 15540 44098
rect 15484 44044 15540 44046
rect 14364 43314 14420 43316
rect 14364 43262 14366 43314
rect 14366 43262 14418 43314
rect 14418 43262 14420 43314
rect 14364 43260 14420 43262
rect 14028 43148 14084 43204
rect 14924 43036 14980 43092
rect 15148 43372 15204 43428
rect 15372 43036 15428 43092
rect 13804 42530 13860 42532
rect 13804 42478 13806 42530
rect 13806 42478 13858 42530
rect 13858 42478 13860 42530
rect 13804 42476 13860 42478
rect 14476 42476 14532 42532
rect 13468 42252 13524 42308
rect 12908 42194 12964 42196
rect 12908 42142 12910 42194
rect 12910 42142 12962 42194
rect 12962 42142 12964 42194
rect 12908 42140 12964 42142
rect 13020 41746 13076 41748
rect 13020 41694 13022 41746
rect 13022 41694 13074 41746
rect 13074 41694 13076 41746
rect 13020 41692 13076 41694
rect 14476 42140 14532 42196
rect 13804 41804 13860 41860
rect 13244 40908 13300 40964
rect 11340 40626 11396 40628
rect 11340 40574 11342 40626
rect 11342 40574 11394 40626
rect 11394 40574 11396 40626
rect 11340 40572 11396 40574
rect 9436 40348 9492 40404
rect 11564 39730 11620 39732
rect 11564 39678 11566 39730
rect 11566 39678 11618 39730
rect 11618 39678 11620 39730
rect 11564 39676 11620 39678
rect 12012 40514 12068 40516
rect 12012 40462 12014 40514
rect 12014 40462 12066 40514
rect 12066 40462 12068 40514
rect 12012 40460 12068 40462
rect 14252 41244 14308 41300
rect 14700 41858 14756 41860
rect 14700 41806 14702 41858
rect 14702 41806 14754 41858
rect 14754 41806 14756 41858
rect 14700 41804 14756 41806
rect 14140 41186 14196 41188
rect 14140 41134 14142 41186
rect 14142 41134 14194 41186
rect 14194 41134 14196 41186
rect 14140 41132 14196 41134
rect 14028 41020 14084 41076
rect 13468 40684 13524 40740
rect 13580 40402 13636 40404
rect 13580 40350 13582 40402
rect 13582 40350 13634 40402
rect 13634 40350 13636 40402
rect 13580 40348 13636 40350
rect 14588 41132 14644 41188
rect 13916 40684 13972 40740
rect 13916 40348 13972 40404
rect 12684 40124 12740 40180
rect 14588 40402 14644 40404
rect 14588 40350 14590 40402
rect 14590 40350 14642 40402
rect 14642 40350 14644 40402
rect 14588 40348 14644 40350
rect 14588 40124 14644 40180
rect 12348 39676 12404 39732
rect 10780 38668 10836 38724
rect 6524 38108 6580 38164
rect 8204 38162 8260 38164
rect 8204 38110 8206 38162
rect 8206 38110 8258 38162
rect 8258 38110 8260 38162
rect 8204 38108 8260 38110
rect 5180 37324 5236 37380
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5292 29426 5348 29428
rect 5292 29374 5294 29426
rect 5294 29374 5346 29426
rect 5346 29374 5348 29426
rect 5292 29372 5348 29374
rect 9660 37100 9716 37156
rect 8540 29426 8596 29428
rect 8540 29374 8542 29426
rect 8542 29374 8594 29426
rect 8594 29374 8596 29426
rect 8540 29372 8596 29374
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 6524 28642 6580 28644
rect 6524 28590 6526 28642
rect 6526 28590 6578 28642
rect 6578 28590 6580 28642
rect 6524 28588 6580 28590
rect 7196 28642 7252 28644
rect 7196 28590 7198 28642
rect 7198 28590 7250 28642
rect 7250 28590 7252 28642
rect 7196 28588 7252 28590
rect 7532 27916 7588 27972
rect 2268 26460 2324 26516
rect 6636 27804 6692 27860
rect 6300 27746 6356 27748
rect 6300 27694 6302 27746
rect 6302 27694 6354 27746
rect 6354 27694 6356 27746
rect 6300 27692 6356 27694
rect 4956 27580 5012 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4844 26908 4900 26964
rect 3500 26460 3556 26516
rect 5628 26962 5684 26964
rect 5628 26910 5630 26962
rect 5630 26910 5682 26962
rect 5682 26910 5684 26962
rect 5628 26908 5684 26910
rect 3500 26124 3556 26180
rect 4172 26124 4228 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 6524 26124 6580 26180
rect 7084 27746 7140 27748
rect 7084 27694 7086 27746
rect 7086 27694 7138 27746
rect 7138 27694 7140 27746
rect 7084 27692 7140 27694
rect 6748 27634 6804 27636
rect 6748 27582 6750 27634
rect 6750 27582 6802 27634
rect 6802 27582 6804 27634
rect 6748 27580 6804 27582
rect 7868 27692 7924 27748
rect 6860 25116 6916 25172
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 3724 23324 3780 23380
rect 5068 22988 5124 23044
rect 4732 22876 4788 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 5404 23378 5460 23380
rect 5404 23326 5406 23378
rect 5406 23326 5458 23378
rect 5458 23326 5460 23378
rect 5404 23324 5460 23326
rect 5740 22988 5796 23044
rect 5740 22540 5796 22596
rect 6076 22876 6132 22932
rect 6412 22652 6468 22708
rect 2828 22316 2884 22372
rect 5740 22370 5796 22372
rect 5740 22318 5742 22370
rect 5742 22318 5794 22370
rect 5794 22318 5796 22370
rect 5740 22316 5796 22318
rect 6524 23154 6580 23156
rect 6524 23102 6526 23154
rect 6526 23102 6578 23154
rect 6578 23102 6580 23154
rect 6524 23100 6580 23102
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3612 20972 3668 21028
rect 5740 21026 5796 21028
rect 5740 20974 5742 21026
rect 5742 20974 5794 21026
rect 5794 20974 5796 21026
rect 5740 20972 5796 20974
rect 4620 20300 4676 20356
rect 2044 17836 2100 17892
rect 2828 20018 2884 20020
rect 2828 19966 2830 20018
rect 2830 19966 2882 20018
rect 2882 19966 2884 20018
rect 2828 19964 2884 19966
rect 5068 20018 5124 20020
rect 5068 19966 5070 20018
rect 5070 19966 5122 20018
rect 5122 19966 5124 20018
rect 5068 19964 5124 19966
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 2156 15820 2212 15876
rect 1820 15036 1876 15092
rect 5404 20300 5460 20356
rect 6076 20076 6132 20132
rect 5964 19964 6020 20020
rect 6860 22092 6916 22148
rect 7420 26178 7476 26180
rect 7420 26126 7422 26178
rect 7422 26126 7474 26178
rect 7474 26126 7476 26178
rect 7420 26124 7476 26126
rect 8428 27970 8484 27972
rect 8428 27918 8430 27970
rect 8430 27918 8482 27970
rect 8482 27918 8484 27970
rect 8428 27916 8484 27918
rect 8316 27634 8372 27636
rect 8316 27582 8318 27634
rect 8318 27582 8370 27634
rect 8370 27582 8372 27634
rect 8316 27580 8372 27582
rect 8092 26908 8148 26964
rect 9548 30098 9604 30100
rect 9548 30046 9550 30098
rect 9550 30046 9602 30098
rect 9602 30046 9604 30098
rect 9548 30044 9604 30046
rect 14812 41692 14868 41748
rect 14812 41244 14868 41300
rect 15708 42866 15764 42868
rect 15708 42814 15710 42866
rect 15710 42814 15762 42866
rect 15762 42814 15764 42866
rect 15708 42812 15764 42814
rect 15932 44044 15988 44100
rect 16156 44210 16212 44212
rect 16156 44158 16158 44210
rect 16158 44158 16210 44210
rect 16210 44158 16212 44210
rect 16156 44156 16212 44158
rect 16380 44828 16436 44884
rect 16716 44828 16772 44884
rect 16380 44322 16436 44324
rect 16380 44270 16382 44322
rect 16382 44270 16434 44322
rect 16434 44270 16436 44322
rect 16380 44268 16436 44270
rect 16156 43596 16212 43652
rect 15932 42812 15988 42868
rect 15372 41746 15428 41748
rect 15372 41694 15374 41746
rect 15374 41694 15426 41746
rect 15426 41694 15428 41746
rect 15372 41692 15428 41694
rect 14252 39618 14308 39620
rect 14252 39566 14254 39618
rect 14254 39566 14306 39618
rect 14306 39566 14308 39618
rect 14252 39564 14308 39566
rect 12908 39452 12964 39508
rect 14924 40402 14980 40404
rect 14924 40350 14926 40402
rect 14926 40350 14978 40402
rect 14978 40350 14980 40402
rect 14924 40348 14980 40350
rect 15148 40348 15204 40404
rect 15036 40236 15092 40292
rect 14924 39618 14980 39620
rect 14924 39566 14926 39618
rect 14926 39566 14978 39618
rect 14978 39566 14980 39618
rect 14924 39564 14980 39566
rect 13020 39228 13076 39284
rect 13356 38834 13412 38836
rect 13356 38782 13358 38834
rect 13358 38782 13410 38834
rect 13410 38782 13412 38834
rect 13356 38780 13412 38782
rect 14364 38220 14420 38276
rect 10108 37100 10164 37156
rect 14028 37772 14084 37828
rect 14812 38946 14868 38948
rect 14812 38894 14814 38946
rect 14814 38894 14866 38946
rect 14866 38894 14868 38946
rect 14812 38892 14868 38894
rect 15148 38610 15204 38612
rect 15148 38558 15150 38610
rect 15150 38558 15202 38610
rect 15202 38558 15204 38610
rect 15148 38556 15204 38558
rect 15036 38220 15092 38276
rect 15036 38050 15092 38052
rect 15036 37998 15038 38050
rect 15038 37998 15090 38050
rect 15090 37998 15092 38050
rect 15036 37996 15092 37998
rect 14140 37548 14196 37604
rect 14812 37660 14868 37716
rect 12908 37154 12964 37156
rect 12908 37102 12910 37154
rect 12910 37102 12962 37154
rect 12962 37102 12964 37154
rect 12908 37100 12964 37102
rect 10332 36988 10388 37044
rect 12012 35308 12068 35364
rect 14476 37154 14532 37156
rect 14476 37102 14478 37154
rect 14478 37102 14530 37154
rect 14530 37102 14532 37154
rect 14476 37100 14532 37102
rect 15260 37884 15316 37940
rect 15484 39506 15540 39508
rect 15484 39454 15486 39506
rect 15486 39454 15538 39506
rect 15538 39454 15540 39506
rect 15484 39452 15540 39454
rect 15708 41916 15764 41972
rect 16716 44044 16772 44100
rect 16828 43596 16884 43652
rect 16828 43426 16884 43428
rect 16828 43374 16830 43426
rect 16830 43374 16882 43426
rect 16882 43374 16884 43426
rect 16828 43372 16884 43374
rect 16380 43314 16436 43316
rect 16380 43262 16382 43314
rect 16382 43262 16434 43314
rect 16434 43262 16436 43314
rect 16380 43260 16436 43262
rect 16380 42978 16436 42980
rect 16380 42926 16382 42978
rect 16382 42926 16434 42978
rect 16434 42926 16436 42978
rect 16380 42924 16436 42926
rect 16492 42642 16548 42644
rect 16492 42590 16494 42642
rect 16494 42590 16546 42642
rect 16546 42590 16548 42642
rect 16492 42588 16548 42590
rect 16044 41692 16100 41748
rect 16044 41186 16100 41188
rect 16044 41134 16046 41186
rect 16046 41134 16098 41186
rect 16098 41134 16100 41186
rect 16044 41132 16100 41134
rect 16492 41692 16548 41748
rect 16268 41580 16324 41636
rect 16492 41186 16548 41188
rect 16492 41134 16494 41186
rect 16494 41134 16546 41186
rect 16546 41134 16548 41186
rect 16492 41132 16548 41134
rect 16380 40962 16436 40964
rect 16380 40910 16382 40962
rect 16382 40910 16434 40962
rect 16434 40910 16436 40962
rect 16380 40908 16436 40910
rect 15932 40572 15988 40628
rect 15932 40236 15988 40292
rect 16268 40348 16324 40404
rect 16828 42140 16884 42196
rect 16716 41916 16772 41972
rect 17724 52220 17780 52276
rect 18284 52274 18340 52276
rect 18284 52222 18286 52274
rect 18286 52222 18338 52274
rect 18338 52222 18340 52274
rect 18284 52220 18340 52222
rect 18732 52162 18788 52164
rect 18732 52110 18734 52162
rect 18734 52110 18786 52162
rect 18786 52110 18788 52162
rect 18732 52108 18788 52110
rect 18172 51884 18228 51940
rect 17612 51490 17668 51492
rect 17612 51438 17614 51490
rect 17614 51438 17666 51490
rect 17666 51438 17668 51490
rect 17612 51436 17668 51438
rect 17612 50988 17668 51044
rect 17948 50876 18004 50932
rect 18172 51324 18228 51380
rect 18396 51436 18452 51492
rect 18732 51266 18788 51268
rect 18732 51214 18734 51266
rect 18734 51214 18786 51266
rect 18786 51214 18788 51266
rect 18732 51212 18788 51214
rect 18732 50988 18788 51044
rect 18396 50540 18452 50596
rect 18508 50370 18564 50372
rect 18508 50318 18510 50370
rect 18510 50318 18562 50370
rect 18562 50318 18564 50370
rect 18508 50316 18564 50318
rect 17052 41804 17108 41860
rect 17164 49026 17220 49028
rect 17164 48974 17166 49026
rect 17166 48974 17218 49026
rect 17218 48974 17220 49026
rect 17164 48972 17220 48974
rect 16940 41468 16996 41524
rect 15708 39058 15764 39060
rect 15708 39006 15710 39058
rect 15710 39006 15762 39058
rect 15762 39006 15764 39058
rect 15708 39004 15764 39006
rect 15596 38722 15652 38724
rect 15596 38670 15598 38722
rect 15598 38670 15650 38722
rect 15650 38670 15652 38722
rect 15596 38668 15652 38670
rect 16156 39564 16212 39620
rect 15932 39340 15988 39396
rect 15820 38668 15876 38724
rect 15484 38556 15540 38612
rect 15596 37772 15652 37828
rect 15036 37548 15092 37604
rect 15036 37378 15092 37380
rect 15036 37326 15038 37378
rect 15038 37326 15090 37378
rect 15090 37326 15092 37378
rect 15036 37324 15092 37326
rect 15260 37436 15316 37492
rect 15820 37660 15876 37716
rect 16268 39900 16324 39956
rect 16156 39004 16212 39060
rect 16716 39394 16772 39396
rect 16716 39342 16718 39394
rect 16718 39342 16770 39394
rect 16770 39342 16772 39394
rect 16716 39340 16772 39342
rect 17052 41356 17108 41412
rect 16940 40796 16996 40852
rect 17052 40012 17108 40068
rect 16604 38892 16660 38948
rect 16044 37436 16100 37492
rect 16156 37548 16212 37604
rect 14812 36988 14868 37044
rect 16492 38556 16548 38612
rect 16380 37996 16436 38052
rect 16268 37212 16324 37268
rect 15260 37100 15316 37156
rect 14924 35756 14980 35812
rect 14812 35644 14868 35700
rect 12908 35308 12964 35364
rect 13804 35420 13860 35476
rect 12684 35084 12740 35140
rect 13468 35138 13524 35140
rect 13468 35086 13470 35138
rect 13470 35086 13522 35138
rect 13522 35086 13524 35138
rect 13468 35084 13524 35086
rect 14588 35196 14644 35252
rect 13580 33628 13636 33684
rect 12348 33292 12404 33348
rect 13580 33346 13636 33348
rect 13580 33294 13582 33346
rect 13582 33294 13634 33346
rect 13634 33294 13636 33346
rect 13580 33292 13636 33294
rect 13020 31836 13076 31892
rect 13468 31666 13524 31668
rect 13468 31614 13470 31666
rect 13470 31614 13522 31666
rect 13522 31614 13524 31666
rect 13468 31612 13524 31614
rect 13692 31890 13748 31892
rect 13692 31838 13694 31890
rect 13694 31838 13746 31890
rect 13746 31838 13748 31890
rect 13692 31836 13748 31838
rect 15708 37100 15764 37156
rect 15484 36652 15540 36708
rect 15484 35698 15540 35700
rect 15484 35646 15486 35698
rect 15486 35646 15538 35698
rect 15538 35646 15540 35698
rect 15484 35644 15540 35646
rect 16604 36988 16660 37044
rect 16492 36876 16548 36932
rect 15596 35586 15652 35588
rect 15596 35534 15598 35586
rect 15598 35534 15650 35586
rect 15650 35534 15652 35586
rect 15596 35532 15652 35534
rect 15820 35196 15876 35252
rect 16156 35868 16212 35924
rect 17052 36204 17108 36260
rect 17500 48412 17556 48468
rect 17276 47068 17332 47124
rect 18620 48972 18676 49028
rect 21868 55244 21924 55300
rect 19964 55074 20020 55076
rect 19964 55022 19966 55074
rect 19966 55022 20018 55074
rect 20018 55022 20020 55074
rect 19964 55020 20020 55022
rect 21420 55074 21476 55076
rect 21420 55022 21422 55074
rect 21422 55022 21474 55074
rect 21474 55022 21476 55074
rect 21420 55020 21476 55022
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19292 54348 19348 54404
rect 19180 53452 19236 53508
rect 20412 54402 20468 54404
rect 20412 54350 20414 54402
rect 20414 54350 20466 54402
rect 20466 54350 20468 54402
rect 20412 54348 20468 54350
rect 19852 54236 19908 54292
rect 19740 53618 19796 53620
rect 19740 53566 19742 53618
rect 19742 53566 19794 53618
rect 19794 53566 19796 53618
rect 19740 53564 19796 53566
rect 19628 53506 19684 53508
rect 19628 53454 19630 53506
rect 19630 53454 19682 53506
rect 19682 53454 19684 53506
rect 19628 53452 19684 53454
rect 19068 52108 19124 52164
rect 19180 52220 19236 52276
rect 19068 51938 19124 51940
rect 19068 51886 19070 51938
rect 19070 51886 19122 51938
rect 19122 51886 19124 51938
rect 19068 51884 19124 51886
rect 19068 51490 19124 51492
rect 19068 51438 19070 51490
rect 19070 51438 19122 51490
rect 19122 51438 19124 51490
rect 19068 51436 19124 51438
rect 20636 53788 20692 53844
rect 20188 53564 20244 53620
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 20636 53506 20692 53508
rect 20636 53454 20638 53506
rect 20638 53454 20690 53506
rect 20690 53454 20692 53506
rect 20636 53452 20692 53454
rect 20524 52220 20580 52276
rect 22316 55020 22372 55076
rect 21420 53506 21476 53508
rect 21420 53454 21422 53506
rect 21422 53454 21474 53506
rect 21474 53454 21476 53506
rect 21420 53452 21476 53454
rect 21868 52892 21924 52948
rect 21532 52220 21588 52276
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19740 51212 19796 51268
rect 20076 51266 20132 51268
rect 20076 51214 20078 51266
rect 20078 51214 20130 51266
rect 20130 51214 20132 51266
rect 20076 51212 20132 51214
rect 19964 51100 20020 51156
rect 19292 50594 19348 50596
rect 19292 50542 19294 50594
rect 19294 50542 19346 50594
rect 19346 50542 19348 50594
rect 19292 50540 19348 50542
rect 19740 50876 19796 50932
rect 19180 50316 19236 50372
rect 19516 50540 19572 50596
rect 18956 49532 19012 49588
rect 18956 49084 19012 49140
rect 18508 48412 18564 48468
rect 18620 48242 18676 48244
rect 18620 48190 18622 48242
rect 18622 48190 18674 48242
rect 18674 48190 18676 48242
rect 18620 48188 18676 48190
rect 17948 47180 18004 47236
rect 18172 47458 18228 47460
rect 18172 47406 18174 47458
rect 18174 47406 18226 47458
rect 18226 47406 18228 47458
rect 18172 47404 18228 47406
rect 17388 46562 17444 46564
rect 17388 46510 17390 46562
rect 17390 46510 17442 46562
rect 17442 46510 17444 46562
rect 17388 46508 17444 46510
rect 17612 46562 17668 46564
rect 17612 46510 17614 46562
rect 17614 46510 17666 46562
rect 17666 46510 17668 46562
rect 17612 46508 17668 46510
rect 17612 44716 17668 44772
rect 17724 45052 17780 45108
rect 17500 44604 17556 44660
rect 17388 44434 17444 44436
rect 17388 44382 17390 44434
rect 17390 44382 17442 44434
rect 17442 44382 17444 44434
rect 17388 44380 17444 44382
rect 17276 43820 17332 43876
rect 17724 43820 17780 43876
rect 17612 43650 17668 43652
rect 17612 43598 17614 43650
rect 17614 43598 17666 43650
rect 17666 43598 17668 43650
rect 17612 43596 17668 43598
rect 17724 43484 17780 43540
rect 18508 46620 18564 46676
rect 18172 45388 18228 45444
rect 18060 45052 18116 45108
rect 17276 42588 17332 42644
rect 17612 42252 17668 42308
rect 17500 41970 17556 41972
rect 17500 41918 17502 41970
rect 17502 41918 17554 41970
rect 17554 41918 17556 41970
rect 17500 41916 17556 41918
rect 17612 41692 17668 41748
rect 17388 41580 17444 41636
rect 17388 41356 17444 41412
rect 17276 41074 17332 41076
rect 17276 41022 17278 41074
rect 17278 41022 17330 41074
rect 17330 41022 17332 41074
rect 17276 41020 17332 41022
rect 17388 40908 17444 40964
rect 17724 41468 17780 41524
rect 17612 40626 17668 40628
rect 17612 40574 17614 40626
rect 17614 40574 17666 40626
rect 17666 40574 17668 40626
rect 17612 40572 17668 40574
rect 18284 44604 18340 44660
rect 18396 44380 18452 44436
rect 18620 45836 18676 45892
rect 18732 44604 18788 44660
rect 18620 44268 18676 44324
rect 18620 44044 18676 44100
rect 18732 43484 18788 43540
rect 18620 43260 18676 43316
rect 18172 42978 18228 42980
rect 18172 42926 18174 42978
rect 18174 42926 18226 42978
rect 18226 42926 18228 42978
rect 18172 42924 18228 42926
rect 17948 41804 18004 41860
rect 18060 41916 18116 41972
rect 17948 40908 18004 40964
rect 17948 40460 18004 40516
rect 17948 40012 18004 40068
rect 17948 39788 18004 39844
rect 17276 37100 17332 37156
rect 17724 39004 17780 39060
rect 18060 38668 18116 38724
rect 17724 37996 17780 38052
rect 17612 37772 17668 37828
rect 17612 37212 17668 37268
rect 17612 36316 17668 36372
rect 17388 35922 17444 35924
rect 17388 35870 17390 35922
rect 17390 35870 17442 35922
rect 17442 35870 17444 35922
rect 17388 35868 17444 35870
rect 18060 37772 18116 37828
rect 17836 37042 17892 37044
rect 17836 36990 17838 37042
rect 17838 36990 17890 37042
rect 17890 36990 17892 37042
rect 17836 36988 17892 36990
rect 18508 42978 18564 42980
rect 18508 42926 18510 42978
rect 18510 42926 18562 42978
rect 18562 42926 18564 42978
rect 18508 42924 18564 42926
rect 18732 42924 18788 42980
rect 19180 47234 19236 47236
rect 19180 47182 19182 47234
rect 19182 47182 19234 47234
rect 19234 47182 19236 47234
rect 19180 47180 19236 47182
rect 20188 50594 20244 50596
rect 20188 50542 20190 50594
rect 20190 50542 20242 50594
rect 20242 50542 20244 50594
rect 20188 50540 20244 50542
rect 19628 50428 19684 50484
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19404 49698 19460 49700
rect 19404 49646 19406 49698
rect 19406 49646 19458 49698
rect 19458 49646 19460 49698
rect 19404 49644 19460 49646
rect 19852 49810 19908 49812
rect 19852 49758 19854 49810
rect 19854 49758 19906 49810
rect 19906 49758 19908 49810
rect 19852 49756 19908 49758
rect 19516 48466 19572 48468
rect 19516 48414 19518 48466
rect 19518 48414 19570 48466
rect 19570 48414 19572 48466
rect 19516 48412 19572 48414
rect 19628 49196 19684 49252
rect 20300 49810 20356 49812
rect 20300 49758 20302 49810
rect 20302 49758 20354 49810
rect 20354 49758 20356 49810
rect 20300 49756 20356 49758
rect 20188 48860 20244 48916
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 20524 49586 20580 49588
rect 20524 49534 20526 49586
rect 20526 49534 20578 49586
rect 20578 49534 20580 49586
rect 20524 49532 20580 49534
rect 20748 50428 20804 50484
rect 22540 53506 22596 53508
rect 22540 53454 22542 53506
rect 22542 53454 22594 53506
rect 22594 53454 22596 53506
rect 22540 53452 22596 53454
rect 22204 52332 22260 52388
rect 22092 51378 22148 51380
rect 22092 51326 22094 51378
rect 22094 51326 22146 51378
rect 22146 51326 22148 51378
rect 22092 51324 22148 51326
rect 21756 51266 21812 51268
rect 21756 51214 21758 51266
rect 21758 51214 21810 51266
rect 21810 51214 21812 51266
rect 21756 51212 21812 51214
rect 21980 50988 22036 51044
rect 20636 48748 20692 48804
rect 20412 48412 20468 48468
rect 20636 48412 20692 48468
rect 19516 47180 19572 47236
rect 19068 45890 19124 45892
rect 19068 45838 19070 45890
rect 19070 45838 19122 45890
rect 19122 45838 19124 45890
rect 19068 45836 19124 45838
rect 19068 45276 19124 45332
rect 18956 45218 19012 45220
rect 18956 45166 18958 45218
rect 18958 45166 19010 45218
rect 19010 45166 19012 45218
rect 18956 45164 19012 45166
rect 18956 44940 19012 44996
rect 19964 48188 20020 48244
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20076 46732 20132 46788
rect 19404 46002 19460 46004
rect 19404 45950 19406 46002
rect 19406 45950 19458 46002
rect 19458 45950 19460 46002
rect 19404 45948 19460 45950
rect 19404 45388 19460 45444
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19404 44828 19460 44884
rect 19740 44604 19796 44660
rect 19292 44322 19348 44324
rect 19292 44270 19294 44322
rect 19294 44270 19346 44322
rect 19346 44270 19348 44322
rect 19292 44268 19348 44270
rect 19068 43148 19124 43204
rect 18732 42530 18788 42532
rect 18732 42478 18734 42530
rect 18734 42478 18786 42530
rect 18786 42478 18788 42530
rect 18732 42476 18788 42478
rect 18396 42252 18452 42308
rect 18396 41916 18452 41972
rect 18284 41580 18340 41636
rect 18284 41410 18340 41412
rect 18284 41358 18286 41410
rect 18286 41358 18338 41410
rect 18338 41358 18340 41410
rect 18284 41356 18340 41358
rect 18284 40908 18340 40964
rect 18844 41804 18900 41860
rect 18956 41580 19012 41636
rect 18956 41074 19012 41076
rect 18956 41022 18958 41074
rect 18958 41022 19010 41074
rect 19010 41022 19012 41074
rect 18956 41020 19012 41022
rect 18620 40572 18676 40628
rect 18284 39788 18340 39844
rect 18396 39676 18452 39732
rect 18284 38892 18340 38948
rect 18284 38668 18340 38724
rect 19292 43372 19348 43428
rect 19516 44380 19572 44436
rect 19516 43596 19572 43652
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19516 43426 19572 43428
rect 19516 43374 19518 43426
rect 19518 43374 19570 43426
rect 19570 43374 19572 43426
rect 19516 43372 19572 43374
rect 20860 48412 20916 48468
rect 20972 48972 21028 49028
rect 21644 49084 21700 49140
rect 21308 48860 21364 48916
rect 21420 48748 21476 48804
rect 21308 48076 21364 48132
rect 20300 45836 20356 45892
rect 20748 45890 20804 45892
rect 20748 45838 20750 45890
rect 20750 45838 20802 45890
rect 20802 45838 20804 45890
rect 20748 45836 20804 45838
rect 20636 44940 20692 44996
rect 20748 45612 20804 45668
rect 20412 44716 20468 44772
rect 21196 46674 21252 46676
rect 21196 46622 21198 46674
rect 21198 46622 21250 46674
rect 21250 46622 21252 46674
rect 21196 46620 21252 46622
rect 20860 45388 20916 45444
rect 20524 44604 20580 44660
rect 20300 43820 20356 43876
rect 20188 43148 20244 43204
rect 19852 42476 19908 42532
rect 20188 42924 20244 42980
rect 19404 42252 19460 42308
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19180 42028 19236 42084
rect 19404 41858 19460 41860
rect 19404 41806 19406 41858
rect 19406 41806 19458 41858
rect 19458 41806 19460 41858
rect 19404 41804 19460 41806
rect 19404 41356 19460 41412
rect 20300 41970 20356 41972
rect 20300 41918 20302 41970
rect 20302 41918 20354 41970
rect 20354 41918 20356 41970
rect 20300 41916 20356 41918
rect 20860 43650 20916 43652
rect 20860 43598 20862 43650
rect 20862 43598 20914 43650
rect 20914 43598 20916 43650
rect 20860 43596 20916 43598
rect 20748 42194 20804 42196
rect 20748 42142 20750 42194
rect 20750 42142 20802 42194
rect 20802 42142 20804 42194
rect 20748 42140 20804 42142
rect 20636 42082 20692 42084
rect 20636 42030 20638 42082
rect 20638 42030 20690 42082
rect 20690 42030 20692 42082
rect 20636 42028 20692 42030
rect 19180 40962 19236 40964
rect 19180 40910 19182 40962
rect 19182 40910 19234 40962
rect 19234 40910 19236 40962
rect 19180 40908 19236 40910
rect 19404 40290 19460 40292
rect 19404 40238 19406 40290
rect 19406 40238 19458 40290
rect 19458 40238 19460 40290
rect 19404 40236 19460 40238
rect 19292 39676 19348 39732
rect 19068 39564 19124 39620
rect 19404 39452 19460 39508
rect 18844 38946 18900 38948
rect 18844 38894 18846 38946
rect 18846 38894 18898 38946
rect 18898 38894 18900 38946
rect 18844 38892 18900 38894
rect 18732 38556 18788 38612
rect 18620 37938 18676 37940
rect 18620 37886 18622 37938
rect 18622 37886 18674 37938
rect 18674 37886 18676 37938
rect 18620 37884 18676 37886
rect 19628 40796 19684 40852
rect 20188 41020 20244 41076
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19964 40402 20020 40404
rect 19964 40350 19966 40402
rect 19966 40350 20018 40402
rect 20018 40350 20020 40402
rect 19964 40348 20020 40350
rect 19628 40178 19684 40180
rect 19628 40126 19630 40178
rect 19630 40126 19682 40178
rect 19682 40126 19684 40178
rect 19628 40124 19684 40126
rect 19628 39564 19684 39620
rect 19516 37548 19572 37604
rect 19964 39506 20020 39508
rect 19964 39454 19966 39506
rect 19966 39454 20018 39506
rect 20018 39454 20020 39506
rect 19964 39452 20020 39454
rect 20076 39394 20132 39396
rect 20076 39342 20078 39394
rect 20078 39342 20130 39394
rect 20130 39342 20132 39394
rect 20076 39340 20132 39342
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19852 38946 19908 38948
rect 19852 38894 19854 38946
rect 19854 38894 19906 38946
rect 19906 38894 19908 38946
rect 19852 38892 19908 38894
rect 20412 41020 20468 41076
rect 20748 41356 20804 41412
rect 20748 40684 20804 40740
rect 20860 40572 20916 40628
rect 20972 40348 21028 40404
rect 20860 40012 20916 40068
rect 20748 39564 20804 39620
rect 20412 38668 20468 38724
rect 19852 38050 19908 38052
rect 19852 37998 19854 38050
rect 19854 37998 19906 38050
rect 19906 37998 19908 38050
rect 19852 37996 19908 37998
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19292 37212 19348 37268
rect 18284 36258 18340 36260
rect 18284 36206 18286 36258
rect 18286 36206 18338 36258
rect 18338 36206 18340 36258
rect 18284 36204 18340 36206
rect 18284 35922 18340 35924
rect 18284 35870 18286 35922
rect 18286 35870 18338 35922
rect 18338 35870 18340 35922
rect 18284 35868 18340 35870
rect 16828 35196 16884 35252
rect 16492 34802 16548 34804
rect 16492 34750 16494 34802
rect 16494 34750 16546 34802
rect 16546 34750 16548 34802
rect 16492 34748 16548 34750
rect 17500 34748 17556 34804
rect 15596 34354 15652 34356
rect 15596 34302 15598 34354
rect 15598 34302 15650 34354
rect 15650 34302 15652 34354
rect 15596 34300 15652 34302
rect 17388 34300 17444 34356
rect 15260 34076 15316 34132
rect 14364 33516 14420 33572
rect 17724 34636 17780 34692
rect 16380 34130 16436 34132
rect 16380 34078 16382 34130
rect 16382 34078 16434 34130
rect 16434 34078 16436 34130
rect 16380 34076 16436 34078
rect 17948 34130 18004 34132
rect 17948 34078 17950 34130
rect 17950 34078 18002 34130
rect 18002 34078 18004 34130
rect 17948 34076 18004 34078
rect 17164 33964 17220 34020
rect 18732 35532 18788 35588
rect 18508 34018 18564 34020
rect 18508 33966 18510 34018
rect 18510 33966 18562 34018
rect 18562 33966 18564 34018
rect 18508 33964 18564 33966
rect 16940 33740 16996 33796
rect 15708 33292 15764 33348
rect 16940 33458 16996 33460
rect 16940 33406 16942 33458
rect 16942 33406 16994 33458
rect 16994 33406 16996 33458
rect 16940 33404 16996 33406
rect 16716 33292 16772 33348
rect 16044 32396 16100 32452
rect 15148 31836 15204 31892
rect 15596 31948 15652 32004
rect 10332 30044 10388 30100
rect 9772 29932 9828 29988
rect 11228 29538 11284 29540
rect 11228 29486 11230 29538
rect 11230 29486 11282 29538
rect 11282 29486 11284 29538
rect 11228 29484 11284 29486
rect 7644 26796 7700 26852
rect 12460 29484 12516 29540
rect 10668 27692 10724 27748
rect 11452 29426 11508 29428
rect 11452 29374 11454 29426
rect 11454 29374 11506 29426
rect 11506 29374 11508 29426
rect 11452 29372 11508 29374
rect 13580 30492 13636 30548
rect 14252 30770 14308 30772
rect 14252 30718 14254 30770
rect 14254 30718 14306 30770
rect 14306 30718 14308 30770
rect 14252 30716 14308 30718
rect 15708 31276 15764 31332
rect 15484 31164 15540 31220
rect 16268 32284 16324 32340
rect 16268 31948 16324 32004
rect 16156 31276 16212 31332
rect 16380 31836 16436 31892
rect 16604 32172 16660 32228
rect 16492 31612 16548 31668
rect 16604 31164 16660 31220
rect 16380 31052 16436 31108
rect 14364 30604 14420 30660
rect 14252 30492 14308 30548
rect 13468 29372 13524 29428
rect 15932 29372 15988 29428
rect 13916 27692 13972 27748
rect 8204 26124 8260 26180
rect 9436 26124 9492 26180
rect 8652 25116 8708 25172
rect 8316 25004 8372 25060
rect 7980 23938 8036 23940
rect 7980 23886 7982 23938
rect 7982 23886 8034 23938
rect 8034 23886 8036 23938
rect 7980 23884 8036 23886
rect 7084 23660 7140 23716
rect 7308 23154 7364 23156
rect 7308 23102 7310 23154
rect 7310 23102 7362 23154
rect 7362 23102 7364 23154
rect 7308 23100 7364 23102
rect 7308 22594 7364 22596
rect 7308 22542 7310 22594
rect 7310 22542 7362 22594
rect 7362 22542 7364 22594
rect 7308 22540 7364 22542
rect 7868 23714 7924 23716
rect 7868 23662 7870 23714
rect 7870 23662 7922 23714
rect 7922 23662 7924 23714
rect 7868 23660 7924 23662
rect 10556 26796 10612 26852
rect 9884 26290 9940 26292
rect 9884 26238 9886 26290
rect 9886 26238 9938 26290
rect 9938 26238 9940 26290
rect 9884 26236 9940 26238
rect 10556 26290 10612 26292
rect 10556 26238 10558 26290
rect 10558 26238 10610 26290
rect 10610 26238 10612 26290
rect 10556 26236 10612 26238
rect 9772 25228 9828 25284
rect 8540 23714 8596 23716
rect 8540 23662 8542 23714
rect 8542 23662 8594 23714
rect 8594 23662 8596 23714
rect 8540 23660 8596 23662
rect 7532 22988 7588 23044
rect 7980 22930 8036 22932
rect 7980 22878 7982 22930
rect 7982 22878 8034 22930
rect 8034 22878 8036 22930
rect 7980 22876 8036 22878
rect 7420 20636 7476 20692
rect 6860 19964 6916 20020
rect 6188 19852 6244 19908
rect 6300 19068 6356 19124
rect 4060 18396 4116 18452
rect 5516 18508 5572 18564
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4620 17778 4676 17780
rect 4620 17726 4622 17778
rect 4622 17726 4674 17778
rect 4674 17726 4676 17778
rect 4620 17724 4676 17726
rect 6300 18508 6356 18564
rect 5964 18450 6020 18452
rect 5964 18398 5966 18450
rect 5966 18398 6018 18450
rect 6018 18398 6020 18450
rect 5964 18396 6020 18398
rect 6524 18508 6580 18564
rect 5740 17890 5796 17892
rect 5740 17838 5742 17890
rect 5742 17838 5794 17890
rect 5794 17838 5796 17890
rect 5740 17836 5796 17838
rect 6076 17890 6132 17892
rect 6076 17838 6078 17890
rect 6078 17838 6130 17890
rect 6130 17838 6132 17890
rect 6076 17836 6132 17838
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4844 16044 4900 16100
rect 4060 15484 4116 15540
rect 2828 15036 2884 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 7756 21810 7812 21812
rect 7756 21758 7758 21810
rect 7758 21758 7810 21810
rect 7810 21758 7812 21810
rect 7756 21756 7812 21758
rect 8764 23042 8820 23044
rect 8764 22990 8766 23042
rect 8766 22990 8818 23042
rect 8818 22990 8820 23042
rect 8764 22988 8820 22990
rect 8316 21868 8372 21924
rect 7756 21586 7812 21588
rect 7756 21534 7758 21586
rect 7758 21534 7810 21586
rect 7810 21534 7812 21586
rect 7756 21532 7812 21534
rect 8204 21532 8260 21588
rect 7084 20130 7140 20132
rect 7084 20078 7086 20130
rect 7086 20078 7138 20130
rect 7138 20078 7140 20130
rect 7084 20076 7140 20078
rect 7308 20130 7364 20132
rect 7308 20078 7310 20130
rect 7310 20078 7362 20130
rect 7362 20078 7364 20130
rect 7308 20076 7364 20078
rect 7868 20690 7924 20692
rect 7868 20638 7870 20690
rect 7870 20638 7922 20690
rect 7922 20638 7924 20690
rect 7868 20636 7924 20638
rect 8092 20578 8148 20580
rect 8092 20526 8094 20578
rect 8094 20526 8146 20578
rect 8146 20526 8148 20578
rect 8092 20524 8148 20526
rect 8204 20412 8260 20468
rect 6972 18620 7028 18676
rect 8652 21586 8708 21588
rect 8652 21534 8654 21586
rect 8654 21534 8706 21586
rect 8706 21534 8708 21586
rect 8652 21532 8708 21534
rect 9212 21868 9268 21924
rect 8876 21196 8932 21252
rect 9100 21026 9156 21028
rect 9100 20974 9102 21026
rect 9102 20974 9154 21026
rect 9154 20974 9156 21026
rect 9100 20972 9156 20974
rect 9324 21532 9380 21588
rect 8652 20412 8708 20468
rect 8764 20300 8820 20356
rect 7756 18844 7812 18900
rect 10892 24892 10948 24948
rect 10892 22316 10948 22372
rect 10892 21698 10948 21700
rect 10892 21646 10894 21698
rect 10894 21646 10946 21698
rect 10946 21646 10948 21698
rect 10892 21644 10948 21646
rect 11452 26290 11508 26292
rect 11452 26238 11454 26290
rect 11454 26238 11506 26290
rect 11506 26238 11508 26290
rect 11452 26236 11508 26238
rect 11676 25564 11732 25620
rect 12572 26236 12628 26292
rect 12236 25228 12292 25284
rect 12348 25618 12404 25620
rect 12348 25566 12350 25618
rect 12350 25566 12402 25618
rect 12402 25566 12404 25618
rect 12348 25564 12404 25566
rect 11676 24946 11732 24948
rect 11676 24894 11678 24946
rect 11678 24894 11730 24946
rect 11730 24894 11732 24946
rect 11676 24892 11732 24894
rect 13916 26460 13972 26516
rect 16828 33068 16884 33124
rect 16828 31836 16884 31892
rect 17052 31666 17108 31668
rect 17052 31614 17054 31666
rect 17054 31614 17106 31666
rect 17106 31614 17108 31666
rect 17052 31612 17108 31614
rect 16828 31500 16884 31556
rect 17276 33570 17332 33572
rect 17276 33518 17278 33570
rect 17278 33518 17330 33570
rect 17330 33518 17332 33570
rect 17276 33516 17332 33518
rect 17724 33122 17780 33124
rect 17724 33070 17726 33122
rect 17726 33070 17778 33122
rect 17778 33070 17780 33122
rect 17724 33068 17780 33070
rect 17276 32732 17332 32788
rect 17724 32562 17780 32564
rect 17724 32510 17726 32562
rect 17726 32510 17778 32562
rect 17778 32510 17780 32562
rect 17724 32508 17780 32510
rect 17612 32396 17668 32452
rect 17500 32284 17556 32340
rect 17836 32172 17892 32228
rect 17388 31500 17444 31556
rect 17388 31218 17444 31220
rect 17388 31166 17390 31218
rect 17390 31166 17442 31218
rect 17442 31166 17444 31218
rect 17388 31164 17444 31166
rect 17500 31106 17556 31108
rect 17500 31054 17502 31106
rect 17502 31054 17554 31106
rect 17554 31054 17556 31106
rect 17500 31052 17556 31054
rect 18060 31500 18116 31556
rect 18172 31612 18228 31668
rect 17948 30940 18004 30996
rect 18620 32396 18676 32452
rect 18396 31948 18452 32004
rect 19404 36988 19460 37044
rect 19068 36876 19124 36932
rect 18956 36764 19012 36820
rect 19516 36428 19572 36484
rect 19068 36316 19124 36372
rect 20076 36652 20132 36708
rect 20300 37826 20356 37828
rect 20300 37774 20302 37826
rect 20302 37774 20354 37826
rect 20354 37774 20356 37826
rect 20300 37772 20356 37774
rect 20188 37212 20244 37268
rect 20076 36482 20132 36484
rect 20076 36430 20078 36482
rect 20078 36430 20130 36482
rect 20130 36430 20132 36482
rect 20076 36428 20132 36430
rect 18956 34690 19012 34692
rect 18956 34638 18958 34690
rect 18958 34638 19010 34690
rect 19010 34638 19012 34690
rect 18956 34636 19012 34638
rect 18844 34242 18900 34244
rect 18844 34190 18846 34242
rect 18846 34190 18898 34242
rect 18898 34190 18900 34242
rect 18844 34188 18900 34190
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20300 36204 20356 36260
rect 19740 35586 19796 35588
rect 19740 35534 19742 35586
rect 19742 35534 19794 35586
rect 19794 35534 19796 35586
rect 19740 35532 19796 35534
rect 19964 34914 20020 34916
rect 19964 34862 19966 34914
rect 19966 34862 20018 34914
rect 20018 34862 20020 34914
rect 19964 34860 20020 34862
rect 20860 39116 20916 39172
rect 21196 43596 21252 43652
rect 21644 46620 21700 46676
rect 21868 49250 21924 49252
rect 21868 49198 21870 49250
rect 21870 49198 21922 49250
rect 21922 49198 21924 49250
rect 21868 49196 21924 49198
rect 21756 45500 21812 45556
rect 21756 45052 21812 45108
rect 21532 43820 21588 43876
rect 21756 43820 21812 43876
rect 21532 43596 21588 43652
rect 21644 43538 21700 43540
rect 21644 43486 21646 43538
rect 21646 43486 21698 43538
rect 21698 43486 21700 43538
rect 21644 43484 21700 43486
rect 21532 43036 21588 43092
rect 21308 42924 21364 42980
rect 21308 42754 21364 42756
rect 21308 42702 21310 42754
rect 21310 42702 21362 42754
rect 21362 42702 21364 42754
rect 21308 42700 21364 42702
rect 21308 42252 21364 42308
rect 21196 41916 21252 41972
rect 21868 42754 21924 42756
rect 21868 42702 21870 42754
rect 21870 42702 21922 42754
rect 21922 42702 21924 42754
rect 21868 42700 21924 42702
rect 21644 42140 21700 42196
rect 20972 38892 21028 38948
rect 21196 39788 21252 39844
rect 20972 38668 21028 38724
rect 20860 38108 20916 38164
rect 21532 40402 21588 40404
rect 21532 40350 21534 40402
rect 21534 40350 21586 40402
rect 21586 40350 21588 40402
rect 21532 40348 21588 40350
rect 22204 50482 22260 50484
rect 22204 50430 22206 50482
rect 22206 50430 22258 50482
rect 22258 50430 22260 50482
rect 22204 50428 22260 50430
rect 23212 56306 23268 56308
rect 23212 56254 23214 56306
rect 23214 56254 23266 56306
rect 23266 56254 23268 56306
rect 23212 56252 23268 56254
rect 24668 56252 24724 56308
rect 23660 54460 23716 54516
rect 23100 53618 23156 53620
rect 23100 53566 23102 53618
rect 23102 53566 23154 53618
rect 23154 53566 23156 53618
rect 23100 53564 23156 53566
rect 22876 53506 22932 53508
rect 22876 53454 22878 53506
rect 22878 53454 22930 53506
rect 22930 53454 22932 53506
rect 22876 53452 22932 53454
rect 22764 52274 22820 52276
rect 22764 52222 22766 52274
rect 22766 52222 22818 52274
rect 22818 52222 22820 52274
rect 22764 52220 22820 52222
rect 22652 52108 22708 52164
rect 22876 51660 22932 51716
rect 22652 51324 22708 51380
rect 22428 51154 22484 51156
rect 22428 51102 22430 51154
rect 22430 51102 22482 51154
rect 22482 51102 22484 51154
rect 22428 51100 22484 51102
rect 23100 51378 23156 51380
rect 23100 51326 23102 51378
rect 23102 51326 23154 51378
rect 23154 51326 23156 51378
rect 23100 51324 23156 51326
rect 23100 50988 23156 51044
rect 22428 50428 22484 50484
rect 23772 53564 23828 53620
rect 24668 55468 24724 55524
rect 24556 54514 24612 54516
rect 24556 54462 24558 54514
rect 24558 54462 24610 54514
rect 24610 54462 24612 54514
rect 24556 54460 24612 54462
rect 23884 53116 23940 53172
rect 23548 52946 23604 52948
rect 23548 52894 23550 52946
rect 23550 52894 23602 52946
rect 23602 52894 23604 52946
rect 23548 52892 23604 52894
rect 23324 52220 23380 52276
rect 23548 51884 23604 51940
rect 23324 50594 23380 50596
rect 23324 50542 23326 50594
rect 23326 50542 23378 50594
rect 23378 50542 23380 50594
rect 23324 50540 23380 50542
rect 23436 50428 23492 50484
rect 24108 53170 24164 53172
rect 24108 53118 24110 53170
rect 24110 53118 24162 53170
rect 24162 53118 24164 53170
rect 24108 53116 24164 53118
rect 25788 55298 25844 55300
rect 25788 55246 25790 55298
rect 25790 55246 25842 55298
rect 25842 55246 25844 55298
rect 25788 55244 25844 55246
rect 26684 55468 26740 55524
rect 25228 54460 25284 54516
rect 24668 53452 24724 53508
rect 25676 53506 25732 53508
rect 25676 53454 25678 53506
rect 25678 53454 25730 53506
rect 25730 53454 25732 53506
rect 25676 53452 25732 53454
rect 24444 52668 24500 52724
rect 24332 52444 24388 52500
rect 23996 52162 24052 52164
rect 23996 52110 23998 52162
rect 23998 52110 24050 52162
rect 24050 52110 24052 52162
rect 23996 52108 24052 52110
rect 25228 52722 25284 52724
rect 25228 52670 25230 52722
rect 25230 52670 25282 52722
rect 25282 52670 25284 52722
rect 25228 52668 25284 52670
rect 25228 52444 25284 52500
rect 24668 52220 24724 52276
rect 23884 51884 23940 51940
rect 23772 51490 23828 51492
rect 23772 51438 23774 51490
rect 23774 51438 23826 51490
rect 23826 51438 23828 51490
rect 23772 51436 23828 51438
rect 23996 51378 24052 51380
rect 23996 51326 23998 51378
rect 23998 51326 24050 51378
rect 24050 51326 24052 51378
rect 23996 51324 24052 51326
rect 24108 51100 24164 51156
rect 24108 50876 24164 50932
rect 23884 50428 23940 50484
rect 23212 49810 23268 49812
rect 23212 49758 23214 49810
rect 23214 49758 23266 49810
rect 23266 49758 23268 49810
rect 23212 49756 23268 49758
rect 23324 49698 23380 49700
rect 23324 49646 23326 49698
rect 23326 49646 23378 49698
rect 23378 49646 23380 49698
rect 23324 49644 23380 49646
rect 23212 49196 23268 49252
rect 22540 48300 22596 48356
rect 22092 47346 22148 47348
rect 22092 47294 22094 47346
rect 22094 47294 22146 47346
rect 22146 47294 22148 47346
rect 22092 47292 22148 47294
rect 22764 48914 22820 48916
rect 22764 48862 22766 48914
rect 22766 48862 22818 48914
rect 22818 48862 22820 48914
rect 22764 48860 22820 48862
rect 24556 51938 24612 51940
rect 24556 51886 24558 51938
rect 24558 51886 24610 51938
rect 24610 51886 24612 51938
rect 24556 51884 24612 51886
rect 24556 51660 24612 51716
rect 24444 51154 24500 51156
rect 24444 51102 24446 51154
rect 24446 51102 24498 51154
rect 24498 51102 24500 51154
rect 24444 51100 24500 51102
rect 24556 50876 24612 50932
rect 24332 50540 24388 50596
rect 23324 48972 23380 49028
rect 23100 48748 23156 48804
rect 23884 49026 23940 49028
rect 23884 48974 23886 49026
rect 23886 48974 23938 49026
rect 23938 48974 23940 49026
rect 23884 48972 23940 48974
rect 25564 52722 25620 52724
rect 25564 52670 25566 52722
rect 25566 52670 25618 52722
rect 25618 52670 25620 52722
rect 25564 52668 25620 52670
rect 27356 55244 27412 55300
rect 29148 55298 29204 55300
rect 29148 55246 29150 55298
rect 29150 55246 29202 55298
rect 29202 55246 29204 55298
rect 29148 55244 29204 55246
rect 28252 54684 28308 54740
rect 29148 54738 29204 54740
rect 29148 54686 29150 54738
rect 29150 54686 29202 54738
rect 29202 54686 29204 54738
rect 29148 54684 29204 54686
rect 30044 56252 30100 56308
rect 30716 56306 30772 56308
rect 30716 56254 30718 56306
rect 30718 56254 30770 56306
rect 30770 56254 30772 56306
rect 30716 56252 30772 56254
rect 31388 56252 31444 56308
rect 30380 55244 30436 55300
rect 28812 53564 28868 53620
rect 32732 57036 32788 57092
rect 32620 56252 32676 56308
rect 34076 56924 34132 56980
rect 34188 57036 34244 57092
rect 33628 56252 33684 56308
rect 34076 55804 34132 55860
rect 30380 53676 30436 53732
rect 27244 52444 27300 52500
rect 27356 52668 27412 52724
rect 26908 51100 26964 51156
rect 24332 49196 24388 49252
rect 26236 50482 26292 50484
rect 26236 50430 26238 50482
rect 26238 50430 26290 50482
rect 26290 50430 26292 50482
rect 26236 50428 26292 50430
rect 23996 48860 24052 48916
rect 23660 48802 23716 48804
rect 23660 48750 23662 48802
rect 23662 48750 23714 48802
rect 23714 48750 23716 48802
rect 23660 48748 23716 48750
rect 23436 48354 23492 48356
rect 23436 48302 23438 48354
rect 23438 48302 23490 48354
rect 23490 48302 23492 48354
rect 23436 48300 23492 48302
rect 22428 48130 22484 48132
rect 22428 48078 22430 48130
rect 22430 48078 22482 48130
rect 22482 48078 22484 48130
rect 22428 48076 22484 48078
rect 22652 48018 22708 48020
rect 22652 47966 22654 48018
rect 22654 47966 22706 48018
rect 22706 47966 22708 48018
rect 22652 47964 22708 47966
rect 22316 47852 22372 47908
rect 22652 47458 22708 47460
rect 22652 47406 22654 47458
rect 22654 47406 22706 47458
rect 22706 47406 22708 47458
rect 22652 47404 22708 47406
rect 23548 47964 23604 48020
rect 23324 47292 23380 47348
rect 22316 46674 22372 46676
rect 22316 46622 22318 46674
rect 22318 46622 22370 46674
rect 22370 46622 22372 46674
rect 22316 46620 22372 46622
rect 22204 46284 22260 46340
rect 22540 46786 22596 46788
rect 22540 46734 22542 46786
rect 22542 46734 22594 46786
rect 22594 46734 22596 46786
rect 22540 46732 22596 46734
rect 22428 46172 22484 46228
rect 22428 45948 22484 46004
rect 22092 45388 22148 45444
rect 22092 44380 22148 44436
rect 21980 42028 22036 42084
rect 22092 43372 22148 43428
rect 22316 44604 22372 44660
rect 22316 42700 22372 42756
rect 23212 46284 23268 46340
rect 22988 45276 23044 45332
rect 23100 46172 23156 46228
rect 22764 44604 22820 44660
rect 23548 47068 23604 47124
rect 23436 45948 23492 46004
rect 22540 43148 22596 43204
rect 22876 43484 22932 43540
rect 23100 43650 23156 43652
rect 23100 43598 23102 43650
rect 23102 43598 23154 43650
rect 23154 43598 23156 43650
rect 23100 43596 23156 43598
rect 23548 45890 23604 45892
rect 23548 45838 23550 45890
rect 23550 45838 23602 45890
rect 23602 45838 23604 45890
rect 23548 45836 23604 45838
rect 23548 44434 23604 44436
rect 23548 44382 23550 44434
rect 23550 44382 23602 44434
rect 23602 44382 23604 44434
rect 23548 44380 23604 44382
rect 23548 43596 23604 43652
rect 23324 43426 23380 43428
rect 23324 43374 23326 43426
rect 23326 43374 23378 43426
rect 23378 43374 23380 43426
rect 23324 43372 23380 43374
rect 23100 43260 23156 43316
rect 22988 42924 23044 42980
rect 23212 43148 23268 43204
rect 22428 42588 22484 42644
rect 22764 42588 22820 42644
rect 22652 42140 22708 42196
rect 22092 41916 22148 41972
rect 22092 41468 22148 41524
rect 22204 41356 22260 41412
rect 22092 41132 22148 41188
rect 21868 40908 21924 40964
rect 21980 40796 22036 40852
rect 21532 39676 21588 39732
rect 21308 39004 21364 39060
rect 21420 39452 21476 39508
rect 21532 39116 21588 39172
rect 21532 36482 21588 36484
rect 21532 36430 21534 36482
rect 21534 36430 21586 36482
rect 21586 36430 21588 36482
rect 21532 36428 21588 36430
rect 20636 34860 20692 34916
rect 19852 34690 19908 34692
rect 19852 34638 19854 34690
rect 19854 34638 19906 34690
rect 19906 34638 19908 34690
rect 19852 34636 19908 34638
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 20188 34076 20244 34132
rect 19180 33516 19236 33572
rect 18956 33346 19012 33348
rect 18956 33294 18958 33346
rect 18958 33294 19010 33346
rect 19010 33294 19012 33346
rect 18956 33292 19012 33294
rect 19628 33346 19684 33348
rect 19628 33294 19630 33346
rect 19630 33294 19682 33346
rect 19682 33294 19684 33346
rect 19628 33292 19684 33294
rect 20412 33628 20468 33684
rect 19628 32844 19684 32900
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20076 32732 20132 32788
rect 20188 32396 20244 32452
rect 19740 32284 19796 32340
rect 18844 31778 18900 31780
rect 18844 31726 18846 31778
rect 18846 31726 18898 31778
rect 18898 31726 18900 31778
rect 18844 31724 18900 31726
rect 16268 29372 16324 29428
rect 16268 27916 16324 27972
rect 16044 27132 16100 27188
rect 12572 25340 12628 25396
rect 12012 24332 12068 24388
rect 11788 22594 11844 22596
rect 11788 22542 11790 22594
rect 11790 22542 11842 22594
rect 11842 22542 11844 22594
rect 11788 22540 11844 22542
rect 11452 22370 11508 22372
rect 11452 22318 11454 22370
rect 11454 22318 11506 22370
rect 11506 22318 11508 22370
rect 11452 22316 11508 22318
rect 12124 21698 12180 21700
rect 12124 21646 12126 21698
rect 12126 21646 12178 21698
rect 12178 21646 12180 21698
rect 12124 21644 12180 21646
rect 10108 21026 10164 21028
rect 10108 20974 10110 21026
rect 10110 20974 10162 21026
rect 10162 20974 10164 21026
rect 10108 20972 10164 20974
rect 8092 19122 8148 19124
rect 8092 19070 8094 19122
rect 8094 19070 8146 19122
rect 8146 19070 8148 19122
rect 8092 19068 8148 19070
rect 9100 19122 9156 19124
rect 9100 19070 9102 19122
rect 9102 19070 9154 19122
rect 9154 19070 9156 19122
rect 9100 19068 9156 19070
rect 7532 18732 7588 18788
rect 7868 18732 7924 18788
rect 6860 17948 6916 18004
rect 6748 17836 6804 17892
rect 7308 18620 7364 18676
rect 6748 17554 6804 17556
rect 6748 17502 6750 17554
rect 6750 17502 6802 17554
rect 6802 17502 6804 17554
rect 6748 17500 6804 17502
rect 6412 16828 6468 16884
rect 6076 16098 6132 16100
rect 6076 16046 6078 16098
rect 6078 16046 6130 16098
rect 6130 16046 6132 16098
rect 6076 16044 6132 16046
rect 5740 15874 5796 15876
rect 5740 15822 5742 15874
rect 5742 15822 5794 15874
rect 5794 15822 5796 15874
rect 5740 15820 5796 15822
rect 6076 15538 6132 15540
rect 6076 15486 6078 15538
rect 6078 15486 6130 15538
rect 6130 15486 6132 15538
rect 6076 15484 6132 15486
rect 7532 18562 7588 18564
rect 7532 18510 7534 18562
rect 7534 18510 7586 18562
rect 7586 18510 7588 18562
rect 7532 18508 7588 18510
rect 7308 17948 7364 18004
rect 8316 18732 8372 18788
rect 9772 19068 9828 19124
rect 9548 18620 9604 18676
rect 8988 18562 9044 18564
rect 8988 18510 8990 18562
rect 8990 18510 9042 18562
rect 9042 18510 9044 18562
rect 8988 18508 9044 18510
rect 10108 19404 10164 19460
rect 12460 24332 12516 24388
rect 14140 25394 14196 25396
rect 14140 25342 14142 25394
rect 14142 25342 14194 25394
rect 14194 25342 14196 25394
rect 14140 25340 14196 25342
rect 15372 26514 15428 26516
rect 15372 26462 15374 26514
rect 15374 26462 15426 26514
rect 15426 26462 15428 26514
rect 15372 26460 15428 26462
rect 15708 26012 15764 26068
rect 12796 25282 12852 25284
rect 12796 25230 12798 25282
rect 12798 25230 12850 25282
rect 12850 25230 12852 25282
rect 12796 25228 12852 25230
rect 13916 25228 13972 25284
rect 12908 24892 12964 24948
rect 13580 24892 13636 24948
rect 13132 24610 13188 24612
rect 13132 24558 13134 24610
rect 13134 24558 13186 24610
rect 13186 24558 13188 24610
rect 13132 24556 13188 24558
rect 13468 24556 13524 24612
rect 12908 23884 12964 23940
rect 13244 24332 13300 24388
rect 12460 22540 12516 22596
rect 13132 22540 13188 22596
rect 12572 22204 12628 22260
rect 12460 22092 12516 22148
rect 12684 21362 12740 21364
rect 12684 21310 12686 21362
rect 12686 21310 12738 21362
rect 12738 21310 12740 21362
rect 12684 21308 12740 21310
rect 12124 21084 12180 21140
rect 10668 20076 10724 20132
rect 10220 19964 10276 20020
rect 9772 18508 9828 18564
rect 8204 18172 8260 18228
rect 9884 18060 9940 18116
rect 10108 18226 10164 18228
rect 10108 18174 10110 18226
rect 10110 18174 10162 18226
rect 10162 18174 10164 18226
rect 10108 18172 10164 18174
rect 10108 17836 10164 17892
rect 8764 17724 8820 17780
rect 9100 17554 9156 17556
rect 9100 17502 9102 17554
rect 9102 17502 9154 17554
rect 9154 17502 9156 17554
rect 9100 17500 9156 17502
rect 9548 17500 9604 17556
rect 8092 17106 8148 17108
rect 8092 17054 8094 17106
rect 8094 17054 8146 17106
rect 8146 17054 8148 17106
rect 8092 17052 8148 17054
rect 8540 17106 8596 17108
rect 8540 17054 8542 17106
rect 8542 17054 8594 17106
rect 8594 17054 8596 17106
rect 8540 17052 8596 17054
rect 6972 16882 7028 16884
rect 6972 16830 6974 16882
rect 6974 16830 7026 16882
rect 7026 16830 7028 16882
rect 6972 16828 7028 16830
rect 5068 15036 5124 15092
rect 5852 15036 5908 15092
rect 6188 14028 6244 14084
rect 6076 13692 6132 13748
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 2940 13132 2996 13188
rect 4620 13074 4676 13076
rect 4620 13022 4622 13074
rect 4622 13022 4674 13074
rect 4674 13022 4676 13074
rect 4620 13020 4676 13022
rect 3724 12908 3780 12964
rect 1820 12124 1876 12180
rect 2380 12178 2436 12180
rect 2380 12126 2382 12178
rect 2382 12126 2434 12178
rect 2434 12126 2436 12178
rect 2380 12124 2436 12126
rect 5068 12908 5124 12964
rect 5404 13244 5460 13300
rect 5068 12124 5124 12180
rect 5740 13186 5796 13188
rect 5740 13134 5742 13186
rect 5742 13134 5794 13186
rect 5794 13134 5796 13186
rect 5740 13132 5796 13134
rect 6076 13074 6132 13076
rect 6076 13022 6078 13074
rect 6078 13022 6130 13074
rect 6130 13022 6132 13074
rect 6076 13020 6132 13022
rect 8652 16940 8708 16996
rect 7420 16716 7476 16772
rect 7868 16604 7924 16660
rect 7868 15708 7924 15764
rect 7980 15372 8036 15428
rect 6972 15036 7028 15092
rect 8428 15426 8484 15428
rect 8428 15374 8430 15426
rect 8430 15374 8482 15426
rect 8482 15374 8484 15426
rect 8428 15372 8484 15374
rect 8540 15148 8596 15204
rect 7084 13692 7140 13748
rect 7980 13692 8036 13748
rect 5628 12178 5684 12180
rect 5628 12126 5630 12178
rect 5630 12126 5682 12178
rect 5682 12126 5684 12178
rect 5628 12124 5684 12126
rect 6188 12178 6244 12180
rect 6188 12126 6190 12178
rect 6190 12126 6242 12178
rect 6242 12126 6244 12178
rect 6188 12124 6244 12126
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 7644 11900 7700 11956
rect 6748 11228 6804 11284
rect 8316 13746 8372 13748
rect 8316 13694 8318 13746
rect 8318 13694 8370 13746
rect 8370 13694 8372 13746
rect 8316 13692 8372 13694
rect 8764 14700 8820 14756
rect 9100 15148 9156 15204
rect 10556 18620 10612 18676
rect 11116 20018 11172 20020
rect 11116 19966 11118 20018
rect 11118 19966 11170 20018
rect 11170 19966 11172 20018
rect 11116 19964 11172 19966
rect 10668 18508 10724 18564
rect 10892 18396 10948 18452
rect 12796 20188 12852 20244
rect 12572 19458 12628 19460
rect 12572 19406 12574 19458
rect 12574 19406 12626 19458
rect 12626 19406 12628 19458
rect 12572 19404 12628 19406
rect 11116 18620 11172 18676
rect 11676 18284 11732 18340
rect 11452 18172 11508 18228
rect 11788 17948 11844 18004
rect 11676 17442 11732 17444
rect 11676 17390 11678 17442
rect 11678 17390 11730 17442
rect 11730 17390 11732 17442
rect 11676 17388 11732 17390
rect 11116 16940 11172 16996
rect 9660 15820 9716 15876
rect 9996 15314 10052 15316
rect 9996 15262 9998 15314
rect 9998 15262 10050 15314
rect 10050 15262 10052 15314
rect 9996 15260 10052 15262
rect 11564 16716 11620 16772
rect 9660 14028 9716 14084
rect 9548 13468 9604 13524
rect 8988 13244 9044 13300
rect 8988 12236 9044 12292
rect 8428 12124 8484 12180
rect 8204 11282 8260 11284
rect 8204 11230 8206 11282
rect 8206 11230 8258 11282
rect 8258 11230 8260 11282
rect 8204 11228 8260 11230
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 5740 9042 5796 9044
rect 5740 8990 5742 9042
rect 5742 8990 5794 9042
rect 5794 8990 5796 9042
rect 5740 8988 5796 8990
rect 8988 12066 9044 12068
rect 8988 12014 8990 12066
rect 8990 12014 9042 12066
rect 9042 12014 9044 12066
rect 8988 12012 9044 12014
rect 9212 12124 9268 12180
rect 9772 13746 9828 13748
rect 9772 13694 9774 13746
rect 9774 13694 9826 13746
rect 9826 13694 9828 13746
rect 9772 13692 9828 13694
rect 11116 14754 11172 14756
rect 11116 14702 11118 14754
rect 11118 14702 11170 14754
rect 11170 14702 11172 14754
rect 11116 14700 11172 14702
rect 9772 12850 9828 12852
rect 9772 12798 9774 12850
rect 9774 12798 9826 12850
rect 9826 12798 9828 12850
rect 9772 12796 9828 12798
rect 10892 14140 10948 14196
rect 10780 13858 10836 13860
rect 10780 13806 10782 13858
rect 10782 13806 10834 13858
rect 10834 13806 10836 13858
rect 10780 13804 10836 13806
rect 10780 12962 10836 12964
rect 10780 12910 10782 12962
rect 10782 12910 10834 12962
rect 10834 12910 10836 12962
rect 10780 12908 10836 12910
rect 11788 16210 11844 16212
rect 11788 16158 11790 16210
rect 11790 16158 11842 16210
rect 11842 16158 11844 16210
rect 11788 16156 11844 16158
rect 11788 15202 11844 15204
rect 11788 15150 11790 15202
rect 11790 15150 11842 15202
rect 11842 15150 11844 15202
rect 11788 15148 11844 15150
rect 12012 17554 12068 17556
rect 12012 17502 12014 17554
rect 12014 17502 12066 17554
rect 12066 17502 12068 17554
rect 12012 17500 12068 17502
rect 12348 18172 12404 18228
rect 12684 18450 12740 18452
rect 12684 18398 12686 18450
rect 12686 18398 12738 18450
rect 12738 18398 12740 18450
rect 12684 18396 12740 18398
rect 12908 19292 12964 19348
rect 13020 18396 13076 18452
rect 12796 18284 12852 18340
rect 12572 18172 12628 18228
rect 12460 17890 12516 17892
rect 12460 17838 12462 17890
rect 12462 17838 12514 17890
rect 12514 17838 12516 17890
rect 12460 17836 12516 17838
rect 12796 17612 12852 17668
rect 12348 17500 12404 17556
rect 12124 16716 12180 16772
rect 12684 16268 12740 16324
rect 12236 15708 12292 15764
rect 12796 16098 12852 16100
rect 12796 16046 12798 16098
rect 12798 16046 12850 16098
rect 12850 16046 12852 16098
rect 12796 16044 12852 16046
rect 12684 15708 12740 15764
rect 12012 14252 12068 14308
rect 11676 13804 11732 13860
rect 11564 12796 11620 12852
rect 11788 13020 11844 13076
rect 9660 11676 9716 11732
rect 11564 12012 11620 12068
rect 11676 11676 11732 11732
rect 11564 10834 11620 10836
rect 11564 10782 11566 10834
rect 11566 10782 11618 10834
rect 11618 10782 11620 10834
rect 11564 10780 11620 10782
rect 10892 10556 10948 10612
rect 8428 8988 8484 9044
rect 8540 9660 8596 9716
rect 7420 8876 7476 8932
rect 8540 8930 8596 8932
rect 8540 8878 8542 8930
rect 8542 8878 8594 8930
rect 8594 8878 8596 8930
rect 8540 8876 8596 8878
rect 8988 9042 9044 9044
rect 8988 8990 8990 9042
rect 8990 8990 9042 9042
rect 9042 8990 9044 9042
rect 8988 8988 9044 8990
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 9884 9042 9940 9044
rect 9884 8990 9886 9042
rect 9886 8990 9938 9042
rect 9938 8990 9940 9042
rect 9884 8988 9940 8990
rect 10444 9042 10500 9044
rect 10444 8990 10446 9042
rect 10446 8990 10498 9042
rect 10498 8990 10500 9042
rect 10444 8988 10500 8990
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 11004 10498 11060 10500
rect 11004 10446 11006 10498
rect 11006 10446 11058 10498
rect 11058 10446 11060 10498
rect 11004 10444 11060 10446
rect 12012 12796 12068 12852
rect 12572 15260 12628 15316
rect 13244 21084 13300 21140
rect 13692 23324 13748 23380
rect 13692 22764 13748 22820
rect 14364 23436 14420 23492
rect 14028 23324 14084 23380
rect 14924 24610 14980 24612
rect 14924 24558 14926 24610
rect 14926 24558 14978 24610
rect 14978 24558 14980 24610
rect 14924 24556 14980 24558
rect 15260 23436 15316 23492
rect 15596 23212 15652 23268
rect 14588 22764 14644 22820
rect 13580 22204 13636 22260
rect 14252 21756 14308 21812
rect 14364 21586 14420 21588
rect 14364 21534 14366 21586
rect 14366 21534 14418 21586
rect 14418 21534 14420 21586
rect 14364 21532 14420 21534
rect 13468 21308 13524 21364
rect 13916 21196 13972 21252
rect 13356 19794 13412 19796
rect 13356 19742 13358 19794
rect 13358 19742 13410 19794
rect 13410 19742 13412 19794
rect 13356 19740 13412 19742
rect 13804 20748 13860 20804
rect 14028 20188 14084 20244
rect 14364 20524 14420 20580
rect 13916 20076 13972 20132
rect 13692 19964 13748 20020
rect 13580 19740 13636 19796
rect 13468 19292 13524 19348
rect 13580 19180 13636 19236
rect 13356 17500 13412 17556
rect 13244 16156 13300 16212
rect 13692 18956 13748 19012
rect 14028 19964 14084 20020
rect 13692 18620 13748 18676
rect 13692 18172 13748 18228
rect 13916 18732 13972 18788
rect 14140 18620 14196 18676
rect 14924 22652 14980 22708
rect 14588 22258 14644 22260
rect 14588 22206 14590 22258
rect 14590 22206 14642 22258
rect 14642 22206 14644 22258
rect 14588 22204 14644 22206
rect 15260 21980 15316 22036
rect 15036 21868 15092 21924
rect 14476 19180 14532 19236
rect 15148 20802 15204 20804
rect 15148 20750 15150 20802
rect 15150 20750 15202 20802
rect 15202 20750 15204 20802
rect 15148 20748 15204 20750
rect 15372 20188 15428 20244
rect 14700 20018 14756 20020
rect 14700 19966 14702 20018
rect 14702 19966 14754 20018
rect 14754 19966 14756 20018
rect 14700 19964 14756 19966
rect 15820 22764 15876 22820
rect 15708 21980 15764 22036
rect 16156 26012 16212 26068
rect 16380 23436 16436 23492
rect 16380 23266 16436 23268
rect 16380 23214 16382 23266
rect 16382 23214 16434 23266
rect 16434 23214 16436 23266
rect 16380 23212 16436 23214
rect 16156 22428 16212 22484
rect 16380 22146 16436 22148
rect 16380 22094 16382 22146
rect 16382 22094 16434 22146
rect 16434 22094 16436 22146
rect 16380 22092 16436 22094
rect 15932 21698 15988 21700
rect 15932 21646 15934 21698
rect 15934 21646 15986 21698
rect 15986 21646 15988 21698
rect 15932 21644 15988 21646
rect 15596 21532 15652 21588
rect 16156 21308 16212 21364
rect 16156 21084 16212 21140
rect 15932 20748 15988 20804
rect 14924 20018 14980 20020
rect 14924 19966 14926 20018
rect 14926 19966 14978 20018
rect 14978 19966 14980 20018
rect 14924 19964 14980 19966
rect 14252 18844 14308 18900
rect 16380 20188 16436 20244
rect 15148 18956 15204 19012
rect 13804 17666 13860 17668
rect 13804 17614 13806 17666
rect 13806 17614 13858 17666
rect 13858 17614 13860 17666
rect 13804 17612 13860 17614
rect 14028 17948 14084 18004
rect 14252 17890 14308 17892
rect 14252 17838 14254 17890
rect 14254 17838 14306 17890
rect 14306 17838 14308 17890
rect 14252 17836 14308 17838
rect 14252 17388 14308 17444
rect 13692 16044 13748 16100
rect 13580 15874 13636 15876
rect 13580 15822 13582 15874
rect 13582 15822 13634 15874
rect 13634 15822 13636 15874
rect 13580 15820 13636 15822
rect 13580 15372 13636 15428
rect 14140 16098 14196 16100
rect 14140 16046 14142 16098
rect 14142 16046 14194 16098
rect 14194 16046 14196 16098
rect 14140 16044 14196 16046
rect 13804 15484 13860 15540
rect 13916 15932 13972 15988
rect 13244 15260 13300 15316
rect 12572 14476 12628 14532
rect 13132 14476 13188 14532
rect 12236 14140 12292 14196
rect 12684 14364 12740 14420
rect 12460 13132 12516 13188
rect 12684 13468 12740 13524
rect 12572 13074 12628 13076
rect 12572 13022 12574 13074
rect 12574 13022 12626 13074
rect 12626 13022 12628 13074
rect 12572 13020 12628 13022
rect 12236 12012 12292 12068
rect 12572 12012 12628 12068
rect 12236 11564 12292 11620
rect 12124 10834 12180 10836
rect 12124 10782 12126 10834
rect 12126 10782 12178 10834
rect 12178 10782 12180 10834
rect 12124 10780 12180 10782
rect 11788 10556 11844 10612
rect 11228 9938 11284 9940
rect 11228 9886 11230 9938
rect 11230 9886 11282 9938
rect 11282 9886 11284 9938
rect 11228 9884 11284 9886
rect 12012 9938 12068 9940
rect 12012 9886 12014 9938
rect 12014 9886 12066 9938
rect 12066 9886 12068 9938
rect 12012 9884 12068 9886
rect 11564 9548 11620 9604
rect 12460 10444 12516 10500
rect 12908 13692 12964 13748
rect 13020 13132 13076 13188
rect 12908 13020 12964 13076
rect 13132 12908 13188 12964
rect 13468 14418 13524 14420
rect 13468 14366 13470 14418
rect 13470 14366 13522 14418
rect 13522 14366 13524 14418
rect 13468 14364 13524 14366
rect 15036 18450 15092 18452
rect 15036 18398 15038 18450
rect 15038 18398 15090 18450
rect 15090 18398 15092 18450
rect 15036 18396 15092 18398
rect 15148 17948 15204 18004
rect 16044 19180 16100 19236
rect 15260 17836 15316 17892
rect 15596 18060 15652 18116
rect 15036 16994 15092 16996
rect 15036 16942 15038 16994
rect 15038 16942 15090 16994
rect 15090 16942 15092 16994
rect 15036 16940 15092 16942
rect 14700 16604 14756 16660
rect 15148 16828 15204 16884
rect 14476 15538 14532 15540
rect 14476 15486 14478 15538
rect 14478 15486 14530 15538
rect 14530 15486 14532 15538
rect 14476 15484 14532 15486
rect 14924 15426 14980 15428
rect 14924 15374 14926 15426
rect 14926 15374 14978 15426
rect 14978 15374 14980 15426
rect 14924 15372 14980 15374
rect 13916 14252 13972 14308
rect 13692 12796 13748 12852
rect 14028 12850 14084 12852
rect 14028 12798 14030 12850
rect 14030 12798 14082 12850
rect 14082 12798 14084 12850
rect 14028 12796 14084 12798
rect 14028 12290 14084 12292
rect 14028 12238 14030 12290
rect 14030 12238 14082 12290
rect 14082 12238 14084 12290
rect 14028 12236 14084 12238
rect 13468 12066 13524 12068
rect 13468 12014 13470 12066
rect 13470 12014 13522 12066
rect 13522 12014 13524 12066
rect 13468 12012 13524 12014
rect 13244 11564 13300 11620
rect 12572 9714 12628 9716
rect 12572 9662 12574 9714
rect 12574 9662 12626 9714
rect 12626 9662 12628 9714
rect 12572 9660 12628 9662
rect 14028 9826 14084 9828
rect 14028 9774 14030 9826
rect 14030 9774 14082 9826
rect 14082 9774 14084 9826
rect 14028 9772 14084 9774
rect 13356 9154 13412 9156
rect 13356 9102 13358 9154
rect 13358 9102 13410 9154
rect 13410 9102 13412 9154
rect 13356 9100 13412 9102
rect 14364 13186 14420 13188
rect 14364 13134 14366 13186
rect 14366 13134 14418 13186
rect 14418 13134 14420 13186
rect 14364 13132 14420 13134
rect 14700 14306 14756 14308
rect 14700 14254 14702 14306
rect 14702 14254 14754 14306
rect 14754 14254 14756 14306
rect 14700 14252 14756 14254
rect 14476 12348 14532 12404
rect 15148 14252 15204 14308
rect 17948 30156 18004 30212
rect 19740 31948 19796 32004
rect 20076 31500 20132 31556
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19068 30994 19124 30996
rect 19068 30942 19070 30994
rect 19070 30942 19122 30994
rect 19122 30942 19124 30994
rect 19068 30940 19124 30942
rect 19516 30492 19572 30548
rect 18396 29484 18452 29540
rect 18060 29260 18116 29316
rect 16716 28754 16772 28756
rect 16716 28702 16718 28754
rect 16718 28702 16770 28754
rect 16770 28702 16772 28754
rect 16716 28700 16772 28702
rect 17948 26236 18004 26292
rect 17836 26178 17892 26180
rect 17836 26126 17838 26178
rect 17838 26126 17890 26178
rect 17890 26126 17892 26178
rect 17836 26124 17892 26126
rect 17500 24610 17556 24612
rect 17500 24558 17502 24610
rect 17502 24558 17554 24610
rect 17554 24558 17556 24610
rect 17500 24556 17556 24558
rect 17948 23436 18004 23492
rect 18620 29260 18676 29316
rect 18956 29314 19012 29316
rect 18956 29262 18958 29314
rect 18958 29262 19010 29314
rect 19010 29262 19012 29314
rect 18956 29260 19012 29262
rect 19740 30210 19796 30212
rect 19740 30158 19742 30210
rect 19742 30158 19794 30210
rect 19794 30158 19796 30210
rect 19740 30156 19796 30158
rect 20972 34860 21028 34916
rect 20748 34300 20804 34356
rect 21868 40572 21924 40628
rect 22876 41356 22932 41412
rect 22316 40908 22372 40964
rect 22092 40236 22148 40292
rect 23100 41746 23156 41748
rect 23100 41694 23102 41746
rect 23102 41694 23154 41746
rect 23154 41694 23156 41746
rect 23100 41692 23156 41694
rect 23100 41132 23156 41188
rect 22540 40402 22596 40404
rect 22540 40350 22542 40402
rect 22542 40350 22594 40402
rect 22594 40350 22596 40402
rect 22540 40348 22596 40350
rect 22092 39340 22148 39396
rect 22204 39004 22260 39060
rect 23100 40572 23156 40628
rect 22988 39564 23044 39620
rect 22764 38668 22820 38724
rect 22876 38780 22932 38836
rect 21868 37436 21924 37492
rect 21980 37042 22036 37044
rect 21980 36990 21982 37042
rect 21982 36990 22034 37042
rect 22034 36990 22036 37042
rect 21980 36988 22036 36990
rect 21868 36316 21924 36372
rect 21980 36540 22036 36596
rect 21420 34636 21476 34692
rect 22652 38050 22708 38052
rect 22652 37998 22654 38050
rect 22654 37998 22706 38050
rect 22706 37998 22708 38050
rect 22652 37996 22708 37998
rect 22204 36764 22260 36820
rect 22988 36988 23044 37044
rect 22092 36428 22148 36484
rect 22652 36370 22708 36372
rect 22652 36318 22654 36370
rect 22654 36318 22706 36370
rect 22706 36318 22708 36370
rect 22652 36316 22708 36318
rect 22204 35868 22260 35924
rect 21980 35756 22036 35812
rect 22316 35756 22372 35812
rect 22204 35532 22260 35588
rect 22876 35810 22932 35812
rect 22876 35758 22878 35810
rect 22878 35758 22930 35810
rect 22930 35758 22932 35810
rect 22876 35756 22932 35758
rect 22428 35698 22484 35700
rect 22428 35646 22430 35698
rect 22430 35646 22482 35698
rect 22482 35646 22484 35698
rect 22428 35644 22484 35646
rect 22764 35644 22820 35700
rect 20748 32172 20804 32228
rect 21196 30604 21252 30660
rect 21980 34636 22036 34692
rect 21980 34188 22036 34244
rect 22092 33292 22148 33348
rect 21756 32284 21812 32340
rect 21420 30492 21476 30548
rect 21868 31666 21924 31668
rect 21868 31614 21870 31666
rect 21870 31614 21922 31666
rect 21922 31614 21924 31666
rect 21868 31612 21924 31614
rect 21980 31554 22036 31556
rect 21980 31502 21982 31554
rect 21982 31502 22034 31554
rect 22034 31502 22036 31554
rect 21980 31500 22036 31502
rect 21644 30716 21700 30772
rect 22204 32060 22260 32116
rect 22652 34914 22708 34916
rect 22652 34862 22654 34914
rect 22654 34862 22706 34914
rect 22706 34862 22708 34914
rect 22652 34860 22708 34862
rect 23436 42364 23492 42420
rect 23436 41916 23492 41972
rect 23324 41468 23380 41524
rect 23884 47740 23940 47796
rect 23772 47516 23828 47572
rect 23884 46786 23940 46788
rect 23884 46734 23886 46786
rect 23886 46734 23938 46786
rect 23938 46734 23940 46786
rect 23884 46732 23940 46734
rect 23772 46508 23828 46564
rect 24332 48242 24388 48244
rect 24332 48190 24334 48242
rect 24334 48190 24386 48242
rect 24386 48190 24388 48242
rect 24332 48188 24388 48190
rect 24108 47628 24164 47684
rect 24220 47404 24276 47460
rect 24556 49810 24612 49812
rect 24556 49758 24558 49810
rect 24558 49758 24610 49810
rect 24610 49758 24612 49810
rect 24556 49756 24612 49758
rect 24668 48354 24724 48356
rect 24668 48302 24670 48354
rect 24670 48302 24722 48354
rect 24722 48302 24724 48354
rect 24668 48300 24724 48302
rect 24332 47180 24388 47236
rect 24220 47068 24276 47124
rect 24108 46620 24164 46676
rect 23996 45164 24052 45220
rect 23884 44604 23940 44660
rect 23996 44380 24052 44436
rect 24444 46562 24500 46564
rect 24444 46510 24446 46562
rect 24446 46510 24498 46562
rect 24498 46510 24500 46562
rect 24444 46508 24500 46510
rect 24332 46396 24388 46452
rect 24444 46060 24500 46116
rect 24668 47068 24724 47124
rect 24556 45724 24612 45780
rect 24556 45218 24612 45220
rect 24556 45166 24558 45218
rect 24558 45166 24610 45218
rect 24610 45166 24612 45218
rect 24556 45164 24612 45166
rect 24444 44322 24500 44324
rect 24444 44270 24446 44322
rect 24446 44270 24498 44322
rect 24498 44270 24500 44322
rect 24444 44268 24500 44270
rect 23884 43372 23940 43428
rect 23772 42924 23828 42980
rect 23884 42754 23940 42756
rect 23884 42702 23886 42754
rect 23886 42702 23938 42754
rect 23938 42702 23940 42754
rect 23884 42700 23940 42702
rect 24220 43650 24276 43652
rect 24220 43598 24222 43650
rect 24222 43598 24274 43650
rect 24274 43598 24276 43650
rect 24220 43596 24276 43598
rect 24444 43260 24500 43316
rect 24444 42642 24500 42644
rect 24444 42590 24446 42642
rect 24446 42590 24498 42642
rect 24498 42590 24500 42642
rect 24444 42588 24500 42590
rect 25004 47234 25060 47236
rect 25004 47182 25006 47234
rect 25006 47182 25058 47234
rect 25058 47182 25060 47234
rect 25004 47180 25060 47182
rect 26796 49644 26852 49700
rect 26460 49532 26516 49588
rect 26012 49138 26068 49140
rect 26012 49086 26014 49138
rect 26014 49086 26066 49138
rect 26066 49086 26068 49138
rect 26012 49084 26068 49086
rect 25564 48972 25620 49028
rect 30716 53116 30772 53172
rect 33180 54402 33236 54404
rect 33180 54350 33182 54402
rect 33182 54350 33234 54402
rect 33234 54350 33236 54402
rect 33180 54348 33236 54350
rect 31164 53730 31220 53732
rect 31164 53678 31166 53730
rect 31166 53678 31218 53730
rect 31218 53678 31220 53730
rect 31164 53676 31220 53678
rect 32284 53676 32340 53732
rect 33292 53676 33348 53732
rect 32508 53058 32564 53060
rect 32508 53006 32510 53058
rect 32510 53006 32562 53058
rect 32562 53006 32564 53058
rect 32508 53004 32564 53006
rect 31276 52050 31332 52052
rect 31276 51998 31278 52050
rect 31278 51998 31330 52050
rect 31330 51998 31332 52050
rect 31276 51996 31332 51998
rect 35420 57036 35476 57092
rect 35308 56306 35364 56308
rect 35308 56254 35310 56306
rect 35310 56254 35362 56306
rect 35362 56254 35364 56306
rect 35308 56252 35364 56254
rect 36316 56252 36372 56308
rect 36428 56924 36484 56980
rect 35756 56028 35812 56084
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35980 55804 36036 55860
rect 37548 56082 37604 56084
rect 37548 56030 37550 56082
rect 37550 56030 37602 56082
rect 37602 56030 37604 56082
rect 37548 56028 37604 56030
rect 37996 57036 38052 57092
rect 38108 56588 38164 56644
rect 39452 56924 39508 56980
rect 39116 56306 39172 56308
rect 39116 56254 39118 56306
rect 39118 56254 39170 56306
rect 39170 56254 39172 56306
rect 39116 56252 39172 56254
rect 34972 55132 35028 55188
rect 36092 55186 36148 55188
rect 36092 55134 36094 55186
rect 36094 55134 36146 55186
rect 36146 55134 36148 55186
rect 36092 55132 36148 55134
rect 34300 54402 34356 54404
rect 34300 54350 34302 54402
rect 34302 54350 34354 54402
rect 34354 54350 34356 54402
rect 34300 54348 34356 54350
rect 34860 54402 34916 54404
rect 34860 54350 34862 54402
rect 34862 54350 34914 54402
rect 34914 54350 34916 54402
rect 34860 54348 34916 54350
rect 35308 54348 35364 54404
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 34748 53228 34804 53284
rect 34636 53170 34692 53172
rect 34636 53118 34638 53170
rect 34638 53118 34690 53170
rect 34690 53118 34692 53170
rect 34636 53116 34692 53118
rect 35308 53506 35364 53508
rect 35308 53454 35310 53506
rect 35310 53454 35362 53506
rect 35362 53454 35364 53506
rect 35308 53452 35364 53454
rect 35532 52946 35588 52948
rect 35532 52894 35534 52946
rect 35534 52894 35586 52946
rect 35586 52894 35588 52946
rect 35532 52892 35588 52894
rect 40348 56812 40404 56868
rect 40348 56588 40404 56644
rect 41692 57036 41748 57092
rect 42028 56924 42084 56980
rect 42140 56252 42196 56308
rect 42924 56812 42980 56868
rect 41468 55186 41524 55188
rect 41468 55134 41470 55186
rect 41470 55134 41522 55186
rect 41522 55134 41524 55186
rect 41468 55132 41524 55134
rect 38668 53842 38724 53844
rect 38668 53790 38670 53842
rect 38670 53790 38722 53842
rect 38722 53790 38724 53842
rect 38668 53788 38724 53790
rect 38108 53452 38164 53508
rect 37212 53058 37268 53060
rect 37212 53006 37214 53058
rect 37214 53006 37266 53058
rect 37266 53006 37268 53058
rect 37212 53004 37268 53006
rect 29260 51212 29316 51268
rect 28140 49868 28196 49924
rect 28140 49698 28196 49700
rect 28140 49646 28142 49698
rect 28142 49646 28194 49698
rect 28194 49646 28196 49698
rect 28140 49644 28196 49646
rect 27020 49084 27076 49140
rect 26684 48914 26740 48916
rect 26684 48862 26686 48914
rect 26686 48862 26738 48914
rect 26738 48862 26740 48914
rect 26684 48860 26740 48862
rect 25788 48300 25844 48356
rect 26012 48242 26068 48244
rect 26012 48190 26014 48242
rect 26014 48190 26066 48242
rect 26066 48190 26068 48242
rect 26012 48188 26068 48190
rect 26460 47628 26516 47684
rect 26572 47740 26628 47796
rect 25452 47068 25508 47124
rect 25340 46732 25396 46788
rect 25676 46956 25732 47012
rect 25788 46620 25844 46676
rect 25340 46396 25396 46452
rect 27356 49026 27412 49028
rect 27356 48974 27358 49026
rect 27358 48974 27410 49026
rect 27410 48974 27412 49026
rect 27356 48972 27412 48974
rect 27244 48914 27300 48916
rect 27244 48862 27246 48914
rect 27246 48862 27298 48914
rect 27298 48862 27300 48914
rect 27244 48860 27300 48862
rect 27580 49084 27636 49140
rect 27468 48636 27524 48692
rect 29036 49868 29092 49924
rect 28364 48972 28420 49028
rect 27804 48636 27860 48692
rect 26684 47292 26740 47348
rect 26124 46732 26180 46788
rect 26348 46956 26404 47012
rect 26124 46396 26180 46452
rect 25228 45500 25284 45556
rect 24780 44268 24836 44324
rect 25004 44380 25060 44436
rect 25452 43820 25508 43876
rect 24892 43596 24948 43652
rect 24780 43484 24836 43540
rect 24668 42700 24724 42756
rect 25116 43036 25172 43092
rect 26012 44828 26068 44884
rect 26796 47068 26852 47124
rect 27356 47068 27412 47124
rect 27132 46956 27188 47012
rect 26572 46732 26628 46788
rect 26572 46396 26628 46452
rect 26684 46508 26740 46564
rect 26460 45836 26516 45892
rect 28252 48130 28308 48132
rect 28252 48078 28254 48130
rect 28254 48078 28306 48130
rect 28306 48078 28308 48130
rect 28252 48076 28308 48078
rect 28140 47964 28196 48020
rect 27692 47068 27748 47124
rect 27020 46508 27076 46564
rect 27132 46060 27188 46116
rect 27244 46396 27300 46452
rect 27692 46450 27748 46452
rect 27692 46398 27694 46450
rect 27694 46398 27746 46450
rect 27746 46398 27748 46450
rect 27692 46396 27748 46398
rect 27804 46172 27860 46228
rect 26236 45052 26292 45108
rect 25788 44380 25844 44436
rect 26572 44044 26628 44100
rect 26012 43820 26068 43876
rect 25676 43538 25732 43540
rect 25676 43486 25678 43538
rect 25678 43486 25730 43538
rect 25730 43486 25732 43538
rect 25676 43484 25732 43486
rect 25564 43260 25620 43316
rect 25340 42700 25396 42756
rect 26012 42924 26068 42980
rect 26348 43820 26404 43876
rect 27356 45890 27412 45892
rect 27356 45838 27358 45890
rect 27358 45838 27410 45890
rect 27410 45838 27412 45890
rect 27356 45836 27412 45838
rect 27804 45890 27860 45892
rect 27804 45838 27806 45890
rect 27806 45838 27858 45890
rect 27858 45838 27860 45890
rect 27804 45836 27860 45838
rect 28140 47516 28196 47572
rect 29148 49196 29204 49252
rect 28924 48860 28980 48916
rect 28700 48524 28756 48580
rect 28700 48300 28756 48356
rect 29036 48076 29092 48132
rect 28140 47180 28196 47236
rect 29484 49026 29540 49028
rect 29484 48974 29486 49026
rect 29486 48974 29538 49026
rect 29538 48974 29540 49026
rect 29484 48972 29540 48974
rect 30044 48972 30100 49028
rect 29372 48748 29428 48804
rect 29708 48802 29764 48804
rect 29708 48750 29710 48802
rect 29710 48750 29762 48802
rect 29762 48750 29764 48802
rect 29708 48748 29764 48750
rect 30604 49586 30660 49588
rect 30604 49534 30606 49586
rect 30606 49534 30658 49586
rect 30658 49534 30660 49586
rect 30604 49532 30660 49534
rect 33628 51772 33684 51828
rect 33516 51436 33572 51492
rect 33852 51490 33908 51492
rect 33852 51438 33854 51490
rect 33854 51438 33906 51490
rect 33906 51438 33908 51490
rect 33852 51436 33908 51438
rect 33740 51266 33796 51268
rect 33740 51214 33742 51266
rect 33742 51214 33794 51266
rect 33794 51214 33796 51266
rect 33740 51212 33796 51214
rect 34300 51884 34356 51940
rect 35084 52834 35140 52836
rect 35084 52782 35086 52834
rect 35086 52782 35138 52834
rect 35138 52782 35140 52834
rect 35084 52780 35140 52782
rect 34860 52668 34916 52724
rect 34412 51548 34468 51604
rect 35308 52722 35364 52724
rect 35308 52670 35310 52722
rect 35310 52670 35362 52722
rect 35362 52670 35364 52722
rect 35308 52668 35364 52670
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34300 51212 34356 51268
rect 35644 52444 35700 52500
rect 36092 52946 36148 52948
rect 36092 52894 36094 52946
rect 36094 52894 36146 52946
rect 36146 52894 36148 52946
rect 36092 52892 36148 52894
rect 38780 53452 38836 53508
rect 35980 52332 36036 52388
rect 35532 51660 35588 51716
rect 37660 52722 37716 52724
rect 37660 52670 37662 52722
rect 37662 52670 37714 52722
rect 37714 52670 37716 52722
rect 37660 52668 37716 52670
rect 37660 52332 37716 52388
rect 37884 52220 37940 52276
rect 37996 52050 38052 52052
rect 37996 51998 37998 52050
rect 37998 51998 38050 52050
rect 38050 51998 38052 52050
rect 37996 51996 38052 51998
rect 35756 51660 35812 51716
rect 36092 51772 36148 51828
rect 35980 51602 36036 51604
rect 35980 51550 35982 51602
rect 35982 51550 36034 51602
rect 36034 51550 36036 51602
rect 35980 51548 36036 51550
rect 34860 51324 34916 51380
rect 35196 51324 35252 51380
rect 36316 51378 36372 51380
rect 36316 51326 36318 51378
rect 36318 51326 36370 51378
rect 36370 51326 36372 51378
rect 36316 51324 36372 51326
rect 34972 51154 35028 51156
rect 34972 51102 34974 51154
rect 34974 51102 35026 51154
rect 35026 51102 35028 51154
rect 34972 51100 35028 51102
rect 34636 50764 34692 50820
rect 34748 50594 34804 50596
rect 34748 50542 34750 50594
rect 34750 50542 34802 50594
rect 34802 50542 34804 50594
rect 34748 50540 34804 50542
rect 30268 48300 30324 48356
rect 30716 48524 30772 48580
rect 29260 47682 29316 47684
rect 29260 47630 29262 47682
rect 29262 47630 29314 47682
rect 29314 47630 29316 47682
rect 29260 47628 29316 47630
rect 28812 47516 28868 47572
rect 28700 46898 28756 46900
rect 28700 46846 28702 46898
rect 28702 46846 28754 46898
rect 28754 46846 28756 46898
rect 28700 46844 28756 46846
rect 28028 45948 28084 46004
rect 28140 46060 28196 46116
rect 27916 45724 27972 45780
rect 27132 45612 27188 45668
rect 26796 45218 26852 45220
rect 26796 45166 26798 45218
rect 26798 45166 26850 45218
rect 26850 45166 26852 45218
rect 26796 45164 26852 45166
rect 27020 45388 27076 45444
rect 27244 44994 27300 44996
rect 27244 44942 27246 44994
rect 27246 44942 27298 44994
rect 27298 44942 27300 44994
rect 27244 44940 27300 44942
rect 28476 45836 28532 45892
rect 27916 45164 27972 45220
rect 27692 45106 27748 45108
rect 27692 45054 27694 45106
rect 27694 45054 27746 45106
rect 27746 45054 27748 45106
rect 27692 45052 27748 45054
rect 28140 45164 28196 45220
rect 27356 44380 27412 44436
rect 26684 43484 26740 43540
rect 27020 44156 27076 44212
rect 27356 44210 27412 44212
rect 27356 44158 27358 44210
rect 27358 44158 27410 44210
rect 27410 44158 27412 44210
rect 27356 44156 27412 44158
rect 26796 42924 26852 42980
rect 26348 42812 26404 42868
rect 26124 42588 26180 42644
rect 24108 42194 24164 42196
rect 24108 42142 24110 42194
rect 24110 42142 24162 42194
rect 24162 42142 24164 42194
rect 24108 42140 24164 42142
rect 25228 42364 25284 42420
rect 24332 42028 24388 42084
rect 23884 41804 23940 41860
rect 23884 41244 23940 41300
rect 23436 40908 23492 40964
rect 23324 40236 23380 40292
rect 23660 38834 23716 38836
rect 23660 38782 23662 38834
rect 23662 38782 23714 38834
rect 23714 38782 23716 38834
rect 23660 38780 23716 38782
rect 23996 41186 24052 41188
rect 23996 41134 23998 41186
rect 23998 41134 24050 41186
rect 24050 41134 24052 41186
rect 23996 41132 24052 41134
rect 24444 41916 24500 41972
rect 23884 40012 23940 40068
rect 23996 40178 24052 40180
rect 23996 40126 23998 40178
rect 23998 40126 24050 40178
rect 24050 40126 24052 40178
rect 23996 40124 24052 40126
rect 23436 38556 23492 38612
rect 23324 36988 23380 37044
rect 23436 35532 23492 35588
rect 24556 41356 24612 41412
rect 25452 42364 25508 42420
rect 25340 42082 25396 42084
rect 25340 42030 25342 42082
rect 25342 42030 25394 42082
rect 25394 42030 25396 42082
rect 25340 42028 25396 42030
rect 25900 42364 25956 42420
rect 26796 42140 26852 42196
rect 26908 42364 26964 42420
rect 28140 43932 28196 43988
rect 28364 45388 28420 45444
rect 28476 45164 28532 45220
rect 28588 45106 28644 45108
rect 28588 45054 28590 45106
rect 28590 45054 28642 45106
rect 28642 45054 28644 45106
rect 28588 45052 28644 45054
rect 29148 47180 29204 47236
rect 29036 47068 29092 47124
rect 29260 46844 29316 46900
rect 30268 48018 30324 48020
rect 30268 47966 30270 48018
rect 30270 47966 30322 48018
rect 30322 47966 30324 48018
rect 30268 47964 30324 47966
rect 30044 47516 30100 47572
rect 29596 46956 29652 47012
rect 29820 46562 29876 46564
rect 29820 46510 29822 46562
rect 29822 46510 29874 46562
rect 29874 46510 29876 46562
rect 29820 46508 29876 46510
rect 29260 45836 29316 45892
rect 29372 45388 29428 45444
rect 29372 45052 29428 45108
rect 28588 43932 28644 43988
rect 28476 43708 28532 43764
rect 28028 43650 28084 43652
rect 28028 43598 28030 43650
rect 28030 43598 28082 43650
rect 28082 43598 28084 43650
rect 28028 43596 28084 43598
rect 27692 43484 27748 43540
rect 27580 43036 27636 43092
rect 27916 43372 27972 43428
rect 27356 42866 27412 42868
rect 27356 42814 27358 42866
rect 27358 42814 27410 42866
rect 27410 42814 27412 42866
rect 27356 42812 27412 42814
rect 28028 43148 28084 43204
rect 27132 42364 27188 42420
rect 25228 41356 25284 41412
rect 25788 41970 25844 41972
rect 25788 41918 25790 41970
rect 25790 41918 25842 41970
rect 25842 41918 25844 41970
rect 25788 41916 25844 41918
rect 26348 41804 26404 41860
rect 24668 41186 24724 41188
rect 24668 41134 24670 41186
rect 24670 41134 24722 41186
rect 24722 41134 24724 41186
rect 24668 41132 24724 41134
rect 25900 41356 25956 41412
rect 25676 41186 25732 41188
rect 25676 41134 25678 41186
rect 25678 41134 25730 41186
rect 25730 41134 25732 41186
rect 25676 41132 25732 41134
rect 24556 40236 24612 40292
rect 24668 40908 24724 40964
rect 24444 38834 24500 38836
rect 24444 38782 24446 38834
rect 24446 38782 24498 38834
rect 24498 38782 24500 38834
rect 24444 38780 24500 38782
rect 23660 38050 23716 38052
rect 23660 37998 23662 38050
rect 23662 37998 23714 38050
rect 23714 37998 23716 38050
rect 23660 37996 23716 37998
rect 24332 37938 24388 37940
rect 24332 37886 24334 37938
rect 24334 37886 24386 37938
rect 24386 37886 24388 37938
rect 24332 37884 24388 37886
rect 25788 40626 25844 40628
rect 25788 40574 25790 40626
rect 25790 40574 25842 40626
rect 25842 40574 25844 40626
rect 25788 40572 25844 40574
rect 25004 40348 25060 40404
rect 25452 40124 25508 40180
rect 26012 41244 26068 41300
rect 26124 41580 26180 41636
rect 25564 40348 25620 40404
rect 25452 39788 25508 39844
rect 25228 39618 25284 39620
rect 25228 39566 25230 39618
rect 25230 39566 25282 39618
rect 25282 39566 25284 39618
rect 25228 39564 25284 39566
rect 25004 38444 25060 38500
rect 25228 38556 25284 38612
rect 25340 38162 25396 38164
rect 25340 38110 25342 38162
rect 25342 38110 25394 38162
rect 25394 38110 25396 38162
rect 25340 38108 25396 38110
rect 25004 37996 25060 38052
rect 24668 37660 24724 37716
rect 24444 36988 24500 37044
rect 24108 36428 24164 36484
rect 25340 37884 25396 37940
rect 25564 37884 25620 37940
rect 25228 37660 25284 37716
rect 23884 35698 23940 35700
rect 23884 35646 23886 35698
rect 23886 35646 23938 35698
rect 23938 35646 23940 35698
rect 23884 35644 23940 35646
rect 23100 34636 23156 34692
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 21308 29820 21364 29876
rect 22092 29820 22148 29876
rect 20044 29764 20100 29766
rect 21308 29260 21364 29316
rect 18956 28418 19012 28420
rect 18956 28366 18958 28418
rect 18958 28366 19010 28418
rect 19010 28366 19012 28418
rect 18956 28364 19012 28366
rect 18844 28028 18900 28084
rect 18732 27186 18788 27188
rect 18732 27134 18734 27186
rect 18734 27134 18786 27186
rect 18786 27134 18788 27186
rect 18732 27132 18788 27134
rect 18620 26908 18676 26964
rect 19068 26684 19124 26740
rect 21308 28530 21364 28532
rect 21308 28478 21310 28530
rect 21310 28478 21362 28530
rect 21362 28478 21364 28530
rect 21308 28476 21364 28478
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19740 28082 19796 28084
rect 19740 28030 19742 28082
rect 19742 28030 19794 28082
rect 19794 28030 19796 28082
rect 19740 28028 19796 28030
rect 20188 27916 20244 27972
rect 20524 27970 20580 27972
rect 20524 27918 20526 27970
rect 20526 27918 20578 27970
rect 20578 27918 20580 27970
rect 20524 27916 20580 27918
rect 20748 27858 20804 27860
rect 20748 27806 20750 27858
rect 20750 27806 20802 27858
rect 20802 27806 20804 27858
rect 20748 27804 20804 27806
rect 19292 26796 19348 26852
rect 18620 26290 18676 26292
rect 18620 26238 18622 26290
rect 18622 26238 18674 26290
rect 18674 26238 18676 26290
rect 18620 26236 18676 26238
rect 18844 26236 18900 26292
rect 18284 25452 18340 25508
rect 18620 25900 18676 25956
rect 18284 25116 18340 25172
rect 18396 24946 18452 24948
rect 18396 24894 18398 24946
rect 18398 24894 18450 24946
rect 18450 24894 18452 24946
rect 18396 24892 18452 24894
rect 17500 23266 17556 23268
rect 17500 23214 17502 23266
rect 17502 23214 17554 23266
rect 17554 23214 17556 23266
rect 17500 23212 17556 23214
rect 16716 22652 16772 22708
rect 16940 22428 16996 22484
rect 16716 22258 16772 22260
rect 16716 22206 16718 22258
rect 16718 22206 16770 22258
rect 16770 22206 16772 22258
rect 16716 22204 16772 22206
rect 17948 22370 18004 22372
rect 17948 22318 17950 22370
rect 17950 22318 18002 22370
rect 18002 22318 18004 22370
rect 17948 22316 18004 22318
rect 17164 22258 17220 22260
rect 17164 22206 17166 22258
rect 17166 22206 17218 22258
rect 17218 22206 17220 22258
rect 17164 22204 17220 22206
rect 18396 23938 18452 23940
rect 18396 23886 18398 23938
rect 18398 23886 18450 23938
rect 18450 23886 18452 23938
rect 18396 23884 18452 23886
rect 16604 19180 16660 19236
rect 16604 19010 16660 19012
rect 16604 18958 16606 19010
rect 16606 18958 16658 19010
rect 16658 18958 16660 19010
rect 16604 18956 16660 18958
rect 16604 18620 16660 18676
rect 16940 18396 16996 18452
rect 16716 17836 16772 17892
rect 15820 17052 15876 17108
rect 15932 16940 15988 16996
rect 16380 17554 16436 17556
rect 16380 17502 16382 17554
rect 16382 17502 16434 17554
rect 16434 17502 16436 17554
rect 16380 17500 16436 17502
rect 16604 17388 16660 17444
rect 16492 17106 16548 17108
rect 16492 17054 16494 17106
rect 16494 17054 16546 17106
rect 16546 17054 16548 17106
rect 16492 17052 16548 17054
rect 16156 16716 16212 16772
rect 16716 17052 16772 17108
rect 16604 16716 16660 16772
rect 16716 16492 16772 16548
rect 16268 15820 16324 15876
rect 16828 16380 16884 16436
rect 17164 16940 17220 16996
rect 18172 19906 18228 19908
rect 18172 19854 18174 19906
rect 18174 19854 18226 19906
rect 18226 19854 18228 19906
rect 18172 19852 18228 19854
rect 17500 18396 17556 18452
rect 18508 23772 18564 23828
rect 18844 25564 18900 25620
rect 18620 21532 18676 21588
rect 18732 25340 18788 25396
rect 18508 20076 18564 20132
rect 20076 27074 20132 27076
rect 20076 27022 20078 27074
rect 20078 27022 20130 27074
rect 20130 27022 20132 27074
rect 20076 27020 20132 27022
rect 22428 31666 22484 31668
rect 22428 31614 22430 31666
rect 22430 31614 22482 31666
rect 22482 31614 22484 31666
rect 22428 31612 22484 31614
rect 21644 28418 21700 28420
rect 21644 28366 21646 28418
rect 21646 28366 21698 28418
rect 21698 28366 21700 28418
rect 21644 28364 21700 28366
rect 22764 33346 22820 33348
rect 22764 33294 22766 33346
rect 22766 33294 22818 33346
rect 22818 33294 22820 33346
rect 22764 33292 22820 33294
rect 23996 34300 24052 34356
rect 24444 34412 24500 34468
rect 23212 33628 23268 33684
rect 23548 33516 23604 33572
rect 23772 33346 23828 33348
rect 23772 33294 23774 33346
rect 23774 33294 23826 33346
rect 23826 33294 23828 33346
rect 23772 33292 23828 33294
rect 23436 33122 23492 33124
rect 23436 33070 23438 33122
rect 23438 33070 23490 33122
rect 23490 33070 23492 33122
rect 23436 33068 23492 33070
rect 24892 33404 24948 33460
rect 23100 32060 23156 32116
rect 23548 32562 23604 32564
rect 23548 32510 23550 32562
rect 23550 32510 23602 32562
rect 23602 32510 23604 32562
rect 23548 32508 23604 32510
rect 23548 32172 23604 32228
rect 24892 32508 24948 32564
rect 23772 32060 23828 32116
rect 23324 31948 23380 32004
rect 22876 31500 22932 31556
rect 22204 28476 22260 28532
rect 22092 28028 22148 28084
rect 21644 27916 21700 27972
rect 21532 27804 21588 27860
rect 19852 26796 19908 26852
rect 19404 26684 19460 26740
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19068 23826 19124 23828
rect 19068 23774 19070 23826
rect 19070 23774 19122 23826
rect 19122 23774 19124 23826
rect 19068 23772 19124 23774
rect 18844 22370 18900 22372
rect 18844 22318 18846 22370
rect 18846 22318 18898 22370
rect 18898 22318 18900 22370
rect 18844 22316 18900 22318
rect 19068 23436 19124 23492
rect 19628 26124 19684 26180
rect 21532 26962 21588 26964
rect 21532 26910 21534 26962
rect 21534 26910 21586 26962
rect 21586 26910 21588 26962
rect 21532 26908 21588 26910
rect 21644 27580 21700 27636
rect 21420 26348 21476 26404
rect 22092 27356 22148 27412
rect 19964 26124 20020 26180
rect 19740 25394 19796 25396
rect 19740 25342 19742 25394
rect 19742 25342 19794 25394
rect 19794 25342 19796 25394
rect 19740 25340 19796 25342
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20076 24780 20132 24836
rect 21420 25506 21476 25508
rect 21420 25454 21422 25506
rect 21422 25454 21474 25506
rect 21474 25454 21476 25506
rect 21420 25452 21476 25454
rect 20188 23884 20244 23940
rect 20636 24780 20692 24836
rect 19628 23772 19684 23828
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19740 23100 19796 23156
rect 19628 23042 19684 23044
rect 19628 22990 19630 23042
rect 19630 22990 19682 23042
rect 19682 22990 19684 23042
rect 19628 22988 19684 22990
rect 21532 25282 21588 25284
rect 21532 25230 21534 25282
rect 21534 25230 21586 25282
rect 21586 25230 21588 25282
rect 21532 25228 21588 25230
rect 20748 25004 20804 25060
rect 20524 23154 20580 23156
rect 20524 23102 20526 23154
rect 20526 23102 20578 23154
rect 20578 23102 20580 23154
rect 20524 23100 20580 23102
rect 20748 24556 20804 24612
rect 20636 22876 20692 22932
rect 19180 22370 19236 22372
rect 19180 22318 19182 22370
rect 19182 22318 19234 22370
rect 19234 22318 19236 22370
rect 19180 22316 19236 22318
rect 20188 22316 20244 22372
rect 19292 22092 19348 22148
rect 19068 21698 19124 21700
rect 19068 21646 19070 21698
rect 19070 21646 19122 21698
rect 19122 21646 19124 21698
rect 19068 21644 19124 21646
rect 19180 20636 19236 20692
rect 18508 19516 18564 19572
rect 18732 19180 18788 19236
rect 19180 19740 19236 19796
rect 18732 18450 18788 18452
rect 18732 18398 18734 18450
rect 18734 18398 18786 18450
rect 18786 18398 18788 18450
rect 18732 18396 18788 18398
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20300 21810 20356 21812
rect 20300 21758 20302 21810
rect 20302 21758 20354 21810
rect 20354 21758 20356 21810
rect 20300 21756 20356 21758
rect 20860 23884 20916 23940
rect 21196 23324 21252 23380
rect 20972 22876 21028 22932
rect 21084 21868 21140 21924
rect 22652 27970 22708 27972
rect 22652 27918 22654 27970
rect 22654 27918 22706 27970
rect 22706 27918 22708 27970
rect 22652 27916 22708 27918
rect 22540 27074 22596 27076
rect 22540 27022 22542 27074
rect 22542 27022 22594 27074
rect 22594 27022 22596 27074
rect 22540 27020 22596 27022
rect 22988 31218 23044 31220
rect 22988 31166 22990 31218
rect 22990 31166 23042 31218
rect 23042 31166 23044 31218
rect 22988 31164 23044 31166
rect 23548 31612 23604 31668
rect 22876 30156 22932 30212
rect 24444 31500 24500 31556
rect 24556 31612 24612 31668
rect 23996 30994 24052 30996
rect 23996 30942 23998 30994
rect 23998 30942 24050 30994
rect 24050 30942 24052 30994
rect 23996 30940 24052 30942
rect 24556 30994 24612 30996
rect 24556 30942 24558 30994
rect 24558 30942 24610 30994
rect 24610 30942 24612 30994
rect 24556 30940 24612 30942
rect 25004 32284 25060 32340
rect 24332 30210 24388 30212
rect 24332 30158 24334 30210
rect 24334 30158 24386 30210
rect 24386 30158 24388 30210
rect 24332 30156 24388 30158
rect 24668 29314 24724 29316
rect 24668 29262 24670 29314
rect 24670 29262 24722 29314
rect 24722 29262 24724 29314
rect 24668 29260 24724 29262
rect 22876 27580 22932 27636
rect 23996 28364 24052 28420
rect 25004 28812 25060 28868
rect 23996 27916 24052 27972
rect 24668 27916 24724 27972
rect 24444 27858 24500 27860
rect 24444 27806 24446 27858
rect 24446 27806 24498 27858
rect 24498 27806 24500 27858
rect 24444 27804 24500 27806
rect 23660 27580 23716 27636
rect 23660 27356 23716 27412
rect 22876 26908 22932 26964
rect 21980 26796 22036 26852
rect 21308 21756 21364 21812
rect 21980 25452 22036 25508
rect 22204 25004 22260 25060
rect 22204 24556 22260 24612
rect 21532 23100 21588 23156
rect 21868 23378 21924 23380
rect 21868 23326 21870 23378
rect 21870 23326 21922 23378
rect 21922 23326 21924 23378
rect 21868 23324 21924 23326
rect 22540 26348 22596 26404
rect 22204 23042 22260 23044
rect 22204 22990 22206 23042
rect 22206 22990 22258 23042
rect 22258 22990 22260 23042
rect 22204 22988 22260 22990
rect 22092 22146 22148 22148
rect 22092 22094 22094 22146
rect 22094 22094 22146 22146
rect 22146 22094 22148 22146
rect 22092 22092 22148 22094
rect 22092 21644 22148 21700
rect 20300 20690 20356 20692
rect 20300 20638 20302 20690
rect 20302 20638 20354 20690
rect 20354 20638 20356 20690
rect 20300 20636 20356 20638
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20524 20578 20580 20580
rect 20524 20526 20526 20578
rect 20526 20526 20578 20578
rect 20578 20526 20580 20578
rect 20524 20524 20580 20526
rect 21420 20578 21476 20580
rect 21420 20526 21422 20578
rect 21422 20526 21474 20578
rect 21474 20526 21476 20578
rect 21420 20524 21476 20526
rect 20188 20076 20244 20132
rect 21084 20412 21140 20468
rect 19852 19234 19908 19236
rect 19852 19182 19854 19234
rect 19854 19182 19906 19234
rect 19906 19182 19908 19234
rect 19852 19180 19908 19182
rect 20300 19794 20356 19796
rect 20300 19742 20302 19794
rect 20302 19742 20354 19794
rect 20354 19742 20356 19794
rect 20300 19740 20356 19742
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 17612 16940 17668 16996
rect 17276 16604 17332 16660
rect 17388 16716 17444 16772
rect 15596 13804 15652 13860
rect 18060 16044 18116 16100
rect 16716 15260 16772 15316
rect 17724 15426 17780 15428
rect 17724 15374 17726 15426
rect 17726 15374 17778 15426
rect 17778 15374 17780 15426
rect 17724 15372 17780 15374
rect 16828 14700 16884 14756
rect 15820 13746 15876 13748
rect 15820 13694 15822 13746
rect 15822 13694 15874 13746
rect 15874 13694 15876 13746
rect 15820 13692 15876 13694
rect 15596 12348 15652 12404
rect 19068 13692 19124 13748
rect 18956 13356 19012 13412
rect 16044 12348 16100 12404
rect 14700 10668 14756 10724
rect 15260 10444 15316 10500
rect 14252 9548 14308 9604
rect 15372 10668 15428 10724
rect 15708 10332 15764 10388
rect 15708 9772 15764 9828
rect 20188 18172 20244 18228
rect 20748 18396 20804 18452
rect 19292 12348 19348 12404
rect 19404 18060 19460 18116
rect 16716 10610 16772 10612
rect 16716 10558 16718 10610
rect 16718 10558 16770 10610
rect 16770 10558 16772 10610
rect 16716 10556 16772 10558
rect 17500 10610 17556 10612
rect 17500 10558 17502 10610
rect 17502 10558 17554 10610
rect 17554 10558 17556 10610
rect 17500 10556 17556 10558
rect 17724 10444 17780 10500
rect 16044 10220 16100 10276
rect 17164 10332 17220 10388
rect 12124 7756 12180 7812
rect 14140 7756 14196 7812
rect 14700 7698 14756 7700
rect 14700 7646 14702 7698
rect 14702 7646 14754 7698
rect 14754 7646 14756 7698
rect 14700 7644 14756 7646
rect 9324 6690 9380 6692
rect 9324 6638 9326 6690
rect 9326 6638 9378 6690
rect 9378 6638 9380 6690
rect 9324 6636 9380 6638
rect 11788 6636 11844 6692
rect 12684 6690 12740 6692
rect 12684 6638 12686 6690
rect 12686 6638 12738 6690
rect 12738 6638 12740 6690
rect 12684 6636 12740 6638
rect 15260 6636 15316 6692
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 16716 7474 16772 7476
rect 16716 7422 16718 7474
rect 16718 7422 16770 7474
rect 16770 7422 16772 7474
rect 16716 7420 16772 7422
rect 18620 10610 18676 10612
rect 18620 10558 18622 10610
rect 18622 10558 18674 10610
rect 18674 10558 18676 10610
rect 18620 10556 18676 10558
rect 17836 10386 17892 10388
rect 17836 10334 17838 10386
rect 17838 10334 17890 10386
rect 17890 10334 17892 10386
rect 17836 10332 17892 10334
rect 17724 9826 17780 9828
rect 17724 9774 17726 9826
rect 17726 9774 17778 9826
rect 17778 9774 17780 9826
rect 17724 9772 17780 9774
rect 17500 7474 17556 7476
rect 17500 7422 17502 7474
rect 17502 7422 17554 7474
rect 17554 7422 17556 7474
rect 17500 7420 17556 7422
rect 19292 9996 19348 10052
rect 18508 9100 18564 9156
rect 18396 8930 18452 8932
rect 18396 8878 18398 8930
rect 18398 8878 18450 8930
rect 18450 8878 18452 8930
rect 18396 8876 18452 8878
rect 18060 7756 18116 7812
rect 19292 8876 19348 8932
rect 19628 17612 19684 17668
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16380 19684 16436
rect 19516 16322 19572 16324
rect 19516 16270 19518 16322
rect 19518 16270 19570 16322
rect 19570 16270 19572 16322
rect 19516 16268 19572 16270
rect 20300 16268 20356 16324
rect 21420 20130 21476 20132
rect 21420 20078 21422 20130
rect 21422 20078 21474 20130
rect 21474 20078 21476 20130
rect 21420 20076 21476 20078
rect 21308 19964 21364 20020
rect 21644 20130 21700 20132
rect 21644 20078 21646 20130
rect 21646 20078 21698 20130
rect 21698 20078 21700 20130
rect 21644 20076 21700 20078
rect 22540 24556 22596 24612
rect 22764 23996 22820 24052
rect 22764 23826 22820 23828
rect 22764 23774 22766 23826
rect 22766 23774 22818 23826
rect 22818 23774 22820 23826
rect 22764 23772 22820 23774
rect 23772 27074 23828 27076
rect 23772 27022 23774 27074
rect 23774 27022 23826 27074
rect 23826 27022 23828 27074
rect 23772 27020 23828 27022
rect 24556 26572 24612 26628
rect 24892 27020 24948 27076
rect 26348 41132 26404 41188
rect 26908 41916 26964 41972
rect 26796 41410 26852 41412
rect 26796 41358 26798 41410
rect 26798 41358 26850 41410
rect 26850 41358 26852 41410
rect 26796 41356 26852 41358
rect 26572 40572 26628 40628
rect 27692 41970 27748 41972
rect 27692 41918 27694 41970
rect 27694 41918 27746 41970
rect 27746 41918 27748 41970
rect 27692 41916 27748 41918
rect 26348 40402 26404 40404
rect 26348 40350 26350 40402
rect 26350 40350 26402 40402
rect 26402 40350 26404 40402
rect 26348 40348 26404 40350
rect 26236 40124 26292 40180
rect 26796 40124 26852 40180
rect 26348 39730 26404 39732
rect 26348 39678 26350 39730
rect 26350 39678 26402 39730
rect 26402 39678 26404 39730
rect 26348 39676 26404 39678
rect 27580 40796 27636 40852
rect 27244 40684 27300 40740
rect 27020 39842 27076 39844
rect 27020 39790 27022 39842
rect 27022 39790 27074 39842
rect 27074 39790 27076 39842
rect 27020 39788 27076 39790
rect 26908 39618 26964 39620
rect 26908 39566 26910 39618
rect 26910 39566 26962 39618
rect 26962 39566 26964 39618
rect 26908 39564 26964 39566
rect 26908 39116 26964 39172
rect 28476 43538 28532 43540
rect 28476 43486 28478 43538
rect 28478 43486 28530 43538
rect 28530 43486 28532 43538
rect 28476 43484 28532 43486
rect 28364 43314 28420 43316
rect 28364 43262 28366 43314
rect 28366 43262 28418 43314
rect 28418 43262 28420 43314
rect 28364 43260 28420 43262
rect 28364 42028 28420 42084
rect 28588 41692 28644 41748
rect 28588 41244 28644 41300
rect 28476 41074 28532 41076
rect 28476 41022 28478 41074
rect 28478 41022 28530 41074
rect 28530 41022 28532 41074
rect 28476 41020 28532 41022
rect 28028 40684 28084 40740
rect 28364 40962 28420 40964
rect 28364 40910 28366 40962
rect 28366 40910 28418 40962
rect 28418 40910 28420 40962
rect 28364 40908 28420 40910
rect 27916 40514 27972 40516
rect 27916 40462 27918 40514
rect 27918 40462 27970 40514
rect 27970 40462 27972 40514
rect 27916 40460 27972 40462
rect 27356 40236 27412 40292
rect 27468 40348 27524 40404
rect 27580 39618 27636 39620
rect 27580 39566 27582 39618
rect 27582 39566 27634 39618
rect 27634 39566 27636 39618
rect 27580 39564 27636 39566
rect 29820 46172 29876 46228
rect 29708 45724 29764 45780
rect 29596 44828 29652 44884
rect 28364 40626 28420 40628
rect 28364 40574 28366 40626
rect 28366 40574 28418 40626
rect 28418 40574 28420 40626
rect 28364 40572 28420 40574
rect 28812 44604 28868 44660
rect 29596 44604 29652 44660
rect 29148 44098 29204 44100
rect 29148 44046 29150 44098
rect 29150 44046 29202 44098
rect 29202 44046 29204 44098
rect 29148 44044 29204 44046
rect 29260 43932 29316 43988
rect 29036 42028 29092 42084
rect 29148 43484 29204 43540
rect 29596 43932 29652 43988
rect 29708 43708 29764 43764
rect 30716 46786 30772 46788
rect 30716 46734 30718 46786
rect 30718 46734 30770 46786
rect 30770 46734 30772 46786
rect 30716 46732 30772 46734
rect 30828 46956 30884 47012
rect 30044 45890 30100 45892
rect 30044 45838 30046 45890
rect 30046 45838 30098 45890
rect 30098 45838 30100 45890
rect 30044 45836 30100 45838
rect 30044 44940 30100 44996
rect 30604 45836 30660 45892
rect 32060 48300 32116 48356
rect 33292 48914 33348 48916
rect 33292 48862 33294 48914
rect 33294 48862 33346 48914
rect 33346 48862 33348 48914
rect 33292 48860 33348 48862
rect 33740 48412 33796 48468
rect 32396 47570 32452 47572
rect 32396 47518 32398 47570
rect 32398 47518 32450 47570
rect 32450 47518 32452 47570
rect 32396 47516 32452 47518
rect 33404 47516 33460 47572
rect 30940 46844 30996 46900
rect 31612 46620 31668 46676
rect 30828 45724 30884 45780
rect 30828 45052 30884 45108
rect 30380 44828 30436 44884
rect 30716 44828 30772 44884
rect 30156 44044 30212 44100
rect 29932 43932 29988 43988
rect 30156 43708 30212 43764
rect 32060 46786 32116 46788
rect 32060 46734 32062 46786
rect 32062 46734 32114 46786
rect 32114 46734 32116 46786
rect 32060 46732 32116 46734
rect 32172 46674 32228 46676
rect 32172 46622 32174 46674
rect 32174 46622 32226 46674
rect 32226 46622 32228 46674
rect 32172 46620 32228 46622
rect 33068 46674 33124 46676
rect 33068 46622 33070 46674
rect 33070 46622 33122 46674
rect 33122 46622 33124 46674
rect 33068 46620 33124 46622
rect 31724 46508 31780 46564
rect 31612 45164 31668 45220
rect 31052 44828 31108 44884
rect 30828 44380 30884 44436
rect 30940 44268 30996 44324
rect 30604 43708 30660 43764
rect 29820 43036 29876 43092
rect 29932 42700 29988 42756
rect 28476 40178 28532 40180
rect 28476 40126 28478 40178
rect 28478 40126 28530 40178
rect 28530 40126 28532 40178
rect 28476 40124 28532 40126
rect 28252 39788 28308 39844
rect 28364 39116 28420 39172
rect 29148 41468 29204 41524
rect 29372 41916 29428 41972
rect 29372 41356 29428 41412
rect 29148 41186 29204 41188
rect 29148 41134 29150 41186
rect 29150 41134 29202 41186
rect 29202 41134 29204 41186
rect 29148 41132 29204 41134
rect 29596 41746 29652 41748
rect 29596 41694 29598 41746
rect 29598 41694 29650 41746
rect 29650 41694 29652 41746
rect 29596 41692 29652 41694
rect 31612 44380 31668 44436
rect 31388 44268 31444 44324
rect 31276 43372 31332 43428
rect 30268 41468 30324 41524
rect 29372 40962 29428 40964
rect 29372 40910 29374 40962
rect 29374 40910 29426 40962
rect 29426 40910 29428 40962
rect 29372 40908 29428 40910
rect 29820 41186 29876 41188
rect 29820 41134 29822 41186
rect 29822 41134 29874 41186
rect 29874 41134 29876 41186
rect 29820 41132 29876 41134
rect 29036 40572 29092 40628
rect 29820 40626 29876 40628
rect 29820 40574 29822 40626
rect 29822 40574 29874 40626
rect 29874 40574 29876 40626
rect 29820 40572 29876 40574
rect 28700 40402 28756 40404
rect 28700 40350 28702 40402
rect 28702 40350 28754 40402
rect 28754 40350 28756 40402
rect 28700 40348 28756 40350
rect 25900 38556 25956 38612
rect 26124 38610 26180 38612
rect 26124 38558 26126 38610
rect 26126 38558 26178 38610
rect 26178 38558 26180 38610
rect 26124 38556 26180 38558
rect 27468 38556 27524 38612
rect 27692 38108 27748 38164
rect 26796 37436 26852 37492
rect 27132 37324 27188 37380
rect 25452 35922 25508 35924
rect 25452 35870 25454 35922
rect 25454 35870 25506 35922
rect 25506 35870 25508 35922
rect 25452 35868 25508 35870
rect 27132 37154 27188 37156
rect 27132 37102 27134 37154
rect 27134 37102 27186 37154
rect 27186 37102 27188 37154
rect 27132 37100 27188 37102
rect 26236 36316 26292 36372
rect 25788 35810 25844 35812
rect 25788 35758 25790 35810
rect 25790 35758 25842 35810
rect 25842 35758 25844 35810
rect 25788 35756 25844 35758
rect 27580 36876 27636 36932
rect 28252 37154 28308 37156
rect 28252 37102 28254 37154
rect 28254 37102 28306 37154
rect 28306 37102 28308 37154
rect 28252 37100 28308 37102
rect 28252 36876 28308 36932
rect 28588 36876 28644 36932
rect 26460 35810 26516 35812
rect 26460 35758 26462 35810
rect 26462 35758 26514 35810
rect 26514 35758 26516 35810
rect 26460 35756 26516 35758
rect 27244 35698 27300 35700
rect 27244 35646 27246 35698
rect 27246 35646 27298 35698
rect 27298 35646 27300 35698
rect 27244 35644 27300 35646
rect 25900 34860 25956 34916
rect 25452 34412 25508 34468
rect 25564 33516 25620 33572
rect 25676 32450 25732 32452
rect 25676 32398 25678 32450
rect 25678 32398 25730 32450
rect 25730 32398 25732 32450
rect 25676 32396 25732 32398
rect 25452 31500 25508 31556
rect 25228 31388 25284 31444
rect 25340 30156 25396 30212
rect 26012 33068 26068 33124
rect 26348 32732 26404 32788
rect 26124 32562 26180 32564
rect 26124 32510 26126 32562
rect 26126 32510 26178 32562
rect 26178 32510 26180 32562
rect 26124 32508 26180 32510
rect 26348 31666 26404 31668
rect 26348 31614 26350 31666
rect 26350 31614 26402 31666
rect 26402 31614 26404 31666
rect 26348 31612 26404 31614
rect 26796 34300 26852 34356
rect 28140 34914 28196 34916
rect 28140 34862 28142 34914
rect 28142 34862 28194 34914
rect 28194 34862 28196 34914
rect 28140 34860 28196 34862
rect 28812 38780 28868 38836
rect 29148 39116 29204 39172
rect 29820 37938 29876 37940
rect 29820 37886 29822 37938
rect 29822 37886 29874 37938
rect 29874 37886 29876 37938
rect 29820 37884 29876 37886
rect 30604 41132 30660 41188
rect 31164 42364 31220 42420
rect 30268 40572 30324 40628
rect 31388 42140 31444 42196
rect 31612 44210 31668 44212
rect 31612 44158 31614 44210
rect 31614 44158 31666 44210
rect 31666 44158 31668 44210
rect 31612 44156 31668 44158
rect 34524 48300 34580 48356
rect 33068 45890 33124 45892
rect 33068 45838 33070 45890
rect 33070 45838 33122 45890
rect 33122 45838 33124 45890
rect 33068 45836 33124 45838
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 36316 51100 36372 51156
rect 35980 50764 36036 50820
rect 35868 50482 35924 50484
rect 35868 50430 35870 50482
rect 35870 50430 35922 50482
rect 35922 50430 35924 50482
rect 35868 50428 35924 50430
rect 36540 50876 36596 50932
rect 36092 50652 36148 50708
rect 36428 50540 36484 50596
rect 37100 51212 37156 51268
rect 37100 50988 37156 51044
rect 35644 49810 35700 49812
rect 35644 49758 35646 49810
rect 35646 49758 35698 49810
rect 35698 49758 35700 49810
rect 35644 49756 35700 49758
rect 36988 50316 37044 50372
rect 37660 50428 37716 50484
rect 36540 50092 36596 50148
rect 36316 50034 36372 50036
rect 36316 49982 36318 50034
rect 36318 49982 36370 50034
rect 36370 49982 36372 50034
rect 36316 49980 36372 49982
rect 37212 49980 37268 50036
rect 37100 49922 37156 49924
rect 37100 49870 37102 49922
rect 37102 49870 37154 49922
rect 37154 49870 37156 49922
rect 37100 49868 37156 49870
rect 36876 49644 36932 49700
rect 37436 50204 37492 50260
rect 38108 51602 38164 51604
rect 38108 51550 38110 51602
rect 38110 51550 38162 51602
rect 38162 51550 38164 51602
rect 38108 51548 38164 51550
rect 37884 50428 37940 50484
rect 37996 51378 38052 51380
rect 37996 51326 37998 51378
rect 37998 51326 38050 51378
rect 38050 51326 38052 51378
rect 37996 51324 38052 51326
rect 38108 51154 38164 51156
rect 38108 51102 38110 51154
rect 38110 51102 38162 51154
rect 38162 51102 38164 51154
rect 38108 51100 38164 51102
rect 38332 52332 38388 52388
rect 38444 53228 38500 53284
rect 38668 53058 38724 53060
rect 38668 53006 38670 53058
rect 38670 53006 38722 53058
rect 38722 53006 38724 53058
rect 38668 53004 38724 53006
rect 38780 52946 38836 52948
rect 38780 52894 38782 52946
rect 38782 52894 38834 52946
rect 38834 52894 38836 52946
rect 38780 52892 38836 52894
rect 38668 52780 38724 52836
rect 38780 52668 38836 52724
rect 38444 51938 38500 51940
rect 38444 51886 38446 51938
rect 38446 51886 38498 51938
rect 38498 51886 38500 51938
rect 38444 51884 38500 51886
rect 38444 51212 38500 51268
rect 38332 50652 38388 50708
rect 38444 50092 38500 50148
rect 37996 49922 38052 49924
rect 37996 49870 37998 49922
rect 37998 49870 38050 49922
rect 38050 49870 38052 49922
rect 37996 49868 38052 49870
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 36092 49026 36148 49028
rect 36092 48974 36094 49026
rect 36094 48974 36146 49026
rect 36146 48974 36148 49026
rect 36092 48972 36148 48974
rect 39116 53004 39172 53060
rect 40124 53452 40180 53508
rect 39676 53170 39732 53172
rect 39676 53118 39678 53170
rect 39678 53118 39730 53170
rect 39730 53118 39732 53170
rect 39676 53116 39732 53118
rect 39116 52444 39172 52500
rect 38892 52162 38948 52164
rect 38892 52110 38894 52162
rect 38894 52110 38946 52162
rect 38946 52110 38948 52162
rect 38892 52108 38948 52110
rect 39452 52332 39508 52388
rect 39564 52274 39620 52276
rect 39564 52222 39566 52274
rect 39566 52222 39618 52274
rect 39618 52222 39620 52274
rect 39564 52220 39620 52222
rect 39004 51884 39060 51940
rect 39340 51996 39396 52052
rect 39116 51548 39172 51604
rect 38668 51324 38724 51380
rect 38892 51212 38948 51268
rect 38668 50988 38724 51044
rect 38892 50652 38948 50708
rect 38780 50428 38836 50484
rect 39004 50594 39060 50596
rect 39004 50542 39006 50594
rect 39006 50542 39058 50594
rect 39058 50542 39060 50594
rect 39004 50540 39060 50542
rect 39228 51490 39284 51492
rect 39228 51438 39230 51490
rect 39230 51438 39282 51490
rect 39282 51438 39284 51490
rect 39228 51436 39284 51438
rect 39676 51996 39732 52052
rect 39340 51324 39396 51380
rect 39564 51436 39620 51492
rect 39452 51154 39508 51156
rect 39452 51102 39454 51154
rect 39454 51102 39506 51154
rect 39506 51102 39508 51154
rect 39452 51100 39508 51102
rect 39228 50988 39284 51044
rect 39564 50988 39620 51044
rect 39340 50764 39396 50820
rect 39228 49980 39284 50036
rect 39116 49644 39172 49700
rect 37436 48972 37492 49028
rect 38668 48860 38724 48916
rect 39452 50370 39508 50372
rect 39452 50318 39454 50370
rect 39454 50318 39506 50370
rect 39506 50318 39508 50370
rect 39452 50316 39508 50318
rect 39452 49196 39508 49252
rect 39004 48802 39060 48804
rect 39004 48750 39006 48802
rect 39006 48750 39058 48802
rect 39058 48750 39060 48802
rect 39004 48748 39060 48750
rect 39228 48860 39284 48916
rect 39676 50428 39732 50484
rect 39676 49644 39732 49700
rect 39900 51548 39956 51604
rect 43036 55916 43092 55972
rect 43596 57036 43652 57092
rect 44044 56306 44100 56308
rect 44044 56254 44046 56306
rect 44046 56254 44098 56306
rect 44098 56254 44100 56306
rect 44044 56252 44100 56254
rect 44492 55970 44548 55972
rect 44492 55918 44494 55970
rect 44494 55918 44546 55970
rect 44546 55918 44548 55970
rect 44492 55916 44548 55918
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 42588 55186 42644 55188
rect 42588 55134 42590 55186
rect 42590 55134 42642 55186
rect 42642 55134 42644 55186
rect 42588 55132 42644 55134
rect 42700 55020 42756 55076
rect 43596 55074 43652 55076
rect 43596 55022 43598 55074
rect 43598 55022 43650 55074
rect 43650 55022 43652 55074
rect 43596 55020 43652 55022
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 44604 54626 44660 54628
rect 44604 54574 44606 54626
rect 44606 54574 44658 54626
rect 44658 54574 44660 54626
rect 44604 54572 44660 54574
rect 45836 54402 45892 54404
rect 45836 54350 45838 54402
rect 45838 54350 45890 54402
rect 45890 54350 45892 54402
rect 45836 54348 45892 54350
rect 42140 53676 42196 53732
rect 42028 53228 42084 53284
rect 40236 52946 40292 52948
rect 40236 52894 40238 52946
rect 40238 52894 40290 52946
rect 40290 52894 40292 52946
rect 40236 52892 40292 52894
rect 40236 52332 40292 52388
rect 40348 52108 40404 52164
rect 40684 52444 40740 52500
rect 41020 52332 41076 52388
rect 41244 53004 41300 53060
rect 40124 51772 40180 51828
rect 40796 51884 40852 51940
rect 40012 51436 40068 51492
rect 40124 51324 40180 51380
rect 39900 50316 39956 50372
rect 39900 49980 39956 50036
rect 40124 50764 40180 50820
rect 40236 50988 40292 51044
rect 40124 50482 40180 50484
rect 40124 50430 40126 50482
rect 40126 50430 40178 50482
rect 40178 50430 40180 50482
rect 40124 50428 40180 50430
rect 40012 49922 40068 49924
rect 40012 49870 40014 49922
rect 40014 49870 40066 49922
rect 40066 49870 40068 49922
rect 40012 49868 40068 49870
rect 40908 51548 40964 51604
rect 41020 51772 41076 51828
rect 41916 53058 41972 53060
rect 41916 53006 41918 53058
rect 41918 53006 41970 53058
rect 41970 53006 41972 53058
rect 41916 53004 41972 53006
rect 41692 52050 41748 52052
rect 41692 51998 41694 52050
rect 41694 51998 41746 52050
rect 41746 51998 41748 52050
rect 41692 51996 41748 51998
rect 40460 50428 40516 50484
rect 41356 51548 41412 51604
rect 42588 53058 42644 53060
rect 42588 53006 42590 53058
rect 42590 53006 42642 53058
rect 42642 53006 42644 53058
rect 42588 53004 42644 53006
rect 42252 52892 42308 52948
rect 43372 52780 43428 52836
rect 44828 53730 44884 53732
rect 44828 53678 44830 53730
rect 44830 53678 44882 53730
rect 44882 53678 44884 53730
rect 44828 53676 44884 53678
rect 48076 54402 48132 54404
rect 48076 54350 48078 54402
rect 48078 54350 48130 54402
rect 48130 54350 48132 54402
rect 48076 54348 48132 54350
rect 45276 53676 45332 53732
rect 43596 52892 43652 52948
rect 43484 52220 43540 52276
rect 42364 51996 42420 52052
rect 42028 51436 42084 51492
rect 41132 50876 41188 50932
rect 40236 50316 40292 50372
rect 40012 49196 40068 49252
rect 40684 49868 40740 49924
rect 40908 49698 40964 49700
rect 40908 49646 40910 49698
rect 40910 49646 40962 49698
rect 40962 49646 40964 49698
rect 40908 49644 40964 49646
rect 41916 50540 41972 50596
rect 42140 50652 42196 50708
rect 41580 50482 41636 50484
rect 41580 50430 41582 50482
rect 41582 50430 41634 50482
rect 41634 50430 41636 50482
rect 41580 50428 41636 50430
rect 42028 50428 42084 50484
rect 41356 49868 41412 49924
rect 42812 52050 42868 52052
rect 42812 51998 42814 52050
rect 42814 51998 42866 52050
rect 42866 51998 42868 52050
rect 42812 51996 42868 51998
rect 43372 51548 43428 51604
rect 43036 51324 43092 51380
rect 42364 50988 42420 51044
rect 42252 50428 42308 50484
rect 42476 50764 42532 50820
rect 44044 52780 44100 52836
rect 43708 51548 43764 51604
rect 43932 51548 43988 51604
rect 43820 51154 43876 51156
rect 43820 51102 43822 51154
rect 43822 51102 43874 51154
rect 43874 51102 43876 51154
rect 43820 51100 43876 51102
rect 43596 50876 43652 50932
rect 43708 50988 43764 51044
rect 42476 50204 42532 50260
rect 41468 49810 41524 49812
rect 41468 49758 41470 49810
rect 41470 49758 41522 49810
rect 41522 49758 41524 49810
rect 41468 49756 41524 49758
rect 42476 49868 42532 49924
rect 43372 50316 43428 50372
rect 43596 50092 43652 50148
rect 43372 49980 43428 50036
rect 43148 49810 43204 49812
rect 43148 49758 43150 49810
rect 43150 49758 43202 49810
rect 43202 49758 43204 49810
rect 43148 49756 43204 49758
rect 42924 49250 42980 49252
rect 42924 49198 42926 49250
rect 42926 49198 42978 49250
rect 42978 49198 42980 49250
rect 42924 49196 42980 49198
rect 43596 49420 43652 49476
rect 43260 49026 43316 49028
rect 43260 48974 43262 49026
rect 43262 48974 43314 49026
rect 43314 48974 43316 49026
rect 43260 48972 43316 48974
rect 41804 48914 41860 48916
rect 41804 48862 41806 48914
rect 41806 48862 41858 48914
rect 41858 48862 41860 48914
rect 41804 48860 41860 48862
rect 42028 48802 42084 48804
rect 42028 48750 42030 48802
rect 42030 48750 42082 48802
rect 42082 48750 42084 48802
rect 42028 48748 42084 48750
rect 41356 48300 41412 48356
rect 36316 48130 36372 48132
rect 36316 48078 36318 48130
rect 36318 48078 36370 48130
rect 36370 48078 36372 48130
rect 36316 48076 36372 48078
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 34412 47346 34468 47348
rect 34412 47294 34414 47346
rect 34414 47294 34466 47346
rect 34466 47294 34468 47346
rect 34412 47292 34468 47294
rect 33852 45836 33908 45892
rect 31948 45218 32004 45220
rect 31948 45166 31950 45218
rect 31950 45166 32002 45218
rect 32002 45166 32004 45218
rect 31948 45164 32004 45166
rect 32284 45106 32340 45108
rect 32284 45054 32286 45106
rect 32286 45054 32338 45106
rect 32338 45054 32340 45106
rect 32284 45052 32340 45054
rect 32060 43820 32116 43876
rect 33516 44828 33572 44884
rect 32396 44492 32452 44548
rect 32284 44210 32340 44212
rect 32284 44158 32286 44210
rect 32286 44158 32338 44210
rect 32338 44158 32340 44210
rect 32284 44156 32340 44158
rect 32396 42812 32452 42868
rect 33740 44604 33796 44660
rect 33628 44492 33684 44548
rect 33628 44210 33684 44212
rect 33628 44158 33630 44210
rect 33630 44158 33682 44210
rect 33682 44158 33684 44210
rect 33628 44156 33684 44158
rect 33964 45218 34020 45220
rect 33964 45166 33966 45218
rect 33966 45166 34018 45218
rect 34018 45166 34020 45218
rect 33964 45164 34020 45166
rect 32172 42364 32228 42420
rect 31724 41970 31780 41972
rect 31724 41918 31726 41970
rect 31726 41918 31778 41970
rect 31778 41918 31780 41970
rect 31724 41916 31780 41918
rect 31948 42194 32004 42196
rect 31948 42142 31950 42194
rect 31950 42142 32002 42194
rect 32002 42142 32004 42194
rect 31948 42140 32004 42142
rect 33404 43484 33460 43540
rect 32620 42140 32676 42196
rect 33292 42082 33348 42084
rect 33292 42030 33294 42082
rect 33294 42030 33346 42082
rect 33346 42030 33348 42082
rect 33292 42028 33348 42030
rect 32508 41916 32564 41972
rect 31836 40908 31892 40964
rect 31612 40572 31668 40628
rect 30492 39900 30548 39956
rect 30492 39004 30548 39060
rect 31724 40796 31780 40852
rect 31724 39676 31780 39732
rect 31948 39564 32004 39620
rect 30156 37996 30212 38052
rect 30156 36370 30212 36372
rect 30156 36318 30158 36370
rect 30158 36318 30210 36370
rect 30210 36318 30212 36370
rect 30156 36316 30212 36318
rect 30380 37938 30436 37940
rect 30380 37886 30382 37938
rect 30382 37886 30434 37938
rect 30434 37886 30436 37938
rect 30380 37884 30436 37886
rect 30828 37548 30884 37604
rect 31276 37884 31332 37940
rect 30828 36876 30884 36932
rect 30268 35308 30324 35364
rect 29708 35084 29764 35140
rect 27580 34354 27636 34356
rect 27580 34302 27582 34354
rect 27582 34302 27634 34354
rect 27634 34302 27636 34354
rect 27580 34300 27636 34302
rect 28588 34300 28644 34356
rect 30156 34690 30212 34692
rect 30156 34638 30158 34690
rect 30158 34638 30210 34690
rect 30210 34638 30212 34690
rect 30156 34636 30212 34638
rect 27132 33740 27188 33796
rect 28700 33516 28756 33572
rect 30044 33516 30100 33572
rect 26684 33458 26740 33460
rect 26684 33406 26686 33458
rect 26686 33406 26738 33458
rect 26738 33406 26740 33458
rect 26684 33404 26740 33406
rect 27020 32396 27076 32452
rect 27244 32732 27300 32788
rect 27468 32508 27524 32564
rect 27804 33122 27860 33124
rect 27804 33070 27806 33122
rect 27806 33070 27858 33122
rect 27858 33070 27860 33122
rect 27804 33068 27860 33070
rect 28812 33068 28868 33124
rect 27580 32844 27636 32900
rect 26572 31612 26628 31668
rect 25900 29820 25956 29876
rect 25452 28588 25508 28644
rect 25340 27970 25396 27972
rect 25340 27918 25342 27970
rect 25342 27918 25394 27970
rect 25394 27918 25396 27970
rect 25340 27916 25396 27918
rect 25452 27804 25508 27860
rect 25452 26908 25508 26964
rect 29932 32284 29988 32340
rect 27804 31836 27860 31892
rect 28364 31890 28420 31892
rect 28364 31838 28366 31890
rect 28366 31838 28418 31890
rect 28418 31838 28420 31890
rect 28364 31836 28420 31838
rect 25564 27132 25620 27188
rect 23324 26178 23380 26180
rect 23324 26126 23326 26178
rect 23326 26126 23378 26178
rect 23378 26126 23380 26178
rect 23324 26124 23380 26126
rect 24108 26124 24164 26180
rect 23100 25506 23156 25508
rect 23100 25454 23102 25506
rect 23102 25454 23154 25506
rect 23154 25454 23156 25506
rect 23100 25452 23156 25454
rect 23772 25340 23828 25396
rect 23660 25116 23716 25172
rect 22988 25004 23044 25060
rect 23436 25004 23492 25060
rect 23436 23996 23492 24052
rect 23212 23938 23268 23940
rect 23212 23886 23214 23938
rect 23214 23886 23266 23938
rect 23266 23886 23268 23938
rect 23212 23884 23268 23886
rect 23100 23436 23156 23492
rect 22316 21698 22372 21700
rect 22316 21646 22318 21698
rect 22318 21646 22370 21698
rect 22370 21646 22372 21698
rect 22316 21644 22372 21646
rect 22204 20524 22260 20580
rect 21420 19852 21476 19908
rect 21308 19180 21364 19236
rect 21084 16156 21140 16212
rect 20300 16098 20356 16100
rect 20300 16046 20302 16098
rect 20302 16046 20354 16098
rect 20354 16046 20356 16098
rect 20300 16044 20356 16046
rect 19516 15932 19572 15988
rect 20076 15986 20132 15988
rect 20076 15934 20078 15986
rect 20078 15934 20130 15986
rect 20130 15934 20132 15986
rect 20076 15932 20132 15934
rect 20188 15820 20244 15876
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 21196 16044 21252 16100
rect 21644 19010 21700 19012
rect 21644 18958 21646 19010
rect 21646 18958 21698 19010
rect 21698 18958 21700 19010
rect 21644 18956 21700 18958
rect 21644 18172 21700 18228
rect 22540 22594 22596 22596
rect 22540 22542 22542 22594
rect 22542 22542 22594 22594
rect 22594 22542 22596 22594
rect 22540 22540 22596 22542
rect 22428 20130 22484 20132
rect 22428 20078 22430 20130
rect 22430 20078 22482 20130
rect 22482 20078 22484 20130
rect 22428 20076 22484 20078
rect 22764 20524 22820 20580
rect 22988 20802 23044 20804
rect 22988 20750 22990 20802
rect 22990 20750 23042 20802
rect 23042 20750 23044 20802
rect 22988 20748 23044 20750
rect 23324 22316 23380 22372
rect 23436 21756 23492 21812
rect 23100 20188 23156 20244
rect 22876 19740 22932 19796
rect 23884 25004 23940 25060
rect 24108 25228 24164 25284
rect 24220 25564 24276 25620
rect 23996 24892 24052 24948
rect 23996 24556 24052 24612
rect 24332 25452 24388 25508
rect 24444 26124 24500 26180
rect 26460 27132 26516 27188
rect 26796 28642 26852 28644
rect 26796 28590 26798 28642
rect 26798 28590 26850 28642
rect 26850 28590 26852 28642
rect 26796 28588 26852 28590
rect 28252 30210 28308 30212
rect 28252 30158 28254 30210
rect 28254 30158 28306 30210
rect 28306 30158 28308 30210
rect 28252 30156 28308 30158
rect 27804 29372 27860 29428
rect 27580 28866 27636 28868
rect 27580 28814 27582 28866
rect 27582 28814 27634 28866
rect 27634 28814 27636 28866
rect 27580 28812 27636 28814
rect 29596 29932 29652 29988
rect 29820 30828 29876 30884
rect 30716 36204 30772 36260
rect 30716 35756 30772 35812
rect 30492 34636 30548 34692
rect 31724 39452 31780 39508
rect 31612 39058 31668 39060
rect 31612 39006 31614 39058
rect 31614 39006 31666 39058
rect 31666 39006 31668 39058
rect 31612 39004 31668 39006
rect 33516 42028 33572 42084
rect 33068 40012 33124 40068
rect 32060 39004 32116 39060
rect 32172 38834 32228 38836
rect 32172 38782 32174 38834
rect 32174 38782 32226 38834
rect 32226 38782 32228 38834
rect 32172 38780 32228 38782
rect 33180 39058 33236 39060
rect 33180 39006 33182 39058
rect 33182 39006 33234 39058
rect 33234 39006 33236 39058
rect 33180 39004 33236 39006
rect 33292 38668 33348 38724
rect 31500 37660 31556 37716
rect 31612 37996 31668 38052
rect 31500 37490 31556 37492
rect 31500 37438 31502 37490
rect 31502 37438 31554 37490
rect 31554 37438 31556 37490
rect 31500 37436 31556 37438
rect 31276 37212 31332 37268
rect 31500 36706 31556 36708
rect 31500 36654 31502 36706
rect 31502 36654 31554 36706
rect 31554 36654 31556 36706
rect 31500 36652 31556 36654
rect 31164 36370 31220 36372
rect 31164 36318 31166 36370
rect 31166 36318 31218 36370
rect 31218 36318 31220 36370
rect 31164 36316 31220 36318
rect 31276 36204 31332 36260
rect 33068 37660 33124 37716
rect 31948 37266 32004 37268
rect 31948 37214 31950 37266
rect 31950 37214 32002 37266
rect 32002 37214 32004 37266
rect 31948 37212 32004 37214
rect 32172 36428 32228 36484
rect 31836 36258 31892 36260
rect 31836 36206 31838 36258
rect 31838 36206 31890 36258
rect 31890 36206 31892 36258
rect 31836 36204 31892 36206
rect 30940 35308 30996 35364
rect 31388 35698 31444 35700
rect 31388 35646 31390 35698
rect 31390 35646 31442 35698
rect 31442 35646 31444 35698
rect 31388 35644 31444 35646
rect 31052 34636 31108 34692
rect 31052 33516 31108 33572
rect 31948 33516 32004 33572
rect 30828 32674 30884 32676
rect 30828 32622 30830 32674
rect 30830 32622 30882 32674
rect 30882 32622 30884 32674
rect 30828 32620 30884 32622
rect 30828 31836 30884 31892
rect 30268 31778 30324 31780
rect 30268 31726 30270 31778
rect 30270 31726 30322 31778
rect 30322 31726 30324 31778
rect 30268 31724 30324 31726
rect 31500 31778 31556 31780
rect 31500 31726 31502 31778
rect 31502 31726 31554 31778
rect 31554 31726 31556 31778
rect 31500 31724 31556 31726
rect 33068 33516 33124 33572
rect 32172 32786 32228 32788
rect 32172 32734 32174 32786
rect 32174 32734 32226 32786
rect 32226 32734 32228 32786
rect 32172 32732 32228 32734
rect 32508 32844 32564 32900
rect 33292 36652 33348 36708
rect 33404 38444 33460 38500
rect 33516 37436 33572 37492
rect 33964 43650 34020 43652
rect 33964 43598 33966 43650
rect 33966 43598 34018 43650
rect 34018 43598 34020 43650
rect 33964 43596 34020 43598
rect 33852 43538 33908 43540
rect 33852 43486 33854 43538
rect 33854 43486 33906 43538
rect 33906 43486 33908 43538
rect 33852 43484 33908 43486
rect 34524 45836 34580 45892
rect 34748 46002 34804 46004
rect 34748 45950 34750 46002
rect 34750 45950 34802 46002
rect 34802 45950 34804 46002
rect 34748 45948 34804 45950
rect 34412 44546 34468 44548
rect 34412 44494 34414 44546
rect 34414 44494 34466 44546
rect 34466 44494 34468 44546
rect 34412 44492 34468 44494
rect 33964 43148 34020 43204
rect 34300 43260 34356 43316
rect 34188 42812 34244 42868
rect 33964 42252 34020 42308
rect 34524 43596 34580 43652
rect 43820 50764 43876 50820
rect 45276 52332 45332 52388
rect 45276 52108 45332 52164
rect 44940 51602 44996 51604
rect 44940 51550 44942 51602
rect 44942 51550 44994 51602
rect 44994 51550 44996 51602
rect 44940 51548 44996 51550
rect 44044 50988 44100 51044
rect 45948 52668 46004 52724
rect 45612 52162 45668 52164
rect 45612 52110 45614 52162
rect 45614 52110 45666 52162
rect 45666 52110 45668 52162
rect 45612 52108 45668 52110
rect 45836 52444 45892 52500
rect 45612 50988 45668 51044
rect 43932 50652 43988 50708
rect 43820 49922 43876 49924
rect 43820 49870 43822 49922
rect 43822 49870 43874 49922
rect 43874 49870 43876 49922
rect 43820 49868 43876 49870
rect 44044 49980 44100 50036
rect 44940 49756 44996 49812
rect 43596 48076 43652 48132
rect 44492 48354 44548 48356
rect 44492 48302 44494 48354
rect 44494 48302 44546 48354
rect 44546 48302 44548 48354
rect 44492 48300 44548 48302
rect 44268 47570 44324 47572
rect 44268 47518 44270 47570
rect 44270 47518 44322 47570
rect 44322 47518 44324 47570
rect 44268 47516 44324 47518
rect 36316 47292 36372 47348
rect 35084 47180 35140 47236
rect 35644 47234 35700 47236
rect 35644 47182 35646 47234
rect 35646 47182 35698 47234
rect 35698 47182 35700 47234
rect 35644 47180 35700 47182
rect 40348 47180 40404 47236
rect 37660 47068 37716 47124
rect 35532 46620 35588 46676
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35644 45948 35700 46004
rect 35532 45890 35588 45892
rect 35532 45838 35534 45890
rect 35534 45838 35586 45890
rect 35586 45838 35588 45890
rect 35532 45836 35588 45838
rect 34972 45164 35028 45220
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34972 44380 35028 44436
rect 36428 43708 36484 43764
rect 35644 43650 35700 43652
rect 35644 43598 35646 43650
rect 35646 43598 35698 43650
rect 35698 43598 35700 43650
rect 35644 43596 35700 43598
rect 34524 42754 34580 42756
rect 34524 42702 34526 42754
rect 34526 42702 34578 42754
rect 34578 42702 34580 42754
rect 34524 42700 34580 42702
rect 34412 42476 34468 42532
rect 34300 42028 34356 42084
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35420 42866 35476 42868
rect 35420 42814 35422 42866
rect 35422 42814 35474 42866
rect 35474 42814 35476 42866
rect 35420 42812 35476 42814
rect 34860 42642 34916 42644
rect 34860 42590 34862 42642
rect 34862 42590 34914 42642
rect 34914 42590 34916 42642
rect 34860 42588 34916 42590
rect 35084 42364 35140 42420
rect 34524 42028 34580 42084
rect 34860 41692 34916 41748
rect 34972 42140 35028 42196
rect 35868 42252 35924 42308
rect 35420 42194 35476 42196
rect 35420 42142 35422 42194
rect 35422 42142 35474 42194
rect 35474 42142 35476 42194
rect 35420 42140 35476 42142
rect 35756 42028 35812 42084
rect 35196 41970 35252 41972
rect 35196 41918 35198 41970
rect 35198 41918 35250 41970
rect 35250 41918 35252 41970
rect 35196 41916 35252 41918
rect 36540 42252 36596 42308
rect 34860 41298 34916 41300
rect 34860 41246 34862 41298
rect 34862 41246 34914 41298
rect 34914 41246 34916 41298
rect 34860 41244 34916 41246
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 34524 40626 34580 40628
rect 34524 40574 34526 40626
rect 34526 40574 34578 40626
rect 34578 40574 34580 40626
rect 34524 40572 34580 40574
rect 33740 40124 33796 40180
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34300 39004 34356 39060
rect 33628 37772 33684 37828
rect 33404 37100 33460 37156
rect 33516 34914 33572 34916
rect 33516 34862 33518 34914
rect 33518 34862 33570 34914
rect 33570 34862 33572 34914
rect 33516 34860 33572 34862
rect 33516 32732 33572 32788
rect 32060 30994 32116 30996
rect 32060 30942 32062 30994
rect 32062 30942 32114 30994
rect 32114 30942 32116 30994
rect 32060 30940 32116 30942
rect 31276 30882 31332 30884
rect 31276 30830 31278 30882
rect 31278 30830 31330 30882
rect 31330 30830 31332 30882
rect 31276 30828 31332 30830
rect 30268 30210 30324 30212
rect 30268 30158 30270 30210
rect 30270 30158 30322 30210
rect 30322 30158 30324 30210
rect 30268 30156 30324 30158
rect 28812 29538 28868 29540
rect 28812 29486 28814 29538
rect 28814 29486 28866 29538
rect 28866 29486 28868 29538
rect 28812 29484 28868 29486
rect 28700 29426 28756 29428
rect 28700 29374 28702 29426
rect 28702 29374 28754 29426
rect 28754 29374 28756 29426
rect 28700 29372 28756 29374
rect 29708 29596 29764 29652
rect 30156 29932 30212 29988
rect 31276 29650 31332 29652
rect 31276 29598 31278 29650
rect 31278 29598 31330 29650
rect 31330 29598 31332 29650
rect 31276 29596 31332 29598
rect 28252 28866 28308 28868
rect 28252 28814 28254 28866
rect 28254 28814 28306 28866
rect 28306 28814 28308 28866
rect 28252 28812 28308 28814
rect 28476 28588 28532 28644
rect 27020 27074 27076 27076
rect 27020 27022 27022 27074
rect 27022 27022 27074 27074
rect 27074 27022 27076 27074
rect 27020 27020 27076 27022
rect 26684 26908 26740 26964
rect 24780 25116 24836 25172
rect 26460 26796 26516 26852
rect 25676 25340 25732 25396
rect 24444 25004 24500 25060
rect 24556 24892 24612 24948
rect 25116 25004 25172 25060
rect 24444 24556 24500 24612
rect 24220 23884 24276 23940
rect 24332 23660 24388 23716
rect 23660 21868 23716 21924
rect 23660 21532 23716 21588
rect 23660 20524 23716 20580
rect 23324 19740 23380 19796
rect 23100 19516 23156 19572
rect 22652 19122 22708 19124
rect 22652 19070 22654 19122
rect 22654 19070 22706 19122
rect 22706 19070 22708 19122
rect 22652 19068 22708 19070
rect 22876 18956 22932 19012
rect 22092 18450 22148 18452
rect 22092 18398 22094 18450
rect 22094 18398 22146 18450
rect 22146 18398 22148 18450
rect 22092 18396 22148 18398
rect 21980 18060 22036 18116
rect 21420 16828 21476 16884
rect 21308 15372 21364 15428
rect 21532 15148 21588 15204
rect 22540 17500 22596 17556
rect 19516 13580 19572 13636
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20412 14028 20468 14084
rect 19628 13356 19684 13412
rect 22316 16828 22372 16884
rect 21196 14028 21252 14084
rect 21868 13746 21924 13748
rect 21868 13694 21870 13746
rect 21870 13694 21922 13746
rect 21922 13694 21924 13746
rect 21868 13692 21924 13694
rect 20300 13580 20356 13636
rect 19740 13020 19796 13076
rect 20300 13186 20356 13188
rect 20300 13134 20302 13186
rect 20302 13134 20354 13186
rect 20354 13134 20356 13186
rect 20300 13132 20356 13134
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19964 12402 20020 12404
rect 19964 12350 19966 12402
rect 19966 12350 20018 12402
rect 20018 12350 20020 12402
rect 19964 12348 20020 12350
rect 21308 13074 21364 13076
rect 21308 13022 21310 13074
rect 21310 13022 21362 13074
rect 21362 13022 21364 13074
rect 21308 13020 21364 13022
rect 19964 11564 20020 11620
rect 20076 11452 20132 11508
rect 21532 12124 21588 12180
rect 20636 11340 20692 11396
rect 20748 11564 20804 11620
rect 20300 11228 20356 11284
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19740 10556 19796 10612
rect 19516 10498 19572 10500
rect 19516 10446 19518 10498
rect 19518 10446 19570 10498
rect 19570 10446 19572 10498
rect 19516 10444 19572 10446
rect 18060 7586 18116 7588
rect 18060 7534 18062 7586
rect 18062 7534 18114 7586
rect 18114 7534 18116 7586
rect 18060 7532 18116 7534
rect 19740 9772 19796 9828
rect 18844 7532 18900 7588
rect 19516 8092 19572 8148
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20076 8146 20132 8148
rect 20076 8094 20078 8146
rect 20078 8094 20130 8146
rect 20130 8094 20132 8146
rect 20076 8092 20132 8094
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 15820 6524 15876 6580
rect 17724 6578 17780 6580
rect 17724 6526 17726 6578
rect 17726 6526 17778 6578
rect 17778 6526 17780 6578
rect 17724 6524 17780 6526
rect 18508 6524 18564 6580
rect 21420 11506 21476 11508
rect 21420 11454 21422 11506
rect 21422 11454 21474 11506
rect 21474 11454 21476 11506
rect 21420 11452 21476 11454
rect 21868 12850 21924 12852
rect 21868 12798 21870 12850
rect 21870 12798 21922 12850
rect 21922 12798 21924 12850
rect 21868 12796 21924 12798
rect 21644 11564 21700 11620
rect 22204 14700 22260 14756
rect 22764 17388 22820 17444
rect 22652 15874 22708 15876
rect 22652 15822 22654 15874
rect 22654 15822 22706 15874
rect 22706 15822 22708 15874
rect 22652 15820 22708 15822
rect 22428 15372 22484 15428
rect 22204 13356 22260 13412
rect 22988 17554 23044 17556
rect 22988 17502 22990 17554
rect 22990 17502 23042 17554
rect 23042 17502 23044 17554
rect 22988 17500 23044 17502
rect 23884 21644 23940 21700
rect 24892 23938 24948 23940
rect 24892 23886 24894 23938
rect 24894 23886 24946 23938
rect 24946 23886 24948 23938
rect 24892 23884 24948 23886
rect 24556 23548 24612 23604
rect 25004 23660 25060 23716
rect 24444 22930 24500 22932
rect 24444 22878 24446 22930
rect 24446 22878 24498 22930
rect 24498 22878 24500 22930
rect 24444 22876 24500 22878
rect 24556 21756 24612 21812
rect 23884 20412 23940 20468
rect 23324 19346 23380 19348
rect 23324 19294 23326 19346
rect 23326 19294 23378 19346
rect 23378 19294 23380 19346
rect 23324 19292 23380 19294
rect 23212 19068 23268 19124
rect 23884 19010 23940 19012
rect 23884 18958 23886 19010
rect 23886 18958 23938 19010
rect 23938 18958 23940 19010
rect 23884 18956 23940 18958
rect 24108 20524 24164 20580
rect 24556 20412 24612 20468
rect 24892 21868 24948 21924
rect 26236 25340 26292 25396
rect 26236 24946 26292 24948
rect 26236 24894 26238 24946
rect 26238 24894 26290 24946
rect 26290 24894 26292 24946
rect 26236 24892 26292 24894
rect 28588 26236 28644 26292
rect 28588 26012 28644 26068
rect 25228 23996 25284 24052
rect 25228 22540 25284 22596
rect 26348 23212 26404 23268
rect 25564 22764 25620 22820
rect 25228 22258 25284 22260
rect 25228 22206 25230 22258
rect 25230 22206 25282 22258
rect 25282 22206 25284 22258
rect 25228 22204 25284 22206
rect 25004 21644 25060 21700
rect 25116 21756 25172 21812
rect 24220 19740 24276 19796
rect 24668 20018 24724 20020
rect 24668 19966 24670 20018
rect 24670 19966 24722 20018
rect 24722 19966 24724 20018
rect 24668 19964 24724 19966
rect 25676 22540 25732 22596
rect 27356 23266 27412 23268
rect 27356 23214 27358 23266
rect 27358 23214 27410 23266
rect 27410 23214 27412 23266
rect 27356 23212 27412 23214
rect 27580 23100 27636 23156
rect 27916 24892 27972 24948
rect 30828 29538 30884 29540
rect 30828 29486 30830 29538
rect 30830 29486 30882 29538
rect 30882 29486 30884 29538
rect 30828 29484 30884 29486
rect 29708 28700 29764 28756
rect 31276 28754 31332 28756
rect 31276 28702 31278 28754
rect 31278 28702 31330 28754
rect 31330 28702 31332 28754
rect 31276 28700 31332 28702
rect 30268 28588 30324 28644
rect 30156 28364 30212 28420
rect 32172 29426 32228 29428
rect 32172 29374 32174 29426
rect 32174 29374 32226 29426
rect 32226 29374 32228 29426
rect 32172 29372 32228 29374
rect 32396 31612 32452 31668
rect 32508 30994 32564 30996
rect 32508 30942 32510 30994
rect 32510 30942 32562 30994
rect 32562 30942 32564 30994
rect 32508 30940 32564 30942
rect 33180 30940 33236 30996
rect 32620 29260 32676 29316
rect 31948 28028 32004 28084
rect 28812 27020 28868 27076
rect 29260 27074 29316 27076
rect 29260 27022 29262 27074
rect 29262 27022 29314 27074
rect 29314 27022 29316 27074
rect 29260 27020 29316 27022
rect 29596 26290 29652 26292
rect 29596 26238 29598 26290
rect 29598 26238 29650 26290
rect 29650 26238 29652 26290
rect 29596 26236 29652 26238
rect 30716 26124 30772 26180
rect 29372 24892 29428 24948
rect 29148 24444 29204 24500
rect 26908 22594 26964 22596
rect 26908 22542 26910 22594
rect 26910 22542 26962 22594
rect 26962 22542 26964 22594
rect 26908 22540 26964 22542
rect 26684 22428 26740 22484
rect 25564 21756 25620 21812
rect 26348 22092 26404 22148
rect 25900 21474 25956 21476
rect 25900 21422 25902 21474
rect 25902 21422 25954 21474
rect 25954 21422 25956 21474
rect 25900 21420 25956 21422
rect 25228 20018 25284 20020
rect 25228 19966 25230 20018
rect 25230 19966 25282 20018
rect 25282 19966 25284 20018
rect 25228 19964 25284 19966
rect 25564 19852 25620 19908
rect 25340 19740 25396 19796
rect 24332 19346 24388 19348
rect 24332 19294 24334 19346
rect 24334 19294 24386 19346
rect 24386 19294 24388 19346
rect 24332 19292 24388 19294
rect 24108 18620 24164 18676
rect 23212 18284 23268 18340
rect 23324 18508 23380 18564
rect 23212 17388 23268 17444
rect 23548 17276 23604 17332
rect 23996 18284 24052 18340
rect 24444 18620 24500 18676
rect 24220 18284 24276 18340
rect 24108 17666 24164 17668
rect 24108 17614 24110 17666
rect 24110 17614 24162 17666
rect 24162 17614 24164 17666
rect 24108 17612 24164 17614
rect 23660 17164 23716 17220
rect 24444 17612 24500 17668
rect 24668 17388 24724 17444
rect 24444 17164 24500 17220
rect 24668 17052 24724 17108
rect 22876 15596 22932 15652
rect 22988 15202 23044 15204
rect 22988 15150 22990 15202
rect 22990 15150 23042 15202
rect 23042 15150 23044 15202
rect 22988 15148 23044 15150
rect 23212 14700 23268 14756
rect 22652 13746 22708 13748
rect 22652 13694 22654 13746
rect 22654 13694 22706 13746
rect 22706 13694 22708 13746
rect 22652 13692 22708 13694
rect 22540 12684 22596 12740
rect 22204 11394 22260 11396
rect 22204 11342 22206 11394
rect 22206 11342 22258 11394
rect 22258 11342 22260 11394
rect 22204 11340 22260 11342
rect 24556 16994 24612 16996
rect 24556 16942 24558 16994
rect 24558 16942 24610 16994
rect 24610 16942 24612 16994
rect 24556 16940 24612 16942
rect 23660 16770 23716 16772
rect 23660 16718 23662 16770
rect 23662 16718 23714 16770
rect 23714 16718 23716 16770
rect 23660 16716 23716 16718
rect 24444 16716 24500 16772
rect 24220 16492 24276 16548
rect 23772 16156 23828 16212
rect 23548 15596 23604 15652
rect 23996 16210 24052 16212
rect 23996 16158 23998 16210
rect 23998 16158 24050 16210
rect 24050 16158 24052 16210
rect 23996 16156 24052 16158
rect 23772 15372 23828 15428
rect 23884 14924 23940 14980
rect 23884 14700 23940 14756
rect 23548 14530 23604 14532
rect 23548 14478 23550 14530
rect 23550 14478 23602 14530
rect 23602 14478 23604 14530
rect 23548 14476 23604 14478
rect 24892 18844 24948 18900
rect 24892 18060 24948 18116
rect 24892 17554 24948 17556
rect 24892 17502 24894 17554
rect 24894 17502 24946 17554
rect 24946 17502 24948 17554
rect 24892 17500 24948 17502
rect 24892 16380 24948 16436
rect 24556 16044 24612 16100
rect 24444 15820 24500 15876
rect 24108 14588 24164 14644
rect 24780 15484 24836 15540
rect 23996 13522 24052 13524
rect 23996 13470 23998 13522
rect 23998 13470 24050 13522
rect 24050 13470 24052 13522
rect 23996 13468 24052 13470
rect 24332 13186 24388 13188
rect 24332 13134 24334 13186
rect 24334 13134 24386 13186
rect 24386 13134 24388 13186
rect 24332 13132 24388 13134
rect 23548 13020 23604 13076
rect 23884 13020 23940 13076
rect 23324 12796 23380 12852
rect 23660 12460 23716 12516
rect 23772 12962 23828 12964
rect 23772 12910 23774 12962
rect 23774 12910 23826 12962
rect 23826 12910 23828 12962
rect 23772 12908 23828 12910
rect 23548 12402 23604 12404
rect 23548 12350 23550 12402
rect 23550 12350 23602 12402
rect 23602 12350 23604 12402
rect 23548 12348 23604 12350
rect 23100 12178 23156 12180
rect 23100 12126 23102 12178
rect 23102 12126 23154 12178
rect 23154 12126 23156 12178
rect 23100 12124 23156 12126
rect 23772 12124 23828 12180
rect 23996 12908 24052 12964
rect 24556 15260 24612 15316
rect 25004 13916 25060 13972
rect 25340 18956 25396 19012
rect 25228 18674 25284 18676
rect 25228 18622 25230 18674
rect 25230 18622 25282 18674
rect 25282 18622 25284 18674
rect 25228 18620 25284 18622
rect 25340 18396 25396 18452
rect 25228 18284 25284 18340
rect 25900 19964 25956 20020
rect 25676 18844 25732 18900
rect 27020 21810 27076 21812
rect 27020 21758 27022 21810
rect 27022 21758 27074 21810
rect 27074 21758 27076 21810
rect 27020 21756 27076 21758
rect 27692 22204 27748 22260
rect 27580 21868 27636 21924
rect 27468 21644 27524 21700
rect 28028 21698 28084 21700
rect 28028 21646 28030 21698
rect 28030 21646 28082 21698
rect 28082 21646 28084 21698
rect 28028 21644 28084 21646
rect 28476 22482 28532 22484
rect 28476 22430 28478 22482
rect 28478 22430 28530 22482
rect 28530 22430 28532 22482
rect 28476 22428 28532 22430
rect 28476 21868 28532 21924
rect 27916 20076 27972 20132
rect 27804 19964 27860 20020
rect 25340 17612 25396 17668
rect 25340 16380 25396 16436
rect 25900 18396 25956 18452
rect 25788 16940 25844 16996
rect 26124 17666 26180 17668
rect 26124 17614 26126 17666
rect 26126 17614 26178 17666
rect 26178 17614 26180 17666
rect 26124 17612 26180 17614
rect 25564 16828 25620 16884
rect 25452 16156 25508 16212
rect 25676 16716 25732 16772
rect 25228 16098 25284 16100
rect 25228 16046 25230 16098
rect 25230 16046 25282 16098
rect 25282 16046 25284 16098
rect 25228 16044 25284 16046
rect 25900 16604 25956 16660
rect 25788 15932 25844 15988
rect 25676 15372 25732 15428
rect 25564 15036 25620 15092
rect 25564 14476 25620 14532
rect 25340 13468 25396 13524
rect 24556 12572 24612 12628
rect 24444 12460 24500 12516
rect 24668 12348 24724 12404
rect 24108 11788 24164 11844
rect 22876 11282 22932 11284
rect 22876 11230 22878 11282
rect 22878 11230 22930 11282
rect 22930 11230 22932 11282
rect 22876 11228 22932 11230
rect 22092 9996 22148 10052
rect 21532 9826 21588 9828
rect 21532 9774 21534 9826
rect 21534 9774 21586 9826
rect 21586 9774 21588 9826
rect 21532 9772 21588 9774
rect 24108 11452 24164 11508
rect 24108 9996 24164 10052
rect 20748 8204 20804 8260
rect 20860 8540 20916 8596
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 21644 9042 21700 9044
rect 21644 8990 21646 9042
rect 21646 8990 21698 9042
rect 21698 8990 21700 9042
rect 21644 8988 21700 8990
rect 22540 8652 22596 8708
rect 21532 8316 21588 8372
rect 21644 8204 21700 8260
rect 21980 8092 22036 8148
rect 21980 7644 22036 7700
rect 22092 6860 22148 6916
rect 22092 6636 22148 6692
rect 21308 5628 21364 5684
rect 21644 5068 21700 5124
rect 20524 4956 20580 5012
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 22316 8316 22372 8372
rect 23212 9154 23268 9156
rect 23212 9102 23214 9154
rect 23214 9102 23266 9154
rect 23266 9102 23268 9154
rect 23212 9100 23268 9102
rect 23324 9042 23380 9044
rect 23324 8990 23326 9042
rect 23326 8990 23378 9042
rect 23378 8990 23380 9042
rect 23324 8988 23380 8990
rect 23100 8652 23156 8708
rect 22876 7698 22932 7700
rect 22876 7646 22878 7698
rect 22878 7646 22930 7698
rect 22930 7646 22932 7698
rect 22876 7644 22932 7646
rect 22540 6690 22596 6692
rect 22540 6638 22542 6690
rect 22542 6638 22594 6690
rect 22594 6638 22596 6690
rect 22540 6636 22596 6638
rect 22204 5964 22260 6020
rect 23100 8370 23156 8372
rect 23100 8318 23102 8370
rect 23102 8318 23154 8370
rect 23154 8318 23156 8370
rect 23100 8316 23156 8318
rect 23324 8204 23380 8260
rect 25228 12796 25284 12852
rect 25452 13074 25508 13076
rect 25452 13022 25454 13074
rect 25454 13022 25506 13074
rect 25506 13022 25508 13074
rect 25452 13020 25508 13022
rect 25900 14252 25956 14308
rect 26796 19180 26852 19236
rect 27692 18396 27748 18452
rect 26348 16940 26404 16996
rect 26460 16828 26516 16884
rect 26572 17164 26628 17220
rect 26684 16828 26740 16884
rect 26684 16322 26740 16324
rect 26684 16270 26686 16322
rect 26686 16270 26738 16322
rect 26738 16270 26740 16322
rect 26684 16268 26740 16270
rect 26572 16156 26628 16212
rect 26236 15932 26292 15988
rect 26908 17388 26964 17444
rect 26236 15596 26292 15652
rect 26236 14812 26292 14868
rect 26236 14588 26292 14644
rect 26124 14364 26180 14420
rect 26236 14306 26292 14308
rect 26236 14254 26238 14306
rect 26238 14254 26290 14306
rect 26290 14254 26292 14306
rect 26236 14252 26292 14254
rect 25788 12684 25844 12740
rect 25788 12402 25844 12404
rect 25788 12350 25790 12402
rect 25790 12350 25842 12402
rect 25842 12350 25844 12402
rect 25788 12348 25844 12350
rect 25676 11506 25732 11508
rect 25676 11454 25678 11506
rect 25678 11454 25730 11506
rect 25730 11454 25732 11506
rect 25676 11452 25732 11454
rect 24668 10220 24724 10276
rect 24332 9100 24388 9156
rect 24780 9212 24836 9268
rect 23996 8204 24052 8260
rect 23660 6860 23716 6916
rect 23324 6018 23380 6020
rect 23324 5966 23326 6018
rect 23326 5966 23378 6018
rect 23378 5966 23380 6018
rect 23324 5964 23380 5966
rect 22764 5682 22820 5684
rect 22764 5630 22766 5682
rect 22766 5630 22818 5682
rect 22818 5630 22820 5682
rect 22764 5628 22820 5630
rect 22764 5122 22820 5124
rect 22764 5070 22766 5122
rect 22766 5070 22818 5122
rect 22818 5070 22820 5122
rect 22764 5068 22820 5070
rect 22092 4956 22148 5012
rect 24668 6690 24724 6692
rect 24668 6638 24670 6690
rect 24670 6638 24722 6690
rect 24722 6638 24724 6690
rect 24668 6636 24724 6638
rect 25564 11228 25620 11284
rect 25564 10220 25620 10276
rect 25340 9266 25396 9268
rect 25340 9214 25342 9266
rect 25342 9214 25394 9266
rect 25394 9214 25396 9266
rect 25340 9212 25396 9214
rect 25340 8428 25396 8484
rect 26124 13020 26180 13076
rect 27132 16492 27188 16548
rect 26572 15708 26628 15764
rect 27020 15708 27076 15764
rect 27916 19068 27972 19124
rect 28364 20076 28420 20132
rect 28028 19010 28084 19012
rect 28028 18958 28030 19010
rect 28030 18958 28082 19010
rect 28082 18958 28084 19010
rect 28028 18956 28084 18958
rect 28364 18450 28420 18452
rect 28364 18398 28366 18450
rect 28366 18398 28418 18450
rect 28418 18398 28420 18450
rect 28364 18396 28420 18398
rect 28028 18226 28084 18228
rect 28028 18174 28030 18226
rect 28030 18174 28082 18226
rect 28082 18174 28084 18226
rect 28028 18172 28084 18174
rect 28364 17836 28420 17892
rect 28588 17612 28644 17668
rect 28364 17388 28420 17444
rect 28140 16994 28196 16996
rect 28140 16942 28142 16994
rect 28142 16942 28194 16994
rect 28194 16942 28196 16994
rect 28140 16940 28196 16942
rect 28700 17164 28756 17220
rect 27468 15986 27524 15988
rect 27468 15934 27470 15986
rect 27470 15934 27522 15986
rect 27522 15934 27524 15986
rect 27468 15932 27524 15934
rect 28588 16882 28644 16884
rect 28588 16830 28590 16882
rect 28590 16830 28642 16882
rect 28642 16830 28644 16882
rect 28588 16828 28644 16830
rect 28252 16770 28308 16772
rect 28252 16718 28254 16770
rect 28254 16718 28306 16770
rect 28306 16718 28308 16770
rect 28252 16716 28308 16718
rect 28140 16268 28196 16324
rect 27244 15538 27300 15540
rect 27244 15486 27246 15538
rect 27246 15486 27298 15538
rect 27298 15486 27300 15538
rect 27244 15484 27300 15486
rect 26460 14364 26516 14420
rect 27132 15148 27188 15204
rect 27580 14924 27636 14980
rect 27020 14700 27076 14756
rect 27244 14812 27300 14868
rect 27020 14418 27076 14420
rect 27020 14366 27022 14418
rect 27022 14366 27074 14418
rect 27074 14366 27076 14418
rect 27020 14364 27076 14366
rect 26460 13746 26516 13748
rect 26460 13694 26462 13746
rect 26462 13694 26514 13746
rect 26514 13694 26516 13746
rect 26460 13692 26516 13694
rect 26460 13522 26516 13524
rect 26460 13470 26462 13522
rect 26462 13470 26514 13522
rect 26514 13470 26516 13522
rect 26460 13468 26516 13470
rect 27020 13970 27076 13972
rect 27020 13918 27022 13970
rect 27022 13918 27074 13970
rect 27074 13918 27076 13970
rect 27020 13916 27076 13918
rect 27468 14700 27524 14756
rect 28028 15036 28084 15092
rect 28588 15426 28644 15428
rect 28588 15374 28590 15426
rect 28590 15374 28642 15426
rect 28642 15374 28644 15426
rect 28588 15372 28644 15374
rect 28252 15314 28308 15316
rect 28252 15262 28254 15314
rect 28254 15262 28306 15314
rect 28306 15262 28308 15314
rect 28252 15260 28308 15262
rect 28476 15036 28532 15092
rect 28252 14700 28308 14756
rect 29484 23212 29540 23268
rect 30716 23266 30772 23268
rect 30716 23214 30718 23266
rect 30718 23214 30770 23266
rect 30770 23214 30772 23266
rect 30716 23212 30772 23214
rect 29596 22482 29652 22484
rect 29596 22430 29598 22482
rect 29598 22430 29650 22482
rect 29650 22430 29652 22482
rect 29596 22428 29652 22430
rect 30044 22316 30100 22372
rect 29820 22258 29876 22260
rect 29820 22206 29822 22258
rect 29822 22206 29874 22258
rect 29874 22206 29876 22258
rect 29820 22204 29876 22206
rect 33516 31724 33572 31780
rect 34188 37826 34244 37828
rect 34188 37774 34190 37826
rect 34190 37774 34242 37826
rect 34242 37774 34244 37826
rect 34188 37772 34244 37774
rect 33964 37660 34020 37716
rect 34412 37548 34468 37604
rect 33740 36482 33796 36484
rect 33740 36430 33742 36482
rect 33742 36430 33794 36482
rect 33794 36430 33796 36482
rect 33740 36428 33796 36430
rect 34748 37436 34804 37492
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35756 41074 35812 41076
rect 35756 41022 35758 41074
rect 35758 41022 35810 41074
rect 35810 41022 35812 41074
rect 35756 41020 35812 41022
rect 36428 41074 36484 41076
rect 36428 41022 36430 41074
rect 36430 41022 36482 41074
rect 36482 41022 36484 41074
rect 36428 41020 36484 41022
rect 36204 40962 36260 40964
rect 36204 40910 36206 40962
rect 36206 40910 36258 40962
rect 36258 40910 36260 40962
rect 36204 40908 36260 40910
rect 36316 40012 36372 40068
rect 36428 39564 36484 39620
rect 37324 45388 37380 45444
rect 37548 43708 37604 43764
rect 36988 42642 37044 42644
rect 36988 42590 36990 42642
rect 36990 42590 37042 42642
rect 37042 42590 37044 42642
rect 36988 42588 37044 42590
rect 37212 42530 37268 42532
rect 37212 42478 37214 42530
rect 37214 42478 37266 42530
rect 37266 42478 37268 42530
rect 37212 42476 37268 42478
rect 37100 42252 37156 42308
rect 37212 42140 37268 42196
rect 37100 41074 37156 41076
rect 37100 41022 37102 41074
rect 37102 41022 37154 41074
rect 37154 41022 37156 41074
rect 37100 41020 37156 41022
rect 37212 40962 37268 40964
rect 37212 40910 37214 40962
rect 37214 40910 37266 40962
rect 37266 40910 37268 40962
rect 37212 40908 37268 40910
rect 37436 40796 37492 40852
rect 37100 39618 37156 39620
rect 37100 39566 37102 39618
rect 37102 39566 37154 39618
rect 37154 39566 37156 39618
rect 37100 39564 37156 39566
rect 38780 46562 38836 46564
rect 38780 46510 38782 46562
rect 38782 46510 38834 46562
rect 38834 46510 38836 46562
rect 38780 46508 38836 46510
rect 38332 45388 38388 45444
rect 37772 44044 37828 44100
rect 38780 45052 38836 45108
rect 38332 44210 38388 44212
rect 38332 44158 38334 44210
rect 38334 44158 38386 44210
rect 38386 44158 38388 44210
rect 38332 44156 38388 44158
rect 38556 44044 38612 44100
rect 37996 43484 38052 43540
rect 39676 45106 39732 45108
rect 39676 45054 39678 45106
rect 39678 45054 39730 45106
rect 39730 45054 39732 45106
rect 39676 45052 39732 45054
rect 40796 45052 40852 45108
rect 39452 44044 39508 44100
rect 39900 43820 39956 43876
rect 39676 43708 39732 43764
rect 38892 43260 38948 43316
rect 39228 43650 39284 43652
rect 39228 43598 39230 43650
rect 39230 43598 39282 43650
rect 39282 43598 39284 43650
rect 39228 43596 39284 43598
rect 39004 43484 39060 43540
rect 39564 43484 39620 43540
rect 38668 42252 38724 42308
rect 38444 41916 38500 41972
rect 38108 41468 38164 41524
rect 38108 40796 38164 40852
rect 37772 40348 37828 40404
rect 38780 40348 38836 40404
rect 37772 40012 37828 40068
rect 37660 39452 37716 39508
rect 36652 38668 36708 38724
rect 36988 38892 37044 38948
rect 36540 38556 36596 38612
rect 35532 37772 35588 37828
rect 36428 37660 36484 37716
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 36204 37266 36260 37268
rect 36204 37214 36206 37266
rect 36206 37214 36258 37266
rect 36258 37214 36260 37266
rect 36204 37212 36260 37214
rect 36876 38444 36932 38500
rect 37324 38556 37380 38612
rect 37884 38610 37940 38612
rect 37884 38558 37886 38610
rect 37886 38558 37938 38610
rect 37938 38558 37940 38610
rect 37884 38556 37940 38558
rect 37772 38444 37828 38500
rect 37100 37660 37156 37716
rect 37212 37548 37268 37604
rect 36652 36988 36708 37044
rect 37212 37212 37268 37268
rect 36092 36482 36148 36484
rect 36092 36430 36094 36482
rect 36094 36430 36146 36482
rect 36146 36430 36148 36482
rect 36092 36428 36148 36430
rect 36988 36482 37044 36484
rect 36988 36430 36990 36482
rect 36990 36430 37042 36482
rect 37042 36430 37044 36482
rect 36988 36428 37044 36430
rect 37212 36482 37268 36484
rect 37212 36430 37214 36482
rect 37214 36430 37266 36482
rect 37266 36430 37268 36482
rect 37212 36428 37268 36430
rect 34636 35756 34692 35812
rect 34076 35644 34132 35700
rect 36988 35756 37044 35812
rect 37996 37996 38052 38052
rect 38444 38946 38500 38948
rect 38444 38894 38446 38946
rect 38446 38894 38498 38946
rect 38498 38894 38500 38946
rect 38444 38892 38500 38894
rect 38332 38834 38388 38836
rect 38332 38782 38334 38834
rect 38334 38782 38386 38834
rect 38386 38782 38388 38834
rect 38332 38780 38388 38782
rect 38108 36764 38164 36820
rect 38780 38780 38836 38836
rect 39788 43314 39844 43316
rect 39788 43262 39790 43314
rect 39790 43262 39842 43314
rect 39842 43262 39844 43314
rect 39788 43260 39844 43262
rect 40124 44322 40180 44324
rect 40124 44270 40126 44322
rect 40126 44270 40178 44322
rect 40178 44270 40180 44322
rect 40124 44268 40180 44270
rect 40236 44156 40292 44212
rect 40236 43484 40292 43540
rect 40348 43820 40404 43876
rect 40348 43372 40404 43428
rect 41244 46450 41300 46452
rect 41244 46398 41246 46450
rect 41246 46398 41298 46450
rect 41298 46398 41300 46450
rect 41244 46396 41300 46398
rect 42140 46844 42196 46900
rect 46620 52444 46676 52500
rect 47404 52444 47460 52500
rect 46620 52274 46676 52276
rect 46620 52222 46622 52274
rect 46622 52222 46674 52274
rect 46674 52222 46676 52274
rect 46620 52220 46676 52222
rect 46508 52162 46564 52164
rect 46508 52110 46510 52162
rect 46510 52110 46562 52162
rect 46562 52110 46564 52162
rect 46508 52108 46564 52110
rect 46060 51324 46116 51380
rect 46620 51602 46676 51604
rect 46620 51550 46622 51602
rect 46622 51550 46674 51602
rect 46674 51550 46676 51602
rect 46620 51548 46676 51550
rect 46956 52108 47012 52164
rect 47068 52050 47124 52052
rect 47068 51998 47070 52050
rect 47070 51998 47122 52050
rect 47122 51998 47124 52050
rect 47068 51996 47124 51998
rect 50092 53788 50148 53844
rect 48188 52162 48244 52164
rect 48188 52110 48190 52162
rect 48190 52110 48242 52162
rect 48242 52110 48244 52162
rect 48188 52108 48244 52110
rect 47180 51324 47236 51380
rect 47740 51324 47796 51380
rect 46060 49084 46116 49140
rect 45388 48300 45444 48356
rect 46172 48130 46228 48132
rect 46172 48078 46174 48130
rect 46174 48078 46226 48130
rect 46226 48078 46228 48130
rect 46172 48076 46228 48078
rect 44604 46620 44660 46676
rect 44828 47570 44884 47572
rect 44828 47518 44830 47570
rect 44830 47518 44882 47570
rect 44882 47518 44884 47570
rect 44828 47516 44884 47518
rect 44380 46562 44436 46564
rect 44380 46510 44382 46562
rect 44382 46510 44434 46562
rect 44434 46510 44436 46562
rect 44380 46508 44436 46510
rect 41804 46396 41860 46452
rect 45052 47234 45108 47236
rect 45052 47182 45054 47234
rect 45054 47182 45106 47234
rect 45106 47182 45108 47234
rect 45052 47180 45108 47182
rect 44940 46674 44996 46676
rect 44940 46622 44942 46674
rect 44942 46622 44994 46674
rect 44994 46622 44996 46674
rect 44940 46620 44996 46622
rect 45052 46508 45108 46564
rect 45164 46844 45220 46900
rect 45500 47516 45556 47572
rect 47068 49810 47124 49812
rect 47068 49758 47070 49810
rect 47070 49758 47122 49810
rect 47122 49758 47124 49810
rect 47068 49756 47124 49758
rect 48076 51324 48132 51380
rect 48300 51996 48356 52052
rect 51324 53842 51380 53844
rect 51324 53790 51326 53842
rect 51326 53790 51378 53842
rect 51378 53790 51380 53842
rect 51324 53788 51380 53790
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 48748 52668 48804 52724
rect 49420 52332 49476 52388
rect 49196 51378 49252 51380
rect 49196 51326 49198 51378
rect 49198 51326 49250 51378
rect 49250 51326 49252 51378
rect 49196 51324 49252 51326
rect 48524 50652 48580 50708
rect 48412 50594 48468 50596
rect 48412 50542 48414 50594
rect 48414 50542 48466 50594
rect 48466 50542 48468 50594
rect 48412 50540 48468 50542
rect 48748 50540 48804 50596
rect 48076 49868 48132 49924
rect 47964 49644 48020 49700
rect 46284 47516 46340 47572
rect 45836 47458 45892 47460
rect 45836 47406 45838 47458
rect 45838 47406 45890 47458
rect 45890 47406 45892 47458
rect 45836 47404 45892 47406
rect 45724 47292 45780 47348
rect 45612 47234 45668 47236
rect 45612 47182 45614 47234
rect 45614 47182 45666 47234
rect 45666 47182 45668 47234
rect 45612 47180 45668 47182
rect 45500 46508 45556 46564
rect 45388 46450 45444 46452
rect 45388 46398 45390 46450
rect 45390 46398 45442 46450
rect 45442 46398 45444 46450
rect 45388 46396 45444 46398
rect 41580 45836 41636 45892
rect 42588 45890 42644 45892
rect 42588 45838 42590 45890
rect 42590 45838 42642 45890
rect 42642 45838 42644 45890
rect 42588 45836 42644 45838
rect 43036 45890 43092 45892
rect 43036 45838 43038 45890
rect 43038 45838 43090 45890
rect 43090 45838 43092 45890
rect 43036 45836 43092 45838
rect 44940 45836 44996 45892
rect 46396 48354 46452 48356
rect 46396 48302 46398 48354
rect 46398 48302 46450 48354
rect 46450 48302 46452 48354
rect 46396 48300 46452 48302
rect 47068 48300 47124 48356
rect 47404 48130 47460 48132
rect 47404 48078 47406 48130
rect 47406 48078 47458 48130
rect 47458 48078 47460 48130
rect 47404 48076 47460 48078
rect 46620 47346 46676 47348
rect 46620 47294 46622 47346
rect 46622 47294 46674 47346
rect 46674 47294 46676 47346
rect 46620 47292 46676 47294
rect 46508 46732 46564 46788
rect 47292 47458 47348 47460
rect 47292 47406 47294 47458
rect 47294 47406 47346 47458
rect 47346 47406 47348 47458
rect 47292 47404 47348 47406
rect 47852 48354 47908 48356
rect 47852 48302 47854 48354
rect 47854 48302 47906 48354
rect 47906 48302 47908 48354
rect 47852 48300 47908 48302
rect 48748 49922 48804 49924
rect 48748 49870 48750 49922
rect 48750 49870 48802 49922
rect 48802 49870 48804 49922
rect 48748 49868 48804 49870
rect 49084 49980 49140 50036
rect 48972 49420 49028 49476
rect 48748 49196 48804 49252
rect 46844 47292 46900 47348
rect 48300 47346 48356 47348
rect 48300 47294 48302 47346
rect 48302 47294 48354 47346
rect 48354 47294 48356 47346
rect 48300 47292 48356 47294
rect 47740 46956 47796 47012
rect 46844 46674 46900 46676
rect 46844 46622 46846 46674
rect 46846 46622 46898 46674
rect 46898 46622 46900 46674
rect 46844 46620 46900 46622
rect 47292 46674 47348 46676
rect 47292 46622 47294 46674
rect 47294 46622 47346 46674
rect 47346 46622 47348 46674
rect 47292 46620 47348 46622
rect 49980 52668 50036 52724
rect 49756 52108 49812 52164
rect 49420 51212 49476 51268
rect 49756 50876 49812 50932
rect 50428 52108 50484 52164
rect 50204 51324 50260 51380
rect 51100 52108 51156 52164
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 51212 51548 51268 51604
rect 50652 51490 50708 51492
rect 50652 51438 50654 51490
rect 50654 51438 50706 51490
rect 50706 51438 50708 51490
rect 50652 51436 50708 51438
rect 53228 51490 53284 51492
rect 53228 51438 53230 51490
rect 53230 51438 53282 51490
rect 53282 51438 53284 51490
rect 53228 51436 53284 51438
rect 50764 51378 50820 51380
rect 50764 51326 50766 51378
rect 50766 51326 50818 51378
rect 50818 51326 50820 51378
rect 50764 51324 50820 51326
rect 50764 51100 50820 51156
rect 50316 50876 50372 50932
rect 50764 50764 50820 50820
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 49868 49980 49924 50036
rect 49756 49868 49812 49924
rect 50764 49922 50820 49924
rect 50764 49870 50766 49922
rect 50766 49870 50818 49922
rect 50818 49870 50820 49922
rect 50764 49868 50820 49870
rect 48972 48636 49028 48692
rect 48860 47570 48916 47572
rect 48860 47518 48862 47570
rect 48862 47518 48914 47570
rect 48914 47518 48916 47570
rect 48860 47516 48916 47518
rect 49196 48412 49252 48468
rect 49644 48802 49700 48804
rect 49644 48750 49646 48802
rect 49646 48750 49698 48802
rect 49698 48750 49700 48802
rect 49644 48748 49700 48750
rect 51100 51266 51156 51268
rect 51100 51214 51102 51266
rect 51102 51214 51154 51266
rect 51154 51214 51156 51266
rect 51100 51212 51156 51214
rect 51996 51212 52052 51268
rect 51996 50764 52052 50820
rect 51660 50706 51716 50708
rect 51660 50654 51662 50706
rect 51662 50654 51714 50706
rect 51714 50654 51716 50706
rect 51660 50652 51716 50654
rect 51884 50540 51940 50596
rect 51548 50428 51604 50484
rect 52108 50706 52164 50708
rect 52108 50654 52110 50706
rect 52110 50654 52162 50706
rect 52162 50654 52164 50706
rect 52108 50652 52164 50654
rect 52668 50652 52724 50708
rect 53900 50652 53956 50708
rect 55580 51212 55636 51268
rect 53452 50482 53508 50484
rect 53452 50430 53454 50482
rect 53454 50430 53506 50482
rect 53506 50430 53508 50482
rect 53452 50428 53508 50430
rect 52220 50034 52276 50036
rect 52220 49982 52222 50034
rect 52222 49982 52274 50034
rect 52274 49982 52276 50034
rect 52220 49980 52276 49982
rect 49980 49698 50036 49700
rect 49980 49646 49982 49698
rect 49982 49646 50034 49698
rect 50034 49646 50036 49698
rect 49980 49644 50036 49646
rect 50316 49084 50372 49140
rect 50092 48972 50148 49028
rect 49980 48636 50036 48692
rect 48972 47068 49028 47124
rect 48748 46956 48804 47012
rect 47964 46732 48020 46788
rect 48076 46674 48132 46676
rect 48076 46622 48078 46674
rect 48078 46622 48130 46674
rect 48130 46622 48132 46674
rect 48076 46620 48132 46622
rect 47740 46450 47796 46452
rect 47740 46398 47742 46450
rect 47742 46398 47794 46450
rect 47794 46398 47796 46450
rect 47740 46396 47796 46398
rect 48860 46674 48916 46676
rect 48860 46622 48862 46674
rect 48862 46622 48914 46674
rect 48914 46622 48916 46674
rect 48860 46620 48916 46622
rect 49084 46674 49140 46676
rect 49084 46622 49086 46674
rect 49086 46622 49138 46674
rect 49138 46622 49140 46674
rect 49084 46620 49140 46622
rect 50204 48860 50260 48916
rect 50876 48972 50932 49028
rect 50540 48860 50596 48916
rect 50428 48748 50484 48804
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50540 48412 50596 48468
rect 50876 48412 50932 48468
rect 51324 49196 51380 49252
rect 51100 48748 51156 48804
rect 53452 48412 53508 48468
rect 49868 47292 49924 47348
rect 50428 47292 50484 47348
rect 49644 47068 49700 47124
rect 49980 46956 50036 47012
rect 44940 45388 44996 45444
rect 47628 45276 47684 45332
rect 41020 44268 41076 44324
rect 40908 44098 40964 44100
rect 40908 44046 40910 44098
rect 40910 44046 40962 44098
rect 40962 44046 40964 44098
rect 40908 44044 40964 44046
rect 40796 43820 40852 43876
rect 41020 43708 41076 43764
rect 40460 43596 40516 43652
rect 40124 42588 40180 42644
rect 40908 42642 40964 42644
rect 40908 42590 40910 42642
rect 40910 42590 40962 42642
rect 40962 42590 40964 42642
rect 40908 42588 40964 42590
rect 39676 41970 39732 41972
rect 39676 41918 39678 41970
rect 39678 41918 39730 41970
rect 39730 41918 39732 41970
rect 39676 41916 39732 41918
rect 39228 41298 39284 41300
rect 39228 41246 39230 41298
rect 39230 41246 39282 41298
rect 39282 41246 39284 41298
rect 39228 41244 39284 41246
rect 39564 41692 39620 41748
rect 39452 40908 39508 40964
rect 39788 41244 39844 41300
rect 39676 40908 39732 40964
rect 40012 40124 40068 40180
rect 39900 39564 39956 39620
rect 40348 39564 40404 39620
rect 41132 42530 41188 42532
rect 41132 42478 41134 42530
rect 41134 42478 41186 42530
rect 41186 42478 41188 42530
rect 41132 42476 41188 42478
rect 41692 44322 41748 44324
rect 41692 44270 41694 44322
rect 41694 44270 41746 44322
rect 41746 44270 41748 44322
rect 41692 44268 41748 44270
rect 41804 44210 41860 44212
rect 41804 44158 41806 44210
rect 41806 44158 41858 44210
rect 41858 44158 41860 44210
rect 41804 44156 41860 44158
rect 42476 44322 42532 44324
rect 42476 44270 42478 44322
rect 42478 44270 42530 44322
rect 42530 44270 42532 44322
rect 42476 44268 42532 44270
rect 42700 44156 42756 44212
rect 41916 44098 41972 44100
rect 41916 44046 41918 44098
rect 41918 44046 41970 44098
rect 41970 44046 41972 44098
rect 41916 44044 41972 44046
rect 42252 43820 42308 43876
rect 41580 43538 41636 43540
rect 41580 43486 41582 43538
rect 41582 43486 41634 43538
rect 41634 43486 41636 43538
rect 41580 43484 41636 43486
rect 41804 43426 41860 43428
rect 41804 43374 41806 43426
rect 41806 43374 41858 43426
rect 41858 43374 41860 43426
rect 41804 43372 41860 43374
rect 49084 45276 49140 45332
rect 50764 47180 50820 47236
rect 51324 47234 51380 47236
rect 51324 47182 51326 47234
rect 51326 47182 51378 47234
rect 51378 47182 51380 47234
rect 51324 47180 51380 47182
rect 51772 47234 51828 47236
rect 51772 47182 51774 47234
rect 51774 47182 51826 47234
rect 51826 47182 51828 47234
rect 51772 47180 51828 47182
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50540 46844 50596 46900
rect 51772 46674 51828 46676
rect 51772 46622 51774 46674
rect 51774 46622 51826 46674
rect 51826 46622 51828 46674
rect 51772 46620 51828 46622
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 44828 44434 44884 44436
rect 44828 44382 44830 44434
rect 44830 44382 44882 44434
rect 44882 44382 44884 44434
rect 44828 44380 44884 44382
rect 44940 43596 44996 43652
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 47068 43650 47124 43652
rect 47068 43598 47070 43650
rect 47070 43598 47122 43650
rect 47122 43598 47124 43650
rect 47068 43596 47124 43598
rect 49980 43596 50036 43652
rect 48188 43484 48244 43540
rect 48860 43538 48916 43540
rect 48860 43486 48862 43538
rect 48862 43486 48914 43538
rect 48914 43486 48916 43538
rect 48860 43484 48916 43486
rect 44380 43372 44436 43428
rect 43484 43260 43540 43316
rect 42252 42754 42308 42756
rect 42252 42702 42254 42754
rect 42254 42702 42306 42754
rect 42306 42702 42308 42754
rect 42252 42700 42308 42702
rect 41804 41746 41860 41748
rect 41804 41694 41806 41746
rect 41806 41694 41858 41746
rect 41858 41694 41860 41746
rect 41804 41692 41860 41694
rect 42476 42530 42532 42532
rect 42476 42478 42478 42530
rect 42478 42478 42530 42530
rect 42530 42478 42532 42530
rect 42476 42476 42532 42478
rect 43372 42530 43428 42532
rect 43372 42478 43374 42530
rect 43374 42478 43426 42530
rect 43426 42478 43428 42530
rect 43372 42476 43428 42478
rect 43372 41692 43428 41748
rect 41580 41074 41636 41076
rect 41580 41022 41582 41074
rect 41582 41022 41634 41074
rect 41634 41022 41636 41074
rect 41580 41020 41636 41022
rect 41692 40962 41748 40964
rect 41692 40910 41694 40962
rect 41694 40910 41746 40962
rect 41746 40910 41748 40962
rect 41692 40908 41748 40910
rect 41916 40572 41972 40628
rect 41468 40402 41524 40404
rect 41468 40350 41470 40402
rect 41470 40350 41522 40402
rect 41522 40350 41524 40402
rect 41468 40348 41524 40350
rect 42588 40908 42644 40964
rect 42812 40460 42868 40516
rect 42140 40348 42196 40404
rect 42700 40402 42756 40404
rect 42700 40350 42702 40402
rect 42702 40350 42754 40402
rect 42754 40350 42756 40402
rect 42700 40348 42756 40350
rect 41356 39618 41412 39620
rect 41356 39566 41358 39618
rect 41358 39566 41410 39618
rect 41410 39566 41412 39618
rect 41356 39564 41412 39566
rect 41468 39452 41524 39508
rect 39228 38050 39284 38052
rect 39228 37998 39230 38050
rect 39230 37998 39282 38050
rect 39282 37998 39284 38050
rect 39228 37996 39284 37998
rect 38780 37548 38836 37604
rect 34972 35644 35028 35700
rect 34860 35532 34916 35588
rect 34860 35308 34916 35364
rect 36764 35644 36820 35700
rect 36652 35532 36708 35588
rect 35532 35474 35588 35476
rect 35532 35422 35534 35474
rect 35534 35422 35586 35474
rect 35586 35422 35588 35474
rect 35532 35420 35588 35422
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 33852 34636 33908 34692
rect 34748 34690 34804 34692
rect 34748 34638 34750 34690
rect 34750 34638 34802 34690
rect 34802 34638 34804 34690
rect 34748 34636 34804 34638
rect 34748 33964 34804 34020
rect 33852 33458 33908 33460
rect 33852 33406 33854 33458
rect 33854 33406 33906 33458
rect 33906 33406 33908 33458
rect 33852 33404 33908 33406
rect 34188 32786 34244 32788
rect 34188 32734 34190 32786
rect 34190 32734 34242 32786
rect 34242 32734 34244 32786
rect 34188 32732 34244 32734
rect 33740 31836 33796 31892
rect 35308 34914 35364 34916
rect 35308 34862 35310 34914
rect 35310 34862 35362 34914
rect 35362 34862 35364 34914
rect 35308 34860 35364 34862
rect 40348 38556 40404 38612
rect 40124 37996 40180 38052
rect 39676 37490 39732 37492
rect 39676 37438 39678 37490
rect 39678 37438 39730 37490
rect 39730 37438 39732 37490
rect 39676 37436 39732 37438
rect 38892 37266 38948 37268
rect 38892 37214 38894 37266
rect 38894 37214 38946 37266
rect 38946 37214 38948 37266
rect 38892 37212 38948 37214
rect 38892 36764 38948 36820
rect 39788 36652 39844 36708
rect 38892 36258 38948 36260
rect 38892 36206 38894 36258
rect 38894 36206 38946 36258
rect 38946 36206 38948 36258
rect 38892 36204 38948 36206
rect 40012 37266 40068 37268
rect 40012 37214 40014 37266
rect 40014 37214 40066 37266
rect 40066 37214 40068 37266
rect 40012 37212 40068 37214
rect 41468 39004 41524 39060
rect 40236 36764 40292 36820
rect 40460 36652 40516 36708
rect 36652 34860 36708 34916
rect 37212 34914 37268 34916
rect 37212 34862 37214 34914
rect 37214 34862 37266 34914
rect 37266 34862 37268 34914
rect 37212 34860 37268 34862
rect 36988 34748 37044 34804
rect 36764 34130 36820 34132
rect 36764 34078 36766 34130
rect 36766 34078 36818 34130
rect 36818 34078 36820 34130
rect 36764 34076 36820 34078
rect 35980 34018 36036 34020
rect 35980 33966 35982 34018
rect 35982 33966 36034 34018
rect 36034 33966 36036 34018
rect 35980 33964 36036 33966
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35084 33404 35140 33460
rect 35532 33346 35588 33348
rect 35532 33294 35534 33346
rect 35534 33294 35586 33346
rect 35586 33294 35588 33346
rect 35532 33292 35588 33294
rect 36652 33964 36708 34020
rect 35980 33292 36036 33348
rect 35420 32844 35476 32900
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 34748 31948 34804 32004
rect 34412 31836 34468 31892
rect 33852 31666 33908 31668
rect 33852 31614 33854 31666
rect 33854 31614 33906 31666
rect 33906 31614 33908 31666
rect 33852 31612 33908 31614
rect 33740 30994 33796 30996
rect 33740 30942 33742 30994
rect 33742 30942 33794 30994
rect 33794 30942 33796 30994
rect 33740 30940 33796 30942
rect 34300 31778 34356 31780
rect 34300 31726 34302 31778
rect 34302 31726 34354 31778
rect 34354 31726 34356 31778
rect 34300 31724 34356 31726
rect 34524 31500 34580 31556
rect 35644 32620 35700 32676
rect 35532 31612 35588 31668
rect 35196 31554 35252 31556
rect 35196 31502 35198 31554
rect 35198 31502 35250 31554
rect 35250 31502 35252 31554
rect 35196 31500 35252 31502
rect 35196 30828 35252 30884
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 33852 30044 33908 30100
rect 33628 29932 33684 29988
rect 33628 29372 33684 29428
rect 33516 29314 33572 29316
rect 33516 29262 33518 29314
rect 33518 29262 33570 29314
rect 33570 29262 33572 29314
rect 33516 29260 33572 29262
rect 33404 28700 33460 28756
rect 32844 28418 32900 28420
rect 32844 28366 32846 28418
rect 32846 28366 32898 28418
rect 32898 28366 32900 28418
rect 32844 28364 32900 28366
rect 32956 27804 33012 27860
rect 32396 27020 32452 27076
rect 33068 27132 33124 27188
rect 32844 26796 32900 26852
rect 32956 26684 33012 26740
rect 33516 28812 33572 28868
rect 33404 27858 33460 27860
rect 33404 27806 33406 27858
rect 33406 27806 33458 27858
rect 33458 27806 33460 27858
rect 33404 27804 33460 27806
rect 33404 27074 33460 27076
rect 33404 27022 33406 27074
rect 33406 27022 33458 27074
rect 33458 27022 33460 27074
rect 33404 27020 33460 27022
rect 33180 26796 33236 26852
rect 33068 26290 33124 26292
rect 33068 26238 33070 26290
rect 33070 26238 33122 26290
rect 33122 26238 33124 26290
rect 33068 26236 33124 26238
rect 33180 26178 33236 26180
rect 33180 26126 33182 26178
rect 33182 26126 33234 26178
rect 33234 26126 33236 26178
rect 33180 26124 33236 26126
rect 33516 25900 33572 25956
rect 33180 24050 33236 24052
rect 33180 23998 33182 24050
rect 33182 23998 33234 24050
rect 33234 23998 33236 24050
rect 33180 23996 33236 23998
rect 34972 30268 35028 30324
rect 34188 29426 34244 29428
rect 34188 29374 34190 29426
rect 34190 29374 34242 29426
rect 34242 29374 34244 29426
rect 34188 29372 34244 29374
rect 34636 29372 34692 29428
rect 35420 29932 35476 29988
rect 35084 29372 35140 29428
rect 35196 29314 35252 29316
rect 35196 29262 35198 29314
rect 35198 29262 35250 29314
rect 35250 29262 35252 29314
rect 35196 29260 35252 29262
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 28866 35252 28868
rect 35196 28814 35198 28866
rect 35198 28814 35250 28866
rect 35250 28814 35252 28866
rect 35196 28812 35252 28814
rect 34412 27804 34468 27860
rect 34860 28028 34916 28084
rect 34188 27020 34244 27076
rect 34636 27074 34692 27076
rect 34636 27022 34638 27074
rect 34638 27022 34690 27074
rect 34690 27022 34692 27074
rect 34636 27020 34692 27022
rect 34300 26908 34356 26964
rect 33740 26290 33796 26292
rect 33740 26238 33742 26290
rect 33742 26238 33794 26290
rect 33794 26238 33796 26290
rect 33740 26236 33796 26238
rect 33964 26124 34020 26180
rect 35196 27804 35252 27860
rect 37548 34076 37604 34132
rect 37100 33964 37156 34020
rect 36988 32844 37044 32900
rect 38892 35644 38948 35700
rect 39564 34636 39620 34692
rect 38556 33516 38612 33572
rect 38556 32844 38612 32900
rect 37436 32674 37492 32676
rect 37436 32622 37438 32674
rect 37438 32622 37490 32674
rect 37490 32622 37492 32674
rect 37436 32620 37492 32622
rect 38444 32620 38500 32676
rect 39340 32508 39396 32564
rect 36204 31836 36260 31892
rect 37548 31836 37604 31892
rect 35980 31554 36036 31556
rect 35980 31502 35982 31554
rect 35982 31502 36034 31554
rect 36034 31502 36036 31554
rect 35980 31500 36036 31502
rect 36428 31554 36484 31556
rect 36428 31502 36430 31554
rect 36430 31502 36482 31554
rect 36482 31502 36484 31554
rect 36428 31500 36484 31502
rect 38108 31836 38164 31892
rect 36092 30434 36148 30436
rect 36092 30382 36094 30434
rect 36094 30382 36146 30434
rect 36146 30382 36148 30434
rect 36092 30380 36148 30382
rect 35756 30322 35812 30324
rect 35756 30270 35758 30322
rect 35758 30270 35810 30322
rect 35810 30270 35812 30322
rect 35756 30268 35812 30270
rect 36540 30156 36596 30212
rect 35980 29986 36036 29988
rect 35980 29934 35982 29986
rect 35982 29934 36034 29986
rect 36034 29934 36036 29986
rect 35980 29932 36036 29934
rect 36092 28700 36148 28756
rect 35980 28588 36036 28644
rect 35644 28028 35700 28084
rect 34860 27132 34916 27188
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35084 27020 35140 27076
rect 35196 27244 35252 27300
rect 35644 27020 35700 27076
rect 35196 26908 35252 26964
rect 34300 26348 34356 26404
rect 34076 25116 34132 25172
rect 33964 24610 34020 24612
rect 33964 24558 33966 24610
rect 33966 24558 34018 24610
rect 34018 24558 34020 24610
rect 33964 24556 34020 24558
rect 33852 23996 33908 24052
rect 33628 23378 33684 23380
rect 33628 23326 33630 23378
rect 33630 23326 33682 23378
rect 33682 23326 33684 23378
rect 33628 23324 33684 23326
rect 34188 23996 34244 24052
rect 34524 25564 34580 25620
rect 35084 26402 35140 26404
rect 35084 26350 35086 26402
rect 35086 26350 35138 26402
rect 35138 26350 35140 26402
rect 35084 26348 35140 26350
rect 35532 26850 35588 26852
rect 35532 26798 35534 26850
rect 35534 26798 35586 26850
rect 35586 26798 35588 26850
rect 35532 26796 35588 26798
rect 34860 26236 34916 26292
rect 35756 26684 35812 26740
rect 35868 27132 35924 27188
rect 34972 26124 35028 26180
rect 34860 25228 34916 25284
rect 34860 24556 34916 24612
rect 34636 23660 34692 23716
rect 32172 22876 32228 22932
rect 29596 19852 29652 19908
rect 29820 19122 29876 19124
rect 29820 19070 29822 19122
rect 29822 19070 29874 19122
rect 29874 19070 29876 19122
rect 29820 19068 29876 19070
rect 29372 18508 29428 18564
rect 29148 17666 29204 17668
rect 29148 17614 29150 17666
rect 29150 17614 29202 17666
rect 29202 17614 29204 17666
rect 29148 17612 29204 17614
rect 29708 18396 29764 18452
rect 29260 16268 29316 16324
rect 29148 16098 29204 16100
rect 29148 16046 29150 16098
rect 29150 16046 29202 16098
rect 29202 16046 29204 16098
rect 29148 16044 29204 16046
rect 29148 15708 29204 15764
rect 29596 17890 29652 17892
rect 29596 17838 29598 17890
rect 29598 17838 29650 17890
rect 29650 17838 29652 17890
rect 29596 17836 29652 17838
rect 29708 16156 29764 16212
rect 29596 15932 29652 15988
rect 29036 15426 29092 15428
rect 29036 15374 29038 15426
rect 29038 15374 29090 15426
rect 29090 15374 29092 15426
rect 29036 15372 29092 15374
rect 29484 15148 29540 15204
rect 27804 13746 27860 13748
rect 27804 13694 27806 13746
rect 27806 13694 27858 13746
rect 27858 13694 27860 13746
rect 27804 13692 27860 13694
rect 27020 13468 27076 13524
rect 26236 12572 26292 12628
rect 26236 12348 26292 12404
rect 26236 11452 26292 11508
rect 25564 8540 25620 8596
rect 26012 8540 26068 8596
rect 25676 7644 25732 7700
rect 23772 5180 23828 5236
rect 27356 12962 27412 12964
rect 27356 12910 27358 12962
rect 27358 12910 27410 12962
rect 27410 12910 27412 12962
rect 27356 12908 27412 12910
rect 27132 12850 27188 12852
rect 27132 12798 27134 12850
rect 27134 12798 27186 12850
rect 27186 12798 27188 12850
rect 27132 12796 27188 12798
rect 28588 12850 28644 12852
rect 28588 12798 28590 12850
rect 28590 12798 28642 12850
rect 28642 12798 28644 12850
rect 28588 12796 28644 12798
rect 28364 12460 28420 12516
rect 27468 12348 27524 12404
rect 28252 12402 28308 12404
rect 28252 12350 28254 12402
rect 28254 12350 28306 12402
rect 28306 12350 28308 12402
rect 28252 12348 28308 12350
rect 28252 12178 28308 12180
rect 28252 12126 28254 12178
rect 28254 12126 28306 12178
rect 28306 12126 28308 12178
rect 28252 12124 28308 12126
rect 28476 11676 28532 11732
rect 26908 11340 26964 11396
rect 26572 10780 26628 10836
rect 29148 12908 29204 12964
rect 29596 12460 29652 12516
rect 29148 12236 29204 12292
rect 28700 11228 28756 11284
rect 27132 10834 27188 10836
rect 27132 10782 27134 10834
rect 27134 10782 27186 10834
rect 27186 10782 27188 10834
rect 27132 10780 27188 10782
rect 26796 10722 26852 10724
rect 26796 10670 26798 10722
rect 26798 10670 26850 10722
rect 26850 10670 26852 10722
rect 26796 10668 26852 10670
rect 28588 10722 28644 10724
rect 28588 10670 28590 10722
rect 28590 10670 28642 10722
rect 28642 10670 28644 10722
rect 28588 10668 28644 10670
rect 26908 9884 26964 9940
rect 27244 9884 27300 9940
rect 27580 9938 27636 9940
rect 27580 9886 27582 9938
rect 27582 9886 27634 9938
rect 27634 9886 27636 9938
rect 27580 9884 27636 9886
rect 28924 9884 28980 9940
rect 28252 9548 28308 9604
rect 27356 8204 27412 8260
rect 26684 7532 26740 7588
rect 26572 6860 26628 6916
rect 27916 8652 27972 8708
rect 30380 19122 30436 19124
rect 30380 19070 30382 19122
rect 30382 19070 30434 19122
rect 30434 19070 30436 19122
rect 30380 19068 30436 19070
rect 33964 22092 34020 22148
rect 34412 22146 34468 22148
rect 34412 22094 34414 22146
rect 34414 22094 34466 22146
rect 34466 22094 34468 22146
rect 34412 22092 34468 22094
rect 34412 21868 34468 21924
rect 34636 21756 34692 21812
rect 34748 22316 34804 22372
rect 34972 23378 35028 23380
rect 34972 23326 34974 23378
rect 34974 23326 35026 23378
rect 35026 23326 35028 23378
rect 34972 23324 35028 23326
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35532 24892 35588 24948
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 23660 35252 23716
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35644 24780 35700 24836
rect 36316 28700 36372 28756
rect 36652 27970 36708 27972
rect 36652 27918 36654 27970
rect 36654 27918 36706 27970
rect 36706 27918 36708 27970
rect 36652 27916 36708 27918
rect 36540 27858 36596 27860
rect 36540 27806 36542 27858
rect 36542 27806 36594 27858
rect 36594 27806 36596 27858
rect 36540 27804 36596 27806
rect 36092 27074 36148 27076
rect 36092 27022 36094 27074
rect 36094 27022 36146 27074
rect 36146 27022 36148 27074
rect 36092 27020 36148 27022
rect 37660 31612 37716 31668
rect 37436 31500 37492 31556
rect 37100 30380 37156 30436
rect 36988 30210 37044 30212
rect 36988 30158 36990 30210
rect 36990 30158 37042 30210
rect 37042 30158 37044 30210
rect 36988 30156 37044 30158
rect 37324 30210 37380 30212
rect 37324 30158 37326 30210
rect 37326 30158 37378 30210
rect 37378 30158 37380 30210
rect 37324 30156 37380 30158
rect 38780 31890 38836 31892
rect 38780 31838 38782 31890
rect 38782 31838 38834 31890
rect 38834 31838 38836 31890
rect 38780 31836 38836 31838
rect 40236 35420 40292 35476
rect 41020 37490 41076 37492
rect 41020 37438 41022 37490
rect 41022 37438 41074 37490
rect 41074 37438 41076 37490
rect 41020 37436 41076 37438
rect 40908 35084 40964 35140
rect 41020 35644 41076 35700
rect 41020 34972 41076 35028
rect 40348 34076 40404 34132
rect 41244 35084 41300 35140
rect 42028 39506 42084 39508
rect 42028 39454 42030 39506
rect 42030 39454 42082 39506
rect 42082 39454 42084 39506
rect 42028 39452 42084 39454
rect 42588 39452 42644 39508
rect 42140 39058 42196 39060
rect 42140 39006 42142 39058
rect 42142 39006 42194 39058
rect 42194 39006 42196 39058
rect 42140 39004 42196 39006
rect 42476 38834 42532 38836
rect 42476 38782 42478 38834
rect 42478 38782 42530 38834
rect 42530 38782 42532 38834
rect 42476 38780 42532 38782
rect 42924 40012 42980 40068
rect 43036 40348 43092 40404
rect 43148 40290 43204 40292
rect 43148 40238 43150 40290
rect 43150 40238 43202 40290
rect 43202 40238 43204 40290
rect 43148 40236 43204 40238
rect 43260 40124 43316 40180
rect 43260 38780 43316 38836
rect 43484 41244 43540 41300
rect 44156 41244 44212 41300
rect 44268 41074 44324 41076
rect 44268 41022 44270 41074
rect 44270 41022 44322 41074
rect 44322 41022 44324 41074
rect 44268 41020 44324 41022
rect 44268 40460 44324 40516
rect 43932 40178 43988 40180
rect 43932 40126 43934 40178
rect 43934 40126 43986 40178
rect 43986 40126 43988 40178
rect 43932 40124 43988 40126
rect 46284 43260 46340 43316
rect 45612 43036 45668 43092
rect 44604 42588 44660 42644
rect 44492 40290 44548 40292
rect 44492 40238 44494 40290
rect 44494 40238 44546 40290
rect 44546 40238 44548 40290
rect 44492 40236 44548 40238
rect 45500 42700 45556 42756
rect 45052 42476 45108 42532
rect 45276 42364 45332 42420
rect 45164 40572 45220 40628
rect 47516 43260 47572 43316
rect 46396 43036 46452 43092
rect 47740 42924 47796 42980
rect 46060 42642 46116 42644
rect 46060 42590 46062 42642
rect 46062 42590 46114 42642
rect 46114 42590 46116 42642
rect 46060 42588 46116 42590
rect 45276 40684 45332 40740
rect 44940 40514 44996 40516
rect 44940 40462 44942 40514
rect 44942 40462 44994 40514
rect 44994 40462 44996 40514
rect 44940 40460 44996 40462
rect 45724 41468 45780 41524
rect 43820 39116 43876 39172
rect 44268 39116 44324 39172
rect 44044 39058 44100 39060
rect 44044 39006 44046 39058
rect 44046 39006 44098 39058
rect 44098 39006 44100 39058
rect 44044 39004 44100 39006
rect 43708 38946 43764 38948
rect 43708 38894 43710 38946
rect 43710 38894 43762 38946
rect 43762 38894 43764 38946
rect 43708 38892 43764 38894
rect 44268 38946 44324 38948
rect 44268 38894 44270 38946
rect 44270 38894 44322 38946
rect 44322 38894 44324 38946
rect 44268 38892 44324 38894
rect 42700 38108 42756 38164
rect 44604 38722 44660 38724
rect 44604 38670 44606 38722
rect 44606 38670 44658 38722
rect 44658 38670 44660 38722
rect 44604 38668 44660 38670
rect 41692 37996 41748 38052
rect 42252 37938 42308 37940
rect 42252 37886 42254 37938
rect 42254 37886 42306 37938
rect 42306 37886 42308 37938
rect 42252 37884 42308 37886
rect 43372 38050 43428 38052
rect 43372 37998 43374 38050
rect 43374 37998 43426 38050
rect 43426 37998 43428 38050
rect 43372 37996 43428 37998
rect 43708 37996 43764 38052
rect 44268 38162 44324 38164
rect 44268 38110 44270 38162
rect 44270 38110 44322 38162
rect 44322 38110 44324 38162
rect 44268 38108 44324 38110
rect 44156 38050 44212 38052
rect 44156 37998 44158 38050
rect 44158 37998 44210 38050
rect 44210 37998 44212 38050
rect 44156 37996 44212 37998
rect 42588 36876 42644 36932
rect 42588 36316 42644 36372
rect 42140 35026 42196 35028
rect 42140 34974 42142 35026
rect 42142 34974 42194 35026
rect 42194 34974 42196 35026
rect 42140 34972 42196 34974
rect 43148 36876 43204 36932
rect 44492 36428 44548 36484
rect 41468 33516 41524 33572
rect 42700 34636 42756 34692
rect 42028 33346 42084 33348
rect 42028 33294 42030 33346
rect 42030 33294 42082 33346
rect 42082 33294 42084 33346
rect 42028 33292 42084 33294
rect 41916 33180 41972 33236
rect 38332 31554 38388 31556
rect 38332 31502 38334 31554
rect 38334 31502 38386 31554
rect 38386 31502 38388 31554
rect 38332 31500 38388 31502
rect 38892 30828 38948 30884
rect 40572 31666 40628 31668
rect 40572 31614 40574 31666
rect 40574 31614 40626 31666
rect 40626 31614 40628 31666
rect 40572 31612 40628 31614
rect 40348 30940 40404 30996
rect 40460 31164 40516 31220
rect 39564 30434 39620 30436
rect 39564 30382 39566 30434
rect 39566 30382 39618 30434
rect 39618 30382 39620 30434
rect 39564 30380 39620 30382
rect 38892 30268 38948 30324
rect 38780 30210 38836 30212
rect 38780 30158 38782 30210
rect 38782 30158 38834 30210
rect 38834 30158 38836 30210
rect 38780 30156 38836 30158
rect 37324 29372 37380 29428
rect 37996 29372 38052 29428
rect 37548 29036 37604 29092
rect 37100 28754 37156 28756
rect 37100 28702 37102 28754
rect 37102 28702 37154 28754
rect 37154 28702 37156 28754
rect 37100 28700 37156 28702
rect 37996 28754 38052 28756
rect 37996 28702 37998 28754
rect 37998 28702 38050 28754
rect 38050 28702 38052 28754
rect 37996 28700 38052 28702
rect 38332 28642 38388 28644
rect 38332 28590 38334 28642
rect 38334 28590 38386 28642
rect 38386 28590 38388 28642
rect 38332 28588 38388 28590
rect 36876 26796 36932 26852
rect 37100 26684 37156 26740
rect 37324 26572 37380 26628
rect 36428 25564 36484 25620
rect 37548 25564 37604 25620
rect 35756 22876 35812 22932
rect 33740 21420 33796 21476
rect 33852 21644 33908 21700
rect 30828 20076 30884 20132
rect 31276 19906 31332 19908
rect 31276 19854 31278 19906
rect 31278 19854 31330 19906
rect 31330 19854 31332 19906
rect 31276 19852 31332 19854
rect 30604 18732 30660 18788
rect 32396 18396 32452 18452
rect 32172 17666 32228 17668
rect 32172 17614 32174 17666
rect 32174 17614 32226 17666
rect 32226 17614 32228 17666
rect 32172 17612 32228 17614
rect 31836 17554 31892 17556
rect 31836 17502 31838 17554
rect 31838 17502 31890 17554
rect 31890 17502 31892 17554
rect 31836 17500 31892 17502
rect 35756 22370 35812 22372
rect 35756 22318 35758 22370
rect 35758 22318 35810 22370
rect 35810 22318 35812 22370
rect 35756 22316 35812 22318
rect 35196 21810 35252 21812
rect 35196 21758 35198 21810
rect 35198 21758 35250 21810
rect 35250 21758 35252 21810
rect 35196 21756 35252 21758
rect 35756 21980 35812 22036
rect 36316 24556 36372 24612
rect 36092 24050 36148 24052
rect 36092 23998 36094 24050
rect 36094 23998 36146 24050
rect 36146 23998 36148 24050
rect 36092 23996 36148 23998
rect 36204 23826 36260 23828
rect 36204 23774 36206 23826
rect 36206 23774 36258 23826
rect 36258 23774 36260 23826
rect 36204 23772 36260 23774
rect 36428 23772 36484 23828
rect 36652 24220 36708 24276
rect 36204 22652 36260 22708
rect 35980 22540 36036 22596
rect 34524 20802 34580 20804
rect 34524 20750 34526 20802
rect 34526 20750 34578 20802
rect 34578 20750 34580 20802
rect 34524 20748 34580 20750
rect 34748 20076 34804 20132
rect 34300 19906 34356 19908
rect 34300 19854 34302 19906
rect 34302 19854 34354 19906
rect 34354 19854 34356 19906
rect 34300 19852 34356 19854
rect 33068 19740 33124 19796
rect 33404 17612 33460 17668
rect 30604 17052 30660 17108
rect 33404 16940 33460 16996
rect 32508 16882 32564 16884
rect 32508 16830 32510 16882
rect 32510 16830 32562 16882
rect 32562 16830 32564 16882
rect 32508 16828 32564 16830
rect 33180 16882 33236 16884
rect 33180 16830 33182 16882
rect 33182 16830 33234 16882
rect 33234 16830 33236 16882
rect 33180 16828 33236 16830
rect 30716 16604 30772 16660
rect 29932 15708 29988 15764
rect 29932 15148 29988 15204
rect 29932 11564 29988 11620
rect 29820 10332 29876 10388
rect 30716 15708 30772 15764
rect 31276 15986 31332 15988
rect 31276 15934 31278 15986
rect 31278 15934 31330 15986
rect 31330 15934 31332 15986
rect 31276 15932 31332 15934
rect 30940 15596 30996 15652
rect 31388 15596 31444 15652
rect 30940 15372 30996 15428
rect 31724 15426 31780 15428
rect 31724 15374 31726 15426
rect 31726 15374 31778 15426
rect 31778 15374 31780 15426
rect 31724 15372 31780 15374
rect 30828 14418 30884 14420
rect 30828 14366 30830 14418
rect 30830 14366 30882 14418
rect 30882 14366 30884 14418
rect 30828 14364 30884 14366
rect 31276 12850 31332 12852
rect 31276 12798 31278 12850
rect 31278 12798 31330 12850
rect 31330 12798 31332 12850
rect 31276 12796 31332 12798
rect 30268 12684 30324 12740
rect 30492 12290 30548 12292
rect 30492 12238 30494 12290
rect 30494 12238 30546 12290
rect 30546 12238 30548 12290
rect 30492 12236 30548 12238
rect 29820 9938 29876 9940
rect 29820 9886 29822 9938
rect 29822 9886 29874 9938
rect 29874 9886 29876 9938
rect 29820 9884 29876 9886
rect 30604 9884 30660 9940
rect 29148 9602 29204 9604
rect 29148 9550 29150 9602
rect 29150 9550 29202 9602
rect 29202 9550 29204 9602
rect 29148 9548 29204 9550
rect 33292 14418 33348 14420
rect 33292 14366 33294 14418
rect 33294 14366 33346 14418
rect 33346 14366 33348 14418
rect 33292 14364 33348 14366
rect 33180 14140 33236 14196
rect 34076 17724 34132 17780
rect 34188 17052 34244 17108
rect 34524 16994 34580 16996
rect 34524 16942 34526 16994
rect 34526 16942 34578 16994
rect 34578 16942 34580 16994
rect 34524 16940 34580 16942
rect 33852 16828 33908 16884
rect 35756 21420 35812 21476
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 20802 35252 20804
rect 35196 20750 35198 20802
rect 35198 20750 35250 20802
rect 35250 20750 35252 20802
rect 35196 20748 35252 20750
rect 35308 20130 35364 20132
rect 35308 20078 35310 20130
rect 35310 20078 35362 20130
rect 35362 20078 35364 20130
rect 35308 20076 35364 20078
rect 34860 19964 34916 20020
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18396 35252 18452
rect 37660 26796 37716 26852
rect 37884 25564 37940 25620
rect 37324 25394 37380 25396
rect 37324 25342 37326 25394
rect 37326 25342 37378 25394
rect 37378 25342 37380 25394
rect 37324 25340 37380 25342
rect 37212 24892 37268 24948
rect 36652 22540 36708 22596
rect 37212 23996 37268 24052
rect 37436 24556 37492 24612
rect 36876 22316 36932 22372
rect 36428 22258 36484 22260
rect 36428 22206 36430 22258
rect 36430 22206 36482 22258
rect 36482 22206 36484 22258
rect 36428 22204 36484 22206
rect 37100 23826 37156 23828
rect 37100 23774 37102 23826
rect 37102 23774 37154 23826
rect 37154 23774 37156 23826
rect 37100 23772 37156 23774
rect 37212 23714 37268 23716
rect 37212 23662 37214 23714
rect 37214 23662 37266 23714
rect 37266 23662 37268 23714
rect 37212 23660 37268 23662
rect 36988 22204 37044 22260
rect 37100 23436 37156 23492
rect 38332 26850 38388 26852
rect 38332 26798 38334 26850
rect 38334 26798 38386 26850
rect 38386 26798 38388 26850
rect 38332 26796 38388 26798
rect 38780 27186 38836 27188
rect 38780 27134 38782 27186
rect 38782 27134 38834 27186
rect 38834 27134 38836 27186
rect 38780 27132 38836 27134
rect 40460 30268 40516 30324
rect 38892 26572 38948 26628
rect 38108 25340 38164 25396
rect 37996 23884 38052 23940
rect 37100 21980 37156 22036
rect 37212 22652 37268 22708
rect 35980 19852 36036 19908
rect 35756 19740 35812 19796
rect 36316 19852 36372 19908
rect 38220 23324 38276 23380
rect 37324 22204 37380 22260
rect 37660 21420 37716 21476
rect 38556 23436 38612 23492
rect 38332 22930 38388 22932
rect 38332 22878 38334 22930
rect 38334 22878 38386 22930
rect 38386 22878 38388 22930
rect 38332 22876 38388 22878
rect 38220 22428 38276 22484
rect 40124 30210 40180 30212
rect 40124 30158 40126 30210
rect 40126 30158 40178 30210
rect 40178 30158 40180 30210
rect 40124 30156 40180 30158
rect 41020 30716 41076 30772
rect 40796 30210 40852 30212
rect 40796 30158 40798 30210
rect 40798 30158 40850 30210
rect 40850 30158 40852 30210
rect 40796 30156 40852 30158
rect 39676 28754 39732 28756
rect 39676 28702 39678 28754
rect 39678 28702 39730 28754
rect 39730 28702 39732 28754
rect 39676 28700 39732 28702
rect 41244 31052 41300 31108
rect 41244 29036 41300 29092
rect 40684 28700 40740 28756
rect 40012 27692 40068 27748
rect 39564 27132 39620 27188
rect 39228 24892 39284 24948
rect 39116 24834 39172 24836
rect 39116 24782 39118 24834
rect 39118 24782 39170 24834
rect 39170 24782 39172 24834
rect 39116 24780 39172 24782
rect 38332 21868 38388 21924
rect 38444 21644 38500 21700
rect 40012 26572 40068 26628
rect 39788 26290 39844 26292
rect 39788 26238 39790 26290
rect 39790 26238 39842 26290
rect 39842 26238 39844 26290
rect 39788 26236 39844 26238
rect 39788 25004 39844 25060
rect 39900 23324 39956 23380
rect 40236 26572 40292 26628
rect 40348 25116 40404 25172
rect 39340 21756 39396 21812
rect 39116 21644 39172 21700
rect 36092 19122 36148 19124
rect 36092 19070 36094 19122
rect 36094 19070 36146 19122
rect 36146 19070 36148 19122
rect 36092 19068 36148 19070
rect 35644 18844 35700 18900
rect 36316 18844 36372 18900
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35532 17778 35588 17780
rect 35532 17726 35534 17778
rect 35534 17726 35586 17778
rect 35586 17726 35588 17778
rect 35532 17724 35588 17726
rect 34636 16828 34692 16884
rect 35532 17052 35588 17108
rect 33964 16658 34020 16660
rect 33964 16606 33966 16658
rect 33966 16606 34018 16658
rect 34018 16606 34020 16658
rect 33964 16604 34020 16606
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 15036 35252 15092
rect 35420 15426 35476 15428
rect 35420 15374 35422 15426
rect 35422 15374 35474 15426
rect 35474 15374 35476 15426
rect 35420 15372 35476 15374
rect 35756 15484 35812 15540
rect 36204 17666 36260 17668
rect 36204 17614 36206 17666
rect 36206 17614 36258 17666
rect 36258 17614 36260 17666
rect 36204 17612 36260 17614
rect 36204 16828 36260 16884
rect 37884 19906 37940 19908
rect 37884 19854 37886 19906
rect 37886 19854 37938 19906
rect 37938 19854 37940 19906
rect 37884 19852 37940 19854
rect 38556 19906 38612 19908
rect 38556 19854 38558 19906
rect 38558 19854 38610 19906
rect 38610 19854 38612 19906
rect 38556 19852 38612 19854
rect 37436 18844 37492 18900
rect 37660 18450 37716 18452
rect 37660 18398 37662 18450
rect 37662 18398 37714 18450
rect 37714 18398 37716 18450
rect 37660 18396 37716 18398
rect 39900 22316 39956 22372
rect 40348 24780 40404 24836
rect 40012 21644 40068 21700
rect 40236 23772 40292 23828
rect 40236 22428 40292 22484
rect 39228 21420 39284 21476
rect 39676 21420 39732 21476
rect 41916 32450 41972 32452
rect 41916 32398 41918 32450
rect 41918 32398 41970 32450
rect 41970 32398 41972 32450
rect 41916 32396 41972 32398
rect 41916 31612 41972 31668
rect 42140 30994 42196 30996
rect 42140 30942 42142 30994
rect 42142 30942 42194 30994
rect 42194 30942 42196 30994
rect 42140 30940 42196 30942
rect 41468 30156 41524 30212
rect 42140 29820 42196 29876
rect 41356 28700 41412 28756
rect 41916 28588 41972 28644
rect 42588 34076 42644 34132
rect 44380 36204 44436 36260
rect 44044 35868 44100 35924
rect 43036 34636 43092 34692
rect 44268 35586 44324 35588
rect 44268 35534 44270 35586
rect 44270 35534 44322 35586
rect 44322 35534 44324 35586
rect 44268 35532 44324 35534
rect 44156 35420 44212 35476
rect 43596 34748 43652 34804
rect 43372 34690 43428 34692
rect 43372 34638 43374 34690
rect 43374 34638 43426 34690
rect 43426 34638 43428 34690
rect 43372 34636 43428 34638
rect 43372 34242 43428 34244
rect 43372 34190 43374 34242
rect 43374 34190 43426 34242
rect 43426 34190 43428 34242
rect 43372 34188 43428 34190
rect 43820 34524 43876 34580
rect 42924 32844 42980 32900
rect 43260 32674 43316 32676
rect 43260 32622 43262 32674
rect 43262 32622 43314 32674
rect 43314 32622 43316 32674
rect 43260 32620 43316 32622
rect 43148 32450 43204 32452
rect 43148 32398 43150 32450
rect 43150 32398 43202 32450
rect 43202 32398 43204 32450
rect 43148 32396 43204 32398
rect 42700 31500 42756 31556
rect 42364 28588 42420 28644
rect 43260 31612 43316 31668
rect 43372 31164 43428 31220
rect 44044 31890 44100 31892
rect 44044 31838 44046 31890
rect 44046 31838 44098 31890
rect 44098 31838 44100 31890
rect 44044 31836 44100 31838
rect 45388 39618 45444 39620
rect 45388 39566 45390 39618
rect 45390 39566 45442 39618
rect 45442 39566 45444 39618
rect 45388 39564 45444 39566
rect 44828 39452 44884 39508
rect 45164 38834 45220 38836
rect 45164 38782 45166 38834
rect 45166 38782 45218 38834
rect 45218 38782 45220 38834
rect 45164 38780 45220 38782
rect 45612 40124 45668 40180
rect 45724 40012 45780 40068
rect 45724 39228 45780 39284
rect 46172 40012 46228 40068
rect 45612 38780 45668 38836
rect 45836 38892 45892 38948
rect 45948 38780 46004 38836
rect 45724 38668 45780 38724
rect 45500 38332 45556 38388
rect 44828 38108 44884 38164
rect 45052 38162 45108 38164
rect 45052 38110 45054 38162
rect 45054 38110 45106 38162
rect 45106 38110 45108 38162
rect 45052 38108 45108 38110
rect 44940 37938 44996 37940
rect 44940 37886 44942 37938
rect 44942 37886 44994 37938
rect 44994 37886 44996 37938
rect 44940 37884 44996 37886
rect 45388 37884 45444 37940
rect 45500 37996 45556 38052
rect 45052 37100 45108 37156
rect 45164 36428 45220 36484
rect 46284 39116 46340 39172
rect 47404 42252 47460 42308
rect 46732 41858 46788 41860
rect 46732 41806 46734 41858
rect 46734 41806 46786 41858
rect 46786 41806 46788 41858
rect 46732 41804 46788 41806
rect 46508 40626 46564 40628
rect 46508 40574 46510 40626
rect 46510 40574 46562 40626
rect 46562 40574 46564 40626
rect 46508 40572 46564 40574
rect 46508 39340 46564 39396
rect 46844 40684 46900 40740
rect 47740 41580 47796 41636
rect 49084 42754 49140 42756
rect 49084 42702 49086 42754
rect 49086 42702 49138 42754
rect 49138 42702 49140 42754
rect 49084 42700 49140 42702
rect 48748 42252 48804 42308
rect 47404 40684 47460 40740
rect 46732 39618 46788 39620
rect 46732 39566 46734 39618
rect 46734 39566 46786 39618
rect 46786 39566 46788 39618
rect 46732 39564 46788 39566
rect 46844 39228 46900 39284
rect 46956 39452 47012 39508
rect 48076 40402 48132 40404
rect 48076 40350 48078 40402
rect 48078 40350 48130 40402
rect 48130 40350 48132 40402
rect 48076 40348 48132 40350
rect 47180 39228 47236 39284
rect 47404 40124 47460 40180
rect 46060 38108 46116 38164
rect 44716 36204 44772 36260
rect 45612 36258 45668 36260
rect 45612 36206 45614 36258
rect 45614 36206 45666 36258
rect 45666 36206 45668 36258
rect 45612 36204 45668 36206
rect 44716 35420 44772 35476
rect 45164 35922 45220 35924
rect 45164 35870 45166 35922
rect 45166 35870 45218 35922
rect 45218 35870 45220 35922
rect 45164 35868 45220 35870
rect 44828 34802 44884 34804
rect 44828 34750 44830 34802
rect 44830 34750 44882 34802
rect 44882 34750 44884 34802
rect 44828 34748 44884 34750
rect 45724 35644 45780 35700
rect 45500 35532 45556 35588
rect 45164 34860 45220 34916
rect 45388 34860 45444 34916
rect 44940 34524 44996 34580
rect 45612 35420 45668 35476
rect 45500 34300 45556 34356
rect 45612 34188 45668 34244
rect 46172 36482 46228 36484
rect 46172 36430 46174 36482
rect 46174 36430 46226 36482
rect 46226 36430 46228 36482
rect 46172 36428 46228 36430
rect 45948 35532 46004 35588
rect 46172 35644 46228 35700
rect 46060 34914 46116 34916
rect 46060 34862 46062 34914
rect 46062 34862 46114 34914
rect 46114 34862 46116 34914
rect 46060 34860 46116 34862
rect 45388 33068 45444 33124
rect 44828 32562 44884 32564
rect 44828 32510 44830 32562
rect 44830 32510 44882 32562
rect 44882 32510 44884 32562
rect 44828 32508 44884 32510
rect 44492 31612 44548 31668
rect 43596 30940 43652 30996
rect 43932 30604 43988 30660
rect 42476 30210 42532 30212
rect 42476 30158 42478 30210
rect 42478 30158 42530 30210
rect 42530 30158 42532 30210
rect 42476 30156 42532 30158
rect 43148 30210 43204 30212
rect 43148 30158 43150 30210
rect 43150 30158 43202 30210
rect 43202 30158 43204 30210
rect 43148 30156 43204 30158
rect 41916 27132 41972 27188
rect 42028 27692 42084 27748
rect 42476 27020 42532 27076
rect 42364 26908 42420 26964
rect 42140 26572 42196 26628
rect 40796 26012 40852 26068
rect 41020 26236 41076 26292
rect 40572 25004 40628 25060
rect 40460 23660 40516 23716
rect 40572 24108 40628 24164
rect 41020 24946 41076 24948
rect 41020 24894 41022 24946
rect 41022 24894 41074 24946
rect 41074 24894 41076 24946
rect 41020 24892 41076 24894
rect 41692 25394 41748 25396
rect 41692 25342 41694 25394
rect 41694 25342 41746 25394
rect 41746 25342 41748 25394
rect 41692 25340 41748 25342
rect 40908 24722 40964 24724
rect 40908 24670 40910 24722
rect 40910 24670 40962 24722
rect 40962 24670 40964 24722
rect 40908 24668 40964 24670
rect 41804 25116 41860 25172
rect 40796 23938 40852 23940
rect 40796 23886 40798 23938
rect 40798 23886 40850 23938
rect 40850 23886 40852 23938
rect 40796 23884 40852 23886
rect 40684 23826 40740 23828
rect 40684 23774 40686 23826
rect 40686 23774 40738 23826
rect 40738 23774 40740 23826
rect 40684 23772 40740 23774
rect 40348 21868 40404 21924
rect 40796 22370 40852 22372
rect 40796 22318 40798 22370
rect 40798 22318 40850 22370
rect 40850 22318 40852 22370
rect 40796 22316 40852 22318
rect 41356 24108 41412 24164
rect 41356 23772 41412 23828
rect 41916 24668 41972 24724
rect 41804 23938 41860 23940
rect 41804 23886 41806 23938
rect 41806 23886 41858 23938
rect 41858 23886 41860 23938
rect 41804 23884 41860 23886
rect 42252 24108 42308 24164
rect 42476 25340 42532 25396
rect 43484 29986 43540 29988
rect 43484 29934 43486 29986
rect 43486 29934 43538 29986
rect 43538 29934 43540 29986
rect 43484 29932 43540 29934
rect 43372 28642 43428 28644
rect 43372 28590 43374 28642
rect 43374 28590 43426 28642
rect 43426 28590 43428 28642
rect 43372 28588 43428 28590
rect 43708 29314 43764 29316
rect 43708 29262 43710 29314
rect 43710 29262 43762 29314
rect 43762 29262 43764 29314
rect 43708 29260 43764 29262
rect 44156 30994 44212 30996
rect 44156 30942 44158 30994
rect 44158 30942 44210 30994
rect 44210 30942 44212 30994
rect 44156 30940 44212 30942
rect 44716 30940 44772 30996
rect 44940 31052 44996 31108
rect 44716 30604 44772 30660
rect 44716 29932 44772 29988
rect 45948 34636 46004 34692
rect 46732 38780 46788 38836
rect 47068 38780 47124 38836
rect 48076 39564 48132 39620
rect 48972 41186 49028 41188
rect 48972 41134 48974 41186
rect 48974 41134 49026 41186
rect 49026 41134 49028 41186
rect 48972 41132 49028 41134
rect 49868 43372 49924 43428
rect 49868 42754 49924 42756
rect 49868 42702 49870 42754
rect 49870 42702 49922 42754
rect 49922 42702 49924 42754
rect 49868 42700 49924 42702
rect 49308 42642 49364 42644
rect 49308 42590 49310 42642
rect 49310 42590 49362 42642
rect 49362 42590 49364 42642
rect 49308 42588 49364 42590
rect 49756 42588 49812 42644
rect 49420 41804 49476 41860
rect 49756 41580 49812 41636
rect 52108 43650 52164 43652
rect 52108 43598 52110 43650
rect 52110 43598 52162 43650
rect 52162 43598 52164 43650
rect 52108 43596 52164 43598
rect 51660 43426 51716 43428
rect 51660 43374 51662 43426
rect 51662 43374 51714 43426
rect 51714 43374 51716 43426
rect 51660 43372 51716 43374
rect 50540 42924 50596 42980
rect 51996 42812 52052 42868
rect 50988 42588 51044 42644
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50316 41186 50372 41188
rect 50316 41134 50318 41186
rect 50318 41134 50370 41186
rect 50370 41134 50372 41186
rect 50316 41132 50372 41134
rect 49420 40572 49476 40628
rect 47740 39116 47796 39172
rect 47628 38722 47684 38724
rect 47628 38670 47630 38722
rect 47630 38670 47682 38722
rect 47682 38670 47684 38722
rect 47628 38668 47684 38670
rect 46620 38332 46676 38388
rect 47628 37490 47684 37492
rect 47628 37438 47630 37490
rect 47630 37438 47682 37490
rect 47682 37438 47684 37490
rect 47628 37436 47684 37438
rect 46620 37100 46676 37156
rect 46508 36652 46564 36708
rect 47628 37212 47684 37268
rect 46956 36428 47012 36484
rect 47068 36764 47124 36820
rect 46732 36204 46788 36260
rect 46732 35698 46788 35700
rect 46732 35646 46734 35698
rect 46734 35646 46786 35698
rect 46786 35646 46788 35698
rect 46732 35644 46788 35646
rect 46620 34802 46676 34804
rect 46620 34750 46622 34802
rect 46622 34750 46674 34802
rect 46674 34750 46676 34802
rect 46620 34748 46676 34750
rect 47292 35644 47348 35700
rect 47068 35532 47124 35588
rect 46732 34130 46788 34132
rect 46732 34078 46734 34130
rect 46734 34078 46786 34130
rect 46786 34078 46788 34130
rect 46732 34076 46788 34078
rect 46060 33292 46116 33348
rect 45836 33068 45892 33124
rect 45724 32508 45780 32564
rect 46508 33234 46564 33236
rect 46508 33182 46510 33234
rect 46510 33182 46562 33234
rect 46562 33182 46564 33234
rect 46508 33180 46564 33182
rect 46620 33122 46676 33124
rect 46620 33070 46622 33122
rect 46622 33070 46674 33122
rect 46674 33070 46676 33122
rect 46620 33068 46676 33070
rect 46060 32338 46116 32340
rect 46060 32286 46062 32338
rect 46062 32286 46114 32338
rect 46114 32286 46116 32338
rect 46060 32284 46116 32286
rect 45612 31724 45668 31780
rect 45276 30492 45332 30548
rect 45388 30380 45444 30436
rect 45500 30268 45556 30324
rect 44828 29596 44884 29652
rect 45164 29932 45220 29988
rect 45052 29820 45108 29876
rect 44156 29426 44212 29428
rect 44156 29374 44158 29426
rect 44158 29374 44210 29426
rect 44210 29374 44212 29426
rect 44156 29372 44212 29374
rect 43932 28642 43988 28644
rect 43932 28590 43934 28642
rect 43934 28590 43986 28642
rect 43986 28590 43988 28642
rect 43932 28588 43988 28590
rect 44940 28924 44996 28980
rect 43036 27692 43092 27748
rect 42924 27244 42980 27300
rect 43036 27132 43092 27188
rect 42700 24668 42756 24724
rect 42812 25900 42868 25956
rect 43260 26962 43316 26964
rect 43260 26910 43262 26962
rect 43262 26910 43314 26962
rect 43314 26910 43316 26962
rect 43260 26908 43316 26910
rect 43148 26236 43204 26292
rect 43148 25506 43204 25508
rect 43148 25454 43150 25506
rect 43150 25454 43202 25506
rect 43202 25454 43204 25506
rect 43148 25452 43204 25454
rect 42364 23884 42420 23940
rect 41916 23548 41972 23604
rect 41468 23324 41524 23380
rect 42924 23884 42980 23940
rect 42028 23266 42084 23268
rect 42028 23214 42030 23266
rect 42030 23214 42082 23266
rect 42082 23214 42084 23266
rect 42028 23212 42084 23214
rect 43036 23660 43092 23716
rect 41804 23154 41860 23156
rect 41804 23102 41806 23154
rect 41806 23102 41858 23154
rect 41858 23102 41860 23154
rect 41804 23100 41860 23102
rect 41692 22316 41748 22372
rect 42588 22764 42644 22820
rect 42364 22092 42420 22148
rect 41580 21868 41636 21924
rect 44828 27244 44884 27300
rect 44156 27074 44212 27076
rect 44156 27022 44158 27074
rect 44158 27022 44210 27074
rect 44210 27022 44212 27074
rect 44156 27020 44212 27022
rect 43820 26460 43876 26516
rect 43484 26348 43540 26404
rect 43932 26348 43988 26404
rect 43820 23996 43876 24052
rect 42476 21868 42532 21924
rect 43484 23212 43540 23268
rect 44268 26572 44324 26628
rect 44716 26572 44772 26628
rect 44380 26290 44436 26292
rect 44380 26238 44382 26290
rect 44382 26238 44434 26290
rect 44434 26238 44436 26290
rect 44380 26236 44436 26238
rect 44716 25228 44772 25284
rect 44940 25116 44996 25172
rect 45836 31388 45892 31444
rect 45836 31164 45892 31220
rect 46284 31164 46340 31220
rect 46396 30492 46452 30548
rect 45836 29260 45892 29316
rect 45276 29148 45332 29204
rect 45164 27692 45220 27748
rect 45500 28924 45556 28980
rect 46060 29148 46116 29204
rect 46620 31052 46676 31108
rect 46620 30380 46676 30436
rect 46844 33346 46900 33348
rect 46844 33294 46846 33346
rect 46846 33294 46898 33346
rect 46898 33294 46900 33346
rect 46844 33292 46900 33294
rect 47180 33068 47236 33124
rect 49196 40402 49252 40404
rect 49196 40350 49198 40402
rect 49198 40350 49250 40402
rect 49250 40350 49252 40402
rect 49196 40348 49252 40350
rect 48748 39340 48804 39396
rect 49980 40124 50036 40180
rect 49868 39618 49924 39620
rect 49868 39566 49870 39618
rect 49870 39566 49922 39618
rect 49922 39566 49924 39618
rect 49868 39564 49924 39566
rect 50092 39564 50148 39620
rect 48524 39228 48580 39284
rect 48076 38946 48132 38948
rect 48076 38894 48078 38946
rect 48078 38894 48130 38946
rect 48130 38894 48132 38946
rect 48076 38892 48132 38894
rect 47964 38834 48020 38836
rect 47964 38782 47966 38834
rect 47966 38782 48018 38834
rect 48018 38782 48020 38834
rect 47964 38780 48020 38782
rect 48748 38892 48804 38948
rect 49308 38834 49364 38836
rect 49308 38782 49310 38834
rect 49310 38782 49362 38834
rect 49362 38782 49364 38834
rect 49308 38780 49364 38782
rect 49532 38834 49588 38836
rect 49532 38782 49534 38834
rect 49534 38782 49586 38834
rect 49586 38782 49588 38834
rect 49532 38780 49588 38782
rect 48524 38668 48580 38724
rect 47628 36764 47684 36820
rect 47516 36428 47572 36484
rect 47516 34412 47572 34468
rect 47740 35980 47796 36036
rect 47852 36204 47908 36260
rect 47740 35756 47796 35812
rect 47852 35532 47908 35588
rect 48188 37042 48244 37044
rect 48188 36990 48190 37042
rect 48190 36990 48242 37042
rect 48242 36990 48244 37042
rect 48188 36988 48244 36990
rect 48076 36482 48132 36484
rect 48076 36430 48078 36482
rect 48078 36430 48130 36482
rect 48130 36430 48132 36482
rect 48076 36428 48132 36430
rect 48188 36316 48244 36372
rect 48076 36092 48132 36148
rect 48076 35644 48132 35700
rect 48076 34242 48132 34244
rect 48076 34190 48078 34242
rect 48078 34190 48130 34242
rect 48130 34190 48132 34242
rect 48076 34188 48132 34190
rect 47516 34130 47572 34132
rect 47516 34078 47518 34130
rect 47518 34078 47570 34130
rect 47570 34078 47572 34130
rect 47516 34076 47572 34078
rect 46732 30268 46788 30324
rect 46956 32396 47012 32452
rect 47180 31948 47236 32004
rect 46956 31724 47012 31780
rect 46956 30828 47012 30884
rect 46508 29372 46564 29428
rect 45724 28812 45780 28868
rect 46284 28700 46340 28756
rect 45948 28252 46004 28308
rect 45836 27580 45892 27636
rect 46620 28812 46676 28868
rect 46508 28418 46564 28420
rect 46508 28366 46510 28418
rect 46510 28366 46562 28418
rect 46562 28366 46564 28418
rect 46508 28364 46564 28366
rect 46508 27020 46564 27076
rect 46620 28028 46676 28084
rect 45388 26402 45444 26404
rect 45388 26350 45390 26402
rect 45390 26350 45442 26402
rect 45442 26350 45444 26402
rect 45388 26348 45444 26350
rect 45500 26124 45556 26180
rect 46396 26514 46452 26516
rect 46396 26462 46398 26514
rect 46398 26462 46450 26514
rect 46450 26462 46452 26514
rect 46396 26460 46452 26462
rect 45724 25788 45780 25844
rect 45836 26348 45892 26404
rect 47180 29372 47236 29428
rect 46956 28700 47012 28756
rect 46844 28028 46900 28084
rect 46844 27356 46900 27412
rect 47404 32674 47460 32676
rect 47404 32622 47406 32674
rect 47406 32622 47458 32674
rect 47458 32622 47460 32674
rect 47404 32620 47460 32622
rect 47516 32450 47572 32452
rect 47516 32398 47518 32450
rect 47518 32398 47570 32450
rect 47570 32398 47572 32450
rect 47516 32396 47572 32398
rect 47628 32060 47684 32116
rect 48076 32508 48132 32564
rect 48188 32172 48244 32228
rect 48076 31948 48132 32004
rect 48524 37212 48580 37268
rect 48860 38556 48916 38612
rect 49868 39058 49924 39060
rect 49868 39006 49870 39058
rect 49870 39006 49922 39058
rect 49922 39006 49924 39058
rect 49868 39004 49924 39006
rect 50204 41020 50260 41076
rect 51660 42642 51716 42644
rect 51660 42590 51662 42642
rect 51662 42590 51714 42642
rect 51714 42590 51716 42642
rect 51660 42588 51716 42590
rect 51548 42476 51604 42532
rect 51884 41804 51940 41860
rect 51996 42028 52052 42084
rect 50764 41020 50820 41076
rect 51548 41356 51604 41412
rect 52220 41916 52276 41972
rect 52668 42754 52724 42756
rect 52668 42702 52670 42754
rect 52670 42702 52722 42754
rect 52722 42702 52724 42754
rect 52668 42700 52724 42702
rect 52780 42530 52836 42532
rect 52780 42478 52782 42530
rect 52782 42478 52834 42530
rect 52834 42478 52836 42530
rect 52780 42476 52836 42478
rect 53788 42476 53844 42532
rect 53004 42082 53060 42084
rect 53004 42030 53006 42082
rect 53006 42030 53058 42082
rect 53058 42030 53060 42082
rect 53004 42028 53060 42030
rect 52780 41804 52836 41860
rect 52668 41356 52724 41412
rect 52780 40962 52836 40964
rect 52780 40910 52782 40962
rect 52782 40910 52834 40962
rect 52834 40910 52836 40962
rect 52780 40908 52836 40910
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50428 40236 50484 40292
rect 50540 40460 50596 40516
rect 50316 40124 50372 40180
rect 52108 40572 52164 40628
rect 50764 40402 50820 40404
rect 50764 40350 50766 40402
rect 50766 40350 50818 40402
rect 50818 40350 50820 40402
rect 50764 40348 50820 40350
rect 52444 40514 52500 40516
rect 52444 40462 52446 40514
rect 52446 40462 52498 40514
rect 52498 40462 52500 40514
rect 52444 40460 52500 40462
rect 51324 40236 51380 40292
rect 51436 40124 51492 40180
rect 51884 40236 51940 40292
rect 51884 39676 51940 39732
rect 50876 39618 50932 39620
rect 50876 39566 50878 39618
rect 50878 39566 50930 39618
rect 50930 39566 50932 39618
rect 50876 39564 50932 39566
rect 50316 39004 50372 39060
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50428 38668 50484 38724
rect 50988 38668 51044 38724
rect 49868 38220 49924 38276
rect 49644 37436 49700 37492
rect 49084 36370 49140 36372
rect 49084 36318 49086 36370
rect 49086 36318 49138 36370
rect 49138 36318 49140 36370
rect 49084 36316 49140 36318
rect 48636 36258 48692 36260
rect 48636 36206 48638 36258
rect 48638 36206 48690 36258
rect 48690 36206 48692 36258
rect 48636 36204 48692 36206
rect 48524 35868 48580 35924
rect 48748 35980 48804 36036
rect 49308 36258 49364 36260
rect 49308 36206 49310 36258
rect 49310 36206 49362 36258
rect 49362 36206 49364 36258
rect 49308 36204 49364 36206
rect 49196 35756 49252 35812
rect 48860 35420 48916 35476
rect 49420 35644 49476 35700
rect 48412 34914 48468 34916
rect 48412 34862 48414 34914
rect 48414 34862 48466 34914
rect 48466 34862 48468 34914
rect 48412 34860 48468 34862
rect 49084 35196 49140 35252
rect 49532 35532 49588 35588
rect 49420 34636 49476 34692
rect 49084 34076 49140 34132
rect 48860 33404 48916 33460
rect 49196 34412 49252 34468
rect 48860 32562 48916 32564
rect 48860 32510 48862 32562
rect 48862 32510 48914 32562
rect 48914 32510 48916 32562
rect 48860 32508 48916 32510
rect 49532 34188 49588 34244
rect 49532 33628 49588 33684
rect 48300 31500 48356 31556
rect 48412 32284 48468 32340
rect 47516 31218 47572 31220
rect 47516 31166 47518 31218
rect 47518 31166 47570 31218
rect 47570 31166 47572 31218
rect 47516 31164 47572 31166
rect 47516 29650 47572 29652
rect 47516 29598 47518 29650
rect 47518 29598 47570 29650
rect 47570 29598 47572 29650
rect 47516 29596 47572 29598
rect 47292 28476 47348 28532
rect 47852 29314 47908 29316
rect 47852 29262 47854 29314
rect 47854 29262 47906 29314
rect 47906 29262 47908 29314
rect 47852 29260 47908 29262
rect 47628 28252 47684 28308
rect 47740 29036 47796 29092
rect 47628 28082 47684 28084
rect 47628 28030 47630 28082
rect 47630 28030 47682 28082
rect 47682 28030 47684 28082
rect 47628 28028 47684 28030
rect 46956 27580 47012 27636
rect 46844 26402 46900 26404
rect 46844 26350 46846 26402
rect 46846 26350 46898 26402
rect 46898 26350 46900 26402
rect 46844 26348 46900 26350
rect 46284 26290 46340 26292
rect 46284 26238 46286 26290
rect 46286 26238 46338 26290
rect 46338 26238 46340 26290
rect 46284 26236 46340 26238
rect 45500 25564 45556 25620
rect 45052 24780 45108 24836
rect 43708 23154 43764 23156
rect 43708 23102 43710 23154
rect 43710 23102 43762 23154
rect 43762 23102 43764 23154
rect 43708 23100 43764 23102
rect 43484 22370 43540 22372
rect 43484 22318 43486 22370
rect 43486 22318 43538 22370
rect 43538 22318 43540 22370
rect 43484 22316 43540 22318
rect 43596 22764 43652 22820
rect 43372 22092 43428 22148
rect 44268 22652 44324 22708
rect 43708 22204 43764 22260
rect 42364 21644 42420 21700
rect 40908 20748 40964 20804
rect 41244 21532 41300 21588
rect 42140 21586 42196 21588
rect 42140 21534 42142 21586
rect 42142 21534 42194 21586
rect 42194 21534 42196 21586
rect 42140 21532 42196 21534
rect 40348 20130 40404 20132
rect 40348 20078 40350 20130
rect 40350 20078 40402 20130
rect 40402 20078 40404 20130
rect 40348 20076 40404 20078
rect 41132 20130 41188 20132
rect 41132 20078 41134 20130
rect 41134 20078 41186 20130
rect 41186 20078 41188 20130
rect 41132 20076 41188 20078
rect 42252 20914 42308 20916
rect 42252 20862 42254 20914
rect 42254 20862 42306 20914
rect 42306 20862 42308 20914
rect 42252 20860 42308 20862
rect 42140 20802 42196 20804
rect 42140 20750 42142 20802
rect 42142 20750 42194 20802
rect 42194 20750 42196 20802
rect 42140 20748 42196 20750
rect 43148 21586 43204 21588
rect 43148 21534 43150 21586
rect 43150 21534 43202 21586
rect 43202 21534 43204 21586
rect 43148 21532 43204 21534
rect 43036 21474 43092 21476
rect 43036 21422 43038 21474
rect 43038 21422 43090 21474
rect 43090 21422 43092 21474
rect 43036 21420 43092 21422
rect 43372 21474 43428 21476
rect 43372 21422 43374 21474
rect 43374 21422 43426 21474
rect 43426 21422 43428 21474
rect 43372 21420 43428 21422
rect 44828 23996 44884 24052
rect 44716 23266 44772 23268
rect 44716 23214 44718 23266
rect 44718 23214 44770 23266
rect 44770 23214 44772 23266
rect 44716 23212 44772 23214
rect 44940 23938 44996 23940
rect 44940 23886 44942 23938
rect 44942 23886 44994 23938
rect 44994 23886 44996 23938
rect 44940 23884 44996 23886
rect 46060 25788 46116 25844
rect 45948 24556 46004 24612
rect 45388 24220 45444 24276
rect 44940 22652 44996 22708
rect 44716 22092 44772 22148
rect 45164 22316 45220 22372
rect 45276 22652 45332 22708
rect 45276 22204 45332 22260
rect 44380 21698 44436 21700
rect 44380 21646 44382 21698
rect 44382 21646 44434 21698
rect 44434 21646 44436 21698
rect 44380 21644 44436 21646
rect 44156 21474 44212 21476
rect 44156 21422 44158 21474
rect 44158 21422 44210 21474
rect 44210 21422 44212 21474
rect 44156 21420 44212 21422
rect 45276 21474 45332 21476
rect 45276 21422 45278 21474
rect 45278 21422 45330 21474
rect 45330 21422 45332 21474
rect 45276 21420 45332 21422
rect 44492 20860 44548 20916
rect 43932 20748 43988 20804
rect 44940 20802 44996 20804
rect 44940 20750 44942 20802
rect 44942 20750 44994 20802
rect 44994 20750 44996 20802
rect 44940 20748 44996 20750
rect 43260 20578 43316 20580
rect 43260 20526 43262 20578
rect 43262 20526 43314 20578
rect 43314 20526 43316 20578
rect 43260 20524 43316 20526
rect 41804 20076 41860 20132
rect 46732 25618 46788 25620
rect 46732 25566 46734 25618
rect 46734 25566 46786 25618
rect 46786 25566 46788 25618
rect 46732 25564 46788 25566
rect 46620 25340 46676 25396
rect 47516 26348 47572 26404
rect 47852 28476 47908 28532
rect 47852 28082 47908 28084
rect 47852 28030 47854 28082
rect 47854 28030 47906 28082
rect 47906 28030 47908 28082
rect 47852 28028 47908 28030
rect 47740 27132 47796 27188
rect 48076 29538 48132 29540
rect 48076 29486 48078 29538
rect 48078 29486 48130 29538
rect 48130 29486 48132 29538
rect 48076 29484 48132 29486
rect 48188 28588 48244 28644
rect 48972 32002 49028 32004
rect 48972 31950 48974 32002
rect 48974 31950 49026 32002
rect 49026 31950 49028 32002
rect 48972 31948 49028 31950
rect 48860 31666 48916 31668
rect 48860 31614 48862 31666
rect 48862 31614 48914 31666
rect 48914 31614 48916 31666
rect 48860 31612 48916 31614
rect 48636 31052 48692 31108
rect 48972 31554 49028 31556
rect 48972 31502 48974 31554
rect 48974 31502 49026 31554
rect 49026 31502 49028 31554
rect 48972 31500 49028 31502
rect 48860 30994 48916 30996
rect 48860 30942 48862 30994
rect 48862 30942 48914 30994
rect 48914 30942 48916 30994
rect 48860 30940 48916 30942
rect 49420 32620 49476 32676
rect 49756 35196 49812 35252
rect 50876 38274 50932 38276
rect 50876 38222 50878 38274
rect 50878 38222 50930 38274
rect 50930 38222 50932 38274
rect 50876 38220 50932 38222
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 49980 36540 50036 36596
rect 49980 36092 50036 36148
rect 49980 35868 50036 35924
rect 50764 36652 50820 36708
rect 50652 36540 50708 36596
rect 50092 35644 50148 35700
rect 50204 36316 50260 36372
rect 50540 36482 50596 36484
rect 50540 36430 50542 36482
rect 50542 36430 50594 36482
rect 50594 36430 50596 36482
rect 50540 36428 50596 36430
rect 51436 39394 51492 39396
rect 51436 39342 51438 39394
rect 51438 39342 51490 39394
rect 51490 39342 51492 39394
rect 51436 39340 51492 39342
rect 52332 40290 52388 40292
rect 52332 40238 52334 40290
rect 52334 40238 52386 40290
rect 52386 40238 52388 40290
rect 52332 40236 52388 40238
rect 52892 40124 52948 40180
rect 52668 39730 52724 39732
rect 52668 39678 52670 39730
rect 52670 39678 52722 39730
rect 52722 39678 52724 39730
rect 52668 39676 52724 39678
rect 50316 36204 50372 36260
rect 50556 36090 50612 36092
rect 50316 35980 50372 36036
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50876 35868 50932 35924
rect 50652 35698 50708 35700
rect 50652 35646 50654 35698
rect 50654 35646 50706 35698
rect 50706 35646 50708 35698
rect 50652 35644 50708 35646
rect 51100 35532 51156 35588
rect 50652 35420 50708 35476
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50316 34130 50372 34132
rect 50316 34078 50318 34130
rect 50318 34078 50370 34130
rect 50370 34078 50372 34130
rect 50316 34076 50372 34078
rect 50316 33628 50372 33684
rect 49868 32508 49924 32564
rect 49532 32172 49588 32228
rect 49420 31778 49476 31780
rect 49420 31726 49422 31778
rect 49422 31726 49474 31778
rect 49474 31726 49476 31778
rect 49420 31724 49476 31726
rect 49644 32060 49700 32116
rect 49084 31164 49140 31220
rect 49196 31388 49252 31444
rect 48412 27916 48468 27972
rect 47964 26908 48020 26964
rect 47180 26236 47236 26292
rect 47516 25564 47572 25620
rect 46956 25340 47012 25396
rect 47404 25452 47460 25508
rect 47292 25282 47348 25284
rect 47292 25230 47294 25282
rect 47294 25230 47346 25282
rect 47346 25230 47348 25282
rect 47292 25228 47348 25230
rect 46620 24834 46676 24836
rect 46620 24782 46622 24834
rect 46622 24782 46674 24834
rect 46674 24782 46676 24834
rect 46620 24780 46676 24782
rect 47292 24780 47348 24836
rect 46284 24050 46340 24052
rect 46284 23998 46286 24050
rect 46286 23998 46338 24050
rect 46338 23998 46340 24050
rect 46284 23996 46340 23998
rect 46508 23938 46564 23940
rect 46508 23886 46510 23938
rect 46510 23886 46562 23938
rect 46562 23886 46564 23938
rect 46508 23884 46564 23886
rect 46060 23324 46116 23380
rect 46396 23154 46452 23156
rect 46396 23102 46398 23154
rect 46398 23102 46450 23154
rect 46450 23102 46452 23154
rect 46396 23100 46452 23102
rect 45948 22876 46004 22932
rect 46508 22876 46564 22932
rect 46732 22540 46788 22596
rect 47068 24610 47124 24612
rect 47068 24558 47070 24610
rect 47070 24558 47122 24610
rect 47122 24558 47124 24610
rect 47068 24556 47124 24558
rect 47180 24050 47236 24052
rect 47180 23998 47182 24050
rect 47182 23998 47234 24050
rect 47234 23998 47236 24050
rect 47180 23996 47236 23998
rect 47852 25788 47908 25844
rect 47740 25340 47796 25396
rect 48188 26460 48244 26516
rect 47740 24108 47796 24164
rect 47516 23938 47572 23940
rect 47516 23886 47518 23938
rect 47518 23886 47570 23938
rect 47570 23886 47572 23938
rect 47516 23884 47572 23886
rect 47404 23772 47460 23828
rect 47068 23436 47124 23492
rect 46844 22428 46900 22484
rect 47516 23100 47572 23156
rect 47180 22482 47236 22484
rect 47180 22430 47182 22482
rect 47182 22430 47234 22482
rect 47234 22430 47236 22482
rect 47180 22428 47236 22430
rect 46060 22370 46116 22372
rect 46060 22318 46062 22370
rect 46062 22318 46114 22370
rect 46114 22318 46116 22370
rect 46060 22316 46116 22318
rect 47292 22316 47348 22372
rect 47740 23154 47796 23156
rect 47740 23102 47742 23154
rect 47742 23102 47794 23154
rect 47794 23102 47796 23154
rect 47740 23100 47796 23102
rect 48076 24668 48132 24724
rect 48300 23938 48356 23940
rect 48300 23886 48302 23938
rect 48302 23886 48354 23938
rect 48354 23886 48356 23938
rect 48300 23884 48356 23886
rect 48076 23212 48132 23268
rect 48188 23378 48244 23380
rect 48188 23326 48190 23378
rect 48190 23326 48242 23378
rect 48242 23326 48244 23378
rect 48188 23324 48244 23326
rect 48188 23100 48244 23156
rect 48188 22428 48244 22484
rect 47404 22092 47460 22148
rect 47852 21980 47908 22036
rect 47628 21420 47684 21476
rect 49532 31388 49588 31444
rect 49084 30380 49140 30436
rect 48860 30044 48916 30100
rect 49308 29596 49364 29652
rect 49308 28642 49364 28644
rect 49308 28590 49310 28642
rect 49310 28590 49362 28642
rect 49362 28590 49364 28642
rect 49308 28588 49364 28590
rect 49420 27186 49476 27188
rect 49420 27134 49422 27186
rect 49422 27134 49474 27186
rect 49474 27134 49476 27186
rect 49420 27132 49476 27134
rect 48524 25788 48580 25844
rect 48748 26908 48804 26964
rect 48860 26348 48916 26404
rect 49308 26348 49364 26404
rect 49420 26460 49476 26516
rect 49084 26290 49140 26292
rect 49084 26238 49086 26290
rect 49086 26238 49138 26290
rect 49138 26238 49140 26290
rect 49084 26236 49140 26238
rect 49644 31164 49700 31220
rect 49644 29596 49700 29652
rect 49980 31948 50036 32004
rect 51324 34860 51380 34916
rect 51436 34076 51492 34132
rect 52220 38220 52276 38276
rect 52556 36652 52612 36708
rect 51996 36428 52052 36484
rect 53676 41970 53732 41972
rect 53676 41918 53678 41970
rect 53678 41918 53730 41970
rect 53730 41918 53732 41970
rect 53676 41916 53732 41918
rect 53340 40962 53396 40964
rect 53340 40910 53342 40962
rect 53342 40910 53394 40962
rect 53394 40910 53396 40962
rect 53340 40908 53396 40910
rect 53788 40626 53844 40628
rect 53788 40574 53790 40626
rect 53790 40574 53842 40626
rect 53842 40574 53844 40626
rect 53788 40572 53844 40574
rect 53452 40402 53508 40404
rect 53452 40350 53454 40402
rect 53454 40350 53506 40402
rect 53506 40350 53508 40402
rect 53452 40348 53508 40350
rect 54012 40348 54068 40404
rect 54796 40236 54852 40292
rect 54012 38834 54068 38836
rect 54012 38782 54014 38834
rect 54014 38782 54066 38834
rect 54066 38782 54068 38834
rect 54012 38780 54068 38782
rect 55468 38780 55524 38836
rect 55580 39340 55636 39396
rect 53228 38722 53284 38724
rect 53228 38670 53230 38722
rect 53230 38670 53282 38722
rect 53282 38670 53284 38722
rect 53228 38668 53284 38670
rect 53116 37436 53172 37492
rect 52108 35084 52164 35140
rect 52108 34636 52164 34692
rect 51212 33404 51268 33460
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50540 32562 50596 32564
rect 50540 32510 50542 32562
rect 50542 32510 50594 32562
rect 50594 32510 50596 32562
rect 50540 32508 50596 32510
rect 50764 32060 50820 32116
rect 51100 32284 51156 32340
rect 50876 31948 50932 32004
rect 52108 33292 52164 33348
rect 53788 37490 53844 37492
rect 53788 37438 53790 37490
rect 53790 37438 53842 37490
rect 53842 37438 53844 37490
rect 53788 37436 53844 37438
rect 54908 37324 54964 37380
rect 53116 37212 53172 37268
rect 53004 36764 53060 36820
rect 53452 37154 53508 37156
rect 53452 37102 53454 37154
rect 53454 37102 53506 37154
rect 53506 37102 53508 37154
rect 53452 37100 53508 37102
rect 54236 36764 54292 36820
rect 54684 37100 54740 37156
rect 55356 37266 55412 37268
rect 55356 37214 55358 37266
rect 55358 37214 55410 37266
rect 55410 37214 55412 37266
rect 55356 37212 55412 37214
rect 54908 36652 54964 36708
rect 55020 36988 55076 37044
rect 53228 36482 53284 36484
rect 53228 36430 53230 36482
rect 53230 36430 53282 36482
rect 53282 36430 53284 36482
rect 53228 36428 53284 36430
rect 53228 35196 53284 35252
rect 53116 35138 53172 35140
rect 53116 35086 53118 35138
rect 53118 35086 53170 35138
rect 53170 35086 53172 35138
rect 53116 35084 53172 35086
rect 52892 35026 52948 35028
rect 52892 34974 52894 35026
rect 52894 34974 52946 35026
rect 52946 34974 52948 35026
rect 52892 34972 52948 34974
rect 52892 34636 52948 34692
rect 53228 33964 53284 34020
rect 54908 36428 54964 36484
rect 53900 36258 53956 36260
rect 53900 36206 53902 36258
rect 53902 36206 53954 36258
rect 53954 36206 53956 36258
rect 53900 36204 53956 36206
rect 54572 35868 54628 35924
rect 53788 34914 53844 34916
rect 53788 34862 53790 34914
rect 53790 34862 53842 34914
rect 53842 34862 53844 34914
rect 53788 34860 53844 34862
rect 54012 34354 54068 34356
rect 54012 34302 54014 34354
rect 54014 34302 54066 34354
rect 54066 34302 54068 34354
rect 54012 34300 54068 34302
rect 54572 35196 54628 35252
rect 54460 35026 54516 35028
rect 54460 34974 54462 35026
rect 54462 34974 54514 35026
rect 54514 34974 54516 35026
rect 54460 34972 54516 34974
rect 55468 36370 55524 36372
rect 55468 36318 55470 36370
rect 55470 36318 55522 36370
rect 55522 36318 55524 36370
rect 55468 36316 55524 36318
rect 54908 35308 54964 35364
rect 55356 35532 55412 35588
rect 55356 35308 55412 35364
rect 54796 34914 54852 34916
rect 54796 34862 54798 34914
rect 54798 34862 54850 34914
rect 54850 34862 54852 34914
rect 54796 34860 54852 34862
rect 55020 34242 55076 34244
rect 55020 34190 55022 34242
rect 55022 34190 55074 34242
rect 55074 34190 55076 34242
rect 55020 34188 55076 34190
rect 52108 32732 52164 32788
rect 52220 33068 52276 33124
rect 50428 31612 50484 31668
rect 49980 31276 50036 31332
rect 49980 30044 50036 30100
rect 49756 29484 49812 29540
rect 50204 31276 50260 31332
rect 50204 30940 50260 30996
rect 49980 29314 50036 29316
rect 49980 29262 49982 29314
rect 49982 29262 50034 29314
rect 50034 29262 50036 29314
rect 49980 29260 50036 29262
rect 50652 31500 50708 31556
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50988 31276 51044 31332
rect 50988 30940 51044 30996
rect 51100 31164 51156 31220
rect 50540 30828 50596 30884
rect 50652 30268 50708 30324
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50428 29426 50484 29428
rect 50428 29374 50430 29426
rect 50430 29374 50482 29426
rect 50482 29374 50484 29426
rect 50428 29372 50484 29374
rect 50316 28642 50372 28644
rect 50316 28590 50318 28642
rect 50318 28590 50370 28642
rect 50370 28590 50372 28642
rect 50316 28588 50372 28590
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50428 27746 50484 27748
rect 50428 27694 50430 27746
rect 50430 27694 50482 27746
rect 50482 27694 50484 27746
rect 50428 27692 50484 27694
rect 49980 27132 50036 27188
rect 49868 27074 49924 27076
rect 49868 27022 49870 27074
rect 49870 27022 49922 27074
rect 49922 27022 49924 27074
rect 49868 27020 49924 27022
rect 50540 27580 50596 27636
rect 50652 27916 50708 27972
rect 50652 27468 50708 27524
rect 51100 29372 51156 29428
rect 50988 28924 51044 28980
rect 51548 32002 51604 32004
rect 51548 31950 51550 32002
rect 51550 31950 51602 32002
rect 51602 31950 51604 32002
rect 51548 31948 51604 31950
rect 51436 30828 51492 30884
rect 52108 32284 52164 32340
rect 52108 31948 52164 32004
rect 52668 31836 52724 31892
rect 51996 31666 52052 31668
rect 51996 31614 51998 31666
rect 51998 31614 52050 31666
rect 52050 31614 52052 31666
rect 51996 31612 52052 31614
rect 52108 31500 52164 31556
rect 51660 31164 51716 31220
rect 51996 31276 52052 31332
rect 51660 30268 51716 30324
rect 51548 30098 51604 30100
rect 51548 30046 51550 30098
rect 51550 30046 51602 30098
rect 51602 30046 51604 30098
rect 51548 30044 51604 30046
rect 52108 30268 52164 30324
rect 53004 30994 53060 30996
rect 53004 30942 53006 30994
rect 53006 30942 53058 30994
rect 53058 30942 53060 30994
rect 53004 30940 53060 30942
rect 52444 30828 52500 30884
rect 53228 31724 53284 31780
rect 53340 31892 53396 31948
rect 55244 34300 55300 34356
rect 57372 38780 57428 38836
rect 55692 37378 55748 37380
rect 55692 37326 55694 37378
rect 55694 37326 55746 37378
rect 55746 37326 55748 37378
rect 55692 37324 55748 37326
rect 55804 37266 55860 37268
rect 55804 37214 55806 37266
rect 55806 37214 55858 37266
rect 55858 37214 55860 37266
rect 55804 37212 55860 37214
rect 55692 37042 55748 37044
rect 55692 36990 55694 37042
rect 55694 36990 55746 37042
rect 55746 36990 55748 37042
rect 55692 36988 55748 36990
rect 56364 36482 56420 36484
rect 56364 36430 56366 36482
rect 56366 36430 56418 36482
rect 56418 36430 56420 36482
rect 56364 36428 56420 36430
rect 55804 36204 55860 36260
rect 55804 34636 55860 34692
rect 55580 34524 55636 34580
rect 53900 34018 53956 34020
rect 53900 33966 53902 34018
rect 53902 33966 53954 34018
rect 53954 33966 53956 34018
rect 53900 33964 53956 33966
rect 54236 33852 54292 33908
rect 54796 33628 54852 33684
rect 54908 33516 54964 33572
rect 55916 34300 55972 34356
rect 55356 33292 55412 33348
rect 56252 34972 56308 35028
rect 57036 36482 57092 36484
rect 57036 36430 57038 36482
rect 57038 36430 57090 36482
rect 57090 36430 57092 36482
rect 57036 36428 57092 36430
rect 56588 36316 56644 36372
rect 56700 35586 56756 35588
rect 56700 35534 56702 35586
rect 56702 35534 56754 35586
rect 56754 35534 56756 35586
rect 56700 35532 56756 35534
rect 57484 36258 57540 36260
rect 57484 36206 57486 36258
rect 57486 36206 57538 36258
rect 57538 36206 57540 36258
rect 57484 36204 57540 36206
rect 57372 35026 57428 35028
rect 57372 34974 57374 35026
rect 57374 34974 57426 35026
rect 57426 34974 57428 35026
rect 57372 34972 57428 34974
rect 56476 34300 56532 34356
rect 57260 34636 57316 34692
rect 56588 34242 56644 34244
rect 56588 34190 56590 34242
rect 56590 34190 56642 34242
rect 56642 34190 56644 34242
rect 56588 34188 56644 34190
rect 57372 34354 57428 34356
rect 57372 34302 57374 34354
rect 57374 34302 57426 34354
rect 57426 34302 57428 34354
rect 57372 34300 57428 34302
rect 56028 33852 56084 33908
rect 56812 33628 56868 33684
rect 57372 33516 57428 33572
rect 56700 33292 56756 33348
rect 53452 31276 53508 31332
rect 53676 31218 53732 31220
rect 53676 31166 53678 31218
rect 53678 31166 53730 31218
rect 53730 31166 53732 31218
rect 53676 31164 53732 31166
rect 56028 31666 56084 31668
rect 56028 31614 56030 31666
rect 56030 31614 56082 31666
rect 56082 31614 56084 31666
rect 56028 31612 56084 31614
rect 54460 31106 54516 31108
rect 54460 31054 54462 31106
rect 54462 31054 54514 31106
rect 54514 31054 54516 31106
rect 54460 31052 54516 31054
rect 56700 31052 56756 31108
rect 58156 33346 58212 33348
rect 58156 33294 58158 33346
rect 58158 33294 58210 33346
rect 58210 33294 58212 33346
rect 58156 33292 58212 33294
rect 52444 29426 52500 29428
rect 52444 29374 52446 29426
rect 52446 29374 52498 29426
rect 52498 29374 52500 29426
rect 52444 29372 52500 29374
rect 52668 29202 52724 29204
rect 52668 29150 52670 29202
rect 52670 29150 52722 29202
rect 52722 29150 52724 29202
rect 52668 29148 52724 29150
rect 52668 28364 52724 28420
rect 51884 27858 51940 27860
rect 51884 27806 51886 27858
rect 51886 27806 51938 27858
rect 51938 27806 51940 27858
rect 51884 27804 51940 27806
rect 51548 27244 51604 27300
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 49644 26348 49700 26404
rect 49644 26178 49700 26180
rect 49644 26126 49646 26178
rect 49646 26126 49698 26178
rect 49698 26126 49700 26178
rect 49644 26124 49700 26126
rect 49532 25900 49588 25956
rect 49980 26236 50036 26292
rect 50764 26290 50820 26292
rect 50764 26238 50766 26290
rect 50766 26238 50818 26290
rect 50818 26238 50820 26290
rect 50764 26236 50820 26238
rect 50876 26178 50932 26180
rect 50876 26126 50878 26178
rect 50878 26126 50930 26178
rect 50930 26126 50932 26178
rect 50876 26124 50932 26126
rect 50988 26012 51044 26068
rect 52108 28082 52164 28084
rect 52108 28030 52110 28082
rect 52110 28030 52162 28082
rect 52162 28030 52164 28082
rect 52108 28028 52164 28030
rect 50876 25900 50932 25956
rect 50764 25564 50820 25620
rect 49420 25340 49476 25396
rect 48636 25282 48692 25284
rect 48636 25230 48638 25282
rect 48638 25230 48690 25282
rect 48690 25230 48692 25282
rect 48636 25228 48692 25230
rect 48860 25116 48916 25172
rect 49084 25282 49140 25284
rect 49084 25230 49086 25282
rect 49086 25230 49138 25282
rect 49138 25230 49140 25282
rect 49084 25228 49140 25230
rect 48972 24780 49028 24836
rect 49084 24722 49140 24724
rect 49084 24670 49086 24722
rect 49086 24670 49138 24722
rect 49138 24670 49140 24722
rect 49084 24668 49140 24670
rect 48748 24108 48804 24164
rect 48748 22540 48804 22596
rect 49084 23212 49140 23268
rect 49196 23436 49252 23492
rect 48300 22258 48356 22260
rect 48300 22206 48302 22258
rect 48302 22206 48354 22258
rect 48354 22206 48356 22258
rect 48300 22204 48356 22206
rect 48524 22092 48580 22148
rect 49196 22258 49252 22260
rect 49196 22206 49198 22258
rect 49198 22206 49250 22258
rect 49250 22206 49252 22258
rect 49196 22204 49252 22206
rect 49532 23938 49588 23940
rect 49532 23886 49534 23938
rect 49534 23886 49586 23938
rect 49586 23886 49588 23938
rect 49532 23884 49588 23886
rect 51436 26290 51492 26292
rect 51436 26238 51438 26290
rect 51438 26238 51490 26290
rect 51490 26238 51492 26290
rect 51436 26236 51492 26238
rect 52332 27692 52388 27748
rect 52332 27020 52388 27076
rect 53340 30156 53396 30212
rect 53900 30994 53956 30996
rect 53900 30942 53902 30994
rect 53902 30942 53954 30994
rect 53954 30942 53956 30994
rect 53900 30940 53956 30942
rect 54348 30604 54404 30660
rect 53564 30268 53620 30324
rect 53788 30210 53844 30212
rect 53788 30158 53790 30210
rect 53790 30158 53842 30210
rect 53842 30158 53844 30210
rect 53788 30156 53844 30158
rect 53676 29426 53732 29428
rect 53676 29374 53678 29426
rect 53678 29374 53730 29426
rect 53730 29374 53732 29426
rect 53676 29372 53732 29374
rect 53228 28924 53284 28980
rect 52780 27858 52836 27860
rect 52780 27806 52782 27858
rect 52782 27806 52834 27858
rect 52834 27806 52836 27858
rect 52780 27804 52836 27806
rect 52668 27692 52724 27748
rect 51996 25900 52052 25956
rect 52220 26012 52276 26068
rect 51548 25452 51604 25508
rect 52108 25676 52164 25732
rect 52108 25506 52164 25508
rect 52108 25454 52110 25506
rect 52110 25454 52162 25506
rect 52162 25454 52164 25506
rect 52108 25452 52164 25454
rect 51436 25228 51492 25284
rect 52108 25228 52164 25284
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50316 24668 50372 24724
rect 50652 23996 50708 24052
rect 50092 23884 50148 23940
rect 51100 23938 51156 23940
rect 51100 23886 51102 23938
rect 51102 23886 51154 23938
rect 51154 23886 51156 23938
rect 51100 23884 51156 23886
rect 51660 23938 51716 23940
rect 51660 23886 51662 23938
rect 51662 23886 51714 23938
rect 51714 23886 51716 23938
rect 51660 23884 51716 23886
rect 49756 23436 49812 23492
rect 51772 23826 51828 23828
rect 51772 23774 51774 23826
rect 51774 23774 51826 23826
rect 51826 23774 51828 23826
rect 51772 23772 51828 23774
rect 51548 23660 51604 23716
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50876 23324 50932 23380
rect 49644 23212 49700 23268
rect 50428 23266 50484 23268
rect 50428 23214 50430 23266
rect 50430 23214 50482 23266
rect 50482 23214 50484 23266
rect 50428 23212 50484 23214
rect 50092 23154 50148 23156
rect 50092 23102 50094 23154
rect 50094 23102 50146 23154
rect 50146 23102 50148 23154
rect 50092 23100 50148 23102
rect 50092 22652 50148 22708
rect 50428 22482 50484 22484
rect 50428 22430 50430 22482
rect 50430 22430 50482 22482
rect 50482 22430 50484 22482
rect 50428 22428 50484 22430
rect 50876 22764 50932 22820
rect 52668 25506 52724 25508
rect 52668 25454 52670 25506
rect 52670 25454 52722 25506
rect 52722 25454 52724 25506
rect 52668 25452 52724 25454
rect 52556 25340 52612 25396
rect 52332 23324 52388 23380
rect 52444 25228 52500 25284
rect 49308 22092 49364 22148
rect 50876 22204 50932 22260
rect 48860 21980 48916 22036
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 48188 20748 48244 20804
rect 39004 19852 39060 19908
rect 39452 19906 39508 19908
rect 39452 19854 39454 19906
rect 39454 19854 39506 19906
rect 39506 19854 39508 19906
rect 39452 19852 39508 19854
rect 52444 22764 52500 22820
rect 51772 22540 51828 22596
rect 51996 22258 52052 22260
rect 51996 22206 51998 22258
rect 51998 22206 52050 22258
rect 52050 22206 52052 22258
rect 51996 22204 52052 22206
rect 53116 28028 53172 28084
rect 53340 28140 53396 28196
rect 53004 27186 53060 27188
rect 53004 27134 53006 27186
rect 53006 27134 53058 27186
rect 53058 27134 53060 27186
rect 53004 27132 53060 27134
rect 53228 27356 53284 27412
rect 53340 26962 53396 26964
rect 53340 26910 53342 26962
rect 53342 26910 53394 26962
rect 53394 26910 53396 26962
rect 53340 26908 53396 26910
rect 54012 28924 54068 28980
rect 53452 26460 53508 26516
rect 53116 25676 53172 25732
rect 53004 25564 53060 25620
rect 52780 25228 52836 25284
rect 53004 23884 53060 23940
rect 52668 23212 52724 23268
rect 53340 25676 53396 25732
rect 53564 27916 53620 27972
rect 54348 27858 54404 27860
rect 54348 27806 54350 27858
rect 54350 27806 54402 27858
rect 54402 27806 54404 27858
rect 54348 27804 54404 27806
rect 53788 27468 53844 27524
rect 53676 27020 53732 27076
rect 53452 25340 53508 25396
rect 54124 27074 54180 27076
rect 54124 27022 54126 27074
rect 54126 27022 54178 27074
rect 54178 27022 54180 27074
rect 54124 27020 54180 27022
rect 54236 25282 54292 25284
rect 54236 25230 54238 25282
rect 54238 25230 54290 25282
rect 54290 25230 54292 25282
rect 54236 25228 54292 25230
rect 57148 30604 57204 30660
rect 54572 29426 54628 29428
rect 54572 29374 54574 29426
rect 54574 29374 54626 29426
rect 54626 29374 54628 29426
rect 54572 29372 54628 29374
rect 57372 29372 57428 29428
rect 55804 29148 55860 29204
rect 55244 28754 55300 28756
rect 55244 28702 55246 28754
rect 55246 28702 55298 28754
rect 55298 28702 55300 28754
rect 55244 28700 55300 28702
rect 55692 28140 55748 28196
rect 55580 28082 55636 28084
rect 55580 28030 55582 28082
rect 55582 28030 55634 28082
rect 55634 28030 55636 28082
rect 55580 28028 55636 28030
rect 55020 27916 55076 27972
rect 54684 27580 54740 27636
rect 54572 27020 54628 27076
rect 54684 25900 54740 25956
rect 54908 27468 54964 27524
rect 54908 26962 54964 26964
rect 54908 26910 54910 26962
rect 54910 26910 54962 26962
rect 54962 26910 54964 26962
rect 54908 26908 54964 26910
rect 55468 27746 55524 27748
rect 55468 27694 55470 27746
rect 55470 27694 55522 27746
rect 55522 27694 55524 27746
rect 55468 27692 55524 27694
rect 55580 26514 55636 26516
rect 55580 26462 55582 26514
rect 55582 26462 55634 26514
rect 55634 26462 55636 26514
rect 55580 26460 55636 26462
rect 54796 25676 54852 25732
rect 53564 23826 53620 23828
rect 53564 23774 53566 23826
rect 53566 23774 53618 23826
rect 53618 23774 53620 23826
rect 53564 23772 53620 23774
rect 53676 23714 53732 23716
rect 53676 23662 53678 23714
rect 53678 23662 53730 23714
rect 53730 23662 53732 23714
rect 53676 23660 53732 23662
rect 52668 22594 52724 22596
rect 52668 22542 52670 22594
rect 52670 22542 52722 22594
rect 52722 22542 52724 22594
rect 52668 22540 52724 22542
rect 56588 28140 56644 28196
rect 56700 27858 56756 27860
rect 56700 27806 56702 27858
rect 56702 27806 56754 27858
rect 56754 27806 56756 27858
rect 56700 27804 56756 27806
rect 55804 23100 55860 23156
rect 52556 22204 52612 22260
rect 50876 20524 50932 20580
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 37100 17666 37156 17668
rect 37100 17614 37102 17666
rect 37102 17614 37154 17666
rect 37154 17614 37156 17666
rect 37100 17612 37156 17614
rect 38556 17612 38612 17668
rect 36316 15484 36372 15540
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 33068 12908 33124 12964
rect 31500 12684 31556 12740
rect 32060 12572 32116 12628
rect 31724 11788 31780 11844
rect 31948 11676 32004 11732
rect 31724 11228 31780 11284
rect 32508 12290 32564 12292
rect 32508 12238 32510 12290
rect 32510 12238 32562 12290
rect 32562 12238 32564 12290
rect 32508 12236 32564 12238
rect 33852 12908 33908 12964
rect 33740 12572 33796 12628
rect 33852 12290 33908 12292
rect 33852 12238 33854 12290
rect 33854 12238 33906 12290
rect 33906 12238 33908 12290
rect 33852 12236 33908 12238
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35644 13746 35700 13748
rect 35644 13694 35646 13746
rect 35646 13694 35698 13746
rect 35698 13694 35700 13746
rect 35644 13692 35700 13694
rect 37884 15426 37940 15428
rect 37884 15374 37886 15426
rect 37886 15374 37938 15426
rect 37938 15374 37940 15426
rect 37884 15372 37940 15374
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 34188 12012 34244 12068
rect 33516 11618 33572 11620
rect 33516 11566 33518 11618
rect 33518 11566 33570 11618
rect 33570 11566 33572 11618
rect 33516 11564 33572 11566
rect 32060 11282 32116 11284
rect 32060 11230 32062 11282
rect 32062 11230 32114 11282
rect 32114 11230 32116 11282
rect 32060 11228 32116 11230
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34300 11228 34356 11284
rect 36316 12962 36372 12964
rect 36316 12910 36318 12962
rect 36318 12910 36370 12962
rect 36370 12910 36372 12962
rect 36316 12908 36372 12910
rect 35868 12738 35924 12740
rect 35868 12686 35870 12738
rect 35870 12686 35922 12738
rect 35922 12686 35924 12738
rect 35868 12684 35924 12686
rect 38444 12684 38500 12740
rect 35980 12066 36036 12068
rect 35980 12014 35982 12066
rect 35982 12014 36034 12066
rect 36034 12014 36036 12066
rect 35980 12012 36036 12014
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 31388 10332 31444 10388
rect 35756 11282 35812 11284
rect 35756 11230 35758 11282
rect 35758 11230 35810 11282
rect 35810 11230 35812 11282
rect 35756 11228 35812 11230
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 35532 10332 35588 10388
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 29932 8258 29988 8260
rect 29932 8206 29934 8258
rect 29934 8206 29986 8258
rect 29986 8206 29988 8258
rect 29932 8204 29988 8206
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 28252 7586 28308 7588
rect 28252 7534 28254 7586
rect 28254 7534 28306 7586
rect 28306 7534 28308 7586
rect 28252 7532 28308 7534
rect 27244 6748 27300 6804
rect 27468 6860 27524 6916
rect 28588 6802 28644 6804
rect 28588 6750 28590 6802
rect 28590 6750 28642 6802
rect 28642 6750 28644 6802
rect 28588 6748 28644 6750
rect 25340 5234 25396 5236
rect 25340 5182 25342 5234
rect 25342 5182 25394 5234
rect 25394 5182 25396 5234
rect 25340 5180 25396 5182
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 26796 5180 26852 5236
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 32722 57036 32732 57092
rect 32788 57036 34188 57092
rect 34244 57036 34254 57092
rect 35410 57036 35420 57092
rect 35476 57036 37996 57092
rect 38052 57036 38062 57092
rect 41682 57036 41692 57092
rect 41748 57036 43596 57092
rect 43652 57036 43662 57092
rect 34066 56924 34076 56980
rect 34132 56924 36428 56980
rect 36484 56924 36494 56980
rect 39442 56924 39452 56980
rect 39508 56924 42028 56980
rect 42084 56924 42094 56980
rect 40338 56812 40348 56868
rect 40404 56812 42924 56868
rect 42980 56812 42990 56868
rect 38098 56588 38108 56644
rect 38164 56588 40348 56644
rect 40404 56588 40414 56644
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4610 56252 4620 56308
rect 4676 56252 5516 56308
rect 5572 56252 5582 56308
rect 23202 56252 23212 56308
rect 23268 56252 24668 56308
rect 24724 56252 24734 56308
rect 30034 56252 30044 56308
rect 30100 56252 30716 56308
rect 30772 56252 30782 56308
rect 31378 56252 31388 56308
rect 31444 56252 32620 56308
rect 32676 56252 32686 56308
rect 33618 56252 33628 56308
rect 33684 56252 35308 56308
rect 35364 56252 35374 56308
rect 36306 56252 36316 56308
rect 36372 56252 39116 56308
rect 39172 56252 39182 56308
rect 42130 56252 42140 56308
rect 42196 56252 44044 56308
rect 44100 56252 44110 56308
rect 5842 56140 5852 56196
rect 5908 56140 8428 56196
rect 8484 56140 8494 56196
rect 15698 56140 15708 56196
rect 15764 56140 17052 56196
rect 17108 56140 17612 56196
rect 17668 56140 17678 56196
rect 17938 56140 17948 56196
rect 18004 56140 18620 56196
rect 18676 56140 18686 56196
rect 20178 56140 20188 56196
rect 20244 56140 21308 56196
rect 21364 56140 21374 56196
rect 17490 56028 17500 56084
rect 17556 56028 19404 56084
rect 19460 56028 19470 56084
rect 35746 56028 35756 56084
rect 35812 56028 37548 56084
rect 37604 56028 37614 56084
rect 43026 55916 43036 55972
rect 43092 55916 44492 55972
rect 44548 55916 44558 55972
rect 18274 55804 18284 55860
rect 18340 55804 18844 55860
rect 18900 55804 18910 55860
rect 34066 55804 34076 55860
rect 34132 55804 35980 55860
rect 36036 55804 36046 55860
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 16818 55468 16828 55524
rect 16884 55468 17500 55524
rect 17556 55468 18396 55524
rect 18452 55468 18462 55524
rect 24658 55468 24668 55524
rect 24724 55468 26684 55524
rect 26740 55468 26750 55524
rect 16930 55356 16940 55412
rect 16996 55356 18844 55412
rect 18900 55356 19852 55412
rect 19908 55356 19918 55412
rect 19170 55244 19180 55300
rect 19236 55244 21868 55300
rect 21924 55244 21934 55300
rect 25778 55244 25788 55300
rect 25844 55244 27356 55300
rect 27412 55244 29148 55300
rect 29204 55244 30380 55300
rect 30436 55244 30446 55300
rect 16258 55132 16268 55188
rect 16324 55132 16828 55188
rect 16884 55132 19068 55188
rect 19124 55132 19134 55188
rect 34962 55132 34972 55188
rect 35028 55132 36092 55188
rect 36148 55132 36158 55188
rect 41458 55132 41468 55188
rect 41524 55132 42588 55188
rect 42644 55132 42654 55188
rect 19954 55020 19964 55076
rect 20020 55020 21420 55076
rect 21476 55020 22316 55076
rect 22372 55020 22382 55076
rect 42690 55020 42700 55076
rect 42756 55020 43596 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 4050 54796 4060 54852
rect 4116 54796 9100 54852
rect 9156 54796 9166 54852
rect 16594 54684 16604 54740
rect 16660 54684 17724 54740
rect 17780 54684 17790 54740
rect 28242 54684 28252 54740
rect 28308 54684 29148 54740
rect 29204 54684 29214 54740
rect 43652 54628 43708 55076
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 2370 54572 2380 54628
rect 2436 54572 6972 54628
rect 7028 54572 7644 54628
rect 7700 54572 7710 54628
rect 43652 54572 44604 54628
rect 44660 54572 44670 54628
rect 17938 54460 17948 54516
rect 18004 54460 18284 54516
rect 18340 54460 18350 54516
rect 23650 54460 23660 54516
rect 23716 54460 24556 54516
rect 24612 54460 25228 54516
rect 25284 54460 25294 54516
rect 19282 54348 19292 54404
rect 19348 54348 20412 54404
rect 20468 54348 20478 54404
rect 33170 54348 33180 54404
rect 33236 54348 34300 54404
rect 34356 54348 34860 54404
rect 34916 54348 35308 54404
rect 35364 54348 35374 54404
rect 45826 54348 45836 54404
rect 45892 54348 48076 54404
rect 48132 54348 48142 54404
rect 16930 54236 16940 54292
rect 16996 54236 17276 54292
rect 17332 54236 19852 54292
rect 19908 54236 19918 54292
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 17490 53900 17500 53956
rect 17556 53900 18172 53956
rect 18228 53900 18238 53956
rect 9650 53788 9660 53844
rect 9716 53788 11452 53844
rect 11508 53788 11518 53844
rect 18386 53788 18396 53844
rect 18452 53788 20636 53844
rect 20692 53788 20702 53844
rect 33516 53788 38668 53844
rect 38724 53788 38734 53844
rect 50082 53788 50092 53844
rect 50148 53788 51324 53844
rect 51380 53788 51390 53844
rect 3602 53676 3612 53732
rect 3668 53676 4956 53732
rect 5012 53676 5022 53732
rect 5170 53676 5180 53732
rect 5236 53676 6748 53732
rect 6804 53676 6814 53732
rect 12898 53676 12908 53732
rect 12964 53676 13468 53732
rect 13524 53676 13534 53732
rect 17266 53676 17276 53732
rect 17332 53676 18620 53732
rect 18676 53676 18686 53732
rect 30370 53676 30380 53732
rect 30436 53676 31164 53732
rect 31220 53676 32284 53732
rect 32340 53676 33292 53732
rect 33348 53676 33358 53732
rect 33516 53620 33572 53788
rect 42130 53676 42140 53732
rect 42196 53676 44828 53732
rect 44884 53676 45276 53732
rect 45332 53676 45342 53732
rect 10770 53564 10780 53620
rect 10836 53564 14364 53620
rect 14420 53564 14430 53620
rect 19730 53564 19740 53620
rect 19796 53564 20188 53620
rect 20244 53564 20254 53620
rect 23090 53564 23100 53620
rect 23156 53564 23772 53620
rect 23828 53564 23838 53620
rect 28802 53564 28812 53620
rect 28868 53564 33572 53620
rect 19170 53452 19180 53508
rect 19236 53452 19628 53508
rect 19684 53452 19694 53508
rect 20626 53452 20636 53508
rect 20692 53452 21420 53508
rect 21476 53452 21486 53508
rect 22530 53452 22540 53508
rect 22596 53452 22876 53508
rect 22932 53452 24668 53508
rect 24724 53452 25676 53508
rect 25732 53452 25742 53508
rect 35298 53452 35308 53508
rect 35364 53452 38108 53508
rect 38164 53452 38174 53508
rect 38770 53452 38780 53508
rect 38836 53452 40124 53508
rect 40180 53452 40190 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 34738 53228 34748 53284
rect 34804 53228 38444 53284
rect 38500 53228 42028 53284
rect 42084 53228 42094 53284
rect 7522 53116 7532 53172
rect 7588 53116 9996 53172
rect 10052 53116 10062 53172
rect 23874 53116 23884 53172
rect 23940 53116 24108 53172
rect 24164 53116 24174 53172
rect 30706 53116 30716 53172
rect 30772 53116 34636 53172
rect 34692 53116 34702 53172
rect 39666 53116 39676 53172
rect 39732 53116 39742 53172
rect 11554 53004 11564 53060
rect 11620 53004 12796 53060
rect 12852 53004 12862 53060
rect 32498 53004 32508 53060
rect 32564 53004 37212 53060
rect 37268 53004 37278 53060
rect 38658 53004 38668 53060
rect 38724 53004 39116 53060
rect 39172 53004 39182 53060
rect 39676 52948 39732 53116
rect 41234 53004 41244 53060
rect 41300 53004 41916 53060
rect 41972 53004 42588 53060
rect 42644 53004 42654 53060
rect 3826 52892 3836 52948
rect 3892 52892 4620 52948
rect 4676 52892 4686 52948
rect 6514 52892 6524 52948
rect 6580 52892 7532 52948
rect 7588 52892 7598 52948
rect 21858 52892 21868 52948
rect 21924 52892 23548 52948
rect 23604 52892 23614 52948
rect 35522 52892 35532 52948
rect 35588 52892 36092 52948
rect 36148 52892 36158 52948
rect 38770 52892 38780 52948
rect 38836 52892 39732 52948
rect 40226 52892 40236 52948
rect 40292 52892 42252 52948
rect 42308 52892 43596 52948
rect 43652 52892 43662 52948
rect 6738 52780 6748 52836
rect 6804 52780 7420 52836
rect 7476 52780 8316 52836
rect 8372 52780 8382 52836
rect 13010 52780 13020 52836
rect 13076 52780 14252 52836
rect 14308 52780 14318 52836
rect 35074 52780 35084 52836
rect 35140 52780 38668 52836
rect 38724 52780 38734 52836
rect 11666 52668 11676 52724
rect 11732 52668 12460 52724
rect 12516 52668 12526 52724
rect 24434 52668 24444 52724
rect 24500 52668 25228 52724
rect 25284 52668 25294 52724
rect 25554 52668 25564 52724
rect 25620 52668 27356 52724
rect 27412 52668 27422 52724
rect 34850 52668 34860 52724
rect 34916 52668 35308 52724
rect 35364 52668 35374 52724
rect 37650 52668 37660 52724
rect 37716 52668 38780 52724
rect 38836 52668 38846 52724
rect 39004 52612 39060 52892
rect 43362 52780 43372 52836
rect 43428 52780 44044 52836
rect 44100 52780 44110 52836
rect 45938 52668 45948 52724
rect 46004 52668 48748 52724
rect 48804 52668 49980 52724
rect 50036 52668 50046 52724
rect 38892 52556 39060 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 38892 52500 38948 52556
rect 5058 52444 5068 52500
rect 5124 52444 6412 52500
rect 6468 52444 6972 52500
rect 7028 52444 7038 52500
rect 10434 52444 10444 52500
rect 10500 52444 10892 52500
rect 10948 52444 12908 52500
rect 12964 52444 13356 52500
rect 13412 52444 13804 52500
rect 13860 52444 13870 52500
rect 24322 52444 24332 52500
rect 24388 52444 25228 52500
rect 25284 52444 27244 52500
rect 27300 52444 27310 52500
rect 35634 52444 35644 52500
rect 35700 52444 38948 52500
rect 39106 52444 39116 52500
rect 39172 52444 40684 52500
rect 40740 52444 40750 52500
rect 45826 52444 45836 52500
rect 45892 52444 46620 52500
rect 46676 52444 47404 52500
rect 47460 52444 47470 52500
rect 5068 52388 5124 52444
rect 38892 52388 38948 52444
rect 4620 52332 5124 52388
rect 22194 52332 22204 52388
rect 22260 52332 23380 52388
rect 35970 52332 35980 52388
rect 36036 52332 37660 52388
rect 37716 52332 38332 52388
rect 38388 52332 38398 52388
rect 38892 52332 39452 52388
rect 39508 52332 39518 52388
rect 40226 52332 40236 52388
rect 40292 52332 41020 52388
rect 41076 52332 41086 52388
rect 45266 52332 45276 52388
rect 45332 52332 49420 52388
rect 49476 52332 49486 52388
rect 4620 52164 4676 52332
rect 23324 52276 23380 52332
rect 4834 52220 4844 52276
rect 4900 52220 7756 52276
rect 7812 52220 7822 52276
rect 12450 52220 12460 52276
rect 12516 52220 15372 52276
rect 15428 52220 15438 52276
rect 17714 52220 17724 52276
rect 17780 52220 18284 52276
rect 18340 52220 19180 52276
rect 19236 52220 19246 52276
rect 20514 52220 20524 52276
rect 20580 52220 21532 52276
rect 21588 52220 22764 52276
rect 22820 52220 22830 52276
rect 23314 52220 23324 52276
rect 23380 52220 24668 52276
rect 24724 52220 24734 52276
rect 37874 52220 37884 52276
rect 37940 52220 39564 52276
rect 39620 52220 39630 52276
rect 43474 52220 43484 52276
rect 43540 52220 46620 52276
rect 46676 52220 46686 52276
rect 4610 52108 4620 52164
rect 4676 52108 4686 52164
rect 4946 52108 4956 52164
rect 5012 52108 5628 52164
rect 5684 52108 5694 52164
rect 10322 52108 10332 52164
rect 10388 52108 11564 52164
rect 11620 52108 11630 52164
rect 12562 52108 12572 52164
rect 12628 52108 14588 52164
rect 14644 52108 14654 52164
rect 15474 52108 15484 52164
rect 15540 52108 18732 52164
rect 18788 52108 19068 52164
rect 19124 52108 19134 52164
rect 22642 52108 22652 52164
rect 22708 52108 23996 52164
rect 24052 52108 24062 52164
rect 38882 52108 38892 52164
rect 38948 52108 40348 52164
rect 40404 52108 40414 52164
rect 45266 52108 45276 52164
rect 45332 52108 45612 52164
rect 45668 52108 45678 52164
rect 46498 52108 46508 52164
rect 46564 52108 46956 52164
rect 47012 52108 48188 52164
rect 48244 52108 48254 52164
rect 49746 52108 49756 52164
rect 49812 52108 50428 52164
rect 50484 52108 51100 52164
rect 51156 52108 51166 52164
rect 38892 52052 38948 52108
rect 2482 51996 2492 52052
rect 2548 51996 4508 52052
rect 4564 51996 4574 52052
rect 31266 51996 31276 52052
rect 31332 51996 31948 52052
rect 37986 51996 37996 52052
rect 38052 51996 38948 52052
rect 39330 51996 39340 52052
rect 39396 51996 39676 52052
rect 39732 51996 39742 52052
rect 41682 51996 41692 52052
rect 41748 51996 42364 52052
rect 42420 51996 42812 52052
rect 42868 51996 42878 52052
rect 47058 51996 47068 52052
rect 47124 51996 48300 52052
rect 48356 51996 48366 52052
rect 3714 51884 3724 51940
rect 3780 51884 5740 51940
rect 5796 51884 5806 51940
rect 11778 51884 11788 51940
rect 11844 51884 12460 51940
rect 12516 51884 12526 51940
rect 13570 51884 13580 51940
rect 13636 51884 13916 51940
rect 13972 51884 14812 51940
rect 14868 51884 14878 51940
rect 18162 51884 18172 51940
rect 18228 51884 19068 51940
rect 19124 51884 19134 51940
rect 23538 51884 23548 51940
rect 23604 51884 23884 51940
rect 23940 51884 24556 51940
rect 24612 51884 24622 51940
rect 31892 51828 31948 51996
rect 34290 51884 34300 51940
rect 34356 51884 38444 51940
rect 38500 51884 38510 51940
rect 38994 51884 39004 51940
rect 39060 51884 40796 51940
rect 40852 51884 40862 51940
rect 31892 51772 33628 51828
rect 33684 51772 33694 51828
rect 36082 51772 36092 51828
rect 36148 51772 40124 51828
rect 40180 51772 41020 51828
rect 41076 51772 41086 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 22866 51660 22876 51716
rect 22932 51660 24556 51716
rect 24612 51660 24622 51716
rect 35522 51660 35532 51716
rect 35588 51660 35756 51716
rect 35812 51660 38164 51716
rect 38108 51604 38164 51660
rect 34402 51548 34412 51604
rect 34468 51548 35980 51604
rect 36036 51548 36046 51604
rect 38098 51548 38108 51604
rect 38164 51548 39116 51604
rect 39172 51548 39900 51604
rect 39956 51548 39966 51604
rect 40898 51548 40908 51604
rect 40964 51548 41356 51604
rect 41412 51548 43372 51604
rect 43428 51548 43708 51604
rect 43764 51548 43774 51604
rect 43922 51548 43932 51604
rect 43988 51548 44940 51604
rect 44996 51548 45006 51604
rect 46610 51548 46620 51604
rect 46676 51548 46686 51604
rect 49196 51548 51212 51604
rect 51268 51548 51278 51604
rect 46620 51492 46676 51548
rect 15362 51436 15372 51492
rect 15428 51436 17612 51492
rect 17668 51436 18396 51492
rect 18452 51436 19068 51492
rect 19124 51436 19134 51492
rect 22652 51436 23772 51492
rect 23828 51436 23838 51492
rect 33506 51436 33516 51492
rect 33572 51436 33852 51492
rect 33908 51436 39228 51492
rect 39284 51436 39294 51492
rect 39554 51436 39564 51492
rect 39620 51436 40012 51492
rect 40068 51436 42028 51492
rect 42084 51436 42094 51492
rect 43036 51436 46676 51492
rect 22652 51380 22708 51436
rect 43036 51380 43092 51436
rect 49196 51380 49252 51548
rect 50642 51436 50652 51492
rect 50708 51436 53228 51492
rect 53284 51436 53294 51492
rect 15250 51324 15260 51380
rect 15316 51324 15326 51380
rect 15586 51324 15596 51380
rect 15652 51324 16492 51380
rect 16548 51324 16558 51380
rect 16818 51324 16828 51380
rect 16884 51324 18172 51380
rect 18228 51324 18238 51380
rect 22082 51324 22092 51380
rect 22148 51324 22652 51380
rect 22708 51324 22718 51380
rect 23090 51324 23100 51380
rect 23156 51324 23996 51380
rect 24052 51324 24062 51380
rect 31892 51324 34860 51380
rect 34916 51324 34926 51380
rect 35186 51324 35196 51380
rect 35252 51324 36316 51380
rect 36372 51324 36382 51380
rect 37986 51324 37996 51380
rect 38052 51324 38668 51380
rect 38724 51324 39340 51380
rect 39396 51324 39406 51380
rect 40114 51324 40124 51380
rect 40180 51324 43036 51380
rect 43092 51324 43102 51380
rect 46050 51324 46060 51380
rect 46116 51324 47180 51380
rect 47236 51324 47740 51380
rect 47796 51324 47806 51380
rect 48066 51324 48076 51380
rect 48132 51324 48142 51380
rect 49186 51324 49196 51380
rect 49252 51324 49262 51380
rect 50194 51324 50204 51380
rect 50260 51324 50764 51380
rect 50820 51324 50830 51380
rect 15260 51268 15316 51324
rect 31892 51268 31948 51324
rect 8082 51212 8092 51268
rect 8148 51212 8764 51268
rect 8820 51212 9660 51268
rect 9716 51212 9726 51268
rect 13794 51212 13804 51268
rect 13860 51212 14252 51268
rect 14308 51212 16044 51268
rect 16100 51212 16110 51268
rect 18722 51212 18732 51268
rect 18788 51212 19740 51268
rect 19796 51212 19806 51268
rect 20066 51212 20076 51268
rect 20132 51212 21756 51268
rect 21812 51212 21822 51268
rect 29250 51212 29260 51268
rect 29316 51212 31948 51268
rect 33730 51212 33740 51268
rect 33796 51212 33806 51268
rect 34290 51212 34300 51268
rect 34356 51212 37100 51268
rect 37156 51212 37166 51268
rect 38434 51212 38444 51268
rect 38500 51212 38892 51268
rect 38948 51212 43708 51268
rect 33740 51156 33796 51212
rect 43652 51156 43708 51212
rect 48076 51156 48132 51324
rect 49410 51212 49420 51268
rect 49476 51212 51100 51268
rect 51156 51212 51166 51268
rect 51986 51212 51996 51268
rect 52052 51212 55580 51268
rect 55636 51212 55646 51268
rect 4834 51100 4844 51156
rect 4900 51100 5740 51156
rect 5796 51100 6636 51156
rect 6692 51100 6702 51156
rect 12898 51100 12908 51156
rect 12964 51100 13580 51156
rect 13636 51100 13646 51156
rect 14578 51100 14588 51156
rect 14644 51100 16268 51156
rect 16324 51100 16334 51156
rect 16482 51100 16492 51156
rect 16548 51100 18788 51156
rect 19954 51100 19964 51156
rect 20020 51100 22428 51156
rect 22484 51100 22494 51156
rect 24098 51100 24108 51156
rect 24164 51100 24444 51156
rect 24500 51100 24510 51156
rect 26898 51100 26908 51156
rect 26964 51100 33796 51156
rect 34962 51100 34972 51156
rect 35028 51100 36316 51156
rect 36372 51100 36382 51156
rect 38098 51100 38108 51156
rect 38164 51100 39452 51156
rect 39508 51100 39518 51156
rect 43652 51100 43820 51156
rect 43876 51100 43886 51156
rect 48076 51100 50764 51156
rect 50820 51100 50830 51156
rect 18732 51044 18788 51100
rect 16034 50988 16044 51044
rect 16100 50988 17612 51044
rect 17668 50988 17678 51044
rect 18722 50988 18732 51044
rect 18788 50988 18798 51044
rect 21970 50988 21980 51044
rect 22036 50988 23100 51044
rect 23156 50988 23166 51044
rect 37090 50988 37100 51044
rect 37156 50988 38668 51044
rect 38724 50988 38734 51044
rect 39218 50988 39228 51044
rect 39284 50988 39564 51044
rect 39620 50988 39630 51044
rect 40226 50988 40236 51044
rect 40292 50988 42364 51044
rect 42420 50988 42430 51044
rect 43698 50988 43708 51044
rect 43764 50988 44044 51044
rect 44100 50988 45612 51044
rect 45668 50988 45678 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 15026 50876 15036 50932
rect 15092 50876 16604 50932
rect 16660 50876 17948 50932
rect 18004 50876 19740 50932
rect 19796 50876 19806 50932
rect 24098 50876 24108 50932
rect 24164 50876 24556 50932
rect 24612 50876 24622 50932
rect 36530 50876 36540 50932
rect 36596 50876 41132 50932
rect 41188 50876 41198 50932
rect 42588 50876 43596 50932
rect 43652 50876 43662 50932
rect 49746 50876 49756 50932
rect 49812 50876 50316 50932
rect 50372 50876 50382 50932
rect 42588 50820 42644 50876
rect 34626 50764 34636 50820
rect 34692 50764 35980 50820
rect 36036 50764 36046 50820
rect 39330 50764 39340 50820
rect 39396 50764 40124 50820
rect 40180 50764 40190 50820
rect 42466 50764 42476 50820
rect 42532 50764 42644 50820
rect 42700 50764 43820 50820
rect 43876 50764 43886 50820
rect 50754 50764 50764 50820
rect 50820 50764 51996 50820
rect 52052 50764 52062 50820
rect 12450 50652 12460 50708
rect 12516 50652 14476 50708
rect 14532 50652 14542 50708
rect 36082 50652 36092 50708
rect 36148 50652 38332 50708
rect 38388 50652 38398 50708
rect 38882 50652 38892 50708
rect 38948 50652 42140 50708
rect 42196 50652 42476 50708
rect 42532 50652 42542 50708
rect 42700 50596 42756 50764
rect 42914 50652 42924 50708
rect 42980 50652 43708 50708
rect 43922 50652 43932 50708
rect 43988 50652 43998 50708
rect 48514 50652 48524 50708
rect 48580 50652 51660 50708
rect 51716 50652 52108 50708
rect 52164 50652 52668 50708
rect 52724 50652 53900 50708
rect 53956 50652 53966 50708
rect 12114 50540 12124 50596
rect 12180 50540 12796 50596
rect 12852 50540 13468 50596
rect 13524 50540 13534 50596
rect 18386 50540 18396 50596
rect 18452 50540 19292 50596
rect 19348 50540 19358 50596
rect 19506 50540 19516 50596
rect 19572 50540 20188 50596
rect 20244 50540 20254 50596
rect 23314 50540 23324 50596
rect 23380 50540 24332 50596
rect 24388 50540 24398 50596
rect 34738 50540 34748 50596
rect 34804 50540 36428 50596
rect 36484 50540 36494 50596
rect 38994 50540 39004 50596
rect 39060 50540 41916 50596
rect 41972 50540 42756 50596
rect 19292 50484 19348 50540
rect 43652 50484 43708 50652
rect 43932 50484 43988 50652
rect 48402 50540 48412 50596
rect 48468 50540 48748 50596
rect 48804 50540 51884 50596
rect 51940 50540 51950 50596
rect 2482 50428 2492 50484
rect 2548 50428 5628 50484
rect 5684 50428 5694 50484
rect 8866 50428 8876 50484
rect 8932 50428 11900 50484
rect 11956 50428 11966 50484
rect 12124 50428 14924 50484
rect 14980 50428 14990 50484
rect 19292 50428 19628 50484
rect 19684 50428 19694 50484
rect 20738 50428 20748 50484
rect 20804 50428 22204 50484
rect 22260 50428 22270 50484
rect 22418 50428 22428 50484
rect 22484 50428 23436 50484
rect 23492 50428 23502 50484
rect 23874 50428 23884 50484
rect 23940 50428 26236 50484
rect 26292 50428 26302 50484
rect 35858 50428 35868 50484
rect 35924 50428 37660 50484
rect 37716 50428 37726 50484
rect 37874 50428 37884 50484
rect 37940 50428 38780 50484
rect 38836 50428 39676 50484
rect 39732 50428 40124 50484
rect 40180 50428 40190 50484
rect 40450 50428 40460 50484
rect 40516 50428 41580 50484
rect 41636 50428 42028 50484
rect 42084 50428 42094 50484
rect 42242 50428 42252 50484
rect 42308 50428 43428 50484
rect 43652 50428 43988 50484
rect 51538 50428 51548 50484
rect 51604 50428 53452 50484
rect 53508 50428 53518 50484
rect 12124 50372 12180 50428
rect 43372 50372 43428 50428
rect 5730 50316 5740 50372
rect 5796 50316 6076 50372
rect 6132 50316 6860 50372
rect 6916 50316 6926 50372
rect 10994 50316 11004 50372
rect 11060 50316 11788 50372
rect 11844 50316 12180 50372
rect 16818 50316 16828 50372
rect 16884 50316 18508 50372
rect 18564 50316 19180 50372
rect 19236 50316 19246 50372
rect 36978 50316 36988 50372
rect 37044 50316 39452 50372
rect 39508 50316 39518 50372
rect 39890 50316 39900 50372
rect 39956 50316 40236 50372
rect 40292 50316 40302 50372
rect 43362 50316 43372 50372
rect 43428 50316 43438 50372
rect 6178 50204 6188 50260
rect 6244 50204 7196 50260
rect 7252 50204 7262 50260
rect 37426 50204 37436 50260
rect 37492 50204 42476 50260
rect 42532 50204 42542 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 36530 50092 36540 50148
rect 36596 50092 38444 50148
rect 38500 50092 43596 50148
rect 43652 50092 43662 50148
rect 36306 49980 36316 50036
rect 36372 49980 37212 50036
rect 37268 49980 37278 50036
rect 39218 49980 39228 50036
rect 39284 49980 39900 50036
rect 39956 49980 39966 50036
rect 43362 49980 43372 50036
rect 43428 49980 44044 50036
rect 44100 49980 49084 50036
rect 49140 49980 49150 50036
rect 49858 49980 49868 50036
rect 49924 49980 52220 50036
rect 52276 49980 52286 50036
rect 28130 49868 28140 49924
rect 28196 49868 29036 49924
rect 29092 49868 29102 49924
rect 37090 49868 37100 49924
rect 37156 49868 37996 49924
rect 38052 49868 40012 49924
rect 40068 49868 40078 49924
rect 40674 49868 40684 49924
rect 40740 49868 41356 49924
rect 41412 49868 42476 49924
rect 42532 49868 43820 49924
rect 43876 49868 43886 49924
rect 48066 49868 48076 49924
rect 48132 49868 48748 49924
rect 48804 49868 48814 49924
rect 49746 49868 49756 49924
rect 49812 49868 50764 49924
rect 50820 49868 50830 49924
rect 5730 49756 5740 49812
rect 5796 49756 7084 49812
rect 7140 49756 7150 49812
rect 12450 49756 12460 49812
rect 12516 49756 13804 49812
rect 13860 49756 14364 49812
rect 14420 49756 14430 49812
rect 19842 49756 19852 49812
rect 19908 49756 20300 49812
rect 20356 49756 20366 49812
rect 23202 49756 23212 49812
rect 23268 49756 24556 49812
rect 24612 49756 24622 49812
rect 35634 49756 35644 49812
rect 35700 49756 35710 49812
rect 41458 49756 41468 49812
rect 41524 49756 43148 49812
rect 43204 49756 43214 49812
rect 44930 49756 44940 49812
rect 44996 49756 47068 49812
rect 47124 49756 47134 49812
rect 35644 49700 35700 49756
rect 4610 49644 4620 49700
rect 4676 49644 5516 49700
rect 5572 49644 7308 49700
rect 7364 49644 7374 49700
rect 19394 49644 19404 49700
rect 19460 49644 23324 49700
rect 23380 49644 23390 49700
rect 26786 49644 26796 49700
rect 26852 49644 28140 49700
rect 28196 49644 28206 49700
rect 35644 49644 36876 49700
rect 36932 49644 39116 49700
rect 39172 49644 39182 49700
rect 39666 49644 39676 49700
rect 39732 49644 40908 49700
rect 40964 49644 40974 49700
rect 47954 49644 47964 49700
rect 48020 49644 49980 49700
rect 50036 49644 50046 49700
rect 14802 49532 14812 49588
rect 14868 49532 15820 49588
rect 15876 49532 15886 49588
rect 18946 49532 18956 49588
rect 19012 49532 20524 49588
rect 20580 49532 20590 49588
rect 26450 49532 26460 49588
rect 26516 49532 30604 49588
rect 30660 49532 30670 49588
rect 12450 49420 12460 49476
rect 12516 49420 13356 49476
rect 13412 49420 13422 49476
rect 43586 49420 43596 49476
rect 43652 49420 48972 49476
rect 49028 49420 49038 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 12786 49196 12796 49252
rect 12852 49196 14812 49252
rect 14868 49196 19628 49252
rect 19684 49196 19694 49252
rect 21858 49196 21868 49252
rect 21924 49196 23212 49252
rect 23268 49196 23278 49252
rect 24322 49196 24332 49252
rect 24388 49196 29148 49252
rect 29204 49196 29214 49252
rect 39442 49196 39452 49252
rect 39508 49196 40012 49252
rect 40068 49196 42924 49252
rect 42980 49196 42990 49252
rect 48738 49196 48748 49252
rect 48804 49196 51324 49252
rect 51380 49196 51390 49252
rect 8082 49084 8092 49140
rect 8148 49084 11340 49140
rect 11396 49084 12348 49140
rect 12404 49084 12414 49140
rect 12898 49084 12908 49140
rect 12964 49084 18956 49140
rect 19012 49084 19022 49140
rect 21634 49084 21644 49140
rect 21700 49084 26012 49140
rect 26068 49084 27020 49140
rect 27076 49084 27580 49140
rect 27636 49084 27646 49140
rect 46050 49084 46060 49140
rect 46116 49084 50316 49140
rect 50372 49084 50382 49140
rect 6066 48972 6076 49028
rect 6132 48972 6636 49028
rect 6692 48972 6702 49028
rect 12674 48972 12684 49028
rect 12740 48972 13916 49028
rect 13972 48972 16380 49028
rect 16436 48972 16446 49028
rect 16594 48972 16604 49028
rect 16660 48972 16670 49028
rect 17154 48972 17164 49028
rect 17220 48972 18620 49028
rect 18676 48972 20972 49028
rect 21028 48972 21038 49028
rect 23314 48972 23324 49028
rect 23380 48972 23884 49028
rect 23940 48972 23950 49028
rect 25554 48972 25564 49028
rect 25620 48972 27356 49028
rect 27412 48972 27422 49028
rect 28354 48972 28364 49028
rect 28420 48972 29484 49028
rect 29540 48972 30044 49028
rect 30100 48972 30110 49028
rect 36082 48972 36092 49028
rect 36148 48972 37436 49028
rect 37492 48972 37502 49028
rect 43250 48972 43260 49028
rect 43316 48972 50092 49028
rect 50148 48972 50876 49028
rect 50932 48972 50942 49028
rect 16604 48916 16660 48972
rect 6178 48860 6188 48916
rect 6244 48860 7420 48916
rect 7476 48860 7486 48916
rect 12114 48860 12124 48916
rect 12180 48860 16660 48916
rect 20178 48860 20188 48916
rect 20244 48860 21308 48916
rect 21364 48860 21374 48916
rect 22754 48860 22764 48916
rect 22820 48860 23996 48916
rect 24052 48860 24062 48916
rect 26674 48860 26684 48916
rect 26740 48860 27244 48916
rect 27300 48860 27310 48916
rect 28914 48860 28924 48916
rect 28980 48860 33292 48916
rect 33348 48860 33358 48916
rect 38658 48860 38668 48916
rect 38724 48860 39228 48916
rect 39284 48860 41804 48916
rect 41860 48860 41870 48916
rect 50194 48860 50204 48916
rect 50260 48860 50540 48916
rect 50596 48860 50606 48916
rect 27244 48804 27300 48860
rect 4722 48748 4732 48804
rect 4788 48748 6076 48804
rect 6132 48748 7084 48804
rect 7140 48748 7150 48804
rect 13682 48748 13692 48804
rect 13748 48748 16156 48804
rect 16212 48748 16828 48804
rect 16884 48748 16894 48804
rect 20626 48748 20636 48804
rect 20692 48748 21420 48804
rect 21476 48748 21486 48804
rect 23090 48748 23100 48804
rect 23156 48748 23660 48804
rect 23716 48748 23726 48804
rect 27244 48748 29372 48804
rect 29428 48748 29708 48804
rect 29764 48748 29774 48804
rect 38994 48748 39004 48804
rect 39060 48748 42028 48804
rect 42084 48748 42094 48804
rect 49634 48748 49644 48804
rect 49700 48748 50428 48804
rect 50484 48748 51100 48804
rect 51156 48748 51166 48804
rect 1810 48636 1820 48692
rect 1876 48636 5068 48692
rect 5124 48636 5134 48692
rect 27458 48636 27468 48692
rect 27524 48636 27804 48692
rect 27860 48636 27870 48692
rect 48962 48636 48972 48692
rect 49028 48636 49980 48692
rect 50036 48636 50046 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 2818 48524 2828 48580
rect 2884 48524 6972 48580
rect 7028 48524 7038 48580
rect 28690 48524 28700 48580
rect 28756 48524 30716 48580
rect 30772 48524 30782 48580
rect 11330 48412 11340 48468
rect 11396 48412 15148 48468
rect 15204 48412 15214 48468
rect 17490 48412 17500 48468
rect 17556 48412 18508 48468
rect 18564 48412 18574 48468
rect 19506 48412 19516 48468
rect 19572 48412 20412 48468
rect 20468 48412 20478 48468
rect 20626 48412 20636 48468
rect 20692 48412 20860 48468
rect 20916 48412 33740 48468
rect 33796 48412 33806 48468
rect 49186 48412 49196 48468
rect 49252 48412 50540 48468
rect 50596 48412 50606 48468
rect 50866 48412 50876 48468
rect 50932 48412 53452 48468
rect 53508 48412 53518 48468
rect 5394 48300 5404 48356
rect 5460 48300 6300 48356
rect 6356 48300 6366 48356
rect 6626 48300 6636 48356
rect 6692 48300 7756 48356
rect 7812 48300 8428 48356
rect 8484 48300 8494 48356
rect 11666 48300 11676 48356
rect 11732 48300 15596 48356
rect 15652 48300 15662 48356
rect 22530 48300 22540 48356
rect 22596 48300 23436 48356
rect 23492 48300 23502 48356
rect 24658 48300 24668 48356
rect 24724 48300 25788 48356
rect 25844 48300 25854 48356
rect 26852 48300 28700 48356
rect 28756 48300 28766 48356
rect 30258 48300 30268 48356
rect 30324 48300 32060 48356
rect 32116 48300 32126 48356
rect 34514 48300 34524 48356
rect 34580 48300 41356 48356
rect 41412 48300 44492 48356
rect 44548 48300 45388 48356
rect 45444 48300 45454 48356
rect 46386 48300 46396 48356
rect 46452 48300 47068 48356
rect 47124 48300 47852 48356
rect 47908 48300 47918 48356
rect 6514 48188 6524 48244
rect 6580 48188 8316 48244
rect 8372 48188 8382 48244
rect 12226 48188 12236 48244
rect 12292 48188 14700 48244
rect 14756 48188 14766 48244
rect 18610 48188 18620 48244
rect 18676 48188 19964 48244
rect 20020 48188 20030 48244
rect 24322 48188 24332 48244
rect 24388 48188 26012 48244
rect 26068 48188 26078 48244
rect 26012 48132 26068 48188
rect 26852 48132 26908 48300
rect 2930 48076 2940 48132
rect 2996 48076 3836 48132
rect 3892 48076 3902 48132
rect 6402 48076 6412 48132
rect 6468 48076 8092 48132
rect 8148 48076 8158 48132
rect 21298 48076 21308 48132
rect 21364 48076 22428 48132
rect 22484 48076 22494 48132
rect 26012 48076 26908 48132
rect 28242 48076 28252 48132
rect 28308 48076 29036 48132
rect 29092 48076 29102 48132
rect 36306 48076 36316 48132
rect 36372 48076 43596 48132
rect 43652 48076 43662 48132
rect 46162 48076 46172 48132
rect 46228 48076 47404 48132
rect 47460 48076 47470 48132
rect 6962 47964 6972 48020
rect 7028 47964 7980 48020
rect 8036 47964 8046 48020
rect 9986 47964 9996 48020
rect 10052 47964 10668 48020
rect 10724 47964 10734 48020
rect 22642 47964 22652 48020
rect 22708 47964 23548 48020
rect 23604 47964 23614 48020
rect 28130 47964 28140 48020
rect 28196 47964 30268 48020
rect 30324 47964 30334 48020
rect 6626 47852 6636 47908
rect 6692 47852 7308 47908
rect 7364 47852 7374 47908
rect 12674 47852 12684 47908
rect 12740 47852 14140 47908
rect 14196 47852 14588 47908
rect 14644 47852 22316 47908
rect 22372 47852 22382 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 15698 47740 15708 47796
rect 15764 47740 23884 47796
rect 23940 47740 26572 47796
rect 26628 47740 26638 47796
rect 15026 47628 15036 47684
rect 15092 47628 24108 47684
rect 24164 47628 24174 47684
rect 26450 47628 26460 47684
rect 26516 47628 29260 47684
rect 29316 47628 29326 47684
rect 23762 47516 23772 47572
rect 23828 47516 28140 47572
rect 28196 47516 28206 47572
rect 28802 47516 28812 47572
rect 28868 47516 30044 47572
rect 30100 47516 30110 47572
rect 32386 47516 32396 47572
rect 32452 47516 33404 47572
rect 33460 47516 33470 47572
rect 44258 47516 44268 47572
rect 44324 47516 44828 47572
rect 44884 47516 45500 47572
rect 45556 47516 45566 47572
rect 46274 47516 46284 47572
rect 46340 47516 48860 47572
rect 48916 47516 48926 47572
rect 16706 47404 16716 47460
rect 16772 47404 18172 47460
rect 18228 47404 18238 47460
rect 22642 47404 22652 47460
rect 22708 47404 24220 47460
rect 24276 47404 24286 47460
rect 45826 47404 45836 47460
rect 45892 47404 47292 47460
rect 47348 47404 47358 47460
rect 13122 47292 13132 47348
rect 13188 47292 13916 47348
rect 13972 47292 13982 47348
rect 14578 47292 14588 47348
rect 14644 47292 16380 47348
rect 16436 47292 16446 47348
rect 16594 47292 16604 47348
rect 16660 47292 22092 47348
rect 22148 47292 22158 47348
rect 23314 47292 23324 47348
rect 23380 47292 26684 47348
rect 26740 47292 27748 47348
rect 34402 47292 34412 47348
rect 34468 47292 36316 47348
rect 36372 47292 36382 47348
rect 45714 47292 45724 47348
rect 45780 47292 46620 47348
rect 46676 47292 46844 47348
rect 46900 47292 46910 47348
rect 48290 47292 48300 47348
rect 48356 47292 49868 47348
rect 49924 47292 50428 47348
rect 50484 47292 50494 47348
rect 16604 47236 16660 47292
rect 13010 47180 13020 47236
rect 13076 47180 16660 47236
rect 17938 47180 17948 47236
rect 18004 47180 18396 47236
rect 18452 47180 19180 47236
rect 19236 47180 19246 47236
rect 19506 47180 19516 47236
rect 19572 47180 24332 47236
rect 24388 47180 25004 47236
rect 25060 47180 25070 47236
rect 27692 47124 27748 47292
rect 28130 47180 28140 47236
rect 28196 47180 29148 47236
rect 29204 47180 29214 47236
rect 35074 47180 35084 47236
rect 35140 47180 35644 47236
rect 35700 47180 40348 47236
rect 40404 47180 40414 47236
rect 45042 47180 45052 47236
rect 45108 47180 45612 47236
rect 45668 47180 45678 47236
rect 50372 47180 50764 47236
rect 50820 47180 51324 47236
rect 51380 47180 51772 47236
rect 51828 47180 51838 47236
rect 50372 47124 50428 47180
rect 15026 47068 15036 47124
rect 15092 47068 17276 47124
rect 17332 47068 17342 47124
rect 23538 47068 23548 47124
rect 23604 47068 24220 47124
rect 24276 47068 24286 47124
rect 24658 47068 24668 47124
rect 24724 47068 25452 47124
rect 25508 47068 26796 47124
rect 26852 47068 27356 47124
rect 27412 47068 27422 47124
rect 27682 47068 27692 47124
rect 27748 47068 29036 47124
rect 29092 47068 29102 47124
rect 37650 47068 37660 47124
rect 37716 47068 48972 47124
rect 49028 47068 49644 47124
rect 49700 47068 50428 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 12674 46956 12684 47012
rect 12740 46956 13692 47012
rect 13748 46956 13758 47012
rect 25666 46956 25676 47012
rect 25732 46956 26348 47012
rect 26404 46956 26414 47012
rect 26852 46956 27132 47012
rect 27188 46956 27198 47012
rect 29586 46956 29596 47012
rect 29652 46956 30828 47012
rect 30884 46956 30894 47012
rect 47730 46956 47740 47012
rect 47796 46956 48748 47012
rect 48804 46956 49980 47012
rect 50036 46956 50428 47012
rect 26852 46900 26908 46956
rect 50372 46900 50428 46956
rect 12338 46844 12348 46900
rect 12404 46844 13468 46900
rect 13524 46844 13534 46900
rect 13682 46844 13692 46900
rect 13748 46844 26908 46900
rect 28690 46844 28700 46900
rect 28756 46844 29260 46900
rect 29316 46844 30940 46900
rect 30996 46844 31006 46900
rect 42130 46844 42140 46900
rect 42196 46844 45164 46900
rect 45220 46844 45230 46900
rect 50372 46844 50540 46900
rect 50596 46844 50606 46900
rect 2258 46732 2268 46788
rect 2324 46732 3276 46788
rect 3332 46732 4508 46788
rect 4564 46732 4574 46788
rect 11554 46732 11564 46788
rect 11620 46732 13916 46788
rect 13972 46732 13982 46788
rect 20066 46732 20076 46788
rect 20132 46732 22540 46788
rect 22596 46732 23884 46788
rect 23940 46732 23950 46788
rect 25302 46732 25340 46788
rect 25396 46732 25406 46788
rect 26114 46732 26124 46788
rect 26180 46732 26572 46788
rect 26628 46732 26638 46788
rect 1586 46620 1596 46676
rect 1652 46620 2156 46676
rect 2212 46620 4172 46676
rect 4228 46620 4238 46676
rect 12002 46620 12012 46676
rect 12068 46620 14028 46676
rect 14084 46620 14094 46676
rect 15810 46620 15820 46676
rect 15876 46620 16156 46676
rect 16212 46620 16222 46676
rect 18498 46620 18508 46676
rect 18564 46620 21196 46676
rect 21252 46620 21644 46676
rect 21700 46620 21710 46676
rect 22306 46620 22316 46676
rect 22372 46620 24108 46676
rect 24164 46620 25788 46676
rect 25844 46620 25854 46676
rect 11218 46508 11228 46564
rect 11284 46508 11900 46564
rect 11956 46508 13692 46564
rect 13748 46508 13758 46564
rect 14242 46508 14252 46564
rect 14308 46508 17388 46564
rect 17444 46508 17454 46564
rect 17602 46508 17612 46564
rect 17668 46508 23772 46564
rect 23828 46508 23838 46564
rect 24434 46508 24444 46564
rect 24500 46508 26684 46564
rect 26740 46508 27020 46564
rect 27076 46508 27086 46564
rect 10098 46396 10108 46452
rect 10164 46396 13468 46452
rect 13524 46396 13534 46452
rect 13906 46396 13916 46452
rect 13972 46396 15708 46452
rect 15764 46396 15774 46452
rect 16370 46396 16380 46452
rect 16436 46396 24332 46452
rect 24388 46396 25340 46452
rect 25396 46396 26124 46452
rect 26180 46396 26190 46452
rect 26562 46396 26572 46452
rect 26628 46396 27244 46452
rect 27300 46396 27692 46452
rect 27748 46396 27758 46452
rect 28700 46340 28756 46844
rect 30706 46732 30716 46788
rect 30772 46732 32060 46788
rect 32116 46732 32126 46788
rect 46498 46732 46508 46788
rect 46564 46732 47964 46788
rect 48020 46732 48030 46788
rect 31602 46620 31612 46676
rect 31668 46620 32172 46676
rect 32228 46620 33068 46676
rect 33124 46620 33134 46676
rect 35522 46620 35532 46676
rect 35588 46620 44604 46676
rect 44660 46620 44670 46676
rect 44930 46620 44940 46676
rect 44996 46620 46844 46676
rect 46900 46620 46910 46676
rect 47282 46620 47292 46676
rect 47348 46620 48076 46676
rect 48132 46620 48860 46676
rect 48916 46620 48926 46676
rect 49074 46620 49084 46676
rect 49140 46620 51772 46676
rect 51828 46620 51838 46676
rect 45500 46564 45556 46620
rect 29810 46508 29820 46564
rect 29876 46508 31724 46564
rect 31780 46508 31790 46564
rect 38770 46508 38780 46564
rect 38836 46508 44380 46564
rect 44436 46508 45052 46564
rect 45108 46508 45118 46564
rect 45490 46508 45500 46564
rect 45556 46508 45566 46564
rect 41234 46396 41244 46452
rect 41300 46396 41804 46452
rect 41860 46396 41870 46452
rect 45378 46396 45388 46452
rect 45444 46396 47740 46452
rect 47796 46396 47806 46452
rect 10434 46284 10444 46340
rect 10500 46284 11228 46340
rect 11284 46284 11294 46340
rect 22194 46284 22204 46340
rect 22260 46284 23212 46340
rect 23268 46284 28756 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 22418 46172 22428 46228
rect 22484 46172 23100 46228
rect 23156 46172 23166 46228
rect 24546 46172 24556 46228
rect 24612 46172 26908 46228
rect 27794 46172 27804 46228
rect 27860 46172 29820 46228
rect 29876 46172 29886 46228
rect 15362 46060 15372 46116
rect 15428 46060 24444 46116
rect 24500 46060 24510 46116
rect 26852 46004 26908 46172
rect 27122 46060 27132 46116
rect 27188 46060 28140 46116
rect 28196 46060 28206 46116
rect 19394 45948 19404 46004
rect 19460 45948 22428 46004
rect 22484 45948 23436 46004
rect 23492 45948 23502 46004
rect 26852 45948 28028 46004
rect 28084 45948 28094 46004
rect 34738 45948 34748 46004
rect 34804 45948 35644 46004
rect 35700 45948 35710 46004
rect 5394 45836 5404 45892
rect 5460 45836 6972 45892
rect 7028 45836 7038 45892
rect 10994 45836 11004 45892
rect 11060 45836 12124 45892
rect 12180 45836 12572 45892
rect 12628 45836 12638 45892
rect 12786 45836 12796 45892
rect 12852 45836 13580 45892
rect 13636 45836 14812 45892
rect 14868 45836 14878 45892
rect 18610 45836 18620 45892
rect 18676 45836 19068 45892
rect 19124 45836 19134 45892
rect 20290 45836 20300 45892
rect 20356 45836 20748 45892
rect 20804 45836 23548 45892
rect 23604 45836 23614 45892
rect 26450 45836 26460 45892
rect 26516 45836 27356 45892
rect 27412 45836 27804 45892
rect 27860 45836 27870 45892
rect 28466 45836 28476 45892
rect 28532 45836 29260 45892
rect 29316 45836 29326 45892
rect 30034 45836 30044 45892
rect 30100 45836 30604 45892
rect 30660 45836 30670 45892
rect 33058 45836 33068 45892
rect 33124 45836 33852 45892
rect 33908 45836 34524 45892
rect 34580 45836 35532 45892
rect 35588 45836 35598 45892
rect 41570 45836 41580 45892
rect 41636 45836 42588 45892
rect 42644 45836 43036 45892
rect 43092 45836 44940 45892
rect 44996 45836 45006 45892
rect 7186 45724 7196 45780
rect 7252 45724 9772 45780
rect 9828 45724 10556 45780
rect 10612 45724 10622 45780
rect 14466 45724 14476 45780
rect 14532 45724 15708 45780
rect 15764 45724 15774 45780
rect 24546 45724 24556 45780
rect 24612 45724 27916 45780
rect 27972 45724 27982 45780
rect 29698 45724 29708 45780
rect 29764 45724 30828 45780
rect 30884 45724 30894 45780
rect 27132 45668 27188 45724
rect 6850 45612 6860 45668
rect 6916 45612 7644 45668
rect 7700 45612 7710 45668
rect 10770 45612 10780 45668
rect 10836 45612 11564 45668
rect 11620 45612 11788 45668
rect 11844 45612 11854 45668
rect 15362 45612 15372 45668
rect 15428 45612 15820 45668
rect 15876 45612 15886 45668
rect 16034 45612 16044 45668
rect 16100 45612 20748 45668
rect 20804 45612 20814 45668
rect 27122 45612 27132 45668
rect 27188 45612 27198 45668
rect 1698 45500 1708 45556
rect 1764 45500 2604 45556
rect 2660 45500 2670 45556
rect 11218 45500 11228 45556
rect 11284 45500 14700 45556
rect 14756 45500 15036 45556
rect 15092 45500 15102 45556
rect 15250 45500 15260 45556
rect 15316 45500 15354 45556
rect 21634 45500 21644 45556
rect 21700 45500 21756 45556
rect 21812 45500 21822 45556
rect 25190 45500 25228 45556
rect 25284 45500 25294 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 2482 45388 2492 45444
rect 2548 45388 3948 45444
rect 4004 45388 4014 45444
rect 11442 45388 11452 45444
rect 11508 45388 12012 45444
rect 12068 45388 12684 45444
rect 12740 45388 13020 45444
rect 13076 45388 13086 45444
rect 14802 45388 14812 45444
rect 14868 45388 15596 45444
rect 15652 45388 15662 45444
rect 18162 45388 18172 45444
rect 18228 45388 19404 45444
rect 19460 45388 19470 45444
rect 20850 45388 20860 45444
rect 20916 45388 22092 45444
rect 22148 45388 22158 45444
rect 27010 45388 27020 45444
rect 27076 45388 28364 45444
rect 28420 45388 29372 45444
rect 29428 45388 29438 45444
rect 37314 45388 37324 45444
rect 37380 45388 38332 45444
rect 38388 45388 38398 45444
rect 44930 45388 44940 45444
rect 44996 45388 47124 45444
rect 47068 45332 47124 45388
rect 5058 45276 5068 45332
rect 5124 45276 5964 45332
rect 6020 45276 8204 45332
rect 8260 45276 9660 45332
rect 9716 45276 10892 45332
rect 10948 45276 11900 45332
rect 11956 45276 11966 45332
rect 13458 45276 13468 45332
rect 13524 45276 15260 45332
rect 15316 45276 15326 45332
rect 19058 45276 19068 45332
rect 19124 45276 20300 45332
rect 20356 45276 22988 45332
rect 23044 45276 23054 45332
rect 47068 45276 47628 45332
rect 47684 45276 49084 45332
rect 49140 45276 49150 45332
rect 11330 45164 11340 45220
rect 11396 45164 11788 45220
rect 11844 45164 11854 45220
rect 18946 45164 18956 45220
rect 19012 45164 23996 45220
rect 24052 45164 24062 45220
rect 24518 45164 24556 45220
rect 24612 45164 24622 45220
rect 26786 45164 26796 45220
rect 26852 45164 27916 45220
rect 27972 45164 27982 45220
rect 28130 45164 28140 45220
rect 28196 45164 28476 45220
rect 28532 45164 28542 45220
rect 31602 45164 31612 45220
rect 31668 45164 31948 45220
rect 32004 45164 32014 45220
rect 33954 45164 33964 45220
rect 34020 45164 34972 45220
rect 35028 45164 35038 45220
rect 2034 45052 2044 45108
rect 2100 45052 3724 45108
rect 3780 45052 3790 45108
rect 10434 45052 10444 45108
rect 10500 45052 11228 45108
rect 11284 45052 12684 45108
rect 12740 45052 14140 45108
rect 14196 45052 14206 45108
rect 17714 45052 17724 45108
rect 17780 45052 18060 45108
rect 18116 45052 21756 45108
rect 21812 45052 21822 45108
rect 26226 45052 26236 45108
rect 26292 45052 27692 45108
rect 27748 45052 27758 45108
rect 28578 45052 28588 45108
rect 28644 45052 29372 45108
rect 29428 45052 30828 45108
rect 30884 45052 32284 45108
rect 32340 45052 32350 45108
rect 38770 45052 38780 45108
rect 38836 45052 39676 45108
rect 39732 45052 40796 45108
rect 40852 45052 40862 45108
rect 7522 44940 7532 44996
rect 7588 44940 8764 44996
rect 8820 44940 8830 44996
rect 18946 44940 18956 44996
rect 19012 44940 20636 44996
rect 20692 44940 20702 44996
rect 27234 44940 27244 44996
rect 27300 44940 30044 44996
rect 30100 44940 30110 44996
rect 16370 44828 16380 44884
rect 16436 44828 16716 44884
rect 16772 44828 19404 44884
rect 19460 44828 26012 44884
rect 26068 44828 29596 44884
rect 29652 44828 29662 44884
rect 30370 44828 30380 44884
rect 30436 44828 30716 44884
rect 30772 44828 31052 44884
rect 31108 44828 33516 44884
rect 33572 44828 33582 44884
rect 17574 44716 17612 44772
rect 17668 44716 20412 44772
rect 20468 44716 20478 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 17490 44604 17500 44660
rect 17556 44604 18284 44660
rect 18340 44604 18732 44660
rect 18788 44604 18798 44660
rect 19730 44604 19740 44660
rect 19796 44604 20524 44660
rect 20580 44604 20590 44660
rect 22306 44604 22316 44660
rect 22372 44604 22764 44660
rect 22820 44604 22830 44660
rect 23874 44604 23884 44660
rect 23940 44604 28812 44660
rect 28868 44604 28878 44660
rect 29586 44604 29596 44660
rect 29652 44604 33740 44660
rect 33796 44604 33806 44660
rect 2370 44492 2380 44548
rect 2436 44492 3276 44548
rect 3332 44492 4172 44548
rect 4228 44492 4238 44548
rect 15922 44492 15932 44548
rect 15988 44492 32396 44548
rect 32452 44492 32462 44548
rect 33618 44492 33628 44548
rect 33684 44492 34412 44548
rect 34468 44492 34478 44548
rect 4610 44380 4620 44436
rect 4676 44380 5684 44436
rect 12674 44380 12684 44436
rect 12740 44380 13804 44436
rect 13860 44380 13870 44436
rect 15092 44380 17388 44436
rect 17444 44380 17454 44436
rect 18386 44380 18396 44436
rect 18452 44380 19516 44436
rect 19572 44380 19582 44436
rect 22082 44380 22092 44436
rect 22148 44380 23548 44436
rect 23604 44380 23614 44436
rect 23986 44380 23996 44436
rect 24052 44380 25004 44436
rect 25060 44380 25788 44436
rect 25844 44380 25854 44436
rect 27346 44380 27356 44436
rect 27412 44380 30436 44436
rect 30818 44380 30828 44436
rect 30884 44380 31612 44436
rect 31668 44380 31678 44436
rect 34962 44380 34972 44436
rect 35028 44380 44828 44436
rect 44884 44380 44894 44436
rect 5628 44324 5684 44380
rect 15092 44324 15148 44380
rect 3826 44268 3836 44324
rect 3892 44268 4956 44324
rect 5012 44268 5022 44324
rect 5618 44268 5628 44324
rect 5684 44268 6300 44324
rect 6356 44268 6366 44324
rect 12450 44268 12460 44324
rect 12516 44268 14476 44324
rect 14532 44268 15148 44324
rect 15810 44268 15820 44324
rect 15876 44268 16380 44324
rect 16436 44268 16446 44324
rect 18610 44268 18620 44324
rect 18676 44268 19292 44324
rect 19348 44268 24444 44324
rect 24500 44268 24510 44324
rect 24770 44268 24780 44324
rect 24836 44268 27412 44324
rect 24444 44212 24500 44268
rect 27356 44212 27412 44268
rect 30380 44212 30436 44380
rect 30930 44268 30940 44324
rect 30996 44268 31388 44324
rect 31444 44268 31454 44324
rect 40114 44268 40124 44324
rect 40180 44268 41020 44324
rect 41076 44268 41692 44324
rect 41748 44268 42476 44324
rect 42532 44268 42542 44324
rect 3042 44156 3052 44212
rect 3108 44156 4284 44212
rect 4340 44156 5740 44212
rect 5796 44156 5806 44212
rect 16146 44156 16156 44212
rect 16212 44156 21476 44212
rect 24444 44156 27020 44212
rect 27076 44156 27086 44212
rect 27346 44156 27356 44212
rect 27412 44156 27422 44212
rect 30380 44156 31612 44212
rect 31668 44156 32284 44212
rect 32340 44156 32350 44212
rect 33618 44156 33628 44212
rect 33684 44156 38332 44212
rect 38388 44156 40236 44212
rect 40292 44156 40302 44212
rect 41794 44156 41804 44212
rect 41860 44156 42700 44212
rect 42756 44156 42766 44212
rect 21420 44100 21476 44156
rect 10658 44044 10668 44100
rect 10724 44044 13692 44100
rect 13748 44044 13758 44100
rect 14914 44044 14924 44100
rect 14980 44044 15484 44100
rect 15540 44044 15932 44100
rect 15988 44044 15998 44100
rect 16706 44044 16716 44100
rect 16772 44044 18620 44100
rect 18676 44044 18686 44100
rect 21420 44044 26572 44100
rect 26628 44044 29148 44100
rect 29204 44044 30156 44100
rect 30212 44044 30222 44100
rect 37762 44044 37772 44100
rect 37828 44044 38556 44100
rect 38612 44044 39452 44100
rect 39508 44044 39518 44100
rect 40898 44044 40908 44100
rect 40964 44044 41916 44100
rect 41972 44044 41982 44100
rect 4050 43932 4060 43988
rect 4116 43932 4732 43988
rect 4788 43932 4798 43988
rect 21532 43932 28140 43988
rect 28196 43932 28588 43988
rect 28644 43932 29260 43988
rect 29316 43932 29596 43988
rect 29652 43932 29932 43988
rect 29988 43932 29998 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 21532 43876 21588 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 1922 43820 1932 43876
rect 1988 43820 3724 43876
rect 3780 43820 3790 43876
rect 17266 43820 17276 43876
rect 17332 43820 17724 43876
rect 17780 43820 17790 43876
rect 20290 43820 20300 43876
rect 20356 43820 21532 43876
rect 21588 43820 21598 43876
rect 21746 43820 21756 43876
rect 21812 43820 25452 43876
rect 25508 43820 26012 43876
rect 26068 43820 26078 43876
rect 26338 43820 26348 43876
rect 26404 43820 32060 43876
rect 32116 43820 32126 43876
rect 39890 43820 39900 43876
rect 39956 43820 40348 43876
rect 40404 43820 40414 43876
rect 40786 43820 40796 43876
rect 40852 43820 42252 43876
rect 42308 43820 42318 43876
rect 10994 43708 11004 43764
rect 11060 43708 11788 43764
rect 11844 43708 11854 43764
rect 12114 43708 12124 43764
rect 12180 43708 14028 43764
rect 14084 43708 14980 43764
rect 28466 43708 28476 43764
rect 28532 43708 29708 43764
rect 29764 43708 29774 43764
rect 30146 43708 30156 43764
rect 30212 43708 30604 43764
rect 30660 43708 30670 43764
rect 36418 43708 36428 43764
rect 36484 43708 37548 43764
rect 37604 43708 37614 43764
rect 39666 43708 39676 43764
rect 39732 43708 41020 43764
rect 41076 43708 41086 43764
rect 4386 43596 4396 43652
rect 4452 43596 5068 43652
rect 5124 43596 5134 43652
rect 8866 43596 8876 43652
rect 8932 43596 10108 43652
rect 10164 43596 10174 43652
rect 4610 43484 4620 43540
rect 4676 43484 6076 43540
rect 6132 43484 6142 43540
rect 10210 43484 10220 43540
rect 10276 43484 11228 43540
rect 11284 43484 11788 43540
rect 11844 43484 12012 43540
rect 12068 43484 12078 43540
rect 3602 43372 3612 43428
rect 3668 43372 4956 43428
rect 5012 43372 5022 43428
rect 5954 43372 5964 43428
rect 6020 43372 11116 43428
rect 11172 43372 11182 43428
rect 12898 43372 12908 43428
rect 12964 43372 13804 43428
rect 13860 43372 13870 43428
rect 14924 43316 14980 43708
rect 16146 43596 16156 43652
rect 16212 43596 16828 43652
rect 16884 43596 17612 43652
rect 17668 43596 17678 43652
rect 19506 43596 19516 43652
rect 19572 43596 20860 43652
rect 20916 43596 20926 43652
rect 21186 43596 21196 43652
rect 21252 43596 21532 43652
rect 21588 43596 21598 43652
rect 23090 43596 23100 43652
rect 23156 43596 23548 43652
rect 23604 43596 24220 43652
rect 24276 43596 24286 43652
rect 24882 43596 24892 43652
rect 24948 43596 28028 43652
rect 28084 43596 28094 43652
rect 33954 43596 33964 43652
rect 34020 43596 34356 43652
rect 34514 43596 34524 43652
rect 34580 43596 35644 43652
rect 35700 43596 35710 43652
rect 39218 43596 39228 43652
rect 39284 43596 40460 43652
rect 40516 43596 40526 43652
rect 44930 43596 44940 43652
rect 44996 43596 47068 43652
rect 47124 43596 47134 43652
rect 49970 43596 49980 43652
rect 50036 43596 52108 43652
rect 52164 43596 52174 43652
rect 34300 43540 34356 43596
rect 17714 43484 17724 43540
rect 17780 43484 18732 43540
rect 18788 43484 18798 43540
rect 21606 43484 21644 43540
rect 21700 43484 22876 43540
rect 22932 43484 24780 43540
rect 24836 43484 24846 43540
rect 25666 43484 25676 43540
rect 25732 43484 26684 43540
rect 26740 43484 27692 43540
rect 27748 43484 27758 43540
rect 28466 43484 28476 43540
rect 28532 43484 29148 43540
rect 29204 43484 29214 43540
rect 33394 43484 33404 43540
rect 33460 43484 33852 43540
rect 33908 43484 33918 43540
rect 34300 43484 37996 43540
rect 38052 43484 39004 43540
rect 39060 43484 39070 43540
rect 39554 43484 39564 43540
rect 39620 43484 40236 43540
rect 40292 43484 41580 43540
rect 41636 43484 41646 43540
rect 48178 43484 48188 43540
rect 48244 43484 48860 43540
rect 48916 43484 48926 43540
rect 15138 43372 15148 43428
rect 15204 43372 16828 43428
rect 16884 43372 16894 43428
rect 19282 43372 19292 43428
rect 19348 43372 19516 43428
rect 19572 43372 22092 43428
rect 22148 43372 22158 43428
rect 23314 43372 23324 43428
rect 23380 43372 23884 43428
rect 23940 43372 23950 43428
rect 27906 43372 27916 43428
rect 27972 43372 31276 43428
rect 31332 43372 31342 43428
rect 40338 43372 40348 43428
rect 40404 43372 41804 43428
rect 41860 43372 44380 43428
rect 44436 43372 44446 43428
rect 49858 43372 49868 43428
rect 49924 43372 51660 43428
rect 51716 43372 51726 43428
rect 4834 43260 4844 43316
rect 4900 43260 5516 43316
rect 5572 43260 5582 43316
rect 8866 43260 8876 43316
rect 8932 43260 14364 43316
rect 14420 43260 14430 43316
rect 14924 43260 16380 43316
rect 16436 43260 18620 43316
rect 18676 43260 18686 43316
rect 23090 43260 23100 43316
rect 23156 43260 24444 43316
rect 24500 43260 25564 43316
rect 25620 43260 25630 43316
rect 28354 43260 28364 43316
rect 28420 43260 34300 43316
rect 34356 43260 34366 43316
rect 38882 43260 38892 43316
rect 38948 43260 39788 43316
rect 39844 43260 43484 43316
rect 43540 43260 43550 43316
rect 46274 43260 46284 43316
rect 46340 43260 47516 43316
rect 47572 43260 47582 43316
rect 13570 43148 13580 43204
rect 13636 43148 14028 43204
rect 14084 43148 14980 43204
rect 19058 43148 19068 43204
rect 19124 43148 20188 43204
rect 20244 43148 20254 43204
rect 22530 43148 22540 43204
rect 22596 43148 23212 43204
rect 23268 43148 23278 43204
rect 28018 43148 28028 43204
rect 28084 43148 33964 43204
rect 34020 43148 34030 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 14924 43092 14980 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 14914 43036 14924 43092
rect 14980 43036 15372 43092
rect 15428 43036 15438 43092
rect 21522 43036 21532 43092
rect 21588 43036 25116 43092
rect 25172 43036 25182 43092
rect 27570 43036 27580 43092
rect 27636 43036 29820 43092
rect 29876 43036 29886 43092
rect 45602 43036 45612 43092
rect 45668 43036 46396 43092
rect 46452 43036 46462 43092
rect 13570 42924 13580 42980
rect 13636 42924 16380 42980
rect 16436 42924 16446 42980
rect 18162 42924 18172 42980
rect 18228 42924 18508 42980
rect 18564 42924 18574 42980
rect 18722 42924 18732 42980
rect 18788 42924 18826 42980
rect 20178 42924 20188 42980
rect 20244 42924 21308 42980
rect 21364 42924 21374 42980
rect 22978 42924 22988 42980
rect 23044 42924 23772 42980
rect 23828 42924 23838 42980
rect 26002 42924 26012 42980
rect 26068 42924 26796 42980
rect 26852 42924 26862 42980
rect 47730 42924 47740 42980
rect 47796 42924 50540 42980
rect 50596 42924 50606 42980
rect 10994 42812 11004 42868
rect 11060 42812 13020 42868
rect 13076 42812 13086 42868
rect 15698 42812 15708 42868
rect 15764 42812 15932 42868
rect 15988 42812 26348 42868
rect 26404 42812 27356 42868
rect 27412 42812 27422 42868
rect 32386 42812 32396 42868
rect 32452 42812 34188 42868
rect 34244 42812 35420 42868
rect 35476 42812 35486 42868
rect 51986 42812 51996 42868
rect 52052 42812 52062 42868
rect 51996 42756 52052 42812
rect 11330 42700 11340 42756
rect 11396 42700 21308 42756
rect 21364 42700 21374 42756
rect 21858 42700 21868 42756
rect 21924 42700 22316 42756
rect 22372 42700 22382 42756
rect 23874 42700 23884 42756
rect 23940 42700 24556 42756
rect 24612 42700 24668 42756
rect 24724 42700 24734 42756
rect 25302 42700 25340 42756
rect 25396 42700 25406 42756
rect 29922 42700 29932 42756
rect 29988 42700 34524 42756
rect 34580 42700 34590 42756
rect 42242 42700 42252 42756
rect 42308 42700 45500 42756
rect 45556 42700 45566 42756
rect 49074 42700 49084 42756
rect 49140 42700 49868 42756
rect 49924 42700 49934 42756
rect 51996 42700 52668 42756
rect 52724 42700 52734 42756
rect 16482 42588 16492 42644
rect 16548 42588 17276 42644
rect 17332 42588 17342 42644
rect 22418 42588 22428 42644
rect 22484 42588 22764 42644
rect 22820 42588 22830 42644
rect 24434 42588 24444 42644
rect 24500 42588 26124 42644
rect 26180 42588 26190 42644
rect 34850 42588 34860 42644
rect 34916 42588 36988 42644
rect 37044 42588 37054 42644
rect 40114 42588 40124 42644
rect 40180 42588 40908 42644
rect 40964 42588 40974 42644
rect 44594 42588 44604 42644
rect 44660 42588 46060 42644
rect 46116 42588 46126 42644
rect 49298 42588 49308 42644
rect 49364 42588 49756 42644
rect 49812 42588 50988 42644
rect 51044 42588 51660 42644
rect 51716 42588 51726 42644
rect 1810 42476 1820 42532
rect 1876 42476 4956 42532
rect 5012 42476 5022 42532
rect 13794 42476 13804 42532
rect 13860 42476 14476 42532
rect 14532 42476 14542 42532
rect 18722 42476 18732 42532
rect 18788 42476 19852 42532
rect 19908 42476 19918 42532
rect 25452 42420 25508 42588
rect 34402 42476 34412 42532
rect 34468 42476 37212 42532
rect 37268 42476 37278 42532
rect 41122 42476 41132 42532
rect 41188 42476 42476 42532
rect 42532 42476 42542 42532
rect 43362 42476 43372 42532
rect 43428 42476 45052 42532
rect 45108 42476 45118 42532
rect 51538 42476 51548 42532
rect 51604 42476 52780 42532
rect 52836 42476 53788 42532
rect 53844 42476 53854 42532
rect 23426 42364 23436 42420
rect 23492 42364 25228 42420
rect 25284 42364 25294 42420
rect 25442 42364 25452 42420
rect 25508 42364 25518 42420
rect 25890 42364 25900 42420
rect 25956 42364 26908 42420
rect 26964 42364 26974 42420
rect 27122 42364 27132 42420
rect 27188 42364 27916 42420
rect 27972 42364 27982 42420
rect 31154 42364 31164 42420
rect 31220 42364 32172 42420
rect 32228 42364 35084 42420
rect 35140 42364 35150 42420
rect 35868 42364 45276 42420
rect 45332 42364 45342 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 35868 42308 35924 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 10210 42252 10220 42308
rect 10276 42252 13468 42308
rect 13524 42252 13534 42308
rect 17602 42252 17612 42308
rect 17668 42252 18396 42308
rect 18452 42252 18462 42308
rect 19366 42252 19404 42308
rect 19460 42252 19470 42308
rect 21298 42252 21308 42308
rect 21364 42252 33964 42308
rect 34020 42252 35868 42308
rect 35924 42252 35934 42308
rect 36530 42252 36540 42308
rect 36596 42252 37100 42308
rect 37156 42252 37166 42308
rect 38658 42252 38668 42308
rect 38724 42252 47404 42308
rect 47460 42252 48748 42308
rect 48804 42252 48814 42308
rect 8978 42140 8988 42196
rect 9044 42140 12908 42196
rect 12964 42140 12974 42196
rect 14466 42140 14476 42196
rect 14532 42140 15260 42196
rect 15316 42140 15326 42196
rect 16818 42140 16828 42196
rect 16884 42140 20748 42196
rect 20804 42140 20814 42196
rect 21634 42140 21644 42196
rect 21700 42140 22652 42196
rect 22708 42140 24108 42196
rect 24164 42140 24174 42196
rect 26786 42140 26796 42196
rect 26852 42140 31388 42196
rect 31444 42140 31454 42196
rect 31938 42140 31948 42196
rect 32004 42140 32620 42196
rect 32676 42140 34972 42196
rect 35028 42140 35038 42196
rect 35410 42140 35420 42196
rect 35476 42140 37212 42196
rect 37268 42140 37278 42196
rect 21644 42084 21700 42140
rect 4946 42028 4956 42084
rect 5012 42028 6076 42084
rect 6132 42028 6142 42084
rect 18060 42028 19180 42084
rect 19236 42028 19246 42084
rect 20626 42028 20636 42084
rect 20692 42028 21700 42084
rect 21942 42028 21980 42084
rect 22036 42028 22046 42084
rect 24322 42028 24332 42084
rect 24388 42028 25340 42084
rect 25396 42028 25406 42084
rect 28354 42028 28364 42084
rect 28420 42028 29036 42084
rect 29092 42028 29102 42084
rect 33282 42028 33292 42084
rect 33348 42028 33516 42084
rect 33572 42028 34300 42084
rect 34356 42028 34366 42084
rect 34514 42028 34524 42084
rect 34580 42028 35756 42084
rect 35812 42028 35822 42084
rect 51986 42028 51996 42084
rect 52052 42028 53004 42084
rect 53060 42028 53070 42084
rect 18060 41972 18116 42028
rect 6850 41916 6860 41972
rect 6916 41916 8428 41972
rect 8484 41916 8876 41972
rect 8932 41916 9660 41972
rect 9716 41916 15708 41972
rect 15764 41916 15774 41972
rect 16706 41916 16716 41972
rect 16772 41916 17500 41972
rect 17556 41916 17566 41972
rect 18050 41916 18060 41972
rect 18116 41916 18126 41972
rect 18386 41916 18396 41972
rect 18452 41916 19460 41972
rect 20290 41916 20300 41972
rect 20356 41916 21196 41972
rect 21252 41916 21262 41972
rect 22082 41916 22092 41972
rect 22148 41916 23436 41972
rect 23492 41916 23502 41972
rect 24434 41916 24444 41972
rect 24500 41916 25788 41972
rect 25844 41916 25854 41972
rect 26898 41916 26908 41972
rect 26964 41916 27692 41972
rect 27748 41916 27758 41972
rect 29362 41916 29372 41972
rect 29428 41916 31724 41972
rect 31780 41916 31790 41972
rect 32498 41916 32508 41972
rect 32564 41916 32574 41972
rect 35186 41916 35196 41972
rect 35252 41916 38444 41972
rect 38500 41916 39676 41972
rect 39732 41916 39742 41972
rect 52210 41916 52220 41972
rect 52276 41916 53676 41972
rect 53732 41916 53742 41972
rect 19404 41860 19460 41916
rect 32508 41860 32564 41916
rect 3938 41804 3948 41860
rect 4004 41804 4172 41860
rect 4228 41804 4956 41860
rect 5012 41804 5964 41860
rect 6020 41804 6030 41860
rect 11554 41804 11564 41860
rect 11620 41804 12236 41860
rect 12292 41804 12572 41860
rect 12628 41804 12638 41860
rect 13794 41804 13804 41860
rect 13860 41804 14700 41860
rect 14756 41804 14766 41860
rect 17014 41804 17052 41860
rect 17108 41804 17118 41860
rect 17938 41804 17948 41860
rect 18004 41804 18844 41860
rect 18900 41804 18910 41860
rect 19394 41804 19404 41860
rect 19460 41804 19470 41860
rect 23874 41804 23884 41860
rect 23940 41804 26348 41860
rect 26404 41804 26414 41860
rect 26852 41804 32564 41860
rect 46722 41804 46732 41860
rect 46788 41804 49420 41860
rect 49476 41804 51884 41860
rect 51940 41804 52780 41860
rect 52836 41804 52846 41860
rect 26852 41748 26908 41804
rect 3826 41692 3836 41748
rect 3892 41692 4620 41748
rect 4676 41692 4686 41748
rect 13010 41692 13020 41748
rect 13076 41692 14812 41748
rect 14868 41692 14878 41748
rect 15362 41692 15372 41748
rect 15428 41692 16044 41748
rect 16100 41692 16110 41748
rect 16482 41692 16492 41748
rect 16548 41692 17612 41748
rect 17668 41692 17678 41748
rect 23090 41692 23100 41748
rect 23156 41692 26908 41748
rect 28578 41692 28588 41748
rect 28644 41692 29596 41748
rect 29652 41692 29662 41748
rect 34850 41692 34860 41748
rect 34916 41692 39564 41748
rect 39620 41692 39630 41748
rect 41794 41692 41804 41748
rect 41860 41692 43372 41748
rect 43428 41692 43438 41748
rect 39564 41636 39620 41692
rect 16258 41580 16268 41636
rect 16324 41580 17388 41636
rect 17444 41580 18284 41636
rect 18340 41580 18350 41636
rect 18722 41580 18732 41636
rect 18788 41580 18956 41636
rect 19012 41580 26124 41636
rect 26180 41580 26190 41636
rect 39564 41580 47740 41636
rect 47796 41580 49756 41636
rect 49812 41580 49822 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 16930 41468 16940 41524
rect 16996 41468 17724 41524
rect 17780 41468 17790 41524
rect 21970 41468 21980 41524
rect 22036 41468 22092 41524
rect 22148 41468 22158 41524
rect 23314 41468 23324 41524
rect 23380 41468 29148 41524
rect 29204 41468 30268 41524
rect 30324 41468 30334 41524
rect 38098 41468 38108 41524
rect 38164 41468 45724 41524
rect 45780 41468 45790 41524
rect 5282 41356 5292 41412
rect 5348 41356 6076 41412
rect 6132 41356 6860 41412
rect 6916 41356 6926 41412
rect 17042 41356 17052 41412
rect 17108 41356 17388 41412
rect 17444 41356 18284 41412
rect 18340 41356 18350 41412
rect 19394 41356 19404 41412
rect 19460 41356 20748 41412
rect 20804 41356 20814 41412
rect 22194 41356 22204 41412
rect 22260 41356 22876 41412
rect 22932 41356 22942 41412
rect 24518 41356 24556 41412
rect 24612 41356 24622 41412
rect 25218 41356 25228 41412
rect 25284 41356 25900 41412
rect 25956 41356 25966 41412
rect 26786 41356 26796 41412
rect 26852 41356 29372 41412
rect 29428 41356 29438 41412
rect 51538 41356 51548 41412
rect 51604 41356 52668 41412
rect 52724 41356 52734 41412
rect 4834 41244 4844 41300
rect 4900 41244 5516 41300
rect 5572 41244 7084 41300
rect 7140 41244 7150 41300
rect 14214 41244 14252 41300
rect 14308 41244 14318 41300
rect 14802 41244 14812 41300
rect 14868 41244 23884 41300
rect 23940 41244 23950 41300
rect 26002 41244 26012 41300
rect 26068 41244 28588 41300
rect 28644 41244 28654 41300
rect 34850 41244 34860 41300
rect 34916 41244 39228 41300
rect 39284 41244 39788 41300
rect 39844 41244 39854 41300
rect 43474 41244 43484 41300
rect 43540 41244 44156 41300
rect 44212 41244 44222 41300
rect 39788 41188 39844 41244
rect 4246 41132 4284 41188
rect 4340 41132 4732 41188
rect 4788 41132 4798 41188
rect 6178 41132 6188 41188
rect 6244 41132 6972 41188
rect 7028 41132 7038 41188
rect 14130 41132 14140 41188
rect 14196 41132 14588 41188
rect 14644 41132 14654 41188
rect 16034 41132 16044 41188
rect 16100 41132 16492 41188
rect 16548 41132 16558 41188
rect 17052 41132 22092 41188
rect 22148 41132 23100 41188
rect 23156 41132 23166 41188
rect 23986 41132 23996 41188
rect 24052 41132 24668 41188
rect 24724 41132 25676 41188
rect 25732 41132 25742 41188
rect 26338 41132 26348 41188
rect 26404 41132 29148 41188
rect 29204 41132 29214 41188
rect 29810 41132 29820 41188
rect 29876 41132 30604 41188
rect 30660 41132 30670 41188
rect 39788 41132 48972 41188
rect 49028 41132 50316 41188
rect 50372 41132 50382 41188
rect 17052 41076 17108 41132
rect 14018 41020 14028 41076
rect 14084 41020 17108 41076
rect 17238 41020 17276 41076
rect 17332 41020 18956 41076
rect 19012 41020 19022 41076
rect 20178 41020 20188 41076
rect 20244 41020 20412 41076
rect 20468 41020 20478 41076
rect 28466 41020 28476 41076
rect 28532 41020 35756 41076
rect 35812 41020 35822 41076
rect 36418 41020 36428 41076
rect 36484 41020 37100 41076
rect 37156 41020 37166 41076
rect 41570 41020 41580 41076
rect 41636 41020 44268 41076
rect 44324 41020 44334 41076
rect 49980 40964 50036 41132
rect 50194 41020 50204 41076
rect 50260 41020 50764 41076
rect 50820 41020 50830 41076
rect 3602 40908 3612 40964
rect 3668 40908 4172 40964
rect 4228 40908 4238 40964
rect 13234 40908 13244 40964
rect 13300 40908 16380 40964
rect 16436 40908 16446 40964
rect 17042 40908 17052 40964
rect 17108 40908 17388 40964
rect 17444 40908 17454 40964
rect 17938 40908 17948 40964
rect 18004 40908 18284 40964
rect 18340 40908 18350 40964
rect 19142 40908 19180 40964
rect 19236 40908 19246 40964
rect 19628 40908 21868 40964
rect 21924 40908 22316 40964
rect 22372 40908 22382 40964
rect 23426 40908 23436 40964
rect 23492 40908 24668 40964
rect 24724 40908 24734 40964
rect 27580 40908 28364 40964
rect 28420 40908 29372 40964
rect 29428 40908 29438 40964
rect 31826 40908 31836 40964
rect 31892 40908 36204 40964
rect 36260 40908 36270 40964
rect 37202 40908 37212 40964
rect 37268 40908 39452 40964
rect 39508 40908 39518 40964
rect 39666 40908 39676 40964
rect 39732 40908 41692 40964
rect 41748 40908 42588 40964
rect 42644 40908 42654 40964
rect 49980 40908 52780 40964
rect 52836 40908 53340 40964
rect 53396 40908 53406 40964
rect 19628 40852 19684 40908
rect 27580 40852 27636 40908
rect 16930 40796 16940 40852
rect 16996 40796 19628 40852
rect 19684 40796 19694 40852
rect 20290 40796 20300 40852
rect 20356 40796 21980 40852
rect 22036 40796 22046 40852
rect 27570 40796 27580 40852
rect 27636 40796 27646 40852
rect 31714 40796 31724 40852
rect 31780 40796 37436 40852
rect 37492 40796 38108 40852
rect 38164 40796 38174 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 13458 40684 13468 40740
rect 13524 40684 13916 40740
rect 13972 40684 19684 40740
rect 20738 40684 20748 40740
rect 20804 40684 27244 40740
rect 27300 40684 28028 40740
rect 28084 40684 28094 40740
rect 45266 40684 45276 40740
rect 45332 40684 46844 40740
rect 46900 40684 47404 40740
rect 47460 40684 47470 40740
rect 2482 40572 2492 40628
rect 2548 40572 4508 40628
rect 4564 40572 4574 40628
rect 8530 40572 8540 40628
rect 8596 40572 11340 40628
rect 11396 40572 11406 40628
rect 14802 40572 14812 40628
rect 14868 40572 15932 40628
rect 15988 40572 15998 40628
rect 17602 40572 17612 40628
rect 17668 40572 18620 40628
rect 18676 40572 18686 40628
rect 19628 40516 19684 40684
rect 20850 40572 20860 40628
rect 20916 40572 21868 40628
rect 21924 40572 23100 40628
rect 23156 40572 23166 40628
rect 25778 40572 25788 40628
rect 25844 40572 26572 40628
rect 26628 40572 26638 40628
rect 28354 40572 28364 40628
rect 28420 40572 29036 40628
rect 29092 40572 29102 40628
rect 29810 40572 29820 40628
rect 29876 40572 30268 40628
rect 30324 40572 30334 40628
rect 31602 40572 31612 40628
rect 31668 40572 34524 40628
rect 34580 40572 34590 40628
rect 41906 40572 41916 40628
rect 41972 40572 45164 40628
rect 45220 40572 46508 40628
rect 46564 40572 46574 40628
rect 49410 40572 49420 40628
rect 49476 40572 52108 40628
rect 52164 40572 53788 40628
rect 53844 40572 53854 40628
rect 6514 40460 6524 40516
rect 6580 40460 7644 40516
rect 7700 40460 7710 40516
rect 12002 40460 12012 40516
rect 12068 40460 17948 40516
rect 18004 40460 18014 40516
rect 19628 40460 25060 40516
rect 27878 40460 27916 40516
rect 27972 40460 27982 40516
rect 42802 40460 42812 40516
rect 42868 40460 44268 40516
rect 44324 40460 44334 40516
rect 44930 40460 44940 40516
rect 44996 40460 45006 40516
rect 50530 40460 50540 40516
rect 50596 40460 52444 40516
rect 52500 40460 52510 40516
rect 25004 40404 25060 40460
rect 44940 40404 44996 40460
rect 4834 40348 4844 40404
rect 4900 40348 5852 40404
rect 5908 40348 6412 40404
rect 6468 40348 6478 40404
rect 9426 40348 9436 40404
rect 9492 40348 13580 40404
rect 13636 40348 13646 40404
rect 13906 40348 13916 40404
rect 13972 40348 14588 40404
rect 14644 40348 14654 40404
rect 14914 40348 14924 40404
rect 14980 40348 15148 40404
rect 15204 40348 15988 40404
rect 16258 40348 16268 40404
rect 16324 40348 16716 40404
rect 16772 40348 16782 40404
rect 19170 40348 19180 40404
rect 19236 40348 19964 40404
rect 20020 40348 20972 40404
rect 21028 40348 21038 40404
rect 21522 40348 21532 40404
rect 21588 40348 22540 40404
rect 22596 40348 22606 40404
rect 24994 40348 25004 40404
rect 25060 40348 25070 40404
rect 25554 40348 25564 40404
rect 25620 40348 26348 40404
rect 26404 40348 26908 40404
rect 27458 40348 27468 40404
rect 27524 40348 28700 40404
rect 28756 40348 28766 40404
rect 37762 40348 37772 40404
rect 37828 40348 38780 40404
rect 38836 40348 41468 40404
rect 41524 40348 41534 40404
rect 42130 40348 42140 40404
rect 42196 40348 42700 40404
rect 42756 40348 42766 40404
rect 43026 40348 43036 40404
rect 43092 40348 44996 40404
rect 48066 40348 48076 40404
rect 48132 40348 49196 40404
rect 49252 40348 49262 40404
rect 50754 40348 50764 40404
rect 50820 40348 53452 40404
rect 53508 40348 54012 40404
rect 54068 40348 54078 40404
rect 15932 40292 15988 40348
rect 26852 40292 26908 40348
rect 14242 40236 14252 40292
rect 14308 40236 15036 40292
rect 15092 40236 15102 40292
rect 15922 40236 15932 40292
rect 15988 40236 19404 40292
rect 19460 40236 22092 40292
rect 22148 40236 22158 40292
rect 23314 40236 23324 40292
rect 23380 40236 24556 40292
rect 24612 40236 24622 40292
rect 26852 40236 27356 40292
rect 27412 40236 27422 40292
rect 43138 40236 43148 40292
rect 43204 40236 44492 40292
rect 44548 40236 44558 40292
rect 50418 40236 50428 40292
rect 50484 40236 51324 40292
rect 51380 40236 51884 40292
rect 51940 40236 51950 40292
rect 52322 40236 52332 40292
rect 52388 40236 54796 40292
rect 54852 40236 54862 40292
rect 4610 40124 4620 40180
rect 4676 40124 6076 40180
rect 6132 40124 6142 40180
rect 12674 40124 12684 40180
rect 12740 40124 14588 40180
rect 14644 40124 19404 40180
rect 19460 40124 19628 40180
rect 19684 40124 19694 40180
rect 23986 40124 23996 40180
rect 24052 40124 25452 40180
rect 25508 40124 26236 40180
rect 26292 40124 26796 40180
rect 26852 40124 26862 40180
rect 28466 40124 28476 40180
rect 28532 40124 33740 40180
rect 33796 40124 33806 40180
rect 40002 40124 40012 40180
rect 40068 40124 43260 40180
rect 43316 40124 43326 40180
rect 43922 40124 43932 40180
rect 43988 40124 45612 40180
rect 45668 40124 47404 40180
rect 47460 40124 47470 40180
rect 49970 40124 49980 40180
rect 50036 40124 50316 40180
rect 50372 40124 51436 40180
rect 51492 40124 52892 40180
rect 52948 40124 52958 40180
rect 17042 40012 17052 40068
rect 17108 40012 17612 40068
rect 17668 40012 17678 40068
rect 17938 40012 17948 40068
rect 18004 40012 20860 40068
rect 20916 40012 20926 40068
rect 23874 40012 23884 40068
rect 23940 40012 33068 40068
rect 33124 40012 33134 40068
rect 36306 40012 36316 40068
rect 36372 40012 37772 40068
rect 37828 40012 37838 40068
rect 42914 40012 42924 40068
rect 42980 40012 45724 40068
rect 45780 40012 46172 40068
rect 46228 40012 46238 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 16258 39900 16268 39956
rect 16324 39900 18396 39956
rect 18452 39900 30492 39956
rect 30548 39900 30558 39956
rect 17938 39788 17948 39844
rect 18004 39788 18284 39844
rect 18340 39788 21196 39844
rect 21252 39788 21262 39844
rect 25442 39788 25452 39844
rect 25508 39788 27020 39844
rect 27076 39788 28252 39844
rect 28308 39788 28318 39844
rect 4610 39676 4620 39732
rect 4676 39676 4956 39732
rect 5012 39676 5516 39732
rect 5572 39676 5582 39732
rect 11554 39676 11564 39732
rect 11620 39676 12348 39732
rect 12404 39676 12414 39732
rect 18386 39676 18396 39732
rect 18452 39676 19292 39732
rect 19348 39676 19358 39732
rect 21522 39676 21532 39732
rect 21588 39676 21598 39732
rect 26338 39676 26348 39732
rect 26404 39676 31724 39732
rect 31780 39676 31790 39732
rect 51874 39676 51884 39732
rect 51940 39676 52668 39732
rect 52724 39676 52734 39732
rect 21532 39620 21588 39676
rect 3938 39564 3948 39620
rect 4004 39564 6636 39620
rect 6692 39564 7196 39620
rect 7252 39564 7262 39620
rect 14214 39564 14252 39620
rect 14308 39564 14318 39620
rect 14914 39564 14924 39620
rect 14980 39564 16156 39620
rect 16212 39564 16222 39620
rect 19058 39564 19068 39620
rect 19124 39564 19628 39620
rect 19684 39564 19694 39620
rect 20738 39564 20748 39620
rect 20804 39564 22988 39620
rect 23044 39564 25228 39620
rect 25284 39564 25294 39620
rect 26898 39564 26908 39620
rect 26964 39564 27580 39620
rect 27636 39564 31948 39620
rect 32004 39564 32014 39620
rect 36418 39564 36428 39620
rect 36484 39564 37100 39620
rect 37156 39564 37166 39620
rect 39890 39564 39900 39620
rect 39956 39564 40348 39620
rect 40404 39564 41356 39620
rect 41412 39564 41422 39620
rect 45350 39564 45388 39620
rect 45444 39564 45454 39620
rect 46722 39564 46732 39620
rect 46788 39564 48076 39620
rect 48132 39564 48142 39620
rect 49858 39564 49868 39620
rect 49924 39564 49934 39620
rect 50082 39564 50092 39620
rect 50148 39564 50876 39620
rect 50932 39564 50942 39620
rect 49868 39508 49924 39564
rect 6290 39452 6300 39508
rect 6356 39452 7532 39508
rect 7588 39452 7598 39508
rect 12898 39452 12908 39508
rect 12964 39452 15484 39508
rect 15540 39452 19404 39508
rect 19460 39452 19470 39508
rect 19954 39452 19964 39508
rect 20020 39452 21420 39508
rect 21476 39452 21486 39508
rect 31714 39452 31724 39508
rect 31780 39452 37660 39508
rect 37716 39452 37726 39508
rect 41458 39452 41468 39508
rect 41524 39452 42028 39508
rect 42084 39452 42588 39508
rect 42644 39452 44828 39508
rect 44884 39452 44894 39508
rect 46946 39452 46956 39508
rect 47012 39452 49924 39508
rect 5058 39340 5068 39396
rect 5124 39340 8316 39396
rect 8372 39340 8382 39396
rect 15922 39340 15932 39396
rect 15988 39340 16716 39396
rect 16772 39340 16782 39396
rect 20066 39340 20076 39396
rect 20132 39340 22092 39396
rect 22148 39340 22158 39396
rect 46498 39340 46508 39396
rect 46564 39340 48748 39396
rect 48804 39340 48814 39396
rect 51426 39340 51436 39396
rect 51492 39340 55580 39396
rect 55636 39340 55646 39396
rect 13010 39228 13020 39284
rect 13076 39228 19684 39284
rect 45714 39228 45724 39284
rect 45780 39228 46844 39284
rect 46900 39228 46910 39284
rect 47170 39228 47180 39284
rect 47236 39228 48524 39284
rect 48580 39228 48590 39284
rect 4834 39116 4844 39172
rect 4900 39116 6860 39172
rect 6916 39116 6926 39172
rect 19628 39060 19684 39228
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 20850 39116 20860 39172
rect 20916 39116 21532 39172
rect 21588 39116 26908 39172
rect 26964 39116 28364 39172
rect 28420 39116 29148 39172
rect 29204 39116 29214 39172
rect 43810 39116 43820 39172
rect 43876 39116 44268 39172
rect 44324 39116 46284 39172
rect 46340 39116 47740 39172
rect 47796 39116 47806 39172
rect 2818 39004 2828 39060
rect 2884 39004 5852 39060
rect 5908 39004 5918 39060
rect 6738 39004 6748 39060
rect 6804 39004 7756 39060
rect 7812 39004 7822 39060
rect 15026 39004 15036 39060
rect 3042 38892 3052 38948
rect 3108 38892 3724 38948
rect 3780 38892 4508 38948
rect 4564 38892 5180 38948
rect 5236 38892 5246 38948
rect 5506 38892 5516 38948
rect 5572 38892 6300 38948
rect 6356 38892 6366 38948
rect 14774 38892 14812 38948
rect 14868 38892 14878 38948
rect 15092 38892 15148 39060
rect 15698 39004 15708 39060
rect 15764 39004 16156 39060
rect 16212 39004 16222 39060
rect 17714 39004 17724 39060
rect 17780 39004 19236 39060
rect 19628 39004 21308 39060
rect 21364 39004 22204 39060
rect 22260 39004 22270 39060
rect 30482 39004 30492 39060
rect 30548 39004 31612 39060
rect 31668 39004 32060 39060
rect 32116 39004 32126 39060
rect 33170 39004 33180 39060
rect 33236 39004 34300 39060
rect 34356 39004 34366 39060
rect 41458 39004 41468 39060
rect 41524 39004 42140 39060
rect 42196 39004 43540 39060
rect 44034 39004 44044 39060
rect 44100 39004 45388 39060
rect 45444 39004 45454 39060
rect 46732 39004 49868 39060
rect 49924 39004 50316 39060
rect 50372 39004 50382 39060
rect 19180 38948 19236 39004
rect 15204 38892 15214 38948
rect 16594 38892 16604 38948
rect 16660 38892 18284 38948
rect 18340 38892 18350 38948
rect 18834 38892 18844 38948
rect 18900 38892 18910 38948
rect 19180 38892 19852 38948
rect 19908 38892 20972 38948
rect 21028 38892 21038 38948
rect 36978 38892 36988 38948
rect 37044 38892 38444 38948
rect 38500 38892 38510 38948
rect 18844 38836 18900 38892
rect 43484 38836 43540 39004
rect 46732 38948 46788 39004
rect 43698 38892 43708 38948
rect 43764 38892 44268 38948
rect 44324 38892 44334 38948
rect 45826 38892 45836 38948
rect 45892 38892 46788 38948
rect 48038 38892 48076 38948
rect 48132 38892 48142 38948
rect 48738 38892 48748 38948
rect 48804 38892 49588 38948
rect 46732 38836 46788 38892
rect 49532 38836 49588 38892
rect 2482 38780 2492 38836
rect 2548 38780 3500 38836
rect 3556 38780 3566 38836
rect 5292 38780 5852 38836
rect 5908 38780 5918 38836
rect 6066 38780 6076 38836
rect 6132 38780 6860 38836
rect 6916 38780 7532 38836
rect 7588 38780 7598 38836
rect 13346 38780 13356 38836
rect 13412 38780 18900 38836
rect 22866 38780 22876 38836
rect 22932 38780 23660 38836
rect 23716 38780 24444 38836
rect 24500 38780 24510 38836
rect 28802 38780 28812 38836
rect 28868 38780 32172 38836
rect 32228 38780 32238 38836
rect 38322 38780 38332 38836
rect 38388 38780 38780 38836
rect 38836 38780 38846 38836
rect 42466 38780 42476 38836
rect 42532 38780 43260 38836
rect 43316 38780 43326 38836
rect 43484 38780 45164 38836
rect 45220 38780 45230 38836
rect 45602 38780 45612 38836
rect 45668 38780 45948 38836
rect 46004 38780 46014 38836
rect 46722 38780 46732 38836
rect 46788 38780 46798 38836
rect 47058 38780 47068 38836
rect 47124 38780 47964 38836
rect 48020 38780 49308 38836
rect 49364 38780 49374 38836
rect 49522 38780 49532 38836
rect 49588 38780 49598 38836
rect 54002 38780 54012 38836
rect 54068 38780 55468 38836
rect 55524 38780 57372 38836
rect 57428 38780 57438 38836
rect 1810 38668 1820 38724
rect 1876 38668 5068 38724
rect 5124 38668 5134 38724
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 5292 38276 5348 38780
rect 10770 38668 10780 38724
rect 10836 38668 15596 38724
rect 15652 38668 15662 38724
rect 15810 38668 15820 38724
rect 15876 38668 18060 38724
rect 18116 38668 18126 38724
rect 18274 38668 18284 38724
rect 18340 38668 18452 38724
rect 20402 38668 20412 38724
rect 20468 38668 20972 38724
rect 21028 38668 21038 38724
rect 22754 38668 22764 38724
rect 22820 38668 23044 38724
rect 33282 38668 33292 38724
rect 33348 38668 36652 38724
rect 36708 38668 36718 38724
rect 44594 38668 44604 38724
rect 44660 38668 45724 38724
rect 45780 38668 47628 38724
rect 47684 38668 47694 38724
rect 48514 38668 48524 38724
rect 48580 38668 50428 38724
rect 50484 38668 50494 38724
rect 50978 38668 50988 38724
rect 51044 38668 53228 38724
rect 53284 38668 53294 38724
rect 18396 38612 18452 38668
rect 22988 38612 23044 38668
rect 47628 38612 47684 38668
rect 15138 38556 15148 38612
rect 15204 38556 15242 38612
rect 15474 38556 15484 38612
rect 15540 38556 16492 38612
rect 16548 38556 16558 38612
rect 18396 38556 18732 38612
rect 18788 38556 18798 38612
rect 22988 38556 23436 38612
rect 23492 38556 23502 38612
rect 25218 38556 25228 38612
rect 25284 38556 25900 38612
rect 25956 38556 25966 38612
rect 26114 38556 26124 38612
rect 26180 38556 27468 38612
rect 27524 38556 27534 38612
rect 36530 38556 36540 38612
rect 36596 38556 37324 38612
rect 37380 38556 37390 38612
rect 37874 38556 37884 38612
rect 37940 38556 40348 38612
rect 40404 38556 40414 38612
rect 47628 38556 48860 38612
rect 48916 38556 48926 38612
rect 24994 38444 25004 38500
rect 25060 38444 33404 38500
rect 33460 38444 33470 38500
rect 36866 38444 36876 38500
rect 36932 38444 37772 38500
rect 37828 38444 37838 38500
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 45490 38332 45500 38388
rect 45556 38332 46620 38388
rect 46676 38332 46686 38388
rect 4610 38220 4620 38276
rect 4676 38220 5348 38276
rect 14354 38220 14364 38276
rect 14420 38220 15036 38276
rect 15092 38220 15102 38276
rect 49858 38220 49868 38276
rect 49924 38220 50876 38276
rect 50932 38220 52220 38276
rect 52276 38220 52286 38276
rect 6514 38108 6524 38164
rect 6580 38108 8204 38164
rect 8260 38108 8270 38164
rect 20850 38108 20860 38164
rect 20916 38108 25340 38164
rect 25396 38108 27692 38164
rect 27748 38108 27758 38164
rect 42690 38108 42700 38164
rect 42756 38108 43764 38164
rect 44258 38108 44268 38164
rect 44324 38108 44828 38164
rect 44884 38108 44894 38164
rect 45042 38108 45052 38164
rect 45108 38108 46060 38164
rect 46116 38108 46126 38164
rect 43708 38052 43764 38108
rect 14802 37996 14812 38052
rect 14868 37996 15036 38052
rect 15092 37996 15102 38052
rect 16370 37996 16380 38052
rect 16436 37996 17724 38052
rect 17780 37996 19852 38052
rect 19908 37996 19918 38052
rect 22642 37996 22652 38052
rect 22708 37996 23660 38052
rect 23716 37996 25004 38052
rect 25060 37996 25070 38052
rect 30146 37996 30156 38052
rect 30212 37996 31612 38052
rect 31668 37996 34244 38052
rect 37986 37996 37996 38052
rect 38052 37996 39228 38052
rect 39284 37996 39294 38052
rect 40114 37996 40124 38052
rect 40180 37996 41692 38052
rect 41748 37996 43372 38052
rect 43428 37996 43438 38052
rect 43698 37996 43708 38052
rect 43764 37996 44156 38052
rect 44212 37996 45500 38052
rect 45556 37996 45566 38052
rect 19852 37940 19908 37996
rect 15250 37884 15260 37940
rect 15316 37884 18620 37940
rect 18676 37884 18686 37940
rect 19852 37884 24332 37940
rect 24388 37884 24398 37940
rect 25330 37884 25340 37940
rect 25396 37884 25564 37940
rect 25620 37884 25630 37940
rect 29810 37884 29820 37940
rect 29876 37884 30380 37940
rect 30436 37884 31276 37940
rect 31332 37884 31342 37940
rect 34188 37828 34244 37996
rect 42242 37884 42252 37940
rect 42308 37884 44940 37940
rect 44996 37884 45006 37940
rect 45350 37884 45388 37940
rect 45444 37884 45454 37940
rect 14018 37772 14028 37828
rect 14084 37772 15596 37828
rect 15652 37772 15662 37828
rect 17602 37772 17612 37828
rect 17668 37772 18060 37828
rect 18116 37772 20300 37828
rect 20356 37772 33628 37828
rect 33684 37772 33694 37828
rect 34178 37772 34188 37828
rect 34244 37772 35532 37828
rect 35588 37772 35598 37828
rect 14802 37660 14812 37716
rect 14868 37660 15820 37716
rect 15876 37660 15886 37716
rect 24658 37660 24668 37716
rect 24724 37660 25228 37716
rect 25284 37660 25294 37716
rect 30828 37660 31500 37716
rect 31556 37660 33068 37716
rect 33124 37660 33134 37716
rect 33954 37660 33964 37716
rect 34020 37660 36428 37716
rect 36484 37660 37100 37716
rect 37156 37660 37166 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 30828 37604 30884 37660
rect 34412 37604 34468 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 14130 37548 14140 37604
rect 14196 37548 15036 37604
rect 15092 37548 16156 37604
rect 16212 37548 16222 37604
rect 19478 37548 19516 37604
rect 19572 37548 19582 37604
rect 30818 37548 30828 37604
rect 30884 37548 30894 37604
rect 34402 37548 34412 37604
rect 34468 37548 34478 37604
rect 37202 37548 37212 37604
rect 37268 37548 38780 37604
rect 38836 37548 38846 37604
rect 15092 37436 15260 37492
rect 15316 37436 15326 37492
rect 16034 37436 16044 37492
rect 16100 37436 21868 37492
rect 21924 37436 21934 37492
rect 26786 37436 26796 37492
rect 26852 37436 26862 37492
rect 31490 37436 31500 37492
rect 31556 37436 33516 37492
rect 33572 37436 34748 37492
rect 34804 37436 34814 37492
rect 38612 37436 39676 37492
rect 39732 37436 41020 37492
rect 41076 37436 41086 37492
rect 47618 37436 47628 37492
rect 47684 37436 49644 37492
rect 49700 37436 49710 37492
rect 53106 37436 53116 37492
rect 53172 37436 53788 37492
rect 53844 37436 53854 37492
rect 15092 37380 15148 37436
rect 26796 37380 26852 37436
rect 38612 37380 38668 37436
rect 4610 37324 4620 37380
rect 4676 37324 5180 37380
rect 5236 37324 5246 37380
rect 15026 37324 15036 37380
rect 15092 37324 26852 37380
rect 27122 37324 27132 37380
rect 27188 37324 38668 37380
rect 54898 37324 54908 37380
rect 54964 37324 55692 37380
rect 55748 37324 55758 37380
rect 16258 37212 16268 37268
rect 16324 37212 17612 37268
rect 17668 37212 17678 37268
rect 19282 37212 19292 37268
rect 19348 37212 20188 37268
rect 20244 37212 20254 37268
rect 31266 37212 31276 37268
rect 31332 37212 31948 37268
rect 32004 37212 32014 37268
rect 36194 37212 36204 37268
rect 36260 37212 37212 37268
rect 37268 37212 37278 37268
rect 38882 37212 38892 37268
rect 38948 37212 40012 37268
rect 40068 37212 40078 37268
rect 47618 37212 47628 37268
rect 47684 37212 48524 37268
rect 48580 37212 48590 37268
rect 53106 37212 53116 37268
rect 53172 37212 55356 37268
rect 55412 37212 55804 37268
rect 55860 37212 55870 37268
rect 9650 37100 9660 37156
rect 9716 37100 10108 37156
rect 10164 37100 12908 37156
rect 12964 37100 12974 37156
rect 14466 37100 14476 37156
rect 14532 37100 15260 37156
rect 15316 37100 15326 37156
rect 15698 37100 15708 37156
rect 15764 37100 17276 37156
rect 17332 37100 17342 37156
rect 27122 37100 27132 37156
rect 27188 37100 28252 37156
rect 28308 37100 28318 37156
rect 33394 37100 33404 37156
rect 33460 37100 45052 37156
rect 45108 37100 46620 37156
rect 46676 37100 46686 37156
rect 53442 37100 53452 37156
rect 53508 37100 54684 37156
rect 54740 37100 54750 37156
rect 10322 36988 10332 37044
rect 10388 36988 14812 37044
rect 14868 36988 14878 37044
rect 16594 36988 16604 37044
rect 16660 36988 17836 37044
rect 17892 36988 17902 37044
rect 19394 36988 19404 37044
rect 19460 36988 21980 37044
rect 22036 36988 22046 37044
rect 22978 36988 22988 37044
rect 23044 36988 23324 37044
rect 23380 36988 24444 37044
rect 24500 36988 24510 37044
rect 36642 36988 36652 37044
rect 36708 36988 37044 37044
rect 48150 36988 48188 37044
rect 48244 36988 48254 37044
rect 55010 36988 55020 37044
rect 55076 36988 55692 37044
rect 55748 36988 55758 37044
rect 36988 36932 37044 36988
rect 16482 36876 16492 36932
rect 16548 36876 19068 36932
rect 19124 36876 19134 36932
rect 27570 36876 27580 36932
rect 27636 36876 28252 36932
rect 28308 36876 28588 36932
rect 28644 36876 30828 36932
rect 30884 36876 30894 36932
rect 36988 36876 42588 36932
rect 42644 36876 43148 36932
rect 43204 36876 43214 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 18946 36764 18956 36820
rect 19012 36764 22204 36820
rect 22260 36764 22270 36820
rect 15474 36652 15484 36708
rect 15540 36652 17276 36708
rect 17332 36652 20076 36708
rect 20132 36652 20142 36708
rect 31490 36652 31500 36708
rect 31556 36652 33292 36708
rect 33348 36652 33358 36708
rect 16706 36540 16716 36596
rect 16772 36540 21980 36596
rect 22036 36540 22046 36596
rect 37212 36484 37268 36876
rect 38098 36764 38108 36820
rect 38164 36764 38892 36820
rect 38948 36764 40236 36820
rect 40292 36764 40302 36820
rect 47058 36764 47068 36820
rect 47124 36764 47628 36820
rect 47684 36764 53004 36820
rect 53060 36764 54236 36820
rect 54292 36764 54302 36820
rect 39778 36652 39788 36708
rect 39844 36652 40460 36708
rect 40516 36652 40526 36708
rect 46498 36652 46508 36708
rect 46564 36652 50764 36708
rect 50820 36652 50830 36708
rect 52546 36652 52556 36708
rect 52612 36652 54908 36708
rect 54964 36652 54974 36708
rect 49970 36540 49980 36596
rect 50036 36540 50652 36596
rect 50708 36540 50718 36596
rect 19478 36428 19516 36484
rect 19572 36428 19582 36484
rect 20066 36428 20076 36484
rect 20132 36428 21532 36484
rect 21588 36428 22092 36484
rect 22148 36428 24108 36484
rect 24164 36428 24174 36484
rect 32162 36428 32172 36484
rect 32228 36428 33740 36484
rect 33796 36428 33806 36484
rect 36082 36428 36092 36484
rect 36148 36428 36988 36484
rect 37044 36428 37054 36484
rect 37202 36428 37212 36484
rect 37268 36428 37278 36484
rect 44482 36428 44492 36484
rect 44548 36428 45164 36484
rect 45220 36428 46172 36484
rect 46228 36428 46238 36484
rect 46946 36428 46956 36484
rect 47012 36428 47022 36484
rect 47506 36428 47516 36484
rect 47572 36428 48076 36484
rect 48132 36428 48142 36484
rect 49532 36428 50540 36484
rect 50596 36428 50606 36484
rect 51986 36428 51996 36484
rect 52052 36428 53228 36484
rect 53284 36428 53294 36484
rect 53900 36428 54908 36484
rect 54964 36428 56364 36484
rect 56420 36428 57036 36484
rect 57092 36428 57102 36484
rect 46956 36372 47012 36428
rect 17602 36316 17612 36372
rect 17668 36316 19068 36372
rect 19124 36316 19134 36372
rect 21858 36316 21868 36372
rect 21924 36316 22652 36372
rect 22708 36316 22718 36372
rect 26226 36316 26236 36372
rect 26292 36316 30156 36372
rect 30212 36316 31164 36372
rect 31220 36316 31230 36372
rect 42578 36316 42588 36372
rect 42644 36316 47012 36372
rect 48150 36316 48188 36372
rect 48244 36316 49084 36372
rect 49140 36316 49150 36372
rect 17042 36204 17052 36260
rect 17108 36204 18284 36260
rect 18340 36204 20300 36260
rect 20356 36204 20366 36260
rect 30706 36204 30716 36260
rect 30772 36204 31276 36260
rect 31332 36204 31836 36260
rect 31892 36204 31902 36260
rect 36988 36204 38892 36260
rect 38948 36204 38958 36260
rect 44370 36204 44380 36260
rect 44436 36204 44716 36260
rect 44772 36204 44782 36260
rect 45602 36204 45612 36260
rect 45668 36204 46732 36260
rect 46788 36204 46798 36260
rect 47842 36204 47852 36260
rect 47908 36204 48636 36260
rect 48692 36204 49308 36260
rect 49364 36204 49374 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 16146 35868 16156 35924
rect 16212 35868 17388 35924
rect 17444 35868 17454 35924
rect 18274 35868 18284 35924
rect 18340 35868 22204 35924
rect 22260 35868 22270 35924
rect 25218 35868 25228 35924
rect 25284 35868 25452 35924
rect 25508 35868 25518 35924
rect 18284 35812 18340 35868
rect 36988 35812 37044 36204
rect 49532 36148 49588 36428
rect 51996 36372 52052 36428
rect 50194 36316 50204 36372
rect 50260 36316 52052 36372
rect 53900 36260 53956 36428
rect 55458 36316 55468 36372
rect 55524 36316 56588 36372
rect 56644 36316 56654 36372
rect 50306 36204 50316 36260
rect 50372 36204 53900 36260
rect 53956 36204 53966 36260
rect 55412 36204 55804 36260
rect 55860 36204 57484 36260
rect 57540 36204 57550 36260
rect 48066 36092 48076 36148
rect 48132 36092 49588 36148
rect 49970 36092 49980 36148
rect 50036 36092 50046 36148
rect 49980 36036 50036 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 47730 35980 47740 36036
rect 47796 35980 48748 36036
rect 48804 35980 48814 36036
rect 49980 35980 50316 36036
rect 50372 35980 50382 36036
rect 55412 35924 55468 36204
rect 44034 35868 44044 35924
rect 44100 35868 45164 35924
rect 45220 35868 48524 35924
rect 48580 35868 48590 35924
rect 49970 35868 49980 35924
rect 50036 35868 50876 35924
rect 50932 35868 54572 35924
rect 54628 35868 55468 35924
rect 14914 35756 14924 35812
rect 14980 35756 18340 35812
rect 21970 35756 21980 35812
rect 22036 35756 22046 35812
rect 22306 35756 22316 35812
rect 22372 35756 22876 35812
rect 22932 35756 22942 35812
rect 25778 35756 25788 35812
rect 25844 35756 26460 35812
rect 26516 35756 30716 35812
rect 30772 35756 30782 35812
rect 34626 35756 34636 35812
rect 34692 35756 36988 35812
rect 37044 35756 37054 35812
rect 47730 35756 47740 35812
rect 47796 35756 49196 35812
rect 49252 35756 49262 35812
rect 21980 35700 22036 35756
rect 14802 35644 14812 35700
rect 14868 35644 15484 35700
rect 15540 35644 15550 35700
rect 21980 35644 22428 35700
rect 22484 35644 22764 35700
rect 22820 35644 23884 35700
rect 23940 35644 27244 35700
rect 27300 35644 27310 35700
rect 31378 35644 31388 35700
rect 31444 35644 34076 35700
rect 34132 35644 34972 35700
rect 35028 35644 35038 35700
rect 36754 35644 36764 35700
rect 36820 35644 38892 35700
rect 38948 35644 41020 35700
rect 41076 35644 41086 35700
rect 45714 35644 45724 35700
rect 45780 35644 46172 35700
rect 46228 35644 46732 35700
rect 46788 35644 47292 35700
rect 47348 35644 47358 35700
rect 48038 35644 48076 35700
rect 48132 35644 48142 35700
rect 49410 35644 49420 35700
rect 49476 35644 50092 35700
rect 50148 35644 50652 35700
rect 50708 35644 50718 35700
rect 15092 35532 15596 35588
rect 15652 35532 15662 35588
rect 18722 35532 18732 35588
rect 18788 35532 19740 35588
rect 19796 35532 19806 35588
rect 22194 35532 22204 35588
rect 22260 35532 23436 35588
rect 23492 35532 23502 35588
rect 34850 35532 34860 35588
rect 34916 35532 36652 35588
rect 36708 35532 36718 35588
rect 44258 35532 44268 35588
rect 44324 35532 45500 35588
rect 45556 35532 45948 35588
rect 46004 35532 46014 35588
rect 47058 35532 47068 35588
rect 47124 35532 47852 35588
rect 47908 35532 47918 35588
rect 49522 35532 49532 35588
rect 49588 35532 51100 35588
rect 51156 35532 51166 35588
rect 55346 35532 55356 35588
rect 55412 35532 56700 35588
rect 56756 35532 56766 35588
rect 15092 35476 15148 35532
rect 13794 35420 13804 35476
rect 13860 35420 15148 35476
rect 35522 35420 35532 35476
rect 35588 35420 40236 35476
rect 40292 35420 40302 35476
rect 44146 35420 44156 35476
rect 44212 35420 44716 35476
rect 44772 35420 45612 35476
rect 45668 35420 48860 35476
rect 48916 35420 50652 35476
rect 50708 35420 50718 35476
rect 12002 35308 12012 35364
rect 12068 35308 12180 35364
rect 12898 35308 12908 35364
rect 12964 35308 12974 35364
rect 30258 35308 30268 35364
rect 30324 35308 30940 35364
rect 30996 35308 34860 35364
rect 34916 35308 34926 35364
rect 54898 35308 54908 35364
rect 54964 35308 55356 35364
rect 55412 35308 55422 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 12124 35252 12180 35308
rect 12908 35252 12964 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 12124 35196 14588 35252
rect 14644 35196 15820 35252
rect 15876 35196 16828 35252
rect 16884 35196 16894 35252
rect 49074 35196 49084 35252
rect 49140 35196 49756 35252
rect 49812 35196 53228 35252
rect 53284 35196 54572 35252
rect 54628 35196 54638 35252
rect 12674 35084 12684 35140
rect 12740 35084 13468 35140
rect 13524 35084 13534 35140
rect 29698 35084 29708 35140
rect 29764 35084 40908 35140
rect 40964 35084 41244 35140
rect 41300 35084 41310 35140
rect 52098 35084 52108 35140
rect 52164 35084 53116 35140
rect 53172 35084 53182 35140
rect 41010 34972 41020 35028
rect 41076 34972 42140 35028
rect 42196 34972 42206 35028
rect 52882 34972 52892 35028
rect 52948 34972 54460 35028
rect 54516 34972 54526 35028
rect 56242 34972 56252 35028
rect 56308 34972 57372 35028
rect 57428 34972 57438 35028
rect 19954 34860 19964 34916
rect 20020 34860 20636 34916
rect 20692 34860 20702 34916
rect 20962 34860 20972 34916
rect 21028 34860 22652 34916
rect 22708 34860 25900 34916
rect 25956 34860 25966 34916
rect 28130 34860 28140 34916
rect 28196 34860 33516 34916
rect 33572 34860 35308 34916
rect 35364 34860 35374 34916
rect 36642 34860 36652 34916
rect 36708 34860 37212 34916
rect 37268 34860 37278 34916
rect 45126 34860 45164 34916
rect 45220 34860 45230 34916
rect 45378 34860 45388 34916
rect 45444 34860 46060 34916
rect 46116 34860 48412 34916
rect 48468 34860 51324 34916
rect 51380 34860 51390 34916
rect 53778 34860 53788 34916
rect 53844 34860 54796 34916
rect 54852 34860 54862 34916
rect 35308 34804 35364 34860
rect 45164 34804 45220 34860
rect 16482 34748 16492 34804
rect 16548 34748 17500 34804
rect 17556 34748 17566 34804
rect 35308 34748 36988 34804
rect 37044 34748 37054 34804
rect 43586 34748 43596 34804
rect 43652 34748 44828 34804
rect 44884 34748 44894 34804
rect 45164 34748 46620 34804
rect 46676 34748 46686 34804
rect 17714 34636 17724 34692
rect 17780 34636 18956 34692
rect 19012 34636 19022 34692
rect 19842 34636 19852 34692
rect 19908 34636 21420 34692
rect 21476 34636 21486 34692
rect 21970 34636 21980 34692
rect 22036 34636 23100 34692
rect 23156 34636 23166 34692
rect 30146 34636 30156 34692
rect 30212 34636 30492 34692
rect 30548 34636 31052 34692
rect 31108 34636 31118 34692
rect 33842 34636 33852 34692
rect 33908 34636 34748 34692
rect 34804 34636 34814 34692
rect 39554 34636 39564 34692
rect 39620 34636 42700 34692
rect 42756 34636 43036 34692
rect 43092 34636 43372 34692
rect 43428 34636 45948 34692
rect 46004 34636 46014 34692
rect 49410 34636 49420 34692
rect 49476 34636 52108 34692
rect 52164 34636 52892 34692
rect 52948 34636 52958 34692
rect 55794 34636 55804 34692
rect 55860 34636 57260 34692
rect 57316 34636 57326 34692
rect 43810 34524 43820 34580
rect 43876 34524 44940 34580
rect 44996 34524 45276 34580
rect 45332 34524 45342 34580
rect 50988 34524 55580 34580
rect 55636 34524 55646 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 24434 34412 24444 34468
rect 24500 34412 25452 34468
rect 25508 34412 25518 34468
rect 47506 34412 47516 34468
rect 47572 34412 49196 34468
rect 49252 34412 49262 34468
rect 50988 34356 51044 34524
rect 15586 34300 15596 34356
rect 15652 34300 17388 34356
rect 17444 34300 20748 34356
rect 20804 34300 20814 34356
rect 23986 34300 23996 34356
rect 24052 34300 26796 34356
rect 26852 34300 27580 34356
rect 27636 34300 28588 34356
rect 28644 34300 28654 34356
rect 45462 34300 45500 34356
rect 45556 34300 45566 34356
rect 46732 34300 51044 34356
rect 54002 34300 54012 34356
rect 54068 34300 55244 34356
rect 55300 34300 55916 34356
rect 55972 34300 55982 34356
rect 56466 34300 56476 34356
rect 56532 34300 57372 34356
rect 57428 34300 57438 34356
rect 18834 34188 18844 34244
rect 18900 34188 21980 34244
rect 22036 34188 22046 34244
rect 43362 34188 43372 34244
rect 43428 34188 45612 34244
rect 45668 34188 45678 34244
rect 46732 34132 46788 34300
rect 48066 34188 48076 34244
rect 48132 34188 49532 34244
rect 49588 34188 49598 34244
rect 55010 34188 55020 34244
rect 55076 34188 56588 34244
rect 56644 34188 56654 34244
rect 15250 34076 15260 34132
rect 15316 34076 16380 34132
rect 16436 34076 17948 34132
rect 18004 34076 20188 34132
rect 20244 34076 20254 34132
rect 36754 34076 36764 34132
rect 36820 34076 37548 34132
rect 37604 34076 40348 34132
rect 40404 34076 40414 34132
rect 42578 34076 42588 34132
rect 42644 34076 46732 34132
rect 46788 34076 46798 34132
rect 47506 34076 47516 34132
rect 47572 34076 49084 34132
rect 49140 34076 49150 34132
rect 50306 34076 50316 34132
rect 50372 34076 51436 34132
rect 51492 34076 51502 34132
rect 17154 33964 17164 34020
rect 17220 33964 18508 34020
rect 18564 33964 18574 34020
rect 34738 33964 34748 34020
rect 34804 33964 35980 34020
rect 36036 33964 36046 34020
rect 36642 33964 36652 34020
rect 36708 33964 37100 34020
rect 37156 33964 37166 34020
rect 53218 33964 53228 34020
rect 53284 33964 53900 34020
rect 53956 33964 53966 34020
rect 54226 33852 54236 33908
rect 54292 33852 56028 33908
rect 56084 33852 56094 33908
rect 16930 33740 16940 33796
rect 16996 33740 27132 33796
rect 27188 33740 27198 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 13570 33628 13580 33684
rect 13636 33628 20412 33684
rect 20468 33628 23212 33684
rect 23268 33628 23278 33684
rect 49522 33628 49532 33684
rect 49588 33628 50316 33684
rect 50372 33628 50382 33684
rect 54786 33628 54796 33684
rect 54852 33628 56812 33684
rect 56868 33628 56878 33684
rect 14354 33516 14364 33572
rect 14420 33516 17276 33572
rect 17332 33516 17342 33572
rect 19170 33516 19180 33572
rect 19236 33516 23548 33572
rect 23604 33516 25564 33572
rect 25620 33516 25630 33572
rect 28690 33516 28700 33572
rect 28756 33516 30044 33572
rect 30100 33516 31052 33572
rect 31108 33516 31948 33572
rect 32004 33516 33068 33572
rect 33124 33516 33134 33572
rect 38546 33516 38556 33572
rect 38612 33516 41468 33572
rect 41524 33516 41534 33572
rect 54898 33516 54908 33572
rect 54964 33516 57372 33572
rect 57428 33516 57438 33572
rect 16902 33404 16940 33460
rect 16996 33404 17006 33460
rect 24882 33404 24892 33460
rect 24948 33404 26684 33460
rect 26740 33404 26750 33460
rect 33842 33404 33852 33460
rect 33908 33404 35084 33460
rect 35140 33404 35150 33460
rect 48850 33404 48860 33460
rect 48916 33404 51212 33460
rect 51268 33404 51278 33460
rect 12338 33292 12348 33348
rect 12404 33292 13580 33348
rect 13636 33292 15708 33348
rect 15764 33292 16716 33348
rect 16772 33292 18956 33348
rect 19012 33292 19628 33348
rect 19684 33292 22092 33348
rect 22148 33292 22764 33348
rect 22820 33292 23772 33348
rect 23828 33292 23838 33348
rect 35522 33292 35532 33348
rect 35588 33292 35980 33348
rect 36036 33292 42028 33348
rect 42084 33292 42094 33348
rect 46050 33292 46060 33348
rect 46116 33292 46844 33348
rect 46900 33292 46910 33348
rect 52098 33292 52108 33348
rect 52164 33292 55356 33348
rect 55412 33292 55422 33348
rect 56690 33292 56700 33348
rect 56756 33292 58156 33348
rect 58212 33292 58222 33348
rect 41906 33180 41916 33236
rect 41972 33180 46508 33236
rect 46564 33180 46574 33236
rect 16818 33068 16828 33124
rect 16884 33068 17724 33124
rect 17780 33068 17790 33124
rect 23426 33068 23436 33124
rect 23492 33068 26012 33124
rect 26068 33068 26078 33124
rect 27794 33068 27804 33124
rect 27860 33068 28812 33124
rect 28868 33068 28878 33124
rect 45378 33068 45388 33124
rect 45444 33068 45836 33124
rect 45892 33068 45902 33124
rect 46610 33068 46620 33124
rect 46676 33068 47180 33124
rect 47236 33068 52220 33124
rect 52276 33068 52286 33124
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 19618 32844 19628 32900
rect 19684 32844 19694 32900
rect 27570 32844 27580 32900
rect 27636 32844 32508 32900
rect 32564 32844 35420 32900
rect 35476 32844 35486 32900
rect 36978 32844 36988 32900
rect 37044 32844 38556 32900
rect 38612 32844 38622 32900
rect 42914 32844 42924 32900
rect 42980 32844 43484 32900
rect 43540 32844 43550 32900
rect 19628 32788 19684 32844
rect 17266 32732 17276 32788
rect 17332 32732 17342 32788
rect 19628 32732 20076 32788
rect 20132 32732 20142 32788
rect 26338 32732 26348 32788
rect 26404 32732 27244 32788
rect 27300 32732 27310 32788
rect 32162 32732 32172 32788
rect 32228 32732 33516 32788
rect 33572 32732 34188 32788
rect 34244 32732 34254 32788
rect 34412 32732 52108 32788
rect 52164 32732 52174 32788
rect 17276 32676 17332 32732
rect 34412 32676 34468 32732
rect 17276 32620 17780 32676
rect 30818 32620 30828 32676
rect 30884 32620 34468 32676
rect 35634 32620 35644 32676
rect 35700 32620 37436 32676
rect 37492 32620 38444 32676
rect 38500 32620 38612 32676
rect 43250 32620 43260 32676
rect 43316 32620 47404 32676
rect 47460 32620 49420 32676
rect 49476 32620 49486 32676
rect 17724 32564 17780 32620
rect 38556 32564 38612 32620
rect 17714 32508 17724 32564
rect 17780 32508 17790 32564
rect 23538 32508 23548 32564
rect 23604 32508 24892 32564
rect 24948 32508 24958 32564
rect 26114 32508 26124 32564
rect 26180 32508 27468 32564
rect 27524 32508 27534 32564
rect 38556 32508 39340 32564
rect 39396 32508 39406 32564
rect 44818 32508 44828 32564
rect 44884 32508 45724 32564
rect 45780 32508 45790 32564
rect 48066 32508 48076 32564
rect 48132 32508 48860 32564
rect 48916 32508 48926 32564
rect 49858 32508 49868 32564
rect 49924 32508 50540 32564
rect 50596 32508 50606 32564
rect 16034 32396 16044 32452
rect 16100 32396 17612 32452
rect 17668 32396 18620 32452
rect 18676 32396 18686 32452
rect 20178 32396 20188 32452
rect 20244 32396 25284 32452
rect 25666 32396 25676 32452
rect 25732 32396 27020 32452
rect 27076 32396 27086 32452
rect 41906 32396 41916 32452
rect 41972 32396 43148 32452
rect 43204 32396 43214 32452
rect 46946 32396 46956 32452
rect 47012 32396 47516 32452
rect 47572 32396 47582 32452
rect 25228 32340 25284 32396
rect 16258 32284 16268 32340
rect 16324 32284 17500 32340
rect 17556 32284 19740 32340
rect 19796 32284 19806 32340
rect 21746 32284 21756 32340
rect 21812 32284 25004 32340
rect 25060 32284 25070 32340
rect 25228 32284 29932 32340
rect 29988 32284 29998 32340
rect 46050 32284 46060 32340
rect 46116 32284 48412 32340
rect 48468 32284 48478 32340
rect 51090 32284 51100 32340
rect 51156 32284 52108 32340
rect 52164 32284 52174 32340
rect 16594 32172 16604 32228
rect 16660 32172 17836 32228
rect 17892 32172 17902 32228
rect 20738 32172 20748 32228
rect 20804 32172 23548 32228
rect 23604 32172 23614 32228
rect 43474 32172 43484 32228
rect 43540 32172 48188 32228
rect 48244 32172 49532 32228
rect 49588 32172 49598 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 17836 32116 17892 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 17836 32060 22204 32116
rect 22260 32060 23100 32116
rect 23156 32060 23772 32116
rect 23828 32060 23838 32116
rect 47618 32060 47628 32116
rect 47684 32060 49644 32116
rect 49700 32060 49710 32116
rect 50754 32060 50764 32116
rect 50820 32060 51156 32116
rect 51100 32004 51156 32060
rect 15586 31948 15596 32004
rect 15652 31948 16268 32004
rect 16324 31948 18396 32004
rect 18452 31948 18462 32004
rect 19730 31948 19740 32004
rect 19796 31948 23324 32004
rect 23380 31948 23390 32004
rect 34738 31948 34748 32004
rect 34804 31948 36652 32004
rect 36708 31948 36718 32004
rect 47170 31948 47180 32004
rect 47236 31948 48076 32004
rect 48132 31948 48142 32004
rect 48962 31948 48972 32004
rect 49028 31948 49980 32004
rect 50036 31948 50876 32004
rect 50932 31948 50942 32004
rect 51100 31948 51548 32004
rect 51604 31948 51614 32004
rect 52098 31948 52108 32004
rect 52164 31948 53396 32004
rect 13010 31836 13020 31892
rect 13076 31836 13692 31892
rect 13748 31836 13758 31892
rect 15138 31836 15148 31892
rect 15204 31836 16380 31892
rect 16436 31836 16446 31892
rect 16818 31836 16828 31892
rect 16884 31836 17108 31892
rect 17052 31668 17108 31836
rect 18806 31724 18844 31780
rect 18900 31724 18910 31780
rect 21868 31668 21924 31948
rect 53330 31892 53340 31948
rect 53396 31892 53406 31948
rect 27794 31836 27804 31892
rect 27860 31836 28364 31892
rect 28420 31836 30828 31892
rect 30884 31836 30894 31892
rect 33730 31836 33740 31892
rect 33796 31836 34412 31892
rect 34468 31836 36204 31892
rect 36260 31836 36270 31892
rect 37538 31836 37548 31892
rect 37604 31836 38108 31892
rect 38164 31836 38780 31892
rect 38836 31836 38846 31892
rect 44034 31836 44044 31892
rect 44100 31836 52668 31892
rect 52724 31836 52734 31892
rect 30258 31724 30268 31780
rect 30324 31724 31500 31780
rect 31556 31724 31566 31780
rect 33506 31724 33516 31780
rect 33572 31724 34300 31780
rect 34356 31724 34366 31780
rect 45602 31724 45612 31780
rect 45668 31724 46956 31780
rect 47012 31724 47022 31780
rect 49410 31724 49420 31780
rect 49476 31724 53228 31780
rect 53284 31724 53294 31780
rect 13458 31612 13468 31668
rect 13524 31612 16492 31668
rect 16548 31612 16558 31668
rect 17042 31612 17052 31668
rect 17108 31612 18172 31668
rect 18228 31612 18238 31668
rect 21858 31612 21868 31668
rect 21924 31612 21934 31668
rect 22418 31612 22428 31668
rect 22484 31612 23548 31668
rect 23604 31612 23614 31668
rect 24546 31612 24556 31668
rect 24612 31612 26348 31668
rect 26404 31612 26572 31668
rect 26628 31612 26638 31668
rect 32386 31612 32396 31668
rect 32452 31612 33852 31668
rect 33908 31612 33918 31668
rect 35522 31612 35532 31668
rect 35588 31612 37660 31668
rect 37716 31612 37726 31668
rect 40562 31612 40572 31668
rect 40628 31612 41916 31668
rect 41972 31612 43260 31668
rect 43316 31612 43326 31668
rect 44454 31612 44492 31668
rect 44548 31612 44558 31668
rect 48850 31612 48860 31668
rect 48916 31612 50428 31668
rect 50484 31612 50494 31668
rect 51986 31612 51996 31668
rect 52052 31612 56028 31668
rect 56084 31612 56094 31668
rect 16818 31500 16828 31556
rect 16884 31500 17388 31556
rect 17444 31500 18060 31556
rect 18116 31500 18126 31556
rect 20066 31500 20076 31556
rect 20132 31500 21812 31556
rect 21970 31500 21980 31556
rect 22036 31500 22876 31556
rect 22932 31500 22942 31556
rect 24434 31500 24444 31556
rect 24500 31500 25452 31556
rect 25508 31500 25518 31556
rect 34514 31500 34524 31556
rect 34580 31500 35196 31556
rect 35252 31500 35262 31556
rect 35970 31500 35980 31556
rect 36036 31500 36428 31556
rect 36484 31500 36494 31556
rect 37426 31500 37436 31556
rect 37492 31500 38332 31556
rect 38388 31500 42700 31556
rect 42756 31500 42766 31556
rect 48290 31500 48300 31556
rect 48356 31500 48972 31556
rect 49028 31500 49038 31556
rect 50642 31500 50652 31556
rect 50708 31500 52108 31556
rect 52164 31500 52174 31556
rect 21756 31444 21812 31500
rect 21756 31388 25228 31444
rect 25284 31388 25294 31444
rect 45826 31388 45836 31444
rect 45892 31388 49196 31444
rect 49252 31388 49532 31444
rect 49588 31388 49598 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 15698 31276 15708 31332
rect 15764 31276 16156 31332
rect 16212 31276 17668 31332
rect 49970 31276 49980 31332
rect 50036 31276 50204 31332
rect 50260 31276 50270 31332
rect 50978 31276 50988 31332
rect 51044 31276 51996 31332
rect 52052 31276 53452 31332
rect 53508 31276 53518 31332
rect 17612 31220 17668 31276
rect 15474 31164 15484 31220
rect 15540 31164 16604 31220
rect 16660 31164 17388 31220
rect 17444 31164 17454 31220
rect 17612 31164 22988 31220
rect 23044 31164 23054 31220
rect 40450 31164 40460 31220
rect 40516 31164 43372 31220
rect 43428 31164 43438 31220
rect 45826 31164 45836 31220
rect 45892 31164 46284 31220
rect 46340 31164 47516 31220
rect 47572 31164 47582 31220
rect 48626 31164 48636 31220
rect 48692 31164 49084 31220
rect 49140 31164 49150 31220
rect 49634 31164 49644 31220
rect 49700 31164 51100 31220
rect 51156 31164 51660 31220
rect 51716 31164 53676 31220
rect 53732 31164 53742 31220
rect 16370 31052 16380 31108
rect 16436 31052 17500 31108
rect 17556 31052 17566 31108
rect 41234 31052 41244 31108
rect 41300 31052 44940 31108
rect 44996 31052 46620 31108
rect 46676 31052 48636 31108
rect 48692 31052 54460 31108
rect 54516 31052 56700 31108
rect 56756 31052 56766 31108
rect 17938 30940 17948 30996
rect 18004 30940 19068 30996
rect 19124 30940 19134 30996
rect 23986 30940 23996 30996
rect 24052 30940 24556 30996
rect 24612 30940 24622 30996
rect 32050 30940 32060 30996
rect 32116 30940 32508 30996
rect 32564 30940 33180 30996
rect 33236 30940 33740 30996
rect 33796 30940 33806 30996
rect 40338 30940 40348 30996
rect 40404 30940 42140 30996
rect 42196 30940 43596 30996
rect 43652 30940 43662 30996
rect 44146 30940 44156 30996
rect 44212 30940 44716 30996
rect 44772 30940 48860 30996
rect 48916 30940 48926 30996
rect 50194 30940 50204 30996
rect 50260 30940 50988 30996
rect 51044 30940 51054 30996
rect 52994 30940 53004 30996
rect 53060 30940 53900 30996
rect 53956 30940 53966 30996
rect 29810 30828 29820 30884
rect 29876 30828 31276 30884
rect 31332 30828 31342 30884
rect 35186 30828 35196 30884
rect 35252 30828 38892 30884
rect 38948 30828 38958 30884
rect 46946 30828 46956 30884
rect 47012 30828 50540 30884
rect 50596 30828 50606 30884
rect 51426 30828 51436 30884
rect 51492 30828 52444 30884
rect 52500 30828 52510 30884
rect 14242 30716 14252 30772
rect 14308 30716 21644 30772
rect 21700 30716 21710 30772
rect 41010 30716 41020 30772
rect 41076 30716 45444 30772
rect 45388 30660 45444 30716
rect 14354 30604 14364 30660
rect 14420 30604 21196 30660
rect 21252 30604 21262 30660
rect 43922 30604 43932 30660
rect 43988 30604 44716 30660
rect 44772 30604 44782 30660
rect 45388 30604 54348 30660
rect 54404 30604 57148 30660
rect 57204 30604 57214 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 13570 30492 13580 30548
rect 13636 30492 14252 30548
rect 14308 30492 14318 30548
rect 19506 30492 19516 30548
rect 19572 30492 21420 30548
rect 21476 30492 21486 30548
rect 45266 30492 45276 30548
rect 45332 30492 46396 30548
rect 46452 30492 46462 30548
rect 36082 30380 36092 30436
rect 36148 30380 37100 30436
rect 37156 30380 37166 30436
rect 39554 30380 39564 30436
rect 39620 30380 45388 30436
rect 45444 30380 46620 30436
rect 46676 30380 46686 30436
rect 49074 30380 49084 30436
rect 49140 30380 49150 30436
rect 34962 30268 34972 30324
rect 35028 30268 35756 30324
rect 35812 30268 35822 30324
rect 38882 30268 38892 30324
rect 38948 30268 40460 30324
rect 40516 30268 40526 30324
rect 45490 30268 45500 30324
rect 45556 30268 46732 30324
rect 46788 30268 46798 30324
rect 49084 30212 49140 30380
rect 50642 30268 50652 30324
rect 50708 30268 51660 30324
rect 51716 30268 51726 30324
rect 52098 30268 52108 30324
rect 52164 30268 53564 30324
rect 53620 30268 53630 30324
rect 17938 30156 17948 30212
rect 18004 30156 19740 30212
rect 19796 30156 22876 30212
rect 22932 30156 22942 30212
rect 24322 30156 24332 30212
rect 24388 30156 25340 30212
rect 25396 30156 25406 30212
rect 26852 30156 28252 30212
rect 28308 30156 30268 30212
rect 30324 30156 30334 30212
rect 36530 30156 36540 30212
rect 36596 30156 36988 30212
rect 37044 30156 37054 30212
rect 37314 30156 37324 30212
rect 37380 30156 38780 30212
rect 38836 30156 38846 30212
rect 40114 30156 40124 30212
rect 40180 30156 40796 30212
rect 40852 30156 41468 30212
rect 41524 30156 41534 30212
rect 42466 30156 42476 30212
rect 42532 30156 43148 30212
rect 43204 30156 43214 30212
rect 49084 30156 50036 30212
rect 53330 30156 53340 30212
rect 53396 30156 53788 30212
rect 53844 30156 53854 30212
rect 9538 30044 9548 30100
rect 9604 30044 10332 30100
rect 10388 30044 10398 30100
rect 26852 29988 26908 30156
rect 49980 30100 50036 30156
rect 33842 30044 33852 30100
rect 33908 30044 48860 30100
rect 48916 30044 48926 30100
rect 49970 30044 49980 30100
rect 50036 30044 51548 30100
rect 51604 30044 51614 30100
rect 9762 29932 9772 29988
rect 9828 29932 26908 29988
rect 29586 29932 29596 29988
rect 29652 29932 30156 29988
rect 30212 29932 30222 29988
rect 33618 29932 33628 29988
rect 33684 29932 35420 29988
rect 35476 29932 35980 29988
rect 36036 29932 36046 29988
rect 43446 29932 43484 29988
rect 43540 29932 43550 29988
rect 44706 29932 44716 29988
rect 44772 29932 45164 29988
rect 45220 29932 46284 29988
rect 46340 29932 46350 29988
rect 21298 29820 21308 29876
rect 21364 29820 22092 29876
rect 22148 29820 25900 29876
rect 25956 29820 25966 29876
rect 42130 29820 42140 29876
rect 42196 29820 44492 29876
rect 44548 29820 45052 29876
rect 45108 29820 45118 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 29698 29596 29708 29652
rect 29764 29596 31276 29652
rect 31332 29596 31342 29652
rect 44818 29596 44828 29652
rect 44884 29596 47516 29652
rect 47572 29596 47582 29652
rect 49298 29596 49308 29652
rect 49364 29596 49644 29652
rect 49700 29596 49710 29652
rect 11218 29484 11228 29540
rect 11284 29484 12460 29540
rect 12516 29484 12526 29540
rect 12684 29484 18396 29540
rect 18452 29484 18462 29540
rect 28802 29484 28812 29540
rect 28868 29484 30828 29540
rect 30884 29484 30894 29540
rect 48066 29484 48076 29540
rect 48132 29484 49756 29540
rect 49812 29484 49822 29540
rect 12684 29428 12740 29484
rect 5282 29372 5292 29428
rect 5348 29372 8540 29428
rect 8596 29372 8606 29428
rect 11442 29372 11452 29428
rect 11508 29372 12740 29428
rect 13458 29372 13468 29428
rect 13524 29372 15932 29428
rect 15988 29372 16268 29428
rect 16324 29372 16334 29428
rect 27794 29372 27804 29428
rect 27860 29372 28700 29428
rect 28756 29372 28766 29428
rect 32162 29372 32172 29428
rect 32228 29372 33628 29428
rect 33684 29372 33694 29428
rect 34178 29372 34188 29428
rect 34244 29372 34636 29428
rect 34692 29372 35084 29428
rect 35140 29372 37324 29428
rect 37380 29372 37390 29428
rect 37986 29372 37996 29428
rect 38052 29372 44156 29428
rect 44212 29372 45500 29428
rect 45556 29372 46508 29428
rect 46564 29372 46574 29428
rect 47170 29372 47180 29428
rect 47236 29372 50428 29428
rect 50484 29372 51100 29428
rect 51156 29372 51166 29428
rect 52434 29372 52444 29428
rect 52500 29372 53676 29428
rect 53732 29372 54572 29428
rect 54628 29372 57372 29428
rect 57428 29372 57438 29428
rect 18050 29260 18060 29316
rect 18116 29260 18620 29316
rect 18676 29260 18956 29316
rect 19012 29260 19022 29316
rect 21298 29260 21308 29316
rect 21364 29260 24668 29316
rect 24724 29260 24734 29316
rect 32610 29260 32620 29316
rect 32676 29260 33516 29316
rect 33572 29260 35196 29316
rect 35252 29260 35262 29316
rect 43670 29260 43708 29316
rect 43764 29260 45164 29316
rect 45220 29260 45836 29316
rect 45892 29260 45902 29316
rect 47842 29260 47852 29316
rect 47908 29260 49980 29316
rect 50036 29260 50046 29316
rect 45238 29148 45276 29204
rect 45332 29148 45342 29204
rect 46050 29148 46060 29204
rect 46116 29148 46508 29204
rect 46564 29148 46574 29204
rect 52658 29148 52668 29204
rect 52724 29148 55804 29204
rect 55860 29148 55870 29204
rect 37538 29036 37548 29092
rect 37604 29036 41244 29092
rect 41300 29036 47740 29092
rect 47796 29036 47806 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 44930 28924 44940 28980
rect 44996 28924 45500 28980
rect 45556 28924 50988 28980
rect 51044 28924 53228 28980
rect 53284 28924 54012 28980
rect 54068 28924 54078 28980
rect 24994 28812 25004 28868
rect 25060 28812 27580 28868
rect 27636 28812 28252 28868
rect 28308 28812 28318 28868
rect 33506 28812 33516 28868
rect 33572 28812 35196 28868
rect 35252 28812 35262 28868
rect 45714 28812 45724 28868
rect 45780 28812 46620 28868
rect 46676 28812 46686 28868
rect 16706 28700 16716 28756
rect 16772 28700 16940 28756
rect 16996 28700 17006 28756
rect 29698 28700 29708 28756
rect 29764 28700 31276 28756
rect 31332 28700 31342 28756
rect 33394 28700 33404 28756
rect 33460 28700 36092 28756
rect 36148 28700 36158 28756
rect 36306 28700 36316 28756
rect 36372 28700 37100 28756
rect 37156 28700 37996 28756
rect 38052 28700 38062 28756
rect 39666 28700 39676 28756
rect 39732 28700 40684 28756
rect 40740 28700 41356 28756
rect 41412 28700 41422 28756
rect 46246 28700 46284 28756
rect 46340 28700 46350 28756
rect 46946 28700 46956 28756
rect 47012 28700 55244 28756
rect 55300 28700 55310 28756
rect 6514 28588 6524 28644
rect 6580 28588 7196 28644
rect 7252 28588 7262 28644
rect 25442 28588 25452 28644
rect 25508 28588 26796 28644
rect 26852 28588 26862 28644
rect 28466 28588 28476 28644
rect 28532 28588 30268 28644
rect 30324 28588 30334 28644
rect 35970 28588 35980 28644
rect 36036 28588 38332 28644
rect 38388 28588 38398 28644
rect 41906 28588 41916 28644
rect 41972 28588 42364 28644
rect 42420 28588 43372 28644
rect 43428 28588 43438 28644
rect 43922 28588 43932 28644
rect 43988 28588 48188 28644
rect 48244 28588 48254 28644
rect 49298 28588 49308 28644
rect 49364 28588 50316 28644
rect 50372 28588 50382 28644
rect 21298 28476 21308 28532
rect 21364 28476 22204 28532
rect 22260 28476 22270 28532
rect 47282 28476 47292 28532
rect 47348 28476 47852 28532
rect 47908 28476 47918 28532
rect 18918 28364 18956 28420
rect 19012 28364 19022 28420
rect 21634 28364 21644 28420
rect 21700 28364 23996 28420
rect 24052 28364 24062 28420
rect 30146 28364 30156 28420
rect 30212 28364 32844 28420
rect 32900 28364 32910 28420
rect 46470 28364 46508 28420
rect 46564 28364 46574 28420
rect 50372 28364 52668 28420
rect 52724 28364 52734 28420
rect 50372 28308 50428 28364
rect 45938 28252 45948 28308
rect 46004 28252 47628 28308
rect 47684 28252 50428 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 53330 28140 53340 28196
rect 53396 28140 55692 28196
rect 55748 28140 56588 28196
rect 56644 28140 56654 28196
rect 18834 28028 18844 28084
rect 18900 28028 19740 28084
rect 19796 28028 22092 28084
rect 22148 28028 22158 28084
rect 31938 28028 31948 28084
rect 32004 28028 34860 28084
rect 34916 28028 35644 28084
rect 35700 28028 38668 28084
rect 46610 28028 46620 28084
rect 46676 28028 46844 28084
rect 46900 28028 47628 28084
rect 47684 28028 47694 28084
rect 47842 28028 47852 28084
rect 47908 28028 52108 28084
rect 52164 28028 52174 28084
rect 53106 28028 53116 28084
rect 53172 28028 55580 28084
rect 55636 28028 55646 28084
rect 7522 27916 7532 27972
rect 7588 27916 8428 27972
rect 8484 27916 8494 27972
rect 16258 27916 16268 27972
rect 16324 27916 20188 27972
rect 20244 27916 20254 27972
rect 20514 27916 20524 27972
rect 20580 27916 21644 27972
rect 21700 27916 22652 27972
rect 22708 27916 22718 27972
rect 23986 27916 23996 27972
rect 24052 27916 24668 27972
rect 24724 27916 25340 27972
rect 25396 27916 25406 27972
rect 34412 27916 36652 27972
rect 36708 27916 36718 27972
rect 34412 27860 34468 27916
rect 6626 27804 6636 27860
rect 6692 27804 7924 27860
rect 20738 27804 20748 27860
rect 20804 27804 21532 27860
rect 21588 27804 21598 27860
rect 24434 27804 24444 27860
rect 24500 27804 25452 27860
rect 25508 27804 25518 27860
rect 32946 27804 32956 27860
rect 33012 27804 33404 27860
rect 33460 27804 33470 27860
rect 34402 27804 34412 27860
rect 34468 27804 34478 27860
rect 35186 27804 35196 27860
rect 35252 27804 36540 27860
rect 36596 27804 36606 27860
rect 7868 27748 7924 27804
rect 6290 27692 6300 27748
rect 6356 27692 7084 27748
rect 7140 27692 7150 27748
rect 7858 27692 7868 27748
rect 7924 27692 10668 27748
rect 10724 27692 13916 27748
rect 13972 27692 13982 27748
rect 4946 27580 4956 27636
rect 5012 27580 6748 27636
rect 6804 27580 6814 27636
rect 8278 27580 8316 27636
rect 8372 27580 8382 27636
rect 21634 27580 21644 27636
rect 21700 27580 22876 27636
rect 22932 27580 23660 27636
rect 23716 27580 23726 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 22082 27356 22092 27412
rect 22148 27356 23660 27412
rect 23716 27356 23726 27412
rect 35532 27300 35588 27804
rect 38612 27748 38668 28028
rect 48402 27916 48412 27972
rect 48468 27916 50652 27972
rect 50708 27916 50718 27972
rect 52780 27916 53564 27972
rect 53620 27916 55020 27972
rect 55076 27916 55086 27972
rect 52780 27860 52836 27916
rect 51874 27804 51884 27860
rect 51940 27804 52780 27860
rect 52836 27804 52846 27860
rect 54338 27804 54348 27860
rect 54404 27804 56700 27860
rect 56756 27804 56766 27860
rect 38612 27692 40012 27748
rect 40068 27692 40078 27748
rect 42018 27692 42028 27748
rect 42084 27692 43036 27748
rect 43092 27692 45164 27748
rect 45220 27692 50428 27748
rect 50484 27692 52332 27748
rect 52388 27692 52398 27748
rect 52658 27692 52668 27748
rect 52724 27692 55468 27748
rect 55524 27692 55534 27748
rect 45826 27580 45836 27636
rect 45892 27580 46956 27636
rect 47012 27580 47022 27636
rect 50530 27580 50540 27636
rect 50596 27580 54684 27636
rect 54740 27580 54750 27636
rect 50642 27468 50652 27524
rect 50708 27468 53788 27524
rect 53844 27468 54908 27524
rect 54964 27468 54974 27524
rect 46834 27356 46844 27412
rect 46900 27356 53228 27412
rect 53284 27356 53294 27412
rect 35186 27244 35196 27300
rect 35252 27244 35588 27300
rect 42914 27244 42924 27300
rect 42980 27244 44828 27300
rect 44884 27244 51548 27300
rect 51604 27244 51614 27300
rect 16034 27132 16044 27188
rect 16100 27132 18732 27188
rect 18788 27132 18798 27188
rect 25554 27132 25564 27188
rect 25620 27132 26460 27188
rect 26516 27132 26526 27188
rect 33058 27132 33068 27188
rect 33124 27132 34860 27188
rect 34916 27132 35868 27188
rect 35924 27132 35934 27188
rect 38770 27132 38780 27188
rect 38836 27132 39564 27188
rect 39620 27132 41916 27188
rect 41972 27132 43036 27188
rect 43092 27132 43102 27188
rect 47730 27132 47740 27188
rect 47796 27132 49420 27188
rect 49476 27132 49486 27188
rect 49970 27132 49980 27188
rect 50036 27132 53004 27188
rect 53060 27132 53070 27188
rect 19180 27020 20076 27076
rect 20132 27020 22540 27076
rect 22596 27020 22606 27076
rect 23762 27020 23772 27076
rect 23828 27020 24892 27076
rect 24948 27020 27020 27076
rect 27076 27020 28812 27076
rect 28868 27020 29260 27076
rect 29316 27020 29326 27076
rect 32386 27020 32396 27076
rect 32452 27020 33404 27076
rect 33460 27020 34188 27076
rect 34244 27020 34254 27076
rect 34626 27020 34636 27076
rect 34692 27020 35084 27076
rect 35140 27020 35150 27076
rect 35634 27020 35644 27076
rect 35700 27020 36092 27076
rect 36148 27020 36158 27076
rect 42466 27020 42476 27076
rect 42532 27020 44156 27076
rect 44212 27020 44222 27076
rect 46498 27020 46508 27076
rect 46564 27020 49868 27076
rect 49924 27020 49934 27076
rect 52322 27020 52332 27076
rect 52388 27020 53676 27076
rect 53732 27020 54124 27076
rect 54180 27020 54572 27076
rect 54628 27020 54638 27076
rect 4834 26908 4844 26964
rect 4900 26908 5628 26964
rect 5684 26908 5694 26964
rect 8082 26908 8092 26964
rect 8148 26908 8428 26964
rect 8484 26908 8494 26964
rect 18610 26908 18620 26964
rect 18676 26908 18900 26964
rect 7634 26796 7644 26852
rect 7700 26796 8428 26852
rect 8484 26796 10556 26852
rect 10612 26796 10622 26852
rect 2258 26460 2268 26516
rect 2324 26460 3500 26516
rect 3556 26460 3566 26516
rect 13906 26460 13916 26516
rect 13972 26460 15372 26516
rect 15428 26460 15438 26516
rect 18844 26292 18900 26908
rect 19180 26852 19236 27020
rect 21522 26908 21532 26964
rect 21588 26908 22876 26964
rect 22932 26908 22942 26964
rect 25442 26908 25452 26964
rect 25508 26908 26684 26964
rect 26740 26908 26750 26964
rect 34290 26908 34300 26964
rect 34356 26908 35196 26964
rect 35252 26908 35262 26964
rect 42354 26908 42364 26964
rect 42420 26908 43260 26964
rect 43316 26908 43326 26964
rect 47954 26908 47964 26964
rect 48020 26908 48748 26964
rect 48804 26908 48814 26964
rect 53330 26908 53340 26964
rect 53396 26908 54908 26964
rect 54964 26908 54974 26964
rect 26460 26852 26516 26908
rect 19180 26796 19292 26852
rect 19348 26796 19358 26852
rect 19842 26796 19852 26852
rect 19908 26796 21980 26852
rect 22036 26796 22046 26852
rect 26450 26796 26460 26852
rect 26516 26796 26526 26852
rect 32834 26796 32844 26852
rect 32900 26796 33180 26852
rect 33236 26796 33246 26852
rect 34412 26740 34468 26908
rect 35522 26796 35532 26852
rect 35588 26796 36876 26852
rect 36932 26796 37660 26852
rect 37716 26796 38332 26852
rect 38388 26796 38398 26852
rect 19058 26684 19068 26740
rect 19124 26684 19404 26740
rect 19460 26684 19470 26740
rect 32946 26684 32956 26740
rect 33012 26684 34468 26740
rect 35746 26684 35756 26740
rect 35812 26684 37100 26740
rect 37156 26684 37166 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 24546 26572 24556 26628
rect 24612 26572 24622 26628
rect 37314 26572 37324 26628
rect 37380 26572 38892 26628
rect 38948 26572 40012 26628
rect 40068 26572 40078 26628
rect 40226 26572 40236 26628
rect 40292 26572 42140 26628
rect 42196 26572 44268 26628
rect 44324 26572 44716 26628
rect 44772 26572 44782 26628
rect 21410 26348 21420 26404
rect 21476 26348 22540 26404
rect 22596 26348 22606 26404
rect 9874 26236 9884 26292
rect 9940 26236 10556 26292
rect 10612 26236 10622 26292
rect 11442 26236 11452 26292
rect 11508 26236 12572 26292
rect 12628 26236 12638 26292
rect 17938 26236 17948 26292
rect 18004 26236 18620 26292
rect 18676 26236 18686 26292
rect 18834 26236 18844 26292
rect 18900 26236 18910 26292
rect 24556 26180 24612 26572
rect 43810 26460 43820 26516
rect 43876 26460 46396 26516
rect 46452 26460 46462 26516
rect 48150 26460 48188 26516
rect 48244 26460 49420 26516
rect 49476 26460 49486 26516
rect 53442 26460 53452 26516
rect 53508 26460 55580 26516
rect 55636 26460 55646 26516
rect 33068 26348 34300 26404
rect 34356 26348 35084 26404
rect 35140 26348 35150 26404
rect 43474 26348 43484 26404
rect 43540 26348 43932 26404
rect 43988 26348 45388 26404
rect 45444 26348 45836 26404
rect 45892 26348 45902 26404
rect 46834 26348 46844 26404
rect 46900 26348 47516 26404
rect 47572 26348 47582 26404
rect 48850 26348 48860 26404
rect 48916 26348 49308 26404
rect 49364 26348 49644 26404
rect 49700 26348 49710 26404
rect 33068 26292 33124 26348
rect 28578 26236 28588 26292
rect 28644 26236 29596 26292
rect 29652 26236 29662 26292
rect 33058 26236 33068 26292
rect 33124 26236 33134 26292
rect 33730 26236 33740 26292
rect 33796 26236 34860 26292
rect 34916 26236 34926 26292
rect 39778 26236 39788 26292
rect 39844 26236 41020 26292
rect 41076 26236 41086 26292
rect 43138 26236 43148 26292
rect 43204 26236 44380 26292
rect 44436 26236 45556 26292
rect 46274 26236 46284 26292
rect 46340 26236 47180 26292
rect 47236 26236 47246 26292
rect 49074 26236 49084 26292
rect 49140 26236 49150 26292
rect 49970 26236 49980 26292
rect 50036 26236 50764 26292
rect 50820 26236 51436 26292
rect 51492 26236 51502 26292
rect 45500 26180 45556 26236
rect 3490 26124 3500 26180
rect 3556 26124 4172 26180
rect 4228 26124 6524 26180
rect 6580 26124 7420 26180
rect 7476 26124 8204 26180
rect 8260 26124 9436 26180
rect 9492 26124 9502 26180
rect 17826 26124 17836 26180
rect 17892 26124 19628 26180
rect 19684 26124 19964 26180
rect 20020 26124 20030 26180
rect 23314 26124 23324 26180
rect 23380 26124 24108 26180
rect 24164 26124 24174 26180
rect 24434 26124 24444 26180
rect 24500 26124 24612 26180
rect 30706 26124 30716 26180
rect 30772 26124 33180 26180
rect 33236 26124 33246 26180
rect 33954 26124 33964 26180
rect 34020 26124 34972 26180
rect 35028 26124 35038 26180
rect 45490 26124 45500 26180
rect 45556 26124 45566 26180
rect 49084 26068 49140 26236
rect 49634 26124 49644 26180
rect 49700 26124 50876 26180
rect 50932 26124 50942 26180
rect 15698 26012 15708 26068
rect 15764 26012 16156 26068
rect 16212 26012 28588 26068
rect 28644 26012 28654 26068
rect 34860 26012 40796 26068
rect 40852 26012 40862 26068
rect 49084 26012 50988 26068
rect 51044 26012 52220 26068
rect 52276 26012 52286 26068
rect 34860 25956 34916 26012
rect 18610 25900 18620 25956
rect 18676 25900 18956 25956
rect 19012 25900 19022 25956
rect 33506 25900 33516 25956
rect 33572 25900 34916 25956
rect 42802 25900 42812 25956
rect 42868 25900 49532 25956
rect 49588 25900 49598 25956
rect 50866 25900 50876 25956
rect 50932 25900 51996 25956
rect 52052 25900 54684 25956
rect 54740 25900 54750 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 45714 25788 45724 25844
rect 45780 25788 46060 25844
rect 46116 25788 46126 25844
rect 47842 25788 47852 25844
rect 47908 25788 48524 25844
rect 48580 25788 48590 25844
rect 52098 25676 52108 25732
rect 52164 25676 53116 25732
rect 53172 25676 53182 25732
rect 53330 25676 53340 25732
rect 53396 25676 54796 25732
rect 54852 25676 54862 25732
rect 11666 25564 11676 25620
rect 11732 25564 12348 25620
rect 12404 25564 12414 25620
rect 18834 25564 18844 25620
rect 18900 25564 24220 25620
rect 24276 25564 24286 25620
rect 34514 25564 34524 25620
rect 34580 25564 36428 25620
rect 36484 25564 37548 25620
rect 37604 25564 37884 25620
rect 37940 25564 37950 25620
rect 45490 25564 45500 25620
rect 45556 25564 46732 25620
rect 46788 25564 47516 25620
rect 47572 25564 47582 25620
rect 50754 25564 50764 25620
rect 50820 25564 53004 25620
rect 53060 25564 53070 25620
rect 18274 25452 18284 25508
rect 18340 25452 21420 25508
rect 21476 25452 21980 25508
rect 22036 25452 22046 25508
rect 23090 25452 23100 25508
rect 23156 25452 24332 25508
rect 24388 25452 24398 25508
rect 43138 25452 43148 25508
rect 43204 25452 47404 25508
rect 47460 25452 47470 25508
rect 51538 25452 51548 25508
rect 51604 25452 52108 25508
rect 52164 25452 52668 25508
rect 52724 25452 52734 25508
rect 12562 25340 12572 25396
rect 12628 25340 14140 25396
rect 14196 25340 14206 25396
rect 18722 25340 18732 25396
rect 18788 25340 19740 25396
rect 19796 25340 19806 25396
rect 23762 25340 23772 25396
rect 23828 25340 25676 25396
rect 25732 25340 26236 25396
rect 26292 25340 26302 25396
rect 37314 25340 37324 25396
rect 37380 25340 38108 25396
rect 38164 25340 38174 25396
rect 41682 25340 41692 25396
rect 41748 25340 42476 25396
rect 42532 25340 42542 25396
rect 46610 25340 46620 25396
rect 46676 25340 46956 25396
rect 47012 25340 47740 25396
rect 47796 25340 47806 25396
rect 48636 25340 49420 25396
rect 49476 25340 49486 25396
rect 52546 25340 52556 25396
rect 52612 25340 53452 25396
rect 53508 25340 53518 25396
rect 48636 25284 48692 25340
rect 9762 25228 9772 25284
rect 9828 25228 12236 25284
rect 12292 25228 12796 25284
rect 12852 25228 13916 25284
rect 13972 25228 13982 25284
rect 18834 25228 18844 25284
rect 18900 25228 21532 25284
rect 21588 25228 21598 25284
rect 24098 25228 24108 25284
rect 24164 25228 25172 25284
rect 6850 25116 6860 25172
rect 6916 25116 8652 25172
rect 8708 25116 18284 25172
rect 18340 25116 18350 25172
rect 23650 25116 23660 25172
rect 23716 25116 24780 25172
rect 24836 25116 24846 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 25116 25060 25172 25228
rect 34076 25228 34860 25284
rect 34916 25228 44716 25284
rect 44772 25228 44782 25284
rect 47282 25228 47292 25284
rect 47348 25228 47358 25284
rect 48598 25228 48636 25284
rect 48692 25228 48702 25284
rect 49074 25228 49084 25284
rect 49140 25228 51436 25284
rect 51492 25228 52108 25284
rect 52164 25228 52174 25284
rect 52434 25228 52444 25284
rect 52500 25228 52780 25284
rect 52836 25228 54236 25284
rect 54292 25228 54302 25284
rect 34076 25172 34132 25228
rect 47292 25172 47348 25228
rect 34066 25116 34076 25172
rect 34132 25116 34142 25172
rect 40338 25116 40348 25172
rect 40404 25116 41804 25172
rect 41860 25116 41870 25172
rect 44930 25116 44940 25172
rect 44996 25116 48860 25172
rect 48916 25116 48926 25172
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 8278 25004 8316 25060
rect 8372 25004 8382 25060
rect 20738 25004 20748 25060
rect 20804 25004 22204 25060
rect 22260 25004 22988 25060
rect 23044 25004 23054 25060
rect 23426 25004 23436 25060
rect 23492 25004 23884 25060
rect 23940 25004 24444 25060
rect 24500 25004 24510 25060
rect 25106 25004 25116 25060
rect 25172 25004 25182 25060
rect 39778 25004 39788 25060
rect 39844 25004 40572 25060
rect 40628 25004 40638 25060
rect 10882 24892 10892 24948
rect 10948 24892 11676 24948
rect 11732 24892 11742 24948
rect 12898 24892 12908 24948
rect 12964 24892 13580 24948
rect 13636 24892 18396 24948
rect 18452 24892 18462 24948
rect 23986 24892 23996 24948
rect 24052 24892 24556 24948
rect 24612 24892 24622 24948
rect 26226 24892 26236 24948
rect 26292 24892 27916 24948
rect 27972 24892 29372 24948
rect 29428 24892 29438 24948
rect 35522 24892 35532 24948
rect 35588 24892 37212 24948
rect 37268 24892 37278 24948
rect 39218 24892 39228 24948
rect 39284 24892 41020 24948
rect 41076 24892 41086 24948
rect 20066 24780 20076 24836
rect 20132 24780 20636 24836
rect 20692 24780 20702 24836
rect 35634 24780 35644 24836
rect 35700 24780 39116 24836
rect 39172 24780 40348 24836
rect 40404 24780 40414 24836
rect 45042 24780 45052 24836
rect 45108 24780 46620 24836
rect 46676 24780 46686 24836
rect 47282 24780 47292 24836
rect 47348 24780 48972 24836
rect 49028 24780 49038 24836
rect 40898 24668 40908 24724
rect 40964 24668 41916 24724
rect 41972 24668 42700 24724
rect 42756 24668 42766 24724
rect 48066 24668 48076 24724
rect 48132 24668 49084 24724
rect 49140 24668 50316 24724
rect 50372 24668 50382 24724
rect 13122 24556 13132 24612
rect 13188 24556 13468 24612
rect 13524 24556 14924 24612
rect 14980 24556 14990 24612
rect 17490 24556 17500 24612
rect 17556 24556 20748 24612
rect 20804 24556 20814 24612
rect 22194 24556 22204 24612
rect 22260 24556 22540 24612
rect 22596 24556 23996 24612
rect 24052 24556 24444 24612
rect 24500 24556 24510 24612
rect 33954 24556 33964 24612
rect 34020 24556 34860 24612
rect 34916 24556 36316 24612
rect 36372 24556 37436 24612
rect 37492 24556 37502 24612
rect 45938 24556 45948 24612
rect 46004 24556 47068 24612
rect 47124 24556 47134 24612
rect 15092 24444 29148 24500
rect 29204 24444 29214 24500
rect 15092 24388 15148 24444
rect 12002 24332 12012 24388
rect 12068 24332 12460 24388
rect 12516 24332 13244 24388
rect 13300 24332 15148 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 36614 24220 36652 24276
rect 36708 24220 43708 24276
rect 43764 24220 45388 24276
rect 45444 24220 45454 24276
rect 40562 24108 40572 24164
rect 40628 24108 41356 24164
rect 41412 24108 42252 24164
rect 42308 24108 42318 24164
rect 47730 24108 47740 24164
rect 47796 24108 48748 24164
rect 48804 24108 48814 24164
rect 22754 23996 22764 24052
rect 22820 23996 23436 24052
rect 23492 23996 25228 24052
rect 25284 23996 25294 24052
rect 33170 23996 33180 24052
rect 33236 23996 33852 24052
rect 33908 23996 34188 24052
rect 34244 23996 34254 24052
rect 36082 23996 36092 24052
rect 36148 23996 37212 24052
rect 37268 23996 37278 24052
rect 43810 23996 43820 24052
rect 43876 23996 44828 24052
rect 44884 23996 46284 24052
rect 46340 23996 46350 24052
rect 47170 23996 47180 24052
rect 47236 23996 50652 24052
rect 50708 23996 50718 24052
rect 7970 23884 7980 23940
rect 8036 23884 12908 23940
rect 12964 23884 12974 23940
rect 18386 23884 18396 23940
rect 18452 23884 20188 23940
rect 20244 23884 20860 23940
rect 20916 23884 23212 23940
rect 23268 23884 23278 23940
rect 24210 23884 24220 23940
rect 24276 23884 24892 23940
rect 24948 23884 24958 23940
rect 37986 23884 37996 23940
rect 38052 23884 40796 23940
rect 40852 23884 41804 23940
rect 41860 23884 42364 23940
rect 42420 23884 42924 23940
rect 42980 23884 42990 23940
rect 44930 23884 44940 23940
rect 44996 23884 46508 23940
rect 46564 23884 47516 23940
rect 47572 23884 47582 23940
rect 48290 23884 48300 23940
rect 48356 23884 49532 23940
rect 49588 23884 49598 23940
rect 50082 23884 50092 23940
rect 50148 23884 51100 23940
rect 51156 23884 51166 23940
rect 51650 23884 51660 23940
rect 51716 23884 53004 23940
rect 53060 23884 53070 23940
rect 48300 23828 48356 23884
rect 18498 23772 18508 23828
rect 18564 23772 18844 23828
rect 18900 23772 19068 23828
rect 19124 23772 19134 23828
rect 19618 23772 19628 23828
rect 19684 23772 22764 23828
rect 22820 23772 22830 23828
rect 36194 23772 36204 23828
rect 36260 23772 36428 23828
rect 36484 23772 37100 23828
rect 37156 23772 37166 23828
rect 40226 23772 40236 23828
rect 40292 23772 40684 23828
rect 40740 23772 41356 23828
rect 41412 23772 41422 23828
rect 47394 23772 47404 23828
rect 47460 23772 48356 23828
rect 51762 23772 51772 23828
rect 51828 23772 53564 23828
rect 53620 23772 53630 23828
rect 7074 23660 7084 23716
rect 7140 23660 7868 23716
rect 7924 23660 8540 23716
rect 8596 23660 8606 23716
rect 24322 23660 24332 23716
rect 24388 23660 25004 23716
rect 25060 23660 25070 23716
rect 34626 23660 34636 23716
rect 34692 23660 35196 23716
rect 35252 23660 37212 23716
rect 37268 23660 37278 23716
rect 40450 23660 40460 23716
rect 40516 23660 43036 23716
rect 43092 23660 43102 23716
rect 51538 23660 51548 23716
rect 51604 23660 53676 23716
rect 53732 23660 53742 23716
rect 23100 23548 24556 23604
rect 24612 23548 24622 23604
rect 41906 23548 41916 23604
rect 41972 23548 45444 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 23100 23492 23156 23548
rect 45388 23492 45444 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 14354 23436 14364 23492
rect 14420 23436 15260 23492
rect 15316 23436 16380 23492
rect 16436 23436 16446 23492
rect 17938 23436 17948 23492
rect 18004 23436 19068 23492
rect 19124 23436 19134 23492
rect 23090 23436 23100 23492
rect 23156 23436 23166 23492
rect 37090 23436 37100 23492
rect 37156 23436 38556 23492
rect 38612 23436 38622 23492
rect 45388 23436 47068 23492
rect 47124 23436 47134 23492
rect 49186 23436 49196 23492
rect 49252 23436 49756 23492
rect 49812 23436 49822 23492
rect 3714 23324 3724 23380
rect 3780 23324 5404 23380
rect 5460 23324 5470 23380
rect 13682 23324 13692 23380
rect 13748 23324 14028 23380
rect 14084 23324 14094 23380
rect 21186 23324 21196 23380
rect 21252 23324 21868 23380
rect 21924 23324 21934 23380
rect 33618 23324 33628 23380
rect 33684 23324 34972 23380
rect 35028 23324 35038 23380
rect 38210 23324 38220 23380
rect 38276 23324 39900 23380
rect 39956 23324 39966 23380
rect 41458 23324 41468 23380
rect 41524 23324 46060 23380
rect 46116 23324 48188 23380
rect 48244 23324 48254 23380
rect 50866 23324 50876 23380
rect 50932 23324 52332 23380
rect 52388 23324 52398 23380
rect 15586 23212 15596 23268
rect 15652 23212 16380 23268
rect 16436 23212 17500 23268
rect 17556 23212 21812 23268
rect 26338 23212 26348 23268
rect 26404 23212 27356 23268
rect 27412 23212 27422 23268
rect 29474 23212 29484 23268
rect 29540 23212 30716 23268
rect 30772 23212 30782 23268
rect 42018 23212 42028 23268
rect 42084 23212 43484 23268
rect 43540 23212 43550 23268
rect 44706 23212 44716 23268
rect 44772 23212 48076 23268
rect 48132 23212 48142 23268
rect 49074 23212 49084 23268
rect 49140 23212 49644 23268
rect 49700 23212 50428 23268
rect 50484 23212 52668 23268
rect 52724 23212 52734 23268
rect 21756 23156 21812 23212
rect 6514 23100 6524 23156
rect 6580 23100 7308 23156
rect 7364 23100 7374 23156
rect 19730 23100 19740 23156
rect 19796 23100 20524 23156
rect 20580 23100 21532 23156
rect 21588 23100 21598 23156
rect 21756 23100 27580 23156
rect 27636 23100 27646 23156
rect 41794 23100 41804 23156
rect 41860 23100 43708 23156
rect 43764 23100 43774 23156
rect 46386 23100 46396 23156
rect 46452 23100 47516 23156
rect 47572 23100 47582 23156
rect 47730 23100 47740 23156
rect 47796 23100 48188 23156
rect 48244 23100 48254 23156
rect 50082 23100 50092 23156
rect 50148 23100 55804 23156
rect 55860 23100 55870 23156
rect 5058 22988 5068 23044
rect 5124 22988 5740 23044
rect 5796 22988 5806 23044
rect 7522 22988 7532 23044
rect 7588 22988 8764 23044
rect 8820 22988 8830 23044
rect 19618 22988 19628 23044
rect 19684 22988 22204 23044
rect 22260 22988 22270 23044
rect 4722 22876 4732 22932
rect 4788 22876 6076 22932
rect 6132 22876 7980 22932
rect 8036 22876 8046 22932
rect 20626 22876 20636 22932
rect 20692 22876 20972 22932
rect 21028 22876 21038 22932
rect 24434 22876 24444 22932
rect 24500 22876 25340 22932
rect 25396 22876 25406 22932
rect 32162 22876 32172 22932
rect 32228 22876 35588 22932
rect 35746 22876 35756 22932
rect 35812 22876 38332 22932
rect 38388 22876 38398 22932
rect 45938 22876 45948 22932
rect 46004 22876 46508 22932
rect 46564 22876 46574 22932
rect 35532 22820 35588 22876
rect 13682 22764 13692 22820
rect 13748 22764 14588 22820
rect 14644 22764 15820 22820
rect 15876 22764 25564 22820
rect 25620 22764 25630 22820
rect 35532 22764 42588 22820
rect 42644 22764 43596 22820
rect 43652 22764 50876 22820
rect 50932 22764 52444 22820
rect 52500 22764 52510 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 6402 22652 6412 22708
rect 6468 22652 14924 22708
rect 14980 22652 16716 22708
rect 16772 22652 16782 22708
rect 36194 22652 36204 22708
rect 36260 22652 37212 22708
rect 37268 22652 44268 22708
rect 44324 22652 44940 22708
rect 44996 22652 45006 22708
rect 45266 22652 45276 22708
rect 45332 22652 50092 22708
rect 50148 22652 50158 22708
rect 5730 22540 5740 22596
rect 5796 22540 7308 22596
rect 7364 22540 7374 22596
rect 11778 22540 11788 22596
rect 11844 22540 12460 22596
rect 12516 22540 12526 22596
rect 13122 22540 13132 22596
rect 13188 22540 14476 22596
rect 14532 22540 22540 22596
rect 22596 22540 22606 22596
rect 25218 22540 25228 22596
rect 25284 22540 25676 22596
rect 25732 22540 26908 22596
rect 26964 22540 26974 22596
rect 35970 22540 35980 22596
rect 36036 22540 36652 22596
rect 36708 22540 46732 22596
rect 46788 22540 46798 22596
rect 47180 22540 48748 22596
rect 48804 22540 48814 22596
rect 51762 22540 51772 22596
rect 51828 22540 52668 22596
rect 52724 22540 52734 22596
rect 47180 22484 47236 22540
rect 16146 22428 16156 22484
rect 16212 22428 16940 22484
rect 16996 22428 26684 22484
rect 26740 22428 26750 22484
rect 28466 22428 28476 22484
rect 28532 22428 29596 22484
rect 29652 22428 29662 22484
rect 38210 22428 38220 22484
rect 38276 22428 40236 22484
rect 40292 22428 40302 22484
rect 46834 22428 46844 22484
rect 46900 22428 47180 22484
rect 47236 22428 47246 22484
rect 48178 22428 48188 22484
rect 48244 22428 50428 22484
rect 50484 22428 50494 22484
rect 2818 22316 2828 22372
rect 2884 22316 5740 22372
rect 5796 22316 5806 22372
rect 10882 22316 10892 22372
rect 10948 22316 11452 22372
rect 11508 22316 11518 22372
rect 17938 22316 17948 22372
rect 18004 22316 18844 22372
rect 18900 22316 18910 22372
rect 19170 22316 19180 22372
rect 19236 22316 20188 22372
rect 20244 22316 23324 22372
rect 23380 22316 23390 22372
rect 23548 22316 30044 22372
rect 30100 22316 30110 22372
rect 34738 22316 34748 22372
rect 34804 22316 35756 22372
rect 35812 22316 36876 22372
rect 36932 22316 36942 22372
rect 39890 22316 39900 22372
rect 39956 22316 40796 22372
rect 40852 22316 41692 22372
rect 41748 22316 41758 22372
rect 43474 22316 43484 22372
rect 43540 22316 45164 22372
rect 45220 22316 45230 22372
rect 46050 22316 46060 22372
rect 46116 22316 47292 22372
rect 47348 22316 47358 22372
rect 23548 22260 23604 22316
rect 12562 22204 12572 22260
rect 12628 22204 13580 22260
rect 13636 22204 14588 22260
rect 14644 22204 14654 22260
rect 16706 22204 16716 22260
rect 16772 22204 17164 22260
rect 17220 22204 23604 22260
rect 25218 22204 25228 22260
rect 25284 22204 27692 22260
rect 27748 22204 29820 22260
rect 29876 22204 29886 22260
rect 36418 22204 36428 22260
rect 36484 22204 36988 22260
rect 37044 22204 37324 22260
rect 37380 22204 37390 22260
rect 43698 22204 43708 22260
rect 43764 22204 45276 22260
rect 45332 22204 45342 22260
rect 48290 22204 48300 22260
rect 48356 22204 49196 22260
rect 49252 22204 49262 22260
rect 50866 22204 50876 22260
rect 50932 22204 51996 22260
rect 52052 22204 52556 22260
rect 52612 22204 52622 22260
rect 6850 22092 6860 22148
rect 6916 22092 12460 22148
rect 12516 22092 16380 22148
rect 16436 22092 19292 22148
rect 19348 22092 19358 22148
rect 22082 22092 22092 22148
rect 22148 22092 26348 22148
rect 26404 22092 26414 22148
rect 33954 22092 33964 22148
rect 34020 22092 34412 22148
rect 34468 22092 34478 22148
rect 42354 22092 42364 22148
rect 42420 22092 43372 22148
rect 43428 22092 44716 22148
rect 44772 22092 44782 22148
rect 47394 22092 47404 22148
rect 47460 22092 48524 22148
rect 48580 22092 49308 22148
rect 49364 22092 49374 22148
rect 10556 21980 15260 22036
rect 15316 21980 15708 22036
rect 15764 21980 15774 22036
rect 35746 21980 35756 22036
rect 35812 21980 37100 22036
rect 37156 21980 37166 22036
rect 47842 21980 47852 22036
rect 47908 21980 48860 22036
rect 48916 21980 48926 22036
rect 10556 21924 10612 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 8306 21868 8316 21924
rect 8372 21868 9212 21924
rect 9268 21868 10612 21924
rect 15026 21868 15036 21924
rect 15092 21812 15148 21924
rect 21074 21868 21084 21924
rect 21140 21868 23660 21924
rect 23716 21868 24892 21924
rect 24948 21868 24958 21924
rect 27570 21868 27580 21924
rect 27636 21868 28476 21924
rect 28532 21868 28542 21924
rect 34402 21868 34412 21924
rect 34468 21868 38332 21924
rect 38388 21868 38398 21924
rect 40338 21868 40348 21924
rect 40404 21868 40414 21924
rect 41570 21868 41580 21924
rect 41636 21868 42476 21924
rect 42532 21868 42542 21924
rect 24892 21812 24948 21868
rect 40348 21812 40404 21868
rect 7746 21756 7756 21812
rect 7812 21756 14252 21812
rect 14308 21756 14318 21812
rect 15092 21756 19124 21812
rect 20290 21756 20300 21812
rect 20356 21756 21308 21812
rect 21364 21756 21374 21812
rect 23426 21756 23436 21812
rect 23492 21756 24556 21812
rect 24612 21756 24622 21812
rect 24892 21756 25116 21812
rect 25172 21756 25182 21812
rect 25554 21756 25564 21812
rect 25620 21756 27020 21812
rect 27076 21756 27086 21812
rect 34626 21756 34636 21812
rect 34692 21756 35196 21812
rect 35252 21756 35262 21812
rect 39330 21756 39340 21812
rect 39396 21756 40404 21812
rect 19068 21700 19124 21756
rect 10882 21644 10892 21700
rect 10948 21644 12124 21700
rect 12180 21644 12190 21700
rect 15092 21644 15932 21700
rect 15988 21644 15998 21700
rect 19058 21644 19068 21700
rect 19124 21644 19134 21700
rect 22082 21644 22092 21700
rect 22148 21644 22316 21700
rect 22372 21644 22382 21700
rect 23874 21644 23884 21700
rect 23940 21644 25004 21700
rect 25060 21644 25070 21700
rect 27458 21644 27468 21700
rect 27524 21644 28028 21700
rect 28084 21644 33852 21700
rect 33908 21644 33918 21700
rect 38434 21644 38444 21700
rect 38500 21644 39116 21700
rect 39172 21644 40012 21700
rect 40068 21644 40078 21700
rect 42354 21644 42364 21700
rect 42420 21644 44380 21700
rect 44436 21644 44446 21700
rect 15092 21588 15148 21644
rect 7746 21532 7756 21588
rect 7812 21532 8204 21588
rect 8260 21532 8652 21588
rect 8708 21532 9324 21588
rect 9380 21532 9390 21588
rect 14354 21532 14364 21588
rect 14420 21532 15148 21588
rect 15586 21532 15596 21588
rect 15652 21532 18620 21588
rect 18676 21532 23660 21588
rect 23716 21532 23726 21588
rect 41234 21532 41244 21588
rect 41300 21532 42140 21588
rect 42196 21532 43148 21588
rect 43204 21532 43214 21588
rect 25890 21420 25900 21476
rect 25956 21420 33740 21476
rect 33796 21420 35756 21476
rect 35812 21420 35822 21476
rect 37650 21420 37660 21476
rect 37716 21420 39228 21476
rect 39284 21420 39294 21476
rect 39666 21420 39676 21476
rect 39732 21420 43036 21476
rect 43092 21420 43102 21476
rect 43362 21420 43372 21476
rect 43428 21420 44156 21476
rect 44212 21420 44222 21476
rect 45266 21420 45276 21476
rect 45332 21420 47628 21476
rect 47684 21420 47694 21476
rect 12674 21308 12684 21364
rect 12740 21308 13468 21364
rect 13524 21308 13534 21364
rect 16118 21308 16156 21364
rect 16212 21308 16222 21364
rect 8866 21196 8876 21252
rect 8932 21196 13916 21252
rect 13972 21196 13982 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 12114 21084 12124 21140
rect 12180 21084 13244 21140
rect 13300 21084 16156 21140
rect 16212 21084 16222 21140
rect 3602 20972 3612 21028
rect 3668 20972 5740 21028
rect 5796 20972 5806 21028
rect 9090 20972 9100 21028
rect 9156 20972 10108 21028
rect 10164 20972 10174 21028
rect 42242 20860 42252 20916
rect 42308 20860 44492 20916
rect 44548 20860 44558 20916
rect 13794 20748 13804 20804
rect 13860 20748 15148 20804
rect 15204 20748 15214 20804
rect 15922 20748 15932 20804
rect 15988 20748 22988 20804
rect 23044 20748 23054 20804
rect 34514 20748 34524 20804
rect 34580 20748 35196 20804
rect 35252 20748 35262 20804
rect 40898 20748 40908 20804
rect 40964 20748 42140 20804
rect 42196 20748 43932 20804
rect 43988 20748 43998 20804
rect 44930 20748 44940 20804
rect 44996 20748 48188 20804
rect 48244 20748 48254 20804
rect 7410 20636 7420 20692
rect 7476 20636 7868 20692
rect 7924 20636 7934 20692
rect 19170 20636 19180 20692
rect 19236 20636 20300 20692
rect 20356 20636 20366 20692
rect 8082 20524 8092 20580
rect 8148 20524 14364 20580
rect 14420 20524 14430 20580
rect 15092 20524 20524 20580
rect 20580 20524 21420 20580
rect 21476 20524 22204 20580
rect 22260 20524 22764 20580
rect 22820 20524 22830 20580
rect 23650 20524 23660 20580
rect 23716 20524 24108 20580
rect 24164 20524 24174 20580
rect 43250 20524 43260 20580
rect 43316 20524 50876 20580
rect 50932 20524 50942 20580
rect 15092 20468 15148 20524
rect 8194 20412 8204 20468
rect 8260 20412 8652 20468
rect 8708 20412 15148 20468
rect 21074 20412 21084 20468
rect 21140 20412 23884 20468
rect 23940 20412 24556 20468
rect 24612 20412 24622 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 4610 20300 4620 20356
rect 4676 20300 5404 20356
rect 5460 20300 8764 20356
rect 8820 20300 8830 20356
rect 12786 20188 12796 20244
rect 12852 20188 14028 20244
rect 14084 20188 14094 20244
rect 15362 20188 15372 20244
rect 15428 20188 15438 20244
rect 16370 20188 16380 20244
rect 16436 20188 23100 20244
rect 23156 20188 23166 20244
rect 15372 20132 15428 20188
rect 6066 20076 6076 20132
rect 6132 20076 7084 20132
rect 7140 20076 7150 20132
rect 7298 20076 7308 20132
rect 7364 20076 10668 20132
rect 10724 20076 10734 20132
rect 13906 20076 13916 20132
rect 13972 20076 15428 20132
rect 18498 20076 18508 20132
rect 18564 20076 20188 20132
rect 20244 20076 21420 20132
rect 21476 20076 21486 20132
rect 21634 20076 21644 20132
rect 21700 20076 21710 20132
rect 22418 20076 22428 20132
rect 22484 20076 27916 20132
rect 27972 20076 27982 20132
rect 28354 20076 28364 20132
rect 28420 20076 30828 20132
rect 30884 20076 30894 20132
rect 34738 20076 34748 20132
rect 34804 20076 35308 20132
rect 35364 20076 35374 20132
rect 40338 20076 40348 20132
rect 40404 20076 41132 20132
rect 41188 20076 41804 20132
rect 41860 20076 41870 20132
rect 21644 20020 21700 20076
rect 2818 19964 2828 20020
rect 2884 19964 5068 20020
rect 5124 19964 5134 20020
rect 5954 19964 5964 20020
rect 6020 19964 6860 20020
rect 6916 19964 6926 20020
rect 10210 19964 10220 20020
rect 10276 19964 11116 20020
rect 11172 19964 11182 20020
rect 13682 19964 13692 20020
rect 13748 19964 14028 20020
rect 14084 19964 14700 20020
rect 14756 19964 14766 20020
rect 14886 19964 14924 20020
rect 14980 19964 14990 20020
rect 21298 19964 21308 20020
rect 21364 19964 21700 20020
rect 24658 19964 24668 20020
rect 24724 19964 25228 20020
rect 25284 19964 25294 20020
rect 25890 19964 25900 20020
rect 25956 19964 26908 20020
rect 27794 19964 27804 20020
rect 27860 19964 34860 20020
rect 34916 19964 34926 20020
rect 6178 19852 6188 19908
rect 6244 19852 18172 19908
rect 18228 19852 18238 19908
rect 21410 19852 21420 19908
rect 21476 19852 25564 19908
rect 25620 19852 25630 19908
rect 26852 19796 26908 19964
rect 29586 19852 29596 19908
rect 29652 19852 31276 19908
rect 31332 19852 31342 19908
rect 34290 19852 34300 19908
rect 34356 19852 35980 19908
rect 36036 19852 36046 19908
rect 36306 19852 36316 19908
rect 36372 19852 37884 19908
rect 37940 19852 38556 19908
rect 38612 19852 39004 19908
rect 39060 19852 39452 19908
rect 39508 19852 39518 19908
rect 13346 19740 13356 19796
rect 13412 19740 13580 19796
rect 13636 19740 13646 19796
rect 19170 19740 19180 19796
rect 19236 19740 20300 19796
rect 20356 19740 20366 19796
rect 22866 19740 22876 19796
rect 22932 19740 23324 19796
rect 23380 19740 23390 19796
rect 24210 19740 24220 19796
rect 24276 19740 25340 19796
rect 25396 19740 25406 19796
rect 26852 19740 33068 19796
rect 33124 19740 35756 19796
rect 35812 19740 35822 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 18498 19516 18508 19572
rect 18564 19516 23100 19572
rect 23156 19516 23166 19572
rect 10098 19404 10108 19460
rect 10164 19404 12572 19460
rect 12628 19404 12638 19460
rect 12898 19292 12908 19348
rect 12964 19292 13468 19348
rect 13524 19292 13534 19348
rect 23314 19292 23324 19348
rect 23380 19292 24332 19348
rect 24388 19292 24398 19348
rect 13570 19180 13580 19236
rect 13636 19180 14476 19236
rect 14532 19180 14542 19236
rect 16034 19180 16044 19236
rect 16100 19180 16604 19236
rect 16660 19180 16670 19236
rect 18722 19180 18732 19236
rect 18788 19180 19404 19236
rect 19460 19180 19852 19236
rect 19908 19180 19918 19236
rect 21298 19180 21308 19236
rect 21364 19180 26796 19236
rect 26852 19180 26862 19236
rect 6290 19068 6300 19124
rect 6356 19068 8092 19124
rect 8148 19068 8158 19124
rect 9090 19068 9100 19124
rect 9156 19068 9772 19124
rect 9828 19068 22652 19124
rect 22708 19068 23212 19124
rect 23268 19068 23278 19124
rect 27906 19068 27916 19124
rect 27972 19068 29820 19124
rect 29876 19068 29886 19124
rect 30370 19068 30380 19124
rect 30436 19068 36092 19124
rect 36148 19068 36158 19124
rect 13682 18956 13692 19012
rect 13748 18956 15148 19012
rect 15204 18956 16604 19012
rect 16660 18956 16670 19012
rect 19628 18956 21644 19012
rect 21700 18956 22876 19012
rect 22932 18956 22942 19012
rect 23874 18956 23884 19012
rect 23940 18956 23950 19012
rect 25330 18956 25340 19012
rect 25396 18956 28028 19012
rect 28084 18956 28094 19012
rect 19628 18900 19684 18956
rect 7746 18844 7756 18900
rect 7812 18844 7868 18900
rect 7924 18844 7934 18900
rect 14242 18844 14252 18900
rect 14308 18844 19684 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 23884 18788 23940 18956
rect 24882 18844 24892 18900
rect 24948 18844 25676 18900
rect 25732 18844 25742 18900
rect 35634 18844 35644 18900
rect 35700 18844 36316 18900
rect 36372 18844 37436 18900
rect 37492 18844 37502 18900
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 7522 18732 7532 18788
rect 7588 18732 7868 18788
rect 7924 18732 7934 18788
rect 8306 18732 8316 18788
rect 8372 18732 13916 18788
rect 13972 18732 13982 18788
rect 23884 18732 30604 18788
rect 30660 18732 30670 18788
rect 6934 18620 6972 18676
rect 7028 18620 7038 18676
rect 7298 18620 7308 18676
rect 7364 18620 9548 18676
rect 9604 18620 9614 18676
rect 10546 18620 10556 18676
rect 10612 18620 11116 18676
rect 11172 18620 11182 18676
rect 13682 18620 13692 18676
rect 13748 18620 14140 18676
rect 14196 18620 14206 18676
rect 16594 18620 16604 18676
rect 16660 18620 24108 18676
rect 24164 18620 24174 18676
rect 24434 18620 24444 18676
rect 24500 18620 25228 18676
rect 25284 18620 25294 18676
rect 5506 18508 5516 18564
rect 5572 18508 6300 18564
rect 6356 18508 6366 18564
rect 6514 18508 6524 18564
rect 6580 18508 7532 18564
rect 7588 18508 7598 18564
rect 8978 18508 8988 18564
rect 9044 18508 9772 18564
rect 9828 18508 10668 18564
rect 10724 18508 10734 18564
rect 23314 18508 23324 18564
rect 23380 18508 29372 18564
rect 29428 18508 29438 18564
rect 4050 18396 4060 18452
rect 4116 18396 5964 18452
rect 6020 18396 6030 18452
rect 10882 18396 10892 18452
rect 10948 18396 12684 18452
rect 12740 18396 12750 18452
rect 13010 18396 13020 18452
rect 13076 18396 15036 18452
rect 15092 18396 15102 18452
rect 16930 18396 16940 18452
rect 16996 18396 17500 18452
rect 17556 18396 18732 18452
rect 18788 18396 20748 18452
rect 20804 18396 22092 18452
rect 22148 18396 25340 18452
rect 25396 18396 25900 18452
rect 25956 18396 25966 18452
rect 27682 18396 27692 18452
rect 27748 18396 28364 18452
rect 28420 18396 29708 18452
rect 29764 18396 32396 18452
rect 32452 18396 32462 18452
rect 35186 18396 35196 18452
rect 35252 18396 37660 18452
rect 37716 18396 37726 18452
rect 11666 18284 11676 18340
rect 11732 18284 12796 18340
rect 12852 18284 12862 18340
rect 23202 18284 23212 18340
rect 23268 18284 23996 18340
rect 24052 18284 24062 18340
rect 24210 18284 24220 18340
rect 24276 18284 25228 18340
rect 25284 18284 25294 18340
rect 8194 18172 8204 18228
rect 8260 18172 10108 18228
rect 10164 18172 10174 18228
rect 11442 18172 11452 18228
rect 11508 18172 12348 18228
rect 12404 18172 12414 18228
rect 12562 18172 12572 18228
rect 12628 18172 13692 18228
rect 13748 18172 15148 18228
rect 20178 18172 20188 18228
rect 20244 18172 21644 18228
rect 21700 18172 28028 18228
rect 28084 18172 28094 18228
rect 15092 18116 15148 18172
rect 9874 18060 9884 18116
rect 9940 18060 14308 18116
rect 15092 18060 15596 18116
rect 15652 18060 15662 18116
rect 19366 18060 19404 18116
rect 19460 18060 19470 18116
rect 21970 18060 21980 18116
rect 22036 18060 24892 18116
rect 24948 18060 24958 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 14252 18004 14308 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 6850 17948 6860 18004
rect 6916 17948 7308 18004
rect 7364 17948 7374 18004
rect 11778 17948 11788 18004
rect 11844 17948 14028 18004
rect 14084 17948 14094 18004
rect 14252 17948 15148 18004
rect 15204 17948 15214 18004
rect 2034 17836 2044 17892
rect 2100 17836 5740 17892
rect 5796 17836 5806 17892
rect 6066 17836 6076 17892
rect 6132 17836 6748 17892
rect 6804 17836 6814 17892
rect 10098 17836 10108 17892
rect 10164 17836 12460 17892
rect 12516 17836 12526 17892
rect 14242 17836 14252 17892
rect 14308 17836 15260 17892
rect 15316 17836 16716 17892
rect 16772 17836 16782 17892
rect 28354 17836 28364 17892
rect 28420 17836 29596 17892
rect 29652 17836 29662 17892
rect 6076 17780 6132 17836
rect 4610 17724 4620 17780
rect 4676 17724 6132 17780
rect 8754 17724 8764 17780
rect 8820 17724 15148 17780
rect 34066 17724 34076 17780
rect 34132 17724 35532 17780
rect 35588 17724 35598 17780
rect 12786 17612 12796 17668
rect 12852 17612 13804 17668
rect 13860 17612 13870 17668
rect 15092 17556 15148 17724
rect 19618 17612 19628 17668
rect 19684 17612 24108 17668
rect 24164 17612 24444 17668
rect 24500 17612 24510 17668
rect 25330 17612 25340 17668
rect 25396 17612 26124 17668
rect 26180 17612 26190 17668
rect 28578 17612 28588 17668
rect 28644 17612 29148 17668
rect 29204 17612 29214 17668
rect 32162 17612 32172 17668
rect 32228 17612 33404 17668
rect 33460 17612 33470 17668
rect 36194 17612 36204 17668
rect 36260 17612 37100 17668
rect 37156 17612 38556 17668
rect 38612 17612 38622 17668
rect 6738 17500 6748 17556
rect 6804 17500 9100 17556
rect 9156 17500 9166 17556
rect 9538 17500 9548 17556
rect 9604 17500 12012 17556
rect 12068 17500 12078 17556
rect 12338 17500 12348 17556
rect 12404 17500 13356 17556
rect 13412 17500 13422 17556
rect 15092 17500 16380 17556
rect 16436 17500 22540 17556
rect 22596 17500 22988 17556
rect 23044 17500 23054 17556
rect 24882 17500 24892 17556
rect 24948 17500 31836 17556
rect 31892 17500 31902 17556
rect 11666 17388 11676 17444
rect 11732 17388 14252 17444
rect 14308 17388 16604 17444
rect 16660 17388 16670 17444
rect 22754 17388 22764 17444
rect 22820 17388 23212 17444
rect 23268 17388 24668 17444
rect 24724 17388 26908 17444
rect 26964 17388 28364 17444
rect 28420 17388 28430 17444
rect 23538 17276 23548 17332
rect 23604 17276 23642 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 23622 17164 23660 17220
rect 23716 17164 23726 17220
rect 24434 17164 24444 17220
rect 24500 17164 26572 17220
rect 26628 17164 28700 17220
rect 28756 17164 28766 17220
rect 8082 17052 8092 17108
rect 8148 17052 8540 17108
rect 8596 17052 15820 17108
rect 15876 17052 15886 17108
rect 16146 17052 16156 17108
rect 16212 17052 16492 17108
rect 16548 17052 16558 17108
rect 16706 17052 16716 17108
rect 16772 17052 24668 17108
rect 24724 17052 24734 17108
rect 30594 17052 30604 17108
rect 30660 17052 34188 17108
rect 34244 17052 35532 17108
rect 35588 17052 35598 17108
rect 8642 16940 8652 16996
rect 8708 16940 11116 16996
rect 11172 16940 11182 16996
rect 14998 16940 15036 16996
rect 15092 16940 15102 16996
rect 15922 16940 15932 16996
rect 15988 16940 17164 16996
rect 17220 16940 17612 16996
rect 17668 16940 17678 16996
rect 24546 16940 24556 16996
rect 24612 16940 25788 16996
rect 25844 16940 25854 16996
rect 26338 16940 26348 16996
rect 26404 16940 28140 16996
rect 28196 16940 28206 16996
rect 33394 16940 33404 16996
rect 33460 16940 34524 16996
rect 34580 16940 34590 16996
rect 6402 16828 6412 16884
rect 6468 16828 6972 16884
rect 7028 16828 7038 16884
rect 15138 16828 15148 16884
rect 15204 16828 21420 16884
rect 21476 16828 21486 16884
rect 22306 16828 22316 16884
rect 22372 16828 25564 16884
rect 25620 16828 26460 16884
rect 26516 16828 26526 16884
rect 26674 16828 26684 16884
rect 26740 16828 28588 16884
rect 28644 16828 28654 16884
rect 32498 16828 32508 16884
rect 32564 16828 33180 16884
rect 33236 16828 33852 16884
rect 33908 16828 34636 16884
rect 34692 16828 36204 16884
rect 36260 16828 36270 16884
rect 6962 16716 6972 16772
rect 7028 16716 7420 16772
rect 7476 16716 7486 16772
rect 11554 16716 11564 16772
rect 11620 16716 12124 16772
rect 12180 16716 12190 16772
rect 16146 16716 16156 16772
rect 16212 16716 16604 16772
rect 16660 16716 17388 16772
rect 17444 16716 17454 16772
rect 23650 16716 23660 16772
rect 23716 16716 24444 16772
rect 24500 16716 24510 16772
rect 25452 16660 25508 16828
rect 25666 16716 25676 16772
rect 25732 16716 28252 16772
rect 28308 16716 28318 16772
rect 7830 16604 7868 16660
rect 7924 16604 14700 16660
rect 14756 16604 17276 16660
rect 17332 16604 17342 16660
rect 25452 16604 25900 16660
rect 25956 16604 25966 16660
rect 30706 16604 30716 16660
rect 30772 16604 33964 16660
rect 34020 16604 34030 16660
rect 16706 16492 16716 16548
rect 16772 16492 24220 16548
rect 24276 16492 27132 16548
rect 27188 16492 27198 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 16818 16380 16828 16436
rect 16884 16380 19628 16436
rect 19684 16380 19694 16436
rect 24882 16380 24892 16436
rect 24948 16380 25340 16436
rect 25396 16380 25406 16436
rect 12674 16268 12684 16324
rect 12740 16268 15148 16324
rect 19506 16268 19516 16324
rect 19572 16268 20300 16324
rect 20356 16268 26684 16324
rect 26740 16268 26750 16324
rect 28130 16268 28140 16324
rect 28196 16268 29260 16324
rect 29316 16268 29326 16324
rect 15092 16212 15148 16268
rect 11778 16156 11788 16212
rect 11844 16156 13244 16212
rect 13300 16156 13310 16212
rect 15092 16156 21084 16212
rect 21140 16156 21150 16212
rect 23650 16156 23660 16212
rect 23716 16156 23772 16212
rect 23828 16156 23838 16212
rect 23986 16156 23996 16212
rect 24052 16156 25452 16212
rect 25508 16156 25518 16212
rect 26562 16156 26572 16212
rect 26628 16156 26638 16212
rect 29148 16156 29708 16212
rect 29764 16156 29774 16212
rect 4834 16044 4844 16100
rect 4900 16044 6076 16100
rect 6132 16044 6142 16100
rect 12786 16044 12796 16100
rect 12852 16044 13692 16100
rect 13748 16044 14140 16100
rect 14196 16044 18060 16100
rect 18116 16044 18126 16100
rect 20290 16044 20300 16100
rect 20356 16044 21196 16100
rect 21252 16044 21262 16100
rect 24546 16044 24556 16100
rect 24612 16044 25228 16100
rect 25284 16044 25294 16100
rect 13906 15932 13916 15988
rect 13972 15932 15036 15988
rect 15092 15932 19516 15988
rect 19572 15932 20076 15988
rect 20132 15932 20142 15988
rect 25778 15932 25788 15988
rect 25844 15932 26236 15988
rect 26292 15932 26302 15988
rect 2146 15820 2156 15876
rect 2212 15820 5740 15876
rect 5796 15820 5806 15876
rect 9650 15820 9660 15876
rect 9716 15820 13580 15876
rect 13636 15820 13646 15876
rect 16146 15820 16156 15876
rect 16212 15820 16268 15876
rect 16324 15820 16334 15876
rect 20178 15820 20188 15876
rect 20244 15820 22652 15876
rect 22708 15820 24444 15876
rect 24500 15820 24510 15876
rect 26572 15764 26628 16156
rect 29148 16100 29204 16156
rect 28242 16044 28252 16100
rect 28308 16044 29148 16100
rect 29204 16044 29214 16100
rect 27458 15932 27468 15988
rect 27524 15932 29596 15988
rect 29652 15932 31276 15988
rect 31332 15932 31342 15988
rect 7858 15708 7868 15764
rect 7924 15708 12236 15764
rect 12292 15708 12684 15764
rect 12740 15708 12750 15764
rect 26562 15708 26572 15764
rect 26628 15708 26796 15764
rect 26852 15708 26862 15764
rect 27010 15708 27020 15764
rect 27076 15708 29148 15764
rect 29204 15708 29214 15764
rect 29922 15708 29932 15764
rect 29988 15708 30716 15764
rect 30772 15708 30782 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 22866 15596 22876 15652
rect 22932 15596 23548 15652
rect 23604 15596 23614 15652
rect 26226 15596 26236 15652
rect 26292 15596 30940 15652
rect 30996 15596 31388 15652
rect 31444 15596 31454 15652
rect 4050 15484 4060 15540
rect 4116 15484 6076 15540
rect 6132 15484 6142 15540
rect 13794 15484 13804 15540
rect 13860 15484 14476 15540
rect 14532 15484 14542 15540
rect 24770 15484 24780 15540
rect 24836 15484 27244 15540
rect 27300 15484 27310 15540
rect 28588 15484 35756 15540
rect 35812 15484 36316 15540
rect 36372 15484 36382 15540
rect 28588 15428 28644 15484
rect 7970 15372 7980 15428
rect 8036 15372 8428 15428
rect 8484 15372 13580 15428
rect 13636 15372 14924 15428
rect 14980 15372 14990 15428
rect 17714 15372 17724 15428
rect 17780 15372 21308 15428
rect 21364 15372 22428 15428
rect 22484 15372 22494 15428
rect 23762 15372 23772 15428
rect 23828 15372 25676 15428
rect 25732 15372 25742 15428
rect 26460 15372 28588 15428
rect 28644 15372 28654 15428
rect 29026 15372 29036 15428
rect 29092 15372 30940 15428
rect 30996 15372 31724 15428
rect 31780 15372 31790 15428
rect 35410 15372 35420 15428
rect 35476 15372 37884 15428
rect 37940 15372 37950 15428
rect 26460 15316 26516 15372
rect 9986 15260 9996 15316
rect 10052 15260 12572 15316
rect 12628 15260 12638 15316
rect 13234 15260 13244 15316
rect 13300 15260 16716 15316
rect 16772 15260 16782 15316
rect 24546 15260 24556 15316
rect 24612 15260 26516 15316
rect 26572 15260 28252 15316
rect 28308 15260 28318 15316
rect 26572 15204 26628 15260
rect 8372 15148 8540 15204
rect 8596 15148 9100 15204
rect 9156 15148 11788 15204
rect 11844 15148 11854 15204
rect 21522 15148 21532 15204
rect 21588 15148 22988 15204
rect 23044 15148 26628 15204
rect 26786 15148 26796 15204
rect 26852 15148 27132 15204
rect 27188 15148 27198 15204
rect 29474 15148 29484 15204
rect 29540 15148 29932 15204
rect 29988 15148 29998 15204
rect 8372 15092 8428 15148
rect 1810 15036 1820 15092
rect 1876 15036 2828 15092
rect 2884 15036 5068 15092
rect 5124 15036 5852 15092
rect 5908 15036 6972 15092
rect 7028 15036 8428 15092
rect 25554 15036 25564 15092
rect 25620 15036 28028 15092
rect 28084 15036 28094 15092
rect 28466 15036 28476 15092
rect 28532 15036 35196 15092
rect 35252 15036 35262 15092
rect 23874 14924 23884 14980
rect 23940 14924 27580 14980
rect 27636 14924 27646 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 26226 14812 26236 14868
rect 26292 14812 27244 14868
rect 27300 14812 27310 14868
rect 8754 14700 8764 14756
rect 8820 14700 11116 14756
rect 11172 14700 11182 14756
rect 16818 14700 16828 14756
rect 16884 14700 22204 14756
rect 22260 14700 22270 14756
rect 23202 14700 23212 14756
rect 23268 14700 23884 14756
rect 23940 14700 27020 14756
rect 27076 14700 27468 14756
rect 27524 14700 28252 14756
rect 28308 14700 28318 14756
rect 22204 14644 22260 14700
rect 22204 14588 24108 14644
rect 24164 14588 26236 14644
rect 26292 14588 26302 14644
rect 12562 14476 12572 14532
rect 12628 14476 13132 14532
rect 13188 14476 23548 14532
rect 23604 14476 25564 14532
rect 25620 14476 25630 14532
rect 12674 14364 12684 14420
rect 12740 14364 13468 14420
rect 13524 14364 13534 14420
rect 26114 14364 26124 14420
rect 26180 14364 26460 14420
rect 26516 14364 26526 14420
rect 27010 14364 27020 14420
rect 27076 14364 27086 14420
rect 30818 14364 30828 14420
rect 30884 14364 33292 14420
rect 33348 14364 33358 14420
rect 12002 14252 12012 14308
rect 12068 14252 13916 14308
rect 13972 14252 13982 14308
rect 14690 14252 14700 14308
rect 14756 14252 15148 14308
rect 15204 14252 15214 14308
rect 25890 14252 25900 14308
rect 25956 14252 26236 14308
rect 26292 14252 26302 14308
rect 27020 14196 27076 14364
rect 10882 14140 10892 14196
rect 10948 14140 12236 14196
rect 12292 14140 12302 14196
rect 27020 14140 33180 14196
rect 33236 14140 33246 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 6178 14028 6188 14084
rect 6244 14028 9660 14084
rect 9716 14028 9726 14084
rect 20402 14028 20412 14084
rect 20468 14028 21196 14084
rect 21252 14028 21262 14084
rect 24994 13916 25004 13972
rect 25060 13916 27020 13972
rect 27076 13916 27086 13972
rect 10770 13804 10780 13860
rect 10836 13804 11676 13860
rect 11732 13804 15596 13860
rect 15652 13804 17220 13860
rect 6066 13692 6076 13748
rect 6132 13692 7084 13748
rect 7140 13692 7980 13748
rect 8036 13692 8046 13748
rect 8306 13692 8316 13748
rect 8372 13692 9772 13748
rect 9828 13692 9838 13748
rect 12898 13692 12908 13748
rect 12964 13692 15820 13748
rect 15876 13692 15886 13748
rect 17164 13636 17220 13804
rect 19058 13692 19068 13748
rect 19124 13692 21868 13748
rect 21924 13692 21934 13748
rect 22642 13692 22652 13748
rect 22708 13692 26460 13748
rect 26516 13692 26526 13748
rect 27794 13692 27804 13748
rect 27860 13692 35644 13748
rect 35700 13692 35710 13748
rect 17164 13580 19516 13636
rect 19572 13580 20300 13636
rect 20356 13580 20366 13636
rect 9538 13468 9548 13524
rect 9604 13468 12684 13524
rect 12740 13468 12750 13524
rect 23958 13468 23996 13524
rect 24052 13468 24062 13524
rect 25302 13468 25340 13524
rect 25396 13468 25406 13524
rect 26450 13468 26460 13524
rect 26516 13468 27020 13524
rect 27076 13468 27086 13524
rect 18946 13356 18956 13412
rect 19012 13356 19628 13412
rect 19684 13356 22204 13412
rect 22260 13356 22270 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 5394 13244 5404 13300
rect 5460 13244 8988 13300
rect 9044 13244 9054 13300
rect 2930 13132 2940 13188
rect 2996 13132 5740 13188
rect 5796 13132 5806 13188
rect 12450 13132 12460 13188
rect 12516 13132 13020 13188
rect 13076 13132 14364 13188
rect 14420 13132 14430 13188
rect 20290 13132 20300 13188
rect 20356 13132 24332 13188
rect 24388 13132 24398 13188
rect 4610 13020 4620 13076
rect 4676 13020 6076 13076
rect 6132 13020 11788 13076
rect 11844 13020 11854 13076
rect 12562 13020 12572 13076
rect 12628 13020 12908 13076
rect 12964 13020 12974 13076
rect 19730 13020 19740 13076
rect 19796 13020 21308 13076
rect 21364 13020 21374 13076
rect 23538 13020 23548 13076
rect 23604 13020 23884 13076
rect 23940 13020 23950 13076
rect 25442 13020 25452 13076
rect 25508 13020 26124 13076
rect 26180 13020 26190 13076
rect 3714 12908 3724 12964
rect 3780 12908 5068 12964
rect 5124 12908 5134 12964
rect 10770 12908 10780 12964
rect 10836 12908 13132 12964
rect 13188 12908 13198 12964
rect 23538 12908 23548 12964
rect 23604 12908 23772 12964
rect 23828 12908 23838 12964
rect 23986 12908 23996 12964
rect 24052 12908 24090 12964
rect 27346 12908 27356 12964
rect 27412 12908 29148 12964
rect 29204 12908 29214 12964
rect 33058 12908 33068 12964
rect 33124 12908 33852 12964
rect 33908 12908 36316 12964
rect 36372 12908 36382 12964
rect 9762 12796 9772 12852
rect 9828 12796 11564 12852
rect 11620 12796 11630 12852
rect 12002 12796 12012 12852
rect 12068 12796 13692 12852
rect 13748 12796 14028 12852
rect 14084 12796 14094 12852
rect 21858 12796 21868 12852
rect 21924 12796 23324 12852
rect 23380 12796 25228 12852
rect 25284 12796 25294 12852
rect 25452 12796 27132 12852
rect 27188 12796 27198 12852
rect 28578 12796 28588 12852
rect 28644 12796 31276 12852
rect 31332 12796 31342 12852
rect 25452 12740 25508 12796
rect 22530 12684 22540 12740
rect 22596 12684 25508 12740
rect 25778 12684 25788 12740
rect 25844 12684 30268 12740
rect 30324 12684 31500 12740
rect 31556 12684 31566 12740
rect 35858 12684 35868 12740
rect 35924 12684 38444 12740
rect 38500 12684 38510 12740
rect 24546 12572 24556 12628
rect 24612 12572 26236 12628
rect 26292 12572 32060 12628
rect 32116 12572 33740 12628
rect 33796 12572 33806 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 23650 12460 23660 12516
rect 23716 12460 24444 12516
rect 24500 12460 24510 12516
rect 28354 12460 28364 12516
rect 28420 12460 29596 12516
rect 29652 12460 29662 12516
rect 14466 12348 14476 12404
rect 14532 12348 15596 12404
rect 15652 12348 16044 12404
rect 16100 12348 16110 12404
rect 19282 12348 19292 12404
rect 19348 12348 19964 12404
rect 20020 12348 20030 12404
rect 23538 12348 23548 12404
rect 23604 12348 24668 12404
rect 24724 12348 24734 12404
rect 25778 12348 25788 12404
rect 25844 12348 26236 12404
rect 26292 12348 26302 12404
rect 27458 12348 27468 12404
rect 27524 12348 28252 12404
rect 28308 12348 28318 12404
rect 8978 12236 8988 12292
rect 9044 12236 14028 12292
rect 14084 12236 14094 12292
rect 29138 12236 29148 12292
rect 29204 12236 30492 12292
rect 30548 12236 30558 12292
rect 32498 12236 32508 12292
rect 32564 12236 33852 12292
rect 33908 12236 33918 12292
rect 1810 12124 1820 12180
rect 1876 12124 2380 12180
rect 2436 12124 5068 12180
rect 5124 12124 5628 12180
rect 5684 12124 6188 12180
rect 6244 12124 8428 12180
rect 8484 12124 9212 12180
rect 9268 12124 9278 12180
rect 21522 12124 21532 12180
rect 21588 12124 23100 12180
rect 23156 12124 23166 12180
rect 23762 12124 23772 12180
rect 23828 12124 28252 12180
rect 28308 12124 28318 12180
rect 8372 12012 8988 12068
rect 9044 12012 9054 12068
rect 11554 12012 11564 12068
rect 11620 12012 12236 12068
rect 12292 12012 12302 12068
rect 12562 12012 12572 12068
rect 12628 12012 13468 12068
rect 13524 12012 13534 12068
rect 34178 12012 34188 12068
rect 34244 12012 35980 12068
rect 36036 12012 36046 12068
rect 8372 11956 8428 12012
rect 7634 11900 7644 11956
rect 7700 11900 8428 11956
rect 24098 11788 24108 11844
rect 24164 11788 31724 11844
rect 31780 11788 31790 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 9650 11676 9660 11732
rect 9716 11676 11676 11732
rect 11732 11676 11742 11732
rect 28466 11676 28476 11732
rect 28532 11676 31948 11732
rect 32004 11676 32014 11732
rect 12226 11564 12236 11620
rect 12292 11564 13244 11620
rect 13300 11564 13310 11620
rect 19954 11564 19964 11620
rect 20020 11564 20748 11620
rect 20804 11564 21644 11620
rect 21700 11564 21710 11620
rect 29922 11564 29932 11620
rect 29988 11564 33516 11620
rect 33572 11564 33582 11620
rect 20066 11452 20076 11508
rect 20132 11452 21420 11508
rect 21476 11452 24108 11508
rect 24164 11452 25676 11508
rect 25732 11452 26236 11508
rect 26292 11452 26302 11508
rect 20626 11340 20636 11396
rect 20692 11340 22204 11396
rect 22260 11340 22270 11396
rect 26898 11340 26908 11396
rect 26964 11340 34356 11396
rect 34300 11284 34356 11340
rect 6738 11228 6748 11284
rect 6804 11228 8204 11284
rect 8260 11228 8270 11284
rect 20290 11228 20300 11284
rect 20356 11228 22876 11284
rect 22932 11228 22942 11284
rect 25554 11228 25564 11284
rect 25620 11228 28700 11284
rect 28756 11228 28766 11284
rect 31714 11228 31724 11284
rect 31780 11228 32060 11284
rect 32116 11228 32126 11284
rect 34290 11228 34300 11284
rect 34356 11228 35756 11284
rect 35812 11228 35822 11284
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 11554 10780 11564 10836
rect 11620 10780 12124 10836
rect 12180 10780 12190 10836
rect 26562 10780 26572 10836
rect 26628 10780 27132 10836
rect 27188 10780 27198 10836
rect 14690 10668 14700 10724
rect 14756 10668 15372 10724
rect 15428 10668 15438 10724
rect 26786 10668 26796 10724
rect 26852 10668 28588 10724
rect 28644 10668 28654 10724
rect 10882 10556 10892 10612
rect 10948 10556 11788 10612
rect 11844 10556 16548 10612
rect 16706 10556 16716 10612
rect 16772 10556 17500 10612
rect 17556 10556 17566 10612
rect 18610 10556 18620 10612
rect 18676 10556 19740 10612
rect 19796 10556 19806 10612
rect 16492 10500 16548 10556
rect 10994 10444 11004 10500
rect 11060 10444 12460 10500
rect 12516 10444 15260 10500
rect 15316 10444 15326 10500
rect 16492 10444 17724 10500
rect 17780 10444 19516 10500
rect 19572 10444 19582 10500
rect 15698 10332 15708 10388
rect 15764 10332 17164 10388
rect 17220 10332 17836 10388
rect 17892 10332 17902 10388
rect 29810 10332 29820 10388
rect 29876 10332 31388 10388
rect 31444 10332 35532 10388
rect 35588 10332 35598 10388
rect 16034 10220 16044 10276
rect 16100 10220 24668 10276
rect 24724 10220 25564 10276
rect 25620 10220 25630 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19282 9996 19292 10052
rect 19348 9996 22092 10052
rect 22148 9996 24108 10052
rect 24164 9996 24174 10052
rect 11218 9884 11228 9940
rect 11284 9884 12012 9940
rect 12068 9884 12078 9940
rect 26898 9884 26908 9940
rect 26964 9884 27244 9940
rect 27300 9884 27580 9940
rect 27636 9884 27646 9940
rect 28914 9884 28924 9940
rect 28980 9884 29820 9940
rect 29876 9884 30604 9940
rect 30660 9884 30670 9940
rect 14018 9772 14028 9828
rect 14084 9772 15708 9828
rect 15764 9772 15774 9828
rect 17714 9772 17724 9828
rect 17780 9772 19740 9828
rect 19796 9772 21532 9828
rect 21588 9772 21598 9828
rect 8530 9660 8540 9716
rect 8596 9660 12572 9716
rect 12628 9660 12638 9716
rect 11554 9548 11564 9604
rect 11620 9548 14252 9604
rect 14308 9548 14318 9604
rect 28242 9548 28252 9604
rect 28308 9548 29148 9604
rect 29204 9548 29214 9604
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 24770 9212 24780 9268
rect 24836 9212 25340 9268
rect 25396 9212 25406 9268
rect 13346 9100 13356 9156
rect 13412 9100 18508 9156
rect 18564 9100 18574 9156
rect 23202 9100 23212 9156
rect 23268 9100 24332 9156
rect 24388 9100 24398 9156
rect 5730 8988 5740 9044
rect 5796 8988 8428 9044
rect 8484 8988 8988 9044
rect 9044 8988 9054 9044
rect 9874 8988 9884 9044
rect 9940 8988 10444 9044
rect 10500 8988 10510 9044
rect 21634 8988 21644 9044
rect 21700 8988 23324 9044
rect 23380 8988 23390 9044
rect 7410 8876 7420 8932
rect 7476 8876 8540 8932
rect 8596 8876 8606 8932
rect 18386 8876 18396 8932
rect 18452 8876 19292 8932
rect 19348 8876 19358 8932
rect 22530 8652 22540 8708
rect 22596 8652 23100 8708
rect 23156 8652 27916 8708
rect 27972 8652 27982 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 20850 8540 20860 8596
rect 20916 8540 25564 8596
rect 25620 8540 26012 8596
rect 26068 8540 26078 8596
rect 25330 8428 25340 8484
rect 25396 8428 27412 8484
rect 21522 8316 21532 8372
rect 21588 8316 22316 8372
rect 22372 8316 23100 8372
rect 23156 8316 23166 8372
rect 27356 8260 27412 8428
rect 20738 8204 20748 8260
rect 20804 8204 21644 8260
rect 21700 8204 23324 8260
rect 23380 8204 23996 8260
rect 24052 8204 24062 8260
rect 27346 8204 27356 8260
rect 27412 8204 29932 8260
rect 29988 8204 29998 8260
rect 19506 8092 19516 8148
rect 19572 8092 20076 8148
rect 20132 8092 21980 8148
rect 22036 8092 22046 8148
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 12114 7756 12124 7812
rect 12180 7756 14140 7812
rect 14196 7756 18060 7812
rect 18116 7756 18126 7812
rect 14662 7644 14700 7700
rect 14756 7644 14766 7700
rect 21970 7644 21980 7700
rect 22036 7644 22876 7700
rect 22932 7644 25676 7700
rect 25732 7644 25742 7700
rect 18050 7532 18060 7588
rect 18116 7532 18844 7588
rect 18900 7532 18910 7588
rect 26674 7532 26684 7588
rect 26740 7532 28252 7588
rect 28308 7532 28318 7588
rect 16706 7420 16716 7476
rect 16772 7420 17500 7476
rect 17556 7420 17566 7476
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 22082 6860 22092 6916
rect 22148 6860 23660 6916
rect 23716 6860 23726 6916
rect 26562 6860 26572 6916
rect 26628 6860 27468 6916
rect 27524 6860 27534 6916
rect 27234 6748 27244 6804
rect 27300 6748 28588 6804
rect 28644 6748 28654 6804
rect 9314 6636 9324 6692
rect 9380 6636 11788 6692
rect 11844 6636 12684 6692
rect 12740 6636 15260 6692
rect 15316 6636 15326 6692
rect 22082 6636 22092 6692
rect 22148 6636 22540 6692
rect 22596 6636 24668 6692
rect 24724 6636 24734 6692
rect 15810 6524 15820 6580
rect 15876 6524 17724 6580
rect 17780 6524 18508 6580
rect 18564 6524 18574 6580
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 22194 5964 22204 6020
rect 22260 5964 23324 6020
rect 23380 5964 23390 6020
rect 21298 5628 21308 5684
rect 21364 5628 22764 5684
rect 22820 5628 22830 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 23762 5180 23772 5236
rect 23828 5180 25340 5236
rect 25396 5180 26796 5236
rect 26852 5180 26862 5236
rect 21634 5068 21644 5124
rect 21700 5068 22764 5124
rect 22820 5068 22830 5124
rect 20514 4956 20524 5012
rect 20580 4956 22092 5012
rect 22148 4956 22158 5012
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 42476 50652 42532 50708
rect 42924 50652 42980 50708
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 18396 47180 18452 47236
rect 15036 47068 15092 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 13692 46844 13748 46900
rect 25340 46732 25396 46788
rect 13692 46508 13748 46564
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 24556 46172 24612 46228
rect 15260 45500 15316 45556
rect 21644 45500 21700 45556
rect 25228 45500 25284 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 20300 45276 20356 45332
rect 24556 45164 24612 45220
rect 17612 44716 17668 44772
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 4284 44156 4340 44212
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 21644 43484 21700 43540
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 18732 42924 18788 42980
rect 24556 42700 24612 42756
rect 25340 42700 25396 42756
rect 27916 42364 27972 42420
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 19404 42252 19460 42308
rect 15260 42140 15316 42196
rect 21980 42028 22036 42084
rect 17052 41804 17108 41860
rect 18732 41580 18788 41636
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 21980 41468 22036 41524
rect 24556 41356 24612 41412
rect 14252 41244 14308 41300
rect 4284 41132 4340 41188
rect 17276 41020 17332 41076
rect 17052 40908 17108 40964
rect 19180 40908 19236 40964
rect 20300 40796 20356 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 14812 40572 14868 40628
rect 27916 40460 27972 40516
rect 16716 40348 16772 40404
rect 19180 40348 19236 40404
rect 14252 40236 14308 40292
rect 19404 40124 19460 40180
rect 17612 40012 17668 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 18396 39900 18452 39956
rect 14252 39564 14308 39620
rect 45388 39564 45444 39620
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 15036 39004 15092 39060
rect 14812 38892 14868 38948
rect 45388 39004 45444 39060
rect 15148 38892 15204 38948
rect 48076 38892 48132 38948
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 15148 38556 15204 38612
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 14812 37996 14868 38052
rect 45388 37884 45444 37940
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 19516 37548 19572 37604
rect 48188 36988 48244 37044
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 17276 36652 17332 36708
rect 16716 36540 16772 36596
rect 19516 36428 19572 36484
rect 48188 36316 48244 36372
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 25228 35868 25284 35924
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 48076 35644 48132 35700
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 45164 34860 45220 34916
rect 45276 34524 45332 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 45500 34300 45556 34356
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 16940 33404 16996 33460
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 43484 32844 43540 32900
rect 43484 32172 43540 32228
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 36652 31948 36708 32004
rect 18844 31724 18900 31780
rect 44492 31612 44548 31668
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 48636 31164 48692 31220
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 43484 29932 43540 29988
rect 46284 29932 46340 29988
rect 44492 29820 44548 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 45500 29372 45556 29428
rect 43708 29260 43764 29316
rect 45164 29260 45220 29316
rect 45276 29148 45332 29204
rect 46508 29148 46564 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 16940 28700 16996 28756
rect 46284 28700 46340 28756
rect 48188 28588 48244 28644
rect 18956 28364 19012 28420
rect 46508 28364 46564 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 8316 27580 8372 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 8428 26908 8484 26964
rect 8428 26796 8484 26852
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 48188 26460 48244 26516
rect 18956 25900 19012 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 18844 25228 18900 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 48636 25228 48692 25284
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 8316 25004 8372 25060
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 36652 24220 36708 24276
rect 43708 24220 43764 24276
rect 18844 23772 18900 23828
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 25340 22876 25396 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 14476 22540 14532 22596
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 16156 21308 16212 21364
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 14924 19964 14980 20020
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19404 19180 19460 19236
rect 7868 18844 7924 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 6972 18620 7028 18676
rect 19404 18060 19460 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 23548 17276 23604 17332
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 23660 17164 23716 17220
rect 16156 17052 16212 17108
rect 15036 16940 15092 16996
rect 6972 16716 7028 16772
rect 7868 16604 7924 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 23660 16156 23716 16212
rect 15036 15932 15092 15988
rect 16156 15820 16212 15876
rect 28252 16044 28308 16100
rect 26796 15708 26852 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 14476 15484 14532 15540
rect 26796 15148 26852 15204
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 23996 13468 24052 13524
rect 25340 13468 25396 13524
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 23548 12908 23604 12964
rect 23996 12908 24052 12964
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 28252 12124 28308 12180
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 14700 7644 14756 7700
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 18396 47236 18452 47246
rect 15036 47124 15092 47134
rect 13692 46900 13748 46910
rect 13692 46564 13748 46844
rect 13692 46498 13748 46508
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4284 44212 4340 44222
rect 4284 41188 4340 44156
rect 4284 41122 4340 41132
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 14252 41300 14308 41310
rect 14252 40292 14308 41244
rect 14252 39620 14308 40236
rect 14252 39554 14308 39564
rect 14812 40628 14868 40638
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 14812 38948 14868 40572
rect 15036 39060 15092 47068
rect 15260 45556 15316 45566
rect 15260 42196 15316 45500
rect 15260 42130 15316 42140
rect 17612 44772 17668 44782
rect 17052 41860 17108 41870
rect 17052 40964 17108 41804
rect 17052 40898 17108 40908
rect 17276 41076 17332 41086
rect 15036 38994 15092 39004
rect 16716 40404 16772 40414
rect 14812 38052 14868 38892
rect 15148 38948 15204 38958
rect 15148 38612 15204 38892
rect 15148 38546 15204 38556
rect 14812 37986 14868 37996
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 16716 36596 16772 40348
rect 17276 36708 17332 41020
rect 17612 40068 17668 44716
rect 17612 40002 17668 40012
rect 18396 39956 18452 47180
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 42476 50708 42532 50718
rect 42924 50708 42980 50718
rect 42532 50652 42924 50698
rect 42476 50642 42980 50652
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 25340 46788 25396 46798
rect 24556 46228 24612 46238
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 21644 45556 21700 45566
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 18732 42980 18788 42990
rect 18732 41636 18788 42924
rect 19808 42364 20128 43876
rect 18732 41570 18788 41580
rect 19404 42308 19460 42318
rect 19180 40964 19236 40974
rect 19180 40404 19236 40908
rect 19180 40338 19236 40348
rect 19404 40180 19460 42252
rect 19404 40114 19460 40124
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 20300 45332 20356 45342
rect 20300 40852 20356 45276
rect 21644 43540 21700 45500
rect 24556 45220 24612 46172
rect 24556 45154 24612 45164
rect 25228 45556 25284 45566
rect 21644 43474 21700 43484
rect 24556 42756 24612 42766
rect 21980 42084 22036 42094
rect 21980 41524 22036 42028
rect 21980 41458 22036 41468
rect 24556 41412 24612 42700
rect 24556 41346 24612 41356
rect 20300 40786 20356 40796
rect 18396 39890 18452 39900
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 17276 36642 17332 36652
rect 19516 37604 19572 37614
rect 16716 36530 16772 36540
rect 19516 36484 19572 37548
rect 19516 36418 19572 36428
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 25228 35924 25284 45500
rect 25340 42756 25396 46732
rect 25340 42690 25396 42700
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 27916 42420 27972 42430
rect 27916 40516 27972 42364
rect 27916 40450 27972 40460
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 25228 35858 25284 35868
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 45388 39620 45444 39630
rect 45388 39060 45444 39564
rect 45388 37940 45444 39004
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 45388 37874 45444 37884
rect 48076 38948 48132 38958
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 16940 33460 16996 33470
rect 16940 28756 16996 33404
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 16940 28690 16996 28700
rect 18844 31780 18900 31790
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 8316 27636 8372 27646
rect 8316 25060 8372 27580
rect 8428 26964 8484 26974
rect 8428 26852 8484 26908
rect 8428 26786 8484 26796
rect 8316 24994 8372 25004
rect 18844 25284 18900 31724
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 18956 28420 19012 28430
rect 18956 25956 19012 28364
rect 18956 25890 19012 25900
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 18844 23828 18900 25228
rect 18844 23762 18900 23772
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 14476 22596 14532 22606
rect 7868 18900 7924 18910
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 6972 18676 7028 18686
rect 6972 16772 7028 18620
rect 6972 16706 7028 16716
rect 7868 16660 7924 18844
rect 7868 16594 7924 16604
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 14476 15540 14532 22540
rect 19808 21980 20128 23492
rect 35168 35308 35488 36820
rect 48076 35700 48132 38892
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 48188 37044 48244 37054
rect 48188 36372 48244 36988
rect 48188 36306 48244 36316
rect 48076 35634 48132 35644
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 45164 34916 45220 34926
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 43484 32900 43540 32910
rect 43484 32228 43540 32844
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 16156 21364 16212 21374
rect 14476 15474 14532 15484
rect 14924 20020 14980 20030
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 14924 8428 14980 19964
rect 16156 17108 16212 21308
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19404 19236 19460 19246
rect 19404 18116 19460 19180
rect 19404 18050 19460 18060
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 15036 16996 15092 17006
rect 15036 15988 15092 16940
rect 15036 15922 15092 15932
rect 16156 15876 16212 17052
rect 16156 15810 16212 15820
rect 19808 17276 20128 18788
rect 25340 22932 25396 22942
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 14700 8372 14980 8428
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 23548 17332 23604 17342
rect 23548 12964 23604 17276
rect 23660 17220 23716 17230
rect 23660 16212 23716 17164
rect 23660 16146 23716 16156
rect 23548 12898 23604 12908
rect 23996 13524 24052 13534
rect 23996 12964 24052 13468
rect 25340 13524 25396 22876
rect 35168 22764 35488 24276
rect 36652 32004 36708 32014
rect 36652 24276 36708 31948
rect 43484 29988 43540 32172
rect 43484 29922 43540 29932
rect 44492 31668 44548 31678
rect 44492 29876 44548 31612
rect 44492 29810 44548 29820
rect 36652 24210 36708 24220
rect 43708 29316 43764 29326
rect 43708 24276 43764 29260
rect 45164 29316 45220 34860
rect 45164 29250 45220 29260
rect 45276 34580 45332 34590
rect 45276 29204 45332 34524
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 45500 34356 45556 34366
rect 45500 29428 45556 34300
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 48636 31220 48692 31230
rect 45500 29362 45556 29372
rect 46284 29988 46340 29998
rect 45276 29138 45332 29148
rect 46284 28756 46340 29932
rect 46284 28690 46340 28700
rect 46508 29204 46564 29214
rect 46508 28420 46564 29148
rect 46508 28354 46564 28364
rect 48188 28644 48244 28654
rect 48188 26516 48244 28588
rect 48188 26450 48244 26460
rect 48636 25284 48692 31164
rect 48636 25218 48692 25228
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 43708 24210 43764 24220
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 28252 16100 28308 16110
rect 26796 15764 26852 15774
rect 26796 15204 26852 15708
rect 26796 15138 26852 15148
rect 25340 13458 25396 13468
rect 23996 12898 24052 12908
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 28252 12180 28308 16044
rect 28252 12114 28308 12124
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 14700 7700 14756 8372
rect 14700 7634 14756 7644
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1287_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42448 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1288_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 52080 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1289_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 47936 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1290_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47824 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1291_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 50624 0 -1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1292_
timestamp 1698431365
transform -1 0 44128 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1293_
timestamp 1698431365
transform 1 0 47936 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1294_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45472 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1295_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46368 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1296_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 49056 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1297_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48048 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1298_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46368 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1299_
timestamp 1698431365
transform -1 0 43456 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1300_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42112 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1301_
timestamp 1698431365
transform 1 0 41888 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1302_
timestamp 1698431365
transform -1 0 39536 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1303_
timestamp 1698431365
transform -1 0 46816 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1304_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42672 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1305_
timestamp 1698431365
transform -1 0 40208 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1306_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41776 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1307_
timestamp 1698431365
transform -1 0 43904 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1308_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42784 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1309_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37520 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1310_
timestamp 1698431365
transform 1 0 44688 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1311_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42784 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1312_
timestamp 1698431365
transform -1 0 41888 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1313_
timestamp 1698431365
transform 1 0 41216 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1314_
timestamp 1698431365
transform -1 0 44128 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1315_
timestamp 1698431365
transform 1 0 42896 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1316_
timestamp 1698431365
transform -1 0 41664 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1317_
timestamp 1698431365
transform -1 0 39536 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1318_
timestamp 1698431365
transform 1 0 41664 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1319_
timestamp 1698431365
transform 1 0 39200 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1320_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38640 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1321_
timestamp 1698431365
transform -1 0 38192 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1322_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40432 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1323_
timestamp 1698431365
transform -1 0 40096 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1324_
timestamp 1698431365
transform -1 0 40320 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1325_
timestamp 1698431365
transform 1 0 39760 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1326_
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1327_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39312 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1698431365
transform 1 0 43568 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1329_
timestamp 1698431365
transform 1 0 37856 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1330_
timestamp 1698431365
transform 1 0 39536 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1331_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39760 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1332_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38304 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1333_
timestamp 1698431365
transform -1 0 32704 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1334_
timestamp 1698431365
transform -1 0 38192 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1335_
timestamp 1698431365
transform -1 0 36176 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1336_
timestamp 1698431365
transform -1 0 35728 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1337_
timestamp 1698431365
transform -1 0 40544 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1338_
timestamp 1698431365
transform -1 0 35952 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1339_
timestamp 1698431365
transform -1 0 41664 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1340_
timestamp 1698431365
transform -1 0 36736 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1341_
timestamp 1698431365
transform -1 0 34608 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1342_
timestamp 1698431365
transform 1 0 34496 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1343_
timestamp 1698431365
transform -1 0 39200 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1344_
timestamp 1698431365
transform -1 0 36288 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1345_
timestamp 1698431365
transform 1 0 36736 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1346_
timestamp 1698431365
transform 1 0 35728 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1347_
timestamp 1698431365
transform -1 0 36400 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1348_
timestamp 1698431365
transform 1 0 11536 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1349_
timestamp 1698431365
transform 1 0 29344 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1350_
timestamp 1698431365
transform 1 0 31696 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1351_
timestamp 1698431365
transform -1 0 34048 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1352_
timestamp 1698431365
transform 1 0 12208 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1353_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14336 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1354_
timestamp 1698431365
transform 1 0 11648 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1355_
timestamp 1698431365
transform 1 0 13552 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1356_
timestamp 1698431365
transform -1 0 19376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1357_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17024 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1358_
timestamp 1698431365
transform 1 0 11088 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1359_
timestamp 1698431365
transform -1 0 11984 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1360_
timestamp 1698431365
transform 1 0 14560 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1361_
timestamp 1698431365
transform 1 0 12432 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1362_
timestamp 1698431365
transform 1 0 10640 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1363_
timestamp 1698431365
transform -1 0 16128 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1364_
timestamp 1698431365
transform 1 0 14448 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1365_
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1366_
timestamp 1698431365
transform 1 0 12544 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1367_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1368_
timestamp 1698431365
transform -1 0 28000 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1369_
timestamp 1698431365
transform 1 0 20048 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1370_
timestamp 1698431365
transform 1 0 20496 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1371_
timestamp 1698431365
transform -1 0 19264 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1372_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19264 0 -1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1373_
timestamp 1698431365
transform 1 0 18368 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1374_
timestamp 1698431365
transform -1 0 18816 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1375_
timestamp 1698431365
transform 1 0 16128 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1376_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13104 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1377_
timestamp 1698431365
transform -1 0 18816 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1378_
timestamp 1698431365
transform -1 0 13104 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1379_
timestamp 1698431365
transform 1 0 11424 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1380_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16912 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1381_
timestamp 1698431365
transform 1 0 12096 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1382_
timestamp 1698431365
transform -1 0 19488 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1383_
timestamp 1698431365
transform 1 0 11088 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1384_
timestamp 1698431365
transform -1 0 12096 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1385_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1386_
timestamp 1698431365
transform 1 0 12544 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1387_
timestamp 1698431365
transform -1 0 32032 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1388_
timestamp 1698431365
transform 1 0 30016 0 -1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1389_
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1390_
timestamp 1698431365
transform -1 0 17024 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1391_
timestamp 1698431365
transform -1 0 19264 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1392_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21840 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1393_
timestamp 1698431365
transform -1 0 17696 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1394_
timestamp 1698431365
transform 1 0 22736 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1395_
timestamp 1698431365
transform -1 0 15904 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1396_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15680 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1397_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24080 0 1 31360
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1398_
timestamp 1698431365
transform 1 0 26208 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1399_
timestamp 1698431365
transform -1 0 27664 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1400_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26880 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1401_
timestamp 1698431365
transform -1 0 24752 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1402_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22624 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1403_
timestamp 1698431365
transform -1 0 24416 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1404_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26320 0 1 29792
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1405_
timestamp 1698431365
transform -1 0 18480 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1406_
timestamp 1698431365
transform 1 0 15904 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1407_
timestamp 1698431365
transform 1 0 18256 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1408_
timestamp 1698431365
transform 1 0 17584 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1409_
timestamp 1698431365
transform -1 0 19488 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1410_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 31360
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1411_
timestamp 1698431365
transform -1 0 18816 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1412_
timestamp 1698431365
transform -1 0 22176 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1413_
timestamp 1698431365
transform 1 0 22736 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1414_
timestamp 1698431365
transform -1 0 17248 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1415_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1416_
timestamp 1698431365
transform 1 0 27664 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1417_
timestamp 1698431365
transform 1 0 15680 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1418_
timestamp 1698431365
transform -1 0 16912 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1419_
timestamp 1698431365
transform 1 0 22848 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1420_
timestamp 1698431365
transform 1 0 29680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1421_
timestamp 1698431365
transform 1 0 26992 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1422_
timestamp 1698431365
transform -1 0 30128 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1423_
timestamp 1698431365
transform 1 0 22176 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1424_
timestamp 1698431365
transform 1 0 23072 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1425_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30128 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1426_
timestamp 1698431365
transform 1 0 16352 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1427_
timestamp 1698431365
transform -1 0 27552 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1428_
timestamp 1698431365
transform 1 0 35392 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1429_
timestamp 1698431365
transform -1 0 29456 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1430_
timestamp 1698431365
transform -1 0 26880 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1431_
timestamp 1698431365
transform -1 0 32480 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1432_
timestamp 1698431365
transform -1 0 29232 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1433_
timestamp 1698431365
transform -1 0 16464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1434_
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1435_
timestamp 1698431365
transform -1 0 28000 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1436_
timestamp 1698431365
transform -1 0 16352 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1437_
timestamp 1698431365
transform -1 0 25200 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1438_
timestamp 1698431365
transform 1 0 34944 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1439_
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1440_
timestamp 1698431365
transform 1 0 27888 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1441_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1442_
timestamp 1698431365
transform -1 0 28672 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1443_
timestamp 1698431365
transform 1 0 23632 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1444_
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1445_
timestamp 1698431365
transform 1 0 24192 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1446_
timestamp 1698431365
transform 1 0 23072 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1447_
timestamp 1698431365
transform 1 0 23408 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1448_
timestamp 1698431365
transform 1 0 16352 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1449_
timestamp 1698431365
transform -1 0 24304 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1450_
timestamp 1698431365
transform -1 0 25648 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1451_
timestamp 1698431365
transform -1 0 13888 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1452_
timestamp 1698431365
transform -1 0 14224 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1453_
timestamp 1698431365
transform 1 0 8400 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1454_
timestamp 1698431365
transform 1 0 8512 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1455_
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1456_
timestamp 1698431365
transform -1 0 16800 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1457_
timestamp 1698431365
transform -1 0 11312 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1458_
timestamp 1698431365
transform 1 0 9520 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1459_
timestamp 1698431365
transform 1 0 10416 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1460_
timestamp 1698431365
transform -1 0 16464 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1461_
timestamp 1698431365
transform 1 0 10976 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1462_
timestamp 1698431365
transform 1 0 11424 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1463_
timestamp 1698431365
transform 1 0 6832 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1464_
timestamp 1698431365
transform -1 0 16240 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1465_
timestamp 1698431365
transform 1 0 7952 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1466_
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1467_
timestamp 1698431365
transform -1 0 16128 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1468_
timestamp 1698431365
transform 1 0 11872 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1469_
timestamp 1698431365
transform 1 0 13664 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1470_
timestamp 1698431365
transform 1 0 11984 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1471_
timestamp 1698431365
transform 1 0 9408 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1472_
timestamp 1698431365
transform 1 0 8624 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1473_
timestamp 1698431365
transform 1 0 9520 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1474_
timestamp 1698431365
transform 1 0 11984 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1475_
timestamp 1698431365
transform -1 0 14560 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1476_
timestamp 1698431365
transform -1 0 12992 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1477_
timestamp 1698431365
transform -1 0 8960 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1478_
timestamp 1698431365
transform -1 0 8624 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1479_
timestamp 1698431365
transform 1 0 7840 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1480_
timestamp 1698431365
transform -1 0 9296 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1481_
timestamp 1698431365
transform 1 0 7952 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1482_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1483_
timestamp 1698431365
transform 1 0 13104 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1484_
timestamp 1698431365
transform -1 0 16464 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1485_
timestamp 1698431365
transform 1 0 22960 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1486_
timestamp 1698431365
transform 1 0 22736 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1487_
timestamp 1698431365
transform 1 0 22736 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1488_
timestamp 1698431365
transform 1 0 26096 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1489_
timestamp 1698431365
transform -1 0 22848 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1490_
timestamp 1698431365
transform -1 0 27440 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1491_
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1492_
timestamp 1698431365
transform -1 0 27216 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1493_
timestamp 1698431365
transform 1 0 23744 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1494_
timestamp 1698431365
transform -1 0 26992 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1495_
timestamp 1698431365
transform 1 0 28000 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1496_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1497_
timestamp 1698431365
transform -1 0 26656 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1498_
timestamp 1698431365
transform -1 0 27552 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1499_
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1500_
timestamp 1698431365
transform -1 0 27216 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1501_
timestamp 1698431365
transform -1 0 26096 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1502_
timestamp 1698431365
transform 1 0 31584 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1503_
timestamp 1698431365
transform 1 0 25536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1504_
timestamp 1698431365
transform 1 0 21280 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1505_
timestamp 1698431365
transform -1 0 26208 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1506_
timestamp 1698431365
transform -1 0 25088 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1507_
timestamp 1698431365
transform 1 0 22512 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1508_
timestamp 1698431365
transform 1 0 18816 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1509_
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1510_
timestamp 1698431365
transform 1 0 21728 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1511_
timestamp 1698431365
transform -1 0 23184 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1512_
timestamp 1698431365
transform 1 0 23408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1513_
timestamp 1698431365
transform 1 0 24304 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1514_
timestamp 1698431365
transform 1 0 11200 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1515_
timestamp 1698431365
transform -1 0 11312 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1516_
timestamp 1698431365
transform -1 0 11872 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1517_
timestamp 1698431365
transform 1 0 10864 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1518_
timestamp 1698431365
transform 1 0 10528 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1519_
timestamp 1698431365
transform 1 0 12096 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1520_
timestamp 1698431365
transform -1 0 15344 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1521_
timestamp 1698431365
transform 1 0 6048 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1522_
timestamp 1698431365
transform 1 0 6720 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1523_
timestamp 1698431365
transform 1 0 7392 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1524_
timestamp 1698431365
transform -1 0 14672 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1525_
timestamp 1698431365
transform 1 0 14672 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1526_
timestamp 1698431365
transform 1 0 14448 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1527_
timestamp 1698431365
transform 1 0 7168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1528_
timestamp 1698431365
transform 1 0 6944 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1529_
timestamp 1698431365
transform 1 0 7504 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1530_
timestamp 1698431365
transform -1 0 15120 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1531_
timestamp 1698431365
transform 1 0 13888 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1532_
timestamp 1698431365
transform -1 0 7280 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1533_
timestamp 1698431365
transform 1 0 7168 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1534_
timestamp 1698431365
transform 1 0 6832 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1535_
timestamp 1698431365
transform 1 0 13664 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1536_
timestamp 1698431365
transform 1 0 14560 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1537_
timestamp 1698431365
transform -1 0 16912 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1538_
timestamp 1698431365
transform 1 0 22848 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1539_
timestamp 1698431365
transform 1 0 22624 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1540_
timestamp 1698431365
transform 1 0 24080 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1541_
timestamp 1698431365
transform -1 0 22288 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1542_
timestamp 1698431365
transform 1 0 11984 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1543_
timestamp 1698431365
transform 1 0 11760 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1544_
timestamp 1698431365
transform -1 0 14224 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1545_
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1546_
timestamp 1698431365
transform 1 0 18032 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1547_
timestamp 1698431365
transform 1 0 18816 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1548_
timestamp 1698431365
transform -1 0 16688 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1549_
timestamp 1698431365
transform 1 0 14672 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1550_
timestamp 1698431365
transform 1 0 30240 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1551_
timestamp 1698431365
transform -1 0 30464 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1552_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1553_
timestamp 1698431365
transform 1 0 21392 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1554_
timestamp 1698431365
transform -1 0 22064 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1555_
timestamp 1698431365
transform 1 0 45136 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1556_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18144 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1557_
timestamp 1698431365
transform 1 0 25872 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1558_
timestamp 1698431365
transform 1 0 20384 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1559_
timestamp 1698431365
transform -1 0 22288 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1560_
timestamp 1698431365
transform -1 0 20048 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1561_
timestamp 1698431365
transform 1 0 19040 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1562_
timestamp 1698431365
transform 1 0 19488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1563_
timestamp 1698431365
transform -1 0 31136 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1564_
timestamp 1698431365
transform 1 0 22064 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1565_
timestamp 1698431365
transform -1 0 15680 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1566_
timestamp 1698431365
transform 1 0 11984 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1567_
timestamp 1698431365
transform 1 0 12880 0 -1 48608
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1568_
timestamp 1698431365
transform 1 0 14000 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1569_
timestamp 1698431365
transform 1 0 14784 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1570_
timestamp 1698431365
transform 1 0 16464 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1571_
timestamp 1698431365
transform -1 0 16128 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1572_
timestamp 1698431365
transform -1 0 32368 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1573_
timestamp 1698431365
transform -1 0 26656 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1574_
timestamp 1698431365
transform 1 0 23968 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1575_
timestamp 1698431365
transform 1 0 23072 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1576_
timestamp 1698431365
transform 1 0 18816 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1577_
timestamp 1698431365
transform 1 0 22736 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1578_
timestamp 1698431365
transform -1 0 18032 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1579_
timestamp 1698431365
transform 1 0 17136 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1580_
timestamp 1698431365
transform -1 0 17136 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1581_
timestamp 1698431365
transform 1 0 16240 0 -1 54880
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1582_
timestamp 1698431365
transform 1 0 17136 0 1 54880
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1583_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17024 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1584_
timestamp 1698431365
transform -1 0 19488 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1585_
timestamp 1698431365
transform 1 0 18816 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1586_
timestamp 1698431365
transform -1 0 25984 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1587_
timestamp 1698431365
transform 1 0 14336 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1588_
timestamp 1698431365
transform 1 0 20272 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1589_
timestamp 1698431365
transform -1 0 19936 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1590_
timestamp 1698431365
transform 1 0 25760 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1591_
timestamp 1698431365
transform -1 0 18928 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1592_
timestamp 1698431365
transform -1 0 15120 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1593_
timestamp 1698431365
transform 1 0 15680 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1594_
timestamp 1698431365
transform -1 0 15344 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1595_
timestamp 1698431365
transform 1 0 14896 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1596_
timestamp 1698431365
transform 1 0 13440 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1597_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14448 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1598_
timestamp 1698431365
transform 1 0 14560 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1599_
timestamp 1698431365
transform 1 0 28224 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1600_
timestamp 1698431365
transform -1 0 23744 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1601_
timestamp 1698431365
transform -1 0 17584 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1602_
timestamp 1698431365
transform -1 0 18144 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1603_
timestamp 1698431365
transform 1 0 15456 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1604_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16576 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1605_
timestamp 1698431365
transform -1 0 14000 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1606_
timestamp 1698431365
transform -1 0 44128 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1607_
timestamp 1698431365
transform 1 0 43120 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1608_
timestamp 1698431365
transform -1 0 42896 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1609_
timestamp 1698431365
transform -1 0 36176 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1610_
timestamp 1698431365
transform -1 0 36736 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1611_
timestamp 1698431365
transform -1 0 36624 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1612_
timestamp 1698431365
transform -1 0 35952 0 -1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1613_
timestamp 1698431365
transform -1 0 35056 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1614_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34720 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1615_
timestamp 1698431365
transform -1 0 41776 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1616_
timestamp 1698431365
transform -1 0 41216 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1617_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 -1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1618_
timestamp 1698431365
transform 1 0 38304 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1619_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39312 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1620_
timestamp 1698431365
transform -1 0 35728 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1621_
timestamp 1698431365
transform -1 0 30912 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1622_
timestamp 1698431365
transform -1 0 34384 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1623_
timestamp 1698431365
transform -1 0 28784 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1624_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18928 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1625_
timestamp 1698431365
transform 1 0 19824 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1626_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19488 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1627_
timestamp 1698431365
transform 1 0 21728 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1628_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17920 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1629_
timestamp 1698431365
transform -1 0 19824 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1630_
timestamp 1698431365
transform -1 0 13440 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1631_
timestamp 1698431365
transform 1 0 18144 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1632_
timestamp 1698431365
transform -1 0 21728 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1633_
timestamp 1698431365
transform -1 0 22064 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1634_
timestamp 1698431365
transform 1 0 27440 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1635_
timestamp 1698431365
transform 1 0 28112 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1636_
timestamp 1698431365
transform -1 0 15904 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1637_
timestamp 1698431365
transform -1 0 25760 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1638_
timestamp 1698431365
transform -1 0 25088 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1639_
timestamp 1698431365
transform -1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1640_
timestamp 1698431365
transform 1 0 18816 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1641_
timestamp 1698431365
transform 1 0 23184 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1642_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23744 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1643_
timestamp 1698431365
transform -1 0 18144 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1644_
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1645_
timestamp 1698431365
transform -1 0 19712 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1646_
timestamp 1698431365
transform 1 0 17360 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1647_
timestamp 1698431365
transform -1 0 19488 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1648_
timestamp 1698431365
transform 1 0 5824 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1649_
timestamp 1698431365
transform -1 0 6160 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1650_
timestamp 1698431365
transform -1 0 31024 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1651_
timestamp 1698431365
transform 1 0 28112 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1652_
timestamp 1698431365
transform -1 0 29792 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1653_
timestamp 1698431365
transform -1 0 12208 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1654_
timestamp 1698431365
transform 1 0 7504 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1655_
timestamp 1698431365
transform -1 0 8512 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1656_
timestamp 1698431365
transform -1 0 28112 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1657_
timestamp 1698431365
transform 1 0 16240 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1658_
timestamp 1698431365
transform 1 0 22736 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1659_
timestamp 1698431365
transform 1 0 22848 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1660_
timestamp 1698431365
transform -1 0 18928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1661_
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1662_
timestamp 1698431365
transform -1 0 3808 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1663_
timestamp 1698431365
transform 1 0 29680 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1664_
timestamp 1698431365
transform -1 0 16912 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1665_
timestamp 1698431365
transform 1 0 4816 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1666_
timestamp 1698431365
transform -1 0 3024 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1667_
timestamp 1698431365
transform -1 0 18480 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1668_
timestamp 1698431365
transform -1 0 21840 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1669_
timestamp 1698431365
transform -1 0 19376 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1670_
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1671_
timestamp 1698431365
transform 1 0 21840 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1672_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1673_
timestamp 1698431365
transform 1 0 22288 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1674_
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1675_
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1676_
timestamp 1698431365
transform -1 0 14000 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1677_
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1678_
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1679_
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1680_
timestamp 1698431365
transform 1 0 24304 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1681_
timestamp 1698431365
transform 1 0 24752 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1682_
timestamp 1698431365
transform -1 0 13888 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1683_
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1684_
timestamp 1698431365
transform 1 0 13552 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1685_
timestamp 1698431365
transform 1 0 11200 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1686_
timestamp 1698431365
transform -1 0 10864 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1687_
timestamp 1698431365
transform 1 0 21728 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1688_
timestamp 1698431365
transform -1 0 19040 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1689_
timestamp 1698431365
transform -1 0 18816 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1690_
timestamp 1698431365
transform 1 0 10080 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1691_
timestamp 1698431365
transform 1 0 9408 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1692_
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1693_
timestamp 1698431365
transform -1 0 10304 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1694_
timestamp 1698431365
transform -1 0 22848 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1695_
timestamp 1698431365
transform 1 0 18480 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1696_
timestamp 1698431365
transform 1 0 20048 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1697_
timestamp 1698431365
transform 1 0 20272 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1698_
timestamp 1698431365
transform -1 0 20832 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1699_
timestamp 1698431365
transform 1 0 17920 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1700_
timestamp 1698431365
transform -1 0 18032 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1701_
timestamp 1698431365
transform -1 0 20608 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1702_
timestamp 1698431365
transform 1 0 18928 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1703_
timestamp 1698431365
transform -1 0 16240 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1704_
timestamp 1698431365
transform -1 0 19040 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1705_
timestamp 1698431365
transform 1 0 12768 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1706_
timestamp 1698431365
transform -1 0 14000 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1707_
timestamp 1698431365
transform -1 0 12320 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1708_
timestamp 1698431365
transform 1 0 10864 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1709_
timestamp 1698431365
transform -1 0 10752 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1710_
timestamp 1698431365
transform -1 0 24752 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1711_
timestamp 1698431365
transform -1 0 19824 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1712_
timestamp 1698431365
transform 1 0 16576 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1713_
timestamp 1698431365
transform -1 0 16912 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1714_
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1715_
timestamp 1698431365
transform -1 0 16912 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1716_
timestamp 1698431365
transform -1 0 7840 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1717_
timestamp 1698431365
transform 1 0 5152 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1718_
timestamp 1698431365
transform -1 0 3920 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1719_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1720_
timestamp 1698431365
transform -1 0 3248 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1721_
timestamp 1698431365
transform 1 0 30912 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1722_
timestamp 1698431365
transform 1 0 49840 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1723_
timestamp 1698431365
transform -1 0 45920 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1724_
timestamp 1698431365
transform -1 0 24192 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1725_
timestamp 1698431365
transform 1 0 22624 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1726_
timestamp 1698431365
transform -1 0 18704 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1727_
timestamp 1698431365
transform -1 0 15344 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1728_
timestamp 1698431365
transform 1 0 13440 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1729_
timestamp 1698431365
transform -1 0 14000 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1730_
timestamp 1698431365
transform 1 0 10192 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1731_
timestamp 1698431365
transform -1 0 10080 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1732_
timestamp 1698431365
transform -1 0 9632 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1733_
timestamp 1698431365
transform 1 0 7728 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1734_
timestamp 1698431365
transform 1 0 7056 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1735_
timestamp 1698431365
transform -1 0 7840 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1736_
timestamp 1698431365
transform -1 0 8288 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1737_
timestamp 1698431365
transform 1 0 6832 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1738_
timestamp 1698431365
transform -1 0 7056 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1739_
timestamp 1698431365
transform 1 0 23632 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1740_
timestamp 1698431365
transform -1 0 7728 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1741_
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1742_
timestamp 1698431365
transform 1 0 1904 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1743_
timestamp 1698431365
transform 1 0 5824 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1744_
timestamp 1698431365
transform -1 0 4256 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1745_
timestamp 1698431365
transform -1 0 7952 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1746_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1747_
timestamp 1698431365
transform 1 0 1792 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1748_
timestamp 1698431365
transform 1 0 5712 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1749_
timestamp 1698431365
transform -1 0 4256 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1750_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18032 0 -1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1751_
timestamp 1698431365
transform -1 0 14336 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1752_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1753_
timestamp 1698431365
transform -1 0 3136 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1754_
timestamp 1698431365
transform 1 0 4816 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1755_
timestamp 1698431365
transform -1 0 3920 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1756_
timestamp 1698431365
transform -1 0 21056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1757_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1758_
timestamp 1698431365
transform -1 0 20496 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1759_
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1760_
timestamp 1698431365
transform -1 0 16912 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1761_
timestamp 1698431365
transform 1 0 18928 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1762_
timestamp 1698431365
transform -1 0 19376 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1763_
timestamp 1698431365
transform -1 0 22064 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1764_
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1765_
timestamp 1698431365
transform -1 0 21840 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1766_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20272 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1767_
timestamp 1698431365
transform 1 0 17472 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1768_
timestamp 1698431365
transform 1 0 25424 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1769_
timestamp 1698431365
transform -1 0 23072 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1770_
timestamp 1698431365
transform 1 0 23072 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1771_
timestamp 1698431365
transform 1 0 25872 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1772_
timestamp 1698431365
transform 1 0 30352 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1773_
timestamp 1698431365
transform 1 0 26880 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1774_
timestamp 1698431365
transform 1 0 19152 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1775_
timestamp 1698431365
transform -1 0 23632 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1776_
timestamp 1698431365
transform -1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1777_
timestamp 1698431365
transform -1 0 24192 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1778_
timestamp 1698431365
transform -1 0 20944 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1779_
timestamp 1698431365
transform -1 0 22624 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1780_
timestamp 1698431365
transform -1 0 14448 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1781_
timestamp 1698431365
transform -1 0 17024 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1782_
timestamp 1698431365
transform 1 0 13104 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1783_
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1784_
timestamp 1698431365
transform -1 0 18256 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1785_
timestamp 1698431365
transform -1 0 17472 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1786_
timestamp 1698431365
transform 1 0 26656 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1787_
timestamp 1698431365
transform 1 0 49504 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1788_
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1789_
timestamp 1698431365
transform 1 0 44240 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1790_
timestamp 1698431365
transform 1 0 45248 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1791_
timestamp 1698431365
transform -1 0 46032 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1792_
timestamp 1698431365
transform -1 0 48384 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1793_
timestamp 1698431365
transform -1 0 49280 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1794_
timestamp 1698431365
transform -1 0 47712 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1795_
timestamp 1698431365
transform -1 0 46816 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1796_
timestamp 1698431365
transform -1 0 46816 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1797_
timestamp 1698431365
transform 1 0 46368 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1798_
timestamp 1698431365
transform -1 0 48384 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1799_
timestamp 1698431365
transform 1 0 45360 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1800_
timestamp 1698431365
transform -1 0 48384 0 1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1801_
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1802_
timestamp 1698431365
transform 1 0 49952 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1803_
timestamp 1698431365
transform 1 0 50512 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1804_
timestamp 1698431365
transform -1 0 50288 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1805_
timestamp 1698431365
transform 1 0 49168 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1806_
timestamp 1698431365
transform 1 0 50176 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1807_
timestamp 1698431365
transform 1 0 49280 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1808_
timestamp 1698431365
transform 1 0 51744 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1809_
timestamp 1698431365
transform 1 0 49952 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1810_
timestamp 1698431365
transform -1 0 50960 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1811_
timestamp 1698431365
transform -1 0 51408 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1812_
timestamp 1698431365
transform -1 0 50624 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1813_
timestamp 1698431365
transform -1 0 49280 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1814_
timestamp 1698431365
transform -1 0 50064 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1815_
timestamp 1698431365
transform 1 0 49056 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1816_
timestamp 1698431365
transform 1 0 50064 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1817_
timestamp 1698431365
transform 1 0 50624 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1818_
timestamp 1698431365
transform -1 0 35616 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1819_
timestamp 1698431365
transform 1 0 27440 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1820_
timestamp 1698431365
transform 1 0 34608 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1821_
timestamp 1698431365
transform 1 0 33712 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1822_
timestamp 1698431365
transform 1 0 34832 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1823_
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1824_
timestamp 1698431365
transform 1 0 37968 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1825_
timestamp 1698431365
transform -1 0 37968 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1826_
timestamp 1698431365
transform -1 0 36960 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1827_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39984 0 -1 34496
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1828_
timestamp 1698431365
transform 1 0 36400 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1829_
timestamp 1698431365
transform 1 0 37744 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1830_
timestamp 1698431365
transform 1 0 39200 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1831_
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1832_
timestamp 1698431365
transform -1 0 36400 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1833_
timestamp 1698431365
transform -1 0 36736 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1834_
timestamp 1698431365
transform 1 0 38192 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1835_
timestamp 1698431365
transform -1 0 39200 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1836_
timestamp 1698431365
transform 1 0 37632 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1837_
timestamp 1698431365
transform -1 0 40544 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1838_
timestamp 1698431365
transform 1 0 37856 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1839_
timestamp 1698431365
transform 1 0 39312 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1840_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1841_
timestamp 1698431365
transform 1 0 36736 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1842_
timestamp 1698431365
transform -1 0 37520 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1843_
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1844_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37296 0 1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1845_
timestamp 1698431365
transform 1 0 38192 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1846_
timestamp 1698431365
transform 1 0 39200 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1847_
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1848_
timestamp 1698431365
transform 1 0 38976 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1849_
timestamp 1698431365
transform -1 0 38528 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1850_
timestamp 1698431365
transform -1 0 39984 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1851_
timestamp 1698431365
transform 1 0 38752 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1852_
timestamp 1698431365
transform -1 0 41216 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1853_
timestamp 1698431365
transform -1 0 42112 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1854_
timestamp 1698431365
transform 1 0 42112 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1855_
timestamp 1698431365
transform 1 0 43232 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1856_
timestamp 1698431365
transform 1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1857_
timestamp 1698431365
transform 1 0 34272 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1858_
timestamp 1698431365
transform 1 0 47264 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1859_
timestamp 1698431365
transform 1 0 39424 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1860_
timestamp 1698431365
transform -1 0 38976 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1861_
timestamp 1698431365
transform -1 0 40544 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1862_
timestamp 1698431365
transform -1 0 38864 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1863_
timestamp 1698431365
transform 1 0 38864 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1864_
timestamp 1698431365
transform 1 0 39984 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1865_
timestamp 1698431365
transform 1 0 40208 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1866_
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1867_
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1868_
timestamp 1698431365
transform -1 0 53536 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1869_
timestamp 1698431365
transform 1 0 48720 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1870_
timestamp 1698431365
transform 1 0 46928 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform -1 0 48720 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1872_
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1873_
timestamp 1698431365
transform -1 0 54208 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1874_
timestamp 1698431365
transform -1 0 46704 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1875_
timestamp 1698431365
transform 1 0 45360 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1876_
timestamp 1698431365
transform 1 0 49728 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1877_
timestamp 1698431365
transform 1 0 50736 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1878_
timestamp 1698431365
transform 1 0 51520 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1879_
timestamp 1698431365
transform -1 0 56112 0 -1 32928
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1880_
timestamp 1698431365
transform 1 0 51184 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1881_
timestamp 1698431365
transform -1 0 50512 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1882_
timestamp 1698431365
transform 1 0 46592 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1883_
timestamp 1698431365
transform -1 0 47824 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1884_
timestamp 1698431365
transform -1 0 56896 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1885_
timestamp 1698431365
transform -1 0 54768 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1886_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1887_
timestamp 1698431365
transform -1 0 47264 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1888_
timestamp 1698431365
transform -1 0 47152 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1889_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45696 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1890_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42784 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1891_
timestamp 1698431365
transform 1 0 46368 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1892_
timestamp 1698431365
transform 1 0 43008 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1893_
timestamp 1698431365
transform -1 0 54544 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1894_
timestamp 1698431365
transform 1 0 45472 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1895_
timestamp 1698431365
transform 1 0 44688 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1896_
timestamp 1698431365
transform 1 0 45696 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1897_
timestamp 1698431365
transform -1 0 39088 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1898_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1899_
timestamp 1698431365
transform -1 0 40544 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1900_
timestamp 1698431365
transform 1 0 38976 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1901_
timestamp 1698431365
transform -1 0 40544 0 -1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1902_
timestamp 1698431365
transform 1 0 37856 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1903_
timestamp 1698431365
transform 1 0 46032 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1904_
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1905_
timestamp 1698431365
transform 1 0 40880 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1906_
timestamp 1698431365
transform 1 0 40656 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1907_
timestamp 1698431365
transform -1 0 40544 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1908_
timestamp 1698431365
transform 1 0 40096 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1909_
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1910_
timestamp 1698431365
transform -1 0 42672 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1911_
timestamp 1698431365
transform 1 0 42224 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1912_
timestamp 1698431365
transform 1 0 43568 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1913_
timestamp 1698431365
transform 1 0 45136 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1914_
timestamp 1698431365
transform 1 0 47376 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1915_
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1916_
timestamp 1698431365
transform 1 0 44128 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1917_
timestamp 1698431365
transform 1 0 40992 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1918_
timestamp 1698431365
transform 1 0 41664 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1919_
timestamp 1698431365
transform -1 0 45920 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1920_
timestamp 1698431365
transform -1 0 45920 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1921_
timestamp 1698431365
transform 1 0 41776 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1922_
timestamp 1698431365
transform 1 0 42448 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1923_
timestamp 1698431365
transform 1 0 51408 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1924_
timestamp 1698431365
transform 1 0 40992 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1925_
timestamp 1698431365
transform 1 0 42336 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1926_
timestamp 1698431365
transform 1 0 44240 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1927_
timestamp 1698431365
transform 1 0 42336 0 -1 40768
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1928_
timestamp 1698431365
transform 1 0 44912 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1929_
timestamp 1698431365
transform 1 0 43008 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1930_
timestamp 1698431365
transform -1 0 43120 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1931_
timestamp 1698431365
transform -1 0 46032 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1932_
timestamp 1698431365
transform 1 0 46256 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1933_
timestamp 1698431365
transform 1 0 48160 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1934_
timestamp 1698431365
transform 1 0 41552 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1935_
timestamp 1698431365
transform 1 0 42672 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1936_
timestamp 1698431365
transform 1 0 41328 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1937_
timestamp 1698431365
transform -1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1938_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44016 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1939_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46928 0 -1 42336
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1940_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 50624 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1941_
timestamp 1698431365
transform 1 0 47824 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1942_
timestamp 1698431365
transform -1 0 47824 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1943_
timestamp 1698431365
transform 1 0 47824 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1944_
timestamp 1698431365
transform 1 0 47824 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1945_
timestamp 1698431365
transform 1 0 46704 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1946_
timestamp 1698431365
transform 1 0 49728 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1947_
timestamp 1698431365
transform 1 0 48832 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1948_
timestamp 1698431365
transform -1 0 46928 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1949_
timestamp 1698431365
transform 1 0 50400 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1950_
timestamp 1698431365
transform -1 0 52192 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1951_
timestamp 1698431365
transform 1 0 50176 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1952_
timestamp 1698431365
transform -1 0 53088 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1953_
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1954_
timestamp 1698431365
transform -1 0 52640 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1955_
timestamp 1698431365
transform 1 0 49392 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1956_
timestamp 1698431365
transform -1 0 51744 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1957_
timestamp 1698431365
transform -1 0 52640 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1958_
timestamp 1698431365
transform 1 0 45920 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1959_
timestamp 1698431365
transform -1 0 49728 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1960_
timestamp 1698431365
transform -1 0 50176 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1961_
timestamp 1698431365
transform 1 0 51856 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1962_
timestamp 1698431365
transform 1 0 51072 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1963_
timestamp 1698431365
transform 1 0 52640 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1964_
timestamp 1698431365
transform 1 0 53648 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1965_
timestamp 1698431365
transform -1 0 47376 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1966_
timestamp 1698431365
transform -1 0 45360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1967_
timestamp 1698431365
transform -1 0 40992 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1968_
timestamp 1698431365
transform -1 0 44464 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1969_
timestamp 1698431365
transform -1 0 44016 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1970_
timestamp 1698431365
transform 1 0 34048 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1971_
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1972_
timestamp 1698431365
transform -1 0 52080 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1973_
timestamp 1698431365
transform -1 0 50512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1974_
timestamp 1698431365
transform 1 0 46032 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1975_
timestamp 1698431365
transform -1 0 48944 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1976_
timestamp 1698431365
transform -1 0 53424 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1977_
timestamp 1698431365
transform -1 0 49504 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1978_
timestamp 1698431365
transform 1 0 46928 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1979_
timestamp 1698431365
transform 1 0 47712 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1980_
timestamp 1698431365
transform 1 0 47712 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1981_
timestamp 1698431365
transform 1 0 48944 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1982_
timestamp 1698431365
transform -1 0 48384 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1983_
timestamp 1698431365
transform -1 0 51184 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1984_
timestamp 1698431365
transform 1 0 54544 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1985_
timestamp 1698431365
transform -1 0 57120 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1986_
timestamp 1698431365
transform -1 0 41664 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1987_
timestamp 1698431365
transform -1 0 53648 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1988_
timestamp 1698431365
transform -1 0 54208 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1989_
timestamp 1698431365
transform -1 0 56000 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1990_
timestamp 1698431365
transform 1 0 47600 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1991_
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1992_
timestamp 1698431365
transform 1 0 47488 0 1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1993_
timestamp 1698431365
transform -1 0 53648 0 -1 37632
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1994_
timestamp 1698431365
transform 1 0 54320 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1995_
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1996_
timestamp 1698431365
transform 1 0 54656 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1997_
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1998_
timestamp 1698431365
transform 1 0 54208 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1999_
timestamp 1698431365
transform -1 0 55440 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2000_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 53424 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2001_
timestamp 1698431365
transform 1 0 57120 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2002_
timestamp 1698431365
transform 1 0 55664 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2003_
timestamp 1698431365
transform -1 0 40320 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2004_
timestamp 1698431365
transform 1 0 39872 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2005_
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2006_
timestamp 1698431365
transform -1 0 53424 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2007_
timestamp 1698431365
transform -1 0 51744 0 -1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2008_
timestamp 1698431365
transform -1 0 52640 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2009_
timestamp 1698431365
transform -1 0 54432 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2010_
timestamp 1698431365
transform -1 0 52304 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2011_
timestamp 1698431365
transform -1 0 53760 0 -1 34496
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2012_
timestamp 1698431365
transform 1 0 48720 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2013_
timestamp 1698431365
transform -1 0 50176 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2014_
timestamp 1698431365
transform -1 0 51072 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2015_
timestamp 1698431365
transform 1 0 31360 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2016_
timestamp 1698431365
transform -1 0 52304 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2017_
timestamp 1698431365
transform 1 0 42336 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2018_
timestamp 1698431365
transform -1 0 46592 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2019_
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2020_
timestamp 1698431365
transform -1 0 50176 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2021_
timestamp 1698431365
transform 1 0 52640 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2022_
timestamp 1698431365
transform -1 0 54096 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2023_
timestamp 1698431365
transform -1 0 51072 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2024_
timestamp 1698431365
transform -1 0 48272 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2025_
timestamp 1698431365
transform -1 0 45024 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2026_
timestamp 1698431365
transform -1 0 44464 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2027_
timestamp 1698431365
transform 1 0 42896 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2028_
timestamp 1698431365
transform -1 0 42112 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2029_
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2030_
timestamp 1698431365
transform -1 0 52640 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2031_
timestamp 1698431365
transform 1 0 50848 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2032_
timestamp 1698431365
transform -1 0 47376 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2033_
timestamp 1698431365
transform 1 0 45808 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2034_
timestamp 1698431365
transform -1 0 45696 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2035_
timestamp 1698431365
transform 1 0 44576 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2036_
timestamp 1698431365
transform -1 0 51408 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2037_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 51184 0 -1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2038_
timestamp 1698431365
transform -1 0 52304 0 1 29792
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2039_
timestamp 1698431365
transform -1 0 49280 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2040_
timestamp 1698431365
transform 1 0 48832 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2041_
timestamp 1698431365
transform -1 0 53648 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2042_
timestamp 1698431365
transform -1 0 54320 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2043_
timestamp 1698431365
transform -1 0 53984 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2044_
timestamp 1698431365
transform -1 0 51744 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2045_
timestamp 1698431365
transform -1 0 49952 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2046_
timestamp 1698431365
transform -1 0 51296 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2047_
timestamp 1698431365
transform 1 0 51520 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2048_
timestamp 1698431365
transform 1 0 50400 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2049_
timestamp 1698431365
transform -1 0 52976 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2050_
timestamp 1698431365
transform -1 0 50400 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2051_
timestamp 1698431365
transform 1 0 54544 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2052_
timestamp 1698431365
transform 1 0 55328 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2053_
timestamp 1698431365
transform -1 0 53872 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2054_
timestamp 1698431365
transform 1 0 49952 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2055_
timestamp 1698431365
transform -1 0 53424 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2056_
timestamp 1698431365
transform 1 0 50624 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2057_
timestamp 1698431365
transform 1 0 53424 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2058_
timestamp 1698431365
transform -1 0 52192 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2059_
timestamp 1698431365
transform -1 0 47824 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2060_
timestamp 1698431365
transform -1 0 36400 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2061_
timestamp 1698431365
transform -1 0 49952 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2062_
timestamp 1698431365
transform -1 0 52304 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2063_
timestamp 1698431365
transform -1 0 49280 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2064_
timestamp 1698431365
transform -1 0 47376 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2065_
timestamp 1698431365
transform -1 0 47376 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2066_
timestamp 1698431365
transform -1 0 46032 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2067_
timestamp 1698431365
transform 1 0 47936 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2068_
timestamp 1698431365
transform 1 0 49392 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2069_
timestamp 1698431365
transform -1 0 48048 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2070_
timestamp 1698431365
transform -1 0 45584 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2071_
timestamp 1698431365
transform 1 0 46032 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2072_
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2073_
timestamp 1698431365
transform -1 0 47488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2074_
timestamp 1698431365
transform -1 0 45696 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2075_
timestamp 1698431365
transform -1 0 46480 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2076_
timestamp 1698431365
transform 1 0 47040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2077_
timestamp 1698431365
transform -1 0 46256 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2078_
timestamp 1698431365
transform 1 0 47488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2079_
timestamp 1698431365
transform -1 0 47936 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2080_
timestamp 1698431365
transform 1 0 47264 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2081_
timestamp 1698431365
transform 1 0 46144 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2082_
timestamp 1698431365
transform -1 0 46592 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2083_
timestamp 1698431365
transform -1 0 48160 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2084_
timestamp 1698431365
transform -1 0 45472 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2085_
timestamp 1698431365
transform -1 0 44240 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2086_
timestamp 1698431365
transform 1 0 47376 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2087_
timestamp 1698431365
transform -1 0 45584 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2088_
timestamp 1698431365
transform 1 0 42224 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2089_
timestamp 1698431365
transform -1 0 44352 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2090_
timestamp 1698431365
transform -1 0 46144 0 -1 26656
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2091_
timestamp 1698431365
transform 1 0 43008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2092_
timestamp 1698431365
transform 1 0 42112 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2093_
timestamp 1698431365
transform -1 0 42560 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2094_
timestamp 1698431365
transform -1 0 41216 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2095_
timestamp 1698431365
transform 1 0 40992 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2096_
timestamp 1698431365
transform -1 0 43904 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2097_
timestamp 1698431365
transform -1 0 42784 0 -1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2098_
timestamp 1698431365
transform 1 0 42000 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2099_
timestamp 1698431365
transform 1 0 43904 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2100_
timestamp 1698431365
transform 1 0 42784 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2101_
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2102_
timestamp 1698431365
transform 1 0 41440 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2103_
timestamp 1698431365
transform -1 0 40544 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2104_
timestamp 1698431365
transform 1 0 40992 0 1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2105_
timestamp 1698431365
transform 1 0 39648 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2106_
timestamp 1698431365
transform -1 0 42224 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2107_
timestamp 1698431365
transform -1 0 46144 0 -1 25088
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2108_
timestamp 1698431365
transform -1 0 34944 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2109_
timestamp 1698431365
transform 1 0 37856 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2110_
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2111_
timestamp 1698431365
transform -1 0 39424 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2112_
timestamp 1698431365
transform -1 0 37856 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2113_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2114_
timestamp 1698431365
transform -1 0 42336 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2115_
timestamp 1698431365
transform -1 0 36064 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2116_
timestamp 1698431365
transform -1 0 35504 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2117_
timestamp 1698431365
transform 1 0 38192 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2118_
timestamp 1698431365
transform -1 0 37520 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2119_
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2120_
timestamp 1698431365
transform -1 0 38864 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2121_
timestamp 1698431365
transform -1 0 40992 0 1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2122_
timestamp 1698431365
transform 1 0 34944 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2123_
timestamp 1698431365
transform -1 0 39760 0 -1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2124_
timestamp 1698431365
transform -1 0 38080 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2125_
timestamp 1698431365
transform 1 0 32032 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2126_
timestamp 1698431365
transform -1 0 36400 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2127_
timestamp 1698431365
transform -1 0 35392 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2128_
timestamp 1698431365
transform -1 0 34944 0 1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2129_
timestamp 1698431365
transform 1 0 34160 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2130_
timestamp 1698431365
transform -1 0 34608 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2131_
timestamp 1698431365
transform 1 0 34608 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2132_
timestamp 1698431365
transform -1 0 33824 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2133_
timestamp 1698431365
transform -1 0 34160 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2134_
timestamp 1698431365
transform 1 0 32368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2135_
timestamp 1698431365
transform -1 0 35504 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2136_
timestamp 1698431365
transform 1 0 32704 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2137_
timestamp 1698431365
transform 1 0 33040 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2138_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2139_
timestamp 1698431365
transform 1 0 34272 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2140_
timestamp 1698431365
transform -1 0 34048 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2141_
timestamp 1698431365
transform -1 0 34832 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2142_
timestamp 1698431365
transform -1 0 34720 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2143_
timestamp 1698431365
transform -1 0 35616 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2144_
timestamp 1698431365
transform -1 0 32704 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2145_
timestamp 1698431365
transform 1 0 33712 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2146_
timestamp 1698431365
transform 1 0 34384 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2147_
timestamp 1698431365
transform 1 0 35616 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2148_
timestamp 1698431365
transform 1 0 36960 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2149_
timestamp 1698431365
transform 1 0 44464 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2150_
timestamp 1698431365
transform 1 0 45808 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2151_
timestamp 1698431365
transform 1 0 19040 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2152_
timestamp 1698431365
transform 1 0 20272 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2153_
timestamp 1698431365
transform 1 0 33712 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2154_
timestamp 1698431365
transform 1 0 34608 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2155_
timestamp 1698431365
transform -1 0 31024 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2156_
timestamp 1698431365
transform 1 0 31024 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2157_
timestamp 1698431365
transform -1 0 23520 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2158_
timestamp 1698431365
transform -1 0 20608 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2159_
timestamp 1698431365
transform 1 0 19488 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2160_
timestamp 1698431365
transform 1 0 22288 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2161_
timestamp 1698431365
transform -1 0 25760 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2162_
timestamp 1698431365
transform -1 0 19264 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2163_
timestamp 1698431365
transform 1 0 18256 0 1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2164_
timestamp 1698431365
transform 1 0 29344 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2165_
timestamp 1698431365
transform 1 0 28560 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2166_
timestamp 1698431365
transform 1 0 30016 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2167_
timestamp 1698431365
transform -1 0 30016 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2168_
timestamp 1698431365
transform -1 0 30576 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2169_
timestamp 1698431365
transform -1 0 31696 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2170_
timestamp 1698431365
transform -1 0 31024 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2171_
timestamp 1698431365
transform -1 0 31360 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2172_
timestamp 1698431365
transform -1 0 26208 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2173_
timestamp 1698431365
transform -1 0 16576 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2174_
timestamp 1698431365
transform -1 0 19600 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2175_
timestamp 1698431365
transform 1 0 17472 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _2176_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14224 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2177_
timestamp 1698431365
transform -1 0 25984 0 1 45472
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2178_
timestamp 1698431365
transform 1 0 19936 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2179_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2180_
timestamp 1698431365
transform 1 0 21056 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2181_
timestamp 1698431365
transform 1 0 28000 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2182_
timestamp 1698431365
transform -1 0 28784 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2183_
timestamp 1698431365
transform 1 0 27664 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2184_
timestamp 1698431365
transform -1 0 29904 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2185_
timestamp 1698431365
transform -1 0 32368 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2186_
timestamp 1698431365
transform 1 0 31248 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2187_
timestamp 1698431365
transform -1 0 28784 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2188_
timestamp 1698431365
transform 1 0 26208 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2189_
timestamp 1698431365
transform -1 0 24864 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2190_
timestamp 1698431365
transform 1 0 24864 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2191_
timestamp 1698431365
transform 1 0 26992 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2192_
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2193_
timestamp 1698431365
transform -1 0 27104 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2194_
timestamp 1698431365
transform 1 0 28000 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2195_
timestamp 1698431365
transform 1 0 29008 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2196_
timestamp 1698431365
transform -1 0 31248 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2197_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29792 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2198_
timestamp 1698431365
transform -1 0 20384 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2199_
timestamp 1698431365
transform -1 0 23744 0 -1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2200_
timestamp 1698431365
transform -1 0 21840 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2201_
timestamp 1698431365
transform 1 0 22400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2202_
timestamp 1698431365
transform 1 0 21840 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2203_
timestamp 1698431365
transform 1 0 22400 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2204_
timestamp 1698431365
transform 1 0 29680 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2205_
timestamp 1698431365
transform -1 0 29008 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2206_
timestamp 1698431365
transform 1 0 29120 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2207_
timestamp 1698431365
transform 1 0 31920 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2208_
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2209_
timestamp 1698431365
transform -1 0 31808 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2210_
timestamp 1698431365
transform 1 0 25648 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2211_
timestamp 1698431365
transform -1 0 27888 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2212_
timestamp 1698431365
transform 1 0 27552 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2213_
timestamp 1698431365
transform 1 0 30128 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2214_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29456 0 -1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2215_
timestamp 1698431365
transform -1 0 31808 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2216_
timestamp 1698431365
transform -1 0 31584 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2217_
timestamp 1698431365
transform 1 0 24976 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2218_
timestamp 1698431365
transform 1 0 28000 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2219_
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2220_
timestamp 1698431365
transform 1 0 23520 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2221_
timestamp 1698431365
transform -1 0 26992 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2222_
timestamp 1698431365
transform 1 0 25648 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2223_
timestamp 1698431365
transform 1 0 25312 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2224_
timestamp 1698431365
transform -1 0 26656 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2225_
timestamp 1698431365
transform 1 0 23744 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2226_
timestamp 1698431365
transform -1 0 11648 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2227_
timestamp 1698431365
transform 1 0 14000 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2228_
timestamp 1698431365
transform 1 0 15568 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2229_
timestamp 1698431365
transform 1 0 25088 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2230_
timestamp 1698431365
transform 1 0 23296 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2231_
timestamp 1698431365
transform -1 0 20272 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2232_
timestamp 1698431365
transform 1 0 31136 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2233_
timestamp 1698431365
transform 1 0 31808 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2234_
timestamp 1698431365
transform -1 0 27664 0 -1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2235_
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2236_
timestamp 1698431365
transform -1 0 30688 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2237_
timestamp 1698431365
transform -1 0 30576 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2238_
timestamp 1698431365
transform 1 0 12544 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2239_
timestamp 1698431365
transform 1 0 21952 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2240_
timestamp 1698431365
transform 1 0 22960 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2241_
timestamp 1698431365
transform -1 0 27776 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2242_
timestamp 1698431365
transform -1 0 29456 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2243_
timestamp 1698431365
transform 1 0 28560 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2244_
timestamp 1698431365
transform 1 0 22400 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2245_
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2246_
timestamp 1698431365
transform -1 0 33488 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2247_
timestamp 1698431365
transform -1 0 32704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2248_
timestamp 1698431365
transform 1 0 31024 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2249_
timestamp 1698431365
transform -1 0 27216 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2250_
timestamp 1698431365
transform 1 0 27440 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2251_
timestamp 1698431365
transform 1 0 16128 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2252_
timestamp 1698431365
transform 1 0 14448 0 1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2253_
timestamp 1698431365
transform 1 0 24080 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2254_
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2255_
timestamp 1698431365
transform -1 0 17024 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2256_
timestamp 1698431365
transform 1 0 19712 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2257_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25312 0 1 43904
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2258_
timestamp 1698431365
transform 1 0 27776 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2259_
timestamp 1698431365
transform -1 0 34384 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2260_
timestamp 1698431365
transform 1 0 34384 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2261_
timestamp 1698431365
transform 1 0 24416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2262_
timestamp 1698431365
transform 1 0 25648 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2263_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2264_
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2265_
timestamp 1698431365
transform 1 0 27552 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2266_
timestamp 1698431365
transform -1 0 29904 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2267_
timestamp 1698431365
transform 1 0 33712 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2268_
timestamp 1698431365
transform -1 0 34272 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2269_
timestamp 1698431365
transform 1 0 25984 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2270_
timestamp 1698431365
transform -1 0 27552 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2271_
timestamp 1698431365
transform 1 0 32144 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2272_
timestamp 1698431365
transform 1 0 33040 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2273_
timestamp 1698431365
transform 1 0 34272 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2274_
timestamp 1698431365
transform 1 0 30240 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2275_
timestamp 1698431365
transform 1 0 31136 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2276_
timestamp 1698431365
transform 1 0 30688 0 -1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2277_
timestamp 1698431365
transform 1 0 30688 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2278_
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2279_
timestamp 1698431365
transform -1 0 36624 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2280_
timestamp 1698431365
transform 1 0 26656 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2281_
timestamp 1698431365
transform 1 0 26432 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2282_
timestamp 1698431365
transform -1 0 29792 0 1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2283_
timestamp 1698431365
transform -1 0 28560 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2284_
timestamp 1698431365
transform -1 0 28784 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2285_
timestamp 1698431365
transform -1 0 36176 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2286_
timestamp 1698431365
transform -1 0 35616 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2287_
timestamp 1698431365
transform -1 0 35952 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2288_
timestamp 1698431365
transform 1 0 29456 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2289_
timestamp 1698431365
transform -1 0 25200 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2290_
timestamp 1698431365
transform -1 0 28112 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2291_
timestamp 1698431365
transform 1 0 27664 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2292_
timestamp 1698431365
transform 1 0 34160 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2293_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2294_
timestamp 1698431365
transform 1 0 29680 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2295_
timestamp 1698431365
transform -1 0 28000 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2296_
timestamp 1698431365
transform -1 0 27552 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2297_
timestamp 1698431365
transform 1 0 29792 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2298_
timestamp 1698431365
transform 1 0 31360 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2299_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2300_
timestamp 1698431365
transform 1 0 14112 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2301_
timestamp 1698431365
transform 1 0 17696 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2302_
timestamp 1698431365
transform 1 0 18368 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2303_
timestamp 1698431365
transform -1 0 20272 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2304_
timestamp 1698431365
transform -1 0 19152 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2305_
timestamp 1698431365
transform -1 0 12544 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2306_
timestamp 1698431365
transform -1 0 7728 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2307_
timestamp 1698431365
transform -1 0 7952 0 1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2308_
timestamp 1698431365
transform 1 0 4256 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2309_
timestamp 1698431365
transform -1 0 9632 0 1 51744
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2310_
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2311_
timestamp 1698431365
transform -1 0 5264 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2312_
timestamp 1698431365
transform 1 0 1792 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2313_
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2314_
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2315_
timestamp 1698431365
transform 1 0 9632 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2316_
timestamp 1698431365
transform 1 0 12320 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2317_
timestamp 1698431365
transform 1 0 11424 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2318_
timestamp 1698431365
transform 1 0 12432 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2319_
timestamp 1698431365
transform -1 0 15232 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2320_
timestamp 1698431365
transform 1 0 12208 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2321_
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2322_
timestamp 1698431365
transform 1 0 20160 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2323_
timestamp 1698431365
transform -1 0 21056 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2324_
timestamp 1698431365
transform -1 0 17136 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2325_
timestamp 1698431365
transform -1 0 13664 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2326_
timestamp 1698431365
transform 1 0 13664 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2327_
timestamp 1698431365
transform 1 0 9968 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2328_
timestamp 1698431365
transform -1 0 14672 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2329_
timestamp 1698431365
transform -1 0 10864 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2330_
timestamp 1698431365
transform -1 0 18368 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2331_
timestamp 1698431365
transform -1 0 17024 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2332_
timestamp 1698431365
transform -1 0 15792 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2333_
timestamp 1698431365
transform 1 0 10416 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2334_
timestamp 1698431365
transform -1 0 10640 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2335_
timestamp 1698431365
transform -1 0 10416 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2336_
timestamp 1698431365
transform -1 0 14896 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2337_
timestamp 1698431365
transform 1 0 13440 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2338_
timestamp 1698431365
transform 1 0 10864 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2339_
timestamp 1698431365
transform -1 0 10864 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2340_
timestamp 1698431365
transform 1 0 11200 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2341_
timestamp 1698431365
transform 1 0 11088 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2342_
timestamp 1698431365
transform 1 0 10192 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2343_
timestamp 1698431365
transform -1 0 10752 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2344_
timestamp 1698431365
transform -1 0 17024 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2345_
timestamp 1698431365
transform 1 0 15232 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2346_
timestamp 1698431365
transform 1 0 11872 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2347_
timestamp 1698431365
transform 1 0 14112 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2348_
timestamp 1698431365
transform 1 0 13216 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2349_
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2350_
timestamp 1698431365
transform -1 0 14000 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2351_
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2352_
timestamp 1698431365
transform 1 0 16016 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2353_
timestamp 1698431365
transform 1 0 15120 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2354_
timestamp 1698431365
transform -1 0 18928 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2355_
timestamp 1698431365
transform 1 0 13888 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2356_
timestamp 1698431365
transform 1 0 14896 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2357_
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2358_
timestamp 1698431365
transform -1 0 16800 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2359_
timestamp 1698431365
transform -1 0 16912 0 -1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2360_
timestamp 1698431365
transform -1 0 11424 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2361_
timestamp 1698431365
transform -1 0 7504 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2362_
timestamp 1698431365
transform 1 0 2576 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2363_
timestamp 1698431365
transform -1 0 4256 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2364_
timestamp 1698431365
transform -1 0 2800 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2365_
timestamp 1698431365
transform -1 0 6832 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2366_
timestamp 1698431365
transform 1 0 4144 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2367_
timestamp 1698431365
transform 1 0 3248 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2368_
timestamp 1698431365
transform 1 0 4256 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2369_
timestamp 1698431365
transform 1 0 5824 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2370_
timestamp 1698431365
transform 1 0 7280 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2371_
timestamp 1698431365
transform -1 0 6944 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2372_
timestamp 1698431365
transform 1 0 6944 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2373_
timestamp 1698431365
transform -1 0 7280 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2374_
timestamp 1698431365
transform 1 0 5376 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2375_
timestamp 1698431365
transform 1 0 6944 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2376_
timestamp 1698431365
transform -1 0 6384 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2377_
timestamp 1698431365
transform 1 0 6272 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2378_
timestamp 1698431365
transform 1 0 5936 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2379_
timestamp 1698431365
transform -1 0 8736 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2380_
timestamp 1698431365
transform -1 0 6160 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2381_
timestamp 1698431365
transform -1 0 7952 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2382_
timestamp 1698431365
transform -1 0 7840 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2383_
timestamp 1698431365
transform -1 0 6944 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2384_
timestamp 1698431365
transform -1 0 7056 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2385_
timestamp 1698431365
transform -1 0 7728 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2386_
timestamp 1698431365
transform -1 0 6048 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2387_
timestamp 1698431365
transform -1 0 7952 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2388_
timestamp 1698431365
transform -1 0 7056 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2389_
timestamp 1698431365
transform 1 0 2576 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2390_
timestamp 1698431365
transform 1 0 4144 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2391_
timestamp 1698431365
transform 1 0 3248 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2392_
timestamp 1698431365
transform 1 0 5040 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2393_
timestamp 1698431365
transform 1 0 4144 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2394_
timestamp 1698431365
transform 1 0 4256 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2395_
timestamp 1698431365
transform 1 0 6720 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2396_
timestamp 1698431365
transform -1 0 5712 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2397_
timestamp 1698431365
transform 1 0 5824 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2398_
timestamp 1698431365
transform -1 0 4368 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2399_
timestamp 1698431365
transform 1 0 3472 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2400_
timestamp 1698431365
transform -1 0 3472 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2401_
timestamp 1698431365
transform 1 0 4816 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2402_
timestamp 1698431365
transform -1 0 4032 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2403_
timestamp 1698431365
transform 1 0 4032 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2404_
timestamp 1698431365
transform 1 0 2240 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2405_
timestamp 1698431365
transform -1 0 4704 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2406_
timestamp 1698431365
transform -1 0 2464 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2407_
timestamp 1698431365
transform -1 0 3808 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2408_
timestamp 1698431365
transform -1 0 3248 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2409_
timestamp 1698431365
transform 1 0 26096 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2410_
timestamp 1698431365
transform -1 0 22848 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2411_
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2412_
timestamp 1698431365
transform 1 0 25200 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2413_
timestamp 1698431365
transform 1 0 26208 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2414_
timestamp 1698431365
transform 1 0 23968 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2415_
timestamp 1698431365
transform -1 0 24416 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2416_
timestamp 1698431365
transform -1 0 24640 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2417_
timestamp 1698431365
transform -1 0 23184 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2418_
timestamp 1698431365
transform -1 0 23296 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2419_
timestamp 1698431365
transform 1 0 21168 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2420_
timestamp 1698431365
transform -1 0 22512 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2421_
timestamp 1698431365
transform -1 0 21168 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2422_
timestamp 1698431365
transform -1 0 20608 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2423_
timestamp 1698431365
transform -1 0 20160 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2424_
timestamp 1698431365
transform -1 0 22960 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2425_
timestamp 1698431365
transform -1 0 20720 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2426_
timestamp 1698431365
transform -1 0 19264 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2427_
timestamp 1698431365
transform 1 0 26880 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2428_
timestamp 1698431365
transform -1 0 25984 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2429_
timestamp 1698431365
transform 1 0 23968 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2430_
timestamp 1698431365
transform -1 0 21840 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2431_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2432_
timestamp 1698431365
transform -1 0 14448 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2433_
timestamp 1698431365
transform -1 0 24752 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2434_
timestamp 1698431365
transform -1 0 22400 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2435_
timestamp 1698431365
transform 1 0 22960 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2436_
timestamp 1698431365
transform -1 0 24304 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2437_
timestamp 1698431365
transform 1 0 18816 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2438_
timestamp 1698431365
transform 1 0 19488 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2439_
timestamp 1698431365
transform -1 0 20384 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2440_
timestamp 1698431365
transform -1 0 20832 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2441_
timestamp 1698431365
transform 1 0 19712 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2442_
timestamp 1698431365
transform -1 0 21280 0 -1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2443_
timestamp 1698431365
transform 1 0 22064 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2444_
timestamp 1698431365
transform -1 0 23296 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2445_
timestamp 1698431365
transform -1 0 24640 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2446_
timestamp 1698431365
transform 1 0 22288 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2447_
timestamp 1698431365
transform 1 0 22736 0 1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2448_
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2449_
timestamp 1698431365
transform 1 0 21504 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2450_
timestamp 1698431365
transform -1 0 25648 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2451_
timestamp 1698431365
transform 1 0 23744 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2452_
timestamp 1698431365
transform 1 0 23856 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2453_
timestamp 1698431365
transform 1 0 23520 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2454_
timestamp 1698431365
transform -1 0 23184 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2455_
timestamp 1698431365
transform 1 0 19152 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2456_
timestamp 1698431365
transform 1 0 22736 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2457_
timestamp 1698431365
transform -1 0 24192 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2458_
timestamp 1698431365
transform -1 0 23296 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2459_
timestamp 1698431365
transform -1 0 23744 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2460_
timestamp 1698431365
transform -1 0 24080 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2461_
timestamp 1698431365
transform 1 0 18032 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2462_
timestamp 1698431365
transform 1 0 19824 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2463_
timestamp 1698431365
transform 1 0 21616 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2464_
timestamp 1698431365
transform 1 0 23408 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2465_
timestamp 1698431365
transform 1 0 24192 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2466_
timestamp 1698431365
transform 1 0 23856 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2467_
timestamp 1698431365
transform 1 0 19712 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2468_
timestamp 1698431365
transform 1 0 22288 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2469_
timestamp 1698431365
transform 1 0 23856 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2470_
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2471_
timestamp 1698431365
transform 1 0 29008 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2472_
timestamp 1698431365
transform 1 0 23184 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2473_
timestamp 1698431365
transform 1 0 33376 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2474_
timestamp 1698431365
transform 1 0 33600 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2475_
timestamp 1698431365
transform 1 0 29344 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2476_
timestamp 1698431365
transform 1 0 34944 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2477_
timestamp 1698431365
transform 1 0 34944 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2478_
timestamp 1698431365
transform -1 0 15568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2479_
timestamp 1698431365
transform -1 0 22064 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2480_
timestamp 1698431365
transform 1 0 18368 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2481_
timestamp 1698431365
transform -1 0 18480 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2482_
timestamp 1698431365
transform -1 0 16016 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2483_
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2484_
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2485_
timestamp 1698431365
transform -1 0 13888 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2486_
timestamp 1698431365
transform -1 0 15008 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2487_
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2488_
timestamp 1698431365
transform 1 0 10976 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2489_
timestamp 1698431365
transform -1 0 10640 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2490_
timestamp 1698431365
transform -1 0 24752 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2491_
timestamp 1698431365
transform 1 0 24864 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2492_
timestamp 1698431365
transform 1 0 29344 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2493_
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2494_
timestamp 1698431365
transform 1 0 30688 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2495_
timestamp 1698431365
transform 1 0 30016 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2496_
timestamp 1698431365
transform -1 0 22624 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2497_
timestamp 1698431365
transform -1 0 21840 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2498_
timestamp 1698431365
transform -1 0 21728 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2499_
timestamp 1698431365
transform 1 0 18928 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2500_
timestamp 1698431365
transform -1 0 18816 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2501_
timestamp 1698431365
transform -1 0 21728 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2502_
timestamp 1698431365
transform 1 0 20160 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2503_
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2504_
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2505_
timestamp 1698431365
transform 1 0 30128 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2506_
timestamp 1698431365
transform 1 0 30240 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2507_
timestamp 1698431365
transform 1 0 30576 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2508_
timestamp 1698431365
transform 1 0 30352 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2509_
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2510_
timestamp 1698431365
transform 1 0 32928 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2511_
timestamp 1698431365
transform 1 0 32032 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2512_
timestamp 1698431365
transform 1 0 34944 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2513_
timestamp 1698431365
transform 1 0 35392 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2514_
timestamp 1698431365
transform -1 0 12992 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2515_
timestamp 1698431365
transform 1 0 10864 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2516_
timestamp 1698431365
transform 1 0 8512 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2517_
timestamp 1698431365
transform 1 0 9520 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2518_
timestamp 1698431365
transform -1 0 8512 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2519_
timestamp 1698431365
transform 1 0 27552 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2520_
timestamp 1698431365
transform 1 0 21952 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2521_
timestamp 1698431365
transform 1 0 26544 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2522_
timestamp 1698431365
transform -1 0 26768 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2523_
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2524_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2525_
timestamp 1698431365
transform -1 0 29680 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2526_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2527_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2528_
timestamp 1698431365
transform -1 0 32592 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2529_
timestamp 1698431365
transform 1 0 34944 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2530_
timestamp 1698431365
transform 1 0 34272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2531_
timestamp 1698431365
transform -1 0 25872 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2532_
timestamp 1698431365
transform 1 0 21392 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2533_
timestamp 1698431365
transform 1 0 20832 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2534_
timestamp 1698431365
transform 1 0 20272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2535_
timestamp 1698431365
transform -1 0 29680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2536_
timestamp 1698431365
transform 1 0 22512 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2537_
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2538_
timestamp 1698431365
transform 1 0 25872 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2539_
timestamp 1698431365
transform 1 0 25424 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2540_
timestamp 1698431365
transform -1 0 25872 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2541_
timestamp 1698431365
transform 1 0 27328 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2542_
timestamp 1698431365
transform 1 0 27664 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2543_
timestamp 1698431365
transform -1 0 24752 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2544_
timestamp 1698431365
transform 1 0 20272 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2545_
timestamp 1698431365
transform -1 0 20944 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2546_
timestamp 1698431365
transform 1 0 21952 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2547_
timestamp 1698431365
transform -1 0 23296 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2548_
timestamp 1698431365
transform 1 0 25872 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2549_
timestamp 1698431365
transform 1 0 25536 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2550_
timestamp 1698431365
transform -1 0 25984 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2551_
timestamp 1698431365
transform 1 0 27664 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2552_
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2553_
timestamp 1698431365
transform 1 0 24752 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2554_
timestamp 1698431365
transform 1 0 26320 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2555_
timestamp 1698431365
transform 1 0 25872 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2556_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2557_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2558_
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2559_
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2560_
timestamp 1698431365
transform 1 0 32256 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2561_
timestamp 1698431365
transform -1 0 32592 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2562_
timestamp 1698431365
transform 1 0 34944 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2563_
timestamp 1698431365
transform 1 0 34720 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2564_
timestamp 1698431365
transform -1 0 8176 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2565_
timestamp 1698431365
transform 1 0 6496 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2566_
timestamp 1698431365
transform -1 0 5152 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2567_
timestamp 1698431365
transform 1 0 6944 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2568_
timestamp 1698431365
transform -1 0 6832 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2569_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3920 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2570_
timestamp 1698431365
transform 1 0 6048 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2571_
timestamp 1698431365
transform 1 0 2128 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2572_
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2573_
timestamp 1698431365
transform 1 0 11984 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2574_
timestamp 1698431365
transform 1 0 9296 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2575_
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2576_
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2577_
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2578_
timestamp 1698431365
transform 1 0 8960 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2579_
timestamp 1698431365
transform 1 0 16688 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2580_
timestamp 1698431365
transform 1 0 18592 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2581_
timestamp 1698431365
transform 1 0 11984 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2582_
timestamp 1698431365
transform 1 0 9184 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2583_
timestamp 1698431365
transform 1 0 15456 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2584_
timestamp 1698431365
transform 1 0 15456 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2585_
timestamp 1698431365
transform 1 0 2016 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2586_
timestamp 1698431365
transform 1 0 1680 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2587_
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2588_
timestamp 1698431365
transform -1 0 28448 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2589_
timestamp 1698431365
transform 1 0 11760 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2590_
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2591_
timestamp 1698431365
transform 1 0 15568 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2592_
timestamp 1698431365
transform 1 0 8512 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2593_
timestamp 1698431365
transform -1 0 27216 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2594_
timestamp 1698431365
transform 1 0 9856 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2595_
timestamp 1698431365
transform -1 0 22400 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2596_
timestamp 1698431365
transform 1 0 12320 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2597_
timestamp 1698431365
transform 1 0 8176 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2598_
timestamp 1698431365
transform 1 0 5936 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2599_
timestamp 1698431365
transform 1 0 5488 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2600_
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2601_
timestamp 1698431365
transform 1 0 2576 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2602_
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2603_
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2604_
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2605_
timestamp 1698431365
transform 1 0 2128 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2606_
timestamp 1698431365
transform 1 0 15456 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2607_
timestamp 1698431365
transform 1 0 17472 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2608_
timestamp 1698431365
transform -1 0 29680 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2609_
timestamp 1698431365
transform 1 0 19488 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2610_
timestamp 1698431365
transform 1 0 12768 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2611_
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2612_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15792 0 1 28224
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2613_
timestamp 1698431365
transform 1 0 25536 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2614_
timestamp 1698431365
transform 1 0 27888 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2615_
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2616_
timestamp 1698431365
transform 1 0 30352 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2617_
timestamp 1698431365
transform 1 0 31024 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2618_
timestamp 1698431365
transform 1 0 32704 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2619_
timestamp 1698431365
transform 1 0 35056 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2620_
timestamp 1698431365
transform -1 0 42448 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2621_
timestamp 1698431365
transform -1 0 45584 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2622_
timestamp 1698431365
transform 1 0 27328 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2623_
timestamp 1698431365
transform 1 0 41216 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2624_
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2625_
timestamp 1698431365
transform -1 0 49280 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2626_
timestamp 1698431365
transform 1 0 49392 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2627_
timestamp 1698431365
transform 1 0 50400 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2628_
timestamp 1698431365
transform -1 0 54208 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2629_
timestamp 1698431365
transform 1 0 48272 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2630_
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2631_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2632_
timestamp 1698431365
transform 1 0 37296 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2633_
timestamp 1698431365
transform 1 0 39088 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2634_
timestamp 1698431365
transform 1 0 39536 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2635_
timestamp 1698431365
transform -1 0 42784 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2636_
timestamp 1698431365
transform 1 0 41216 0 -1 45472
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2637_
timestamp 1698431365
transform -1 0 43232 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2638_
timestamp 1698431365
transform -1 0 48272 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2639_
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2640_
timestamp 1698431365
transform -1 0 55776 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2641_
timestamp 1698431365
transform 1 0 42448 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2642_
timestamp 1698431365
transform -1 0 54208 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2643_
timestamp 1698431365
transform -1 0 58352 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2644_
timestamp 1698431365
transform -1 0 58352 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2645_
timestamp 1698431365
transform -1 0 57008 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2646_
timestamp 1698431365
transform 1 0 40992 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2647_
timestamp 1698431365
transform 1 0 54320 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2648_
timestamp 1698431365
transform 1 0 53984 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2649_
timestamp 1698431365
transform 1 0 52080 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2650_
timestamp 1698431365
transform 1 0 50624 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2651_
timestamp 1698431365
transform 1 0 44688 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2652_
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2653_
timestamp 1698431365
transform 1 0 42784 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2654_
timestamp 1698431365
transform -1 0 41888 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2655_
timestamp 1698431365
transform 1 0 38752 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2656_
timestamp 1698431365
transform 1 0 37520 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2657_
timestamp 1698431365
transform 1 0 36064 0 -1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2658_
timestamp 1698431365
transform 1 0 35504 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2659_
timestamp 1698431365
transform 1 0 29792 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2660_
timestamp 1698431365
transform 1 0 29232 0 -1 28224
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2661_
timestamp 1698431365
transform 1 0 33488 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2662_
timestamp 1698431365
transform 1 0 36736 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2663_
timestamp 1698431365
transform -1 0 47936 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2664_
timestamp 1698431365
transform 1 0 33264 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2665_
timestamp 1698431365
transform 1 0 35728 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2666_
timestamp 1698431365
transform 1 0 19264 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2667_
timestamp 1698431365
transform 1 0 19488 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2668_
timestamp 1698431365
transform -1 0 32256 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2669_
timestamp 1698431365
transform -1 0 32256 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2670_
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2671_
timestamp 1698431365
transform 1 0 27216 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2672_
timestamp 1698431365
transform -1 0 34272 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2673_
timestamp 1698431365
transform 1 0 30800 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2674_
timestamp 1698431365
transform 1 0 28448 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2675_
timestamp 1698431365
transform 1 0 31248 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2676_
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2677_
timestamp 1698431365
transform 1 0 34272 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2678_
timestamp 1698431365
transform 1 0 34720 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2679_
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2680_
timestamp 1698431365
transform 1 0 34720 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2681_
timestamp 1698431365
transform 1 0 35616 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2682_
timestamp 1698431365
transform 1 0 31808 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2683_
timestamp 1698431365
transform 1 0 8064 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2684_
timestamp 1698431365
transform 1 0 7952 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2685_
timestamp 1698431365
transform 1 0 7952 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2686_
timestamp 1698431365
transform 1 0 8064 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2687_
timestamp 1698431365
transform 1 0 7952 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2688_
timestamp 1698431365
transform 1 0 6608 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2689_
timestamp 1698431365
transform 1 0 9856 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2690_
timestamp 1698431365
transform 1 0 12096 0 -1 54880
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2691_
timestamp 1698431365
transform 1 0 16912 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2692_
timestamp 1698431365
transform 1 0 15232 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2693_
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2694_
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2695_
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2696_
timestamp 1698431365
transform -1 0 9072 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2697_
timestamp 1698431365
transform 1 0 5264 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2698_
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2699_
timestamp 1698431365
transform -1 0 7840 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2700_
timestamp 1698431365
transform 1 0 5712 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2701_
timestamp 1698431365
transform -1 0 9184 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2702_
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2703_
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2704_
timestamp 1698431365
transform -1 0 8624 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2705_
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2706_
timestamp 1698431365
transform -1 0 4816 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2707_
timestamp 1698431365
transform -1 0 4816 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2708_
timestamp 1698431365
transform -1 0 4816 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2709_
timestamp 1698431365
transform -1 0 29120 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2710_
timestamp 1698431365
transform 1 0 23520 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2711_
timestamp 1698431365
transform 1 0 21056 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2712_
timestamp 1698431365
transform 1 0 15344 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2713_
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2714_
timestamp 1698431365
transform -1 0 29792 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2715_
timestamp 1698431365
transform 1 0 23632 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2716_
timestamp 1698431365
transform 1 0 19824 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2717_
timestamp 1698431365
transform 1 0 12096 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2718_
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2719_
timestamp 1698431365
transform -1 0 27216 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2720_
timestamp 1698431365
transform 1 0 22176 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2721_
timestamp 1698431365
transform -1 0 27664 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2722_
timestamp 1698431365
transform -1 0 28336 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2723_
timestamp 1698431365
transform -1 0 36512 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2724_
timestamp 1698431365
transform -1 0 38864 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2725_
timestamp 1698431365
transform 1 0 16800 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2726_
timestamp 1698431365
transform -1 0 23296 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2727_
timestamp 1698431365
transform -1 0 16128 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2728_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2729_
timestamp 1698431365
transform -1 0 32256 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2730_
timestamp 1698431365
transform 1 0 30128 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2731_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2732_
timestamp 1698431365
transform 1 0 19936 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2733_
timestamp 1698431365
transform -1 0 32704 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2734_
timestamp 1698431365
transform -1 0 34272 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2735_
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2736_
timestamp 1698431365
transform -1 0 39424 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2737_
timestamp 1698431365
transform 1 0 8288 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2738_
timestamp 1698431365
transform 1 0 6720 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2739_
timestamp 1698431365
transform 1 0 24864 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2740_
timestamp 1698431365
transform 1 0 28224 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2741_
timestamp 1698431365
transform 1 0 31024 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2742_
timestamp 1698431365
transform 1 0 34384 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2743_
timestamp 1698431365
transform 1 0 20272 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2744_
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2745_
timestamp 1698431365
transform 1 0 24416 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2746_
timestamp 1698431365
transform 1 0 27104 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2747_
timestamp 1698431365
transform 1 0 19264 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2748_
timestamp 1698431365
transform 1 0 21280 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2749_
timestamp 1698431365
transform 1 0 24528 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2750_
timestamp 1698431365
transform 1 0 27552 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2751_
timestamp 1698431365
transform -1 0 28336 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2752_
timestamp 1698431365
transform -1 0 31696 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2753_
timestamp 1698431365
transform 1 0 31024 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2754_
timestamp 1698431365
transform -1 0 38640 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2755_
timestamp 1698431365
transform 1 0 3248 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2756_
timestamp 1698431365
transform 1 0 5040 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__I asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__I
timestamp 1698431365
transform 1 0 29120 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A3
timestamp 1698431365
transform -1 0 14000 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1374__A1
timestamp 1698431365
transform 1 0 17920 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A1
timestamp 1698431365
transform -1 0 16128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A2
timestamp 1698431365
transform -1 0 17696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A1
timestamp 1698431365
transform 1 0 14560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A1
timestamp 1698431365
transform -1 0 11312 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__I
timestamp 1698431365
transform 1 0 17472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__I
timestamp 1698431365
transform 1 0 17136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A1
timestamp 1698431365
transform -1 0 10640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1464__I
timestamp 1698431365
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1476__S
timestamp 1698431365
transform 1 0 13216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__A2
timestamp 1698431365
transform -1 0 22736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__S
timestamp 1698431365
transform 1 0 15568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__S
timestamp 1698431365
transform -1 0 16352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__A2
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A2
timestamp 1698431365
transform -1 0 15680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__B
timestamp 1698431365
transform 1 0 16352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1553__I
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__I
timestamp 1698431365
transform 1 0 47600 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A1
timestamp 1698431365
transform 1 0 19376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A1
timestamp 1698431365
transform 1 0 26320 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A1
timestamp 1698431365
transform -1 0 20832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__B
timestamp 1698431365
transform 1 0 20160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__A1
timestamp 1698431365
transform 1 0 16128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__A1
timestamp 1698431365
transform -1 0 25200 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__B
timestamp 1698431365
transform -1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A1
timestamp 1698431365
transform -1 0 14896 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__B
timestamp 1698431365
transform -1 0 14560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__I
timestamp 1698431365
transform 1 0 26880 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__I
timestamp 1698431365
transform 1 0 23968 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A1
timestamp 1698431365
transform 1 0 11648 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__I
timestamp 1698431365
transform 1 0 16128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__A1
timestamp 1698431365
transform -1 0 18816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__A2
timestamp 1698431365
transform 1 0 19712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__I
timestamp 1698431365
transform 1 0 12432 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A1
timestamp 1698431365
transform 1 0 19824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__I
timestamp 1698431365
transform 1 0 17136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__I
timestamp 1698431365
transform 1 0 22624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A2
timestamp 1698431365
transform 1 0 13104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A2
timestamp 1698431365
transform 1 0 15792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A1
timestamp 1698431365
transform 1 0 19712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__A1
timestamp 1698431365
transform 1 0 21392 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__I
timestamp 1698431365
transform -1 0 16464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__A1
timestamp 1698431365
transform 1 0 19712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__A2
timestamp 1698431365
transform 1 0 19264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__I
timestamp 1698431365
transform -1 0 11648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__A1
timestamp 1698431365
transform 1 0 19824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__A2
timestamp 1698431365
transform 1 0 20048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__A1
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__I
timestamp 1698431365
transform -1 0 49168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A1
timestamp 1698431365
transform -1 0 15568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__I
timestamp 1698431365
transform 1 0 9856 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__A1
timestamp 1698431365
transform -1 0 8512 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__I
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A1
timestamp 1698431365
transform -1 0 7952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__A1
timestamp 1698431365
transform 1 0 7952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__A1
timestamp 1698431365
transform -1 0 14560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A1
timestamp 1698431365
transform 1 0 21392 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A2
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1773__C
timestamp 1698431365
transform -1 0 28448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__I
timestamp 1698431365
transform -1 0 27664 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__A1
timestamp 1698431365
transform -1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__A1
timestamp 1698431365
transform 1 0 26432 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__I
timestamp 1698431365
transform 1 0 51296 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__A1
timestamp 1698431365
transform 1 0 51744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__I
timestamp 1698431365
transform 1 0 27216 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__B
timestamp 1698431365
transform 1 0 33488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__B
timestamp 1698431365
transform -1 0 37072 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__A1
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__A1
timestamp 1698431365
transform 1 0 40992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__I
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__A1
timestamp 1698431365
transform 1 0 40320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__B
timestamp 1698431365
transform -1 0 41216 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__A1
timestamp 1698431365
transform 1 0 39200 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A1
timestamp 1698431365
transform -1 0 44352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__I
timestamp 1698431365
transform 1 0 44240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A2
timestamp 1698431365
transform 1 0 46144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__C
timestamp 1698431365
transform 1 0 46592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__I
timestamp 1698431365
transform 1 0 43120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__A2
timestamp 1698431365
transform 1 0 47040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__B
timestamp 1698431365
transform 1 0 42112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A1
timestamp 1698431365
transform 1 0 48048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__I
timestamp 1698431365
transform 1 0 47152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A2
timestamp 1698431365
transform 1 0 49952 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A1
timestamp 1698431365
transform -1 0 49616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A1
timestamp 1698431365
transform -1 0 47600 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__A1
timestamp 1698431365
transform 1 0 48944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A1
timestamp 1698431365
transform 1 0 53312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1956__A2
timestamp 1698431365
transform 1 0 52864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__A1
timestamp 1698431365
transform 1 0 53760 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__A1
timestamp 1698431365
transform -1 0 43344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A2
timestamp 1698431365
transform 1 0 44240 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__C
timestamp 1698431365
transform 1 0 46592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__B
timestamp 1698431365
transform 1 0 47040 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__B
timestamp 1698431365
transform -1 0 47712 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A2
timestamp 1698431365
transform -1 0 50064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__C
timestamp 1698431365
transform 1 0 53872 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__A1
timestamp 1698431365
transform 1 0 57792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A2
timestamp 1698431365
transform 1 0 58016 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__C
timestamp 1698431365
transform 1 0 52080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A1
timestamp 1698431365
transform 1 0 57120 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A2
timestamp 1698431365
transform 1 0 57456 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__C
timestamp 1698431365
transform 1 0 57008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__B
timestamp 1698431365
transform 1 0 48160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__A2
timestamp 1698431365
transform -1 0 51184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__C
timestamp 1698431365
transform -1 0 51520 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2027__A2
timestamp 1698431365
transform 1 0 42672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__A1
timestamp 1698431365
transform 1 0 41216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__A2
timestamp 1698431365
transform 1 0 44128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__C
timestamp 1698431365
transform 1 0 43680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A2
timestamp 1698431365
transform 1 0 55552 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__C
timestamp 1698431365
transform 1 0 54208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A1
timestamp 1698431365
transform -1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2048__A1
timestamp 1698431365
transform 1 0 54656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2057__A1
timestamp 1698431365
transform 1 0 54320 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__A2
timestamp 1698431365
transform 1 0 50848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__C
timestamp 1698431365
transform 1 0 50848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__B
timestamp 1698431365
transform 1 0 49616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2066__A2
timestamp 1698431365
transform 1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2066__C
timestamp 1698431365
transform 1 0 46704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__A2
timestamp 1698431365
transform -1 0 46928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__B
timestamp 1698431365
transform 1 0 48160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__B
timestamp 1698431365
transform 1 0 43904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2093__A2
timestamp 1698431365
transform 1 0 43344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2094__A1
timestamp 1698431365
transform 1 0 39648 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__B
timestamp 1698431365
transform 1 0 43568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__A2
timestamp 1698431365
transform -1 0 43344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__C
timestamp 1698431365
transform 1 0 42560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2109__A1
timestamp 1698431365
transform -1 0 39200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A2
timestamp 1698431365
transform 1 0 41888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__B
timestamp 1698431365
transform -1 0 41440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__A1
timestamp 1698431365
transform 1 0 39984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__A2
timestamp 1698431365
transform -1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__C
timestamp 1698431365
transform -1 0 34384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__A2
timestamp 1698431365
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__A1
timestamp 1698431365
transform -1 0 33712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2133__A2
timestamp 1698431365
transform 1 0 35056 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2133__C
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__A2
timestamp 1698431365
transform 1 0 35728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__C
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__A2
timestamp 1698431365
transform 1 0 35168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__C
timestamp 1698431365
transform 1 0 33488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2148__A1
timestamp 1698431365
transform 1 0 38304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__A1
timestamp 1698431365
transform -1 0 47152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__A2
timestamp 1698431365
transform 1 0 46032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A1
timestamp 1698431365
transform 1 0 45584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A2
timestamp 1698431365
transform -1 0 47600 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__A1
timestamp 1698431365
transform 1 0 34048 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__A1
timestamp 1698431365
transform -1 0 35728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__A2
timestamp 1698431365
transform 1 0 30128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2158__A2
timestamp 1698431365
transform 1 0 19824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2159__A2
timestamp 1698431365
transform 1 0 21392 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__A3
timestamp 1698431365
transform 1 0 20608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2167__B
timestamp 1698431365
transform 1 0 31248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__A1
timestamp 1698431365
transform -1 0 27104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__A2
timestamp 1698431365
transform 1 0 25536 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__B2
timestamp 1698431365
transform 1 0 25984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2211__A1
timestamp 1698431365
transform -1 0 27216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__B2
timestamp 1698431365
transform 1 0 29232 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2219__I
timestamp 1698431365
transform 1 0 25872 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2220__I
timestamp 1698431365
transform -1 0 23520 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2247__B
timestamp 1698431365
transform 1 0 31584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2264__A1
timestamp 1698431365
transform 1 0 23856 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A1
timestamp 1698431365
transform -1 0 28448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2268__B
timestamp 1698431365
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__A1
timestamp 1698431365
transform 1 0 26544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2278__B
timestamp 1698431365
transform -1 0 38192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2285__I
timestamp 1698431365
transform 1 0 33936 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2286__B
timestamp 1698431365
transform -1 0 34272 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A1
timestamp 1698431365
transform 1 0 27328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__B2
timestamp 1698431365
transform 1 0 28560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__A1
timestamp 1698431365
transform -1 0 32704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2316__A1
timestamp 1698431365
transform 1 0 11648 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2317__A1
timestamp 1698431365
transform 1 0 12208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2318__C
timestamp 1698431365
transform -1 0 14784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__A1
timestamp 1698431365
transform -1 0 15456 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A1
timestamp 1698431365
transform 1 0 17472 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A2
timestamp 1698431365
transform -1 0 18592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__A1
timestamp 1698431365
transform -1 0 9968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2332__A1
timestamp 1698431365
transform -1 0 16016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2337__B
timestamp 1698431365
transform 1 0 15008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2338__A1
timestamp 1698431365
transform 1 0 11760 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2345__A2
timestamp 1698431365
transform 1 0 15680 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2345__B
timestamp 1698431365
transform -1 0 16352 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2357__B
timestamp 1698431365
transform 1 0 19152 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A1
timestamp 1698431365
transform -1 0 11648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2409__I
timestamp 1698431365
transform 1 0 25872 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2410__B
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2415__B
timestamp 1698431365
transform 1 0 22624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__A1
timestamp 1698431365
transform -1 0 23520 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2429__A1
timestamp 1698431365
transform -1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__A1
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2431__A1
timestamp 1698431365
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2432__A1
timestamp 1698431365
transform 1 0 14672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__C
timestamp 1698431365
transform 1 0 24304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2458__A1
timestamp 1698431365
transform -1 0 22624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2465__A1
timestamp 1698431365
transform -1 0 25760 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A1
timestamp 1698431365
transform 1 0 25984 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2471__I
timestamp 1698431365
transform 1 0 28784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2472__A1
timestamp 1698431365
transform 1 0 24304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2475__I
timestamp 1698431365
transform 1 0 29232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2478__I
timestamp 1698431365
transform -1 0 14896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A2
timestamp 1698431365
transform -1 0 20048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__I
timestamp 1698431365
transform -1 0 16240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__A1
timestamp 1698431365
transform -1 0 15008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A1
timestamp 1698431365
transform 1 0 21952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A1
timestamp 1698431365
transform 1 0 23744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2509__A1
timestamp 1698431365
transform 1 0 25760 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__A1
timestamp 1698431365
transform 1 0 12208 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__I
timestamp 1698431365
transform 1 0 28448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A1
timestamp 1698431365
transform 1 0 22736 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2523__I
timestamp 1698431365
transform 1 0 30240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__A1
timestamp 1698431365
transform 1 0 26992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__I
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A1
timestamp 1698431365
transform -1 0 22960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A2
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__I
timestamp 1698431365
transform 1 0 29680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A1
timestamp 1698431365
transform 1 0 25648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__A1
timestamp 1698431365
transform 1 0 24416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__A2
timestamp 1698431365
transform -1 0 23408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__A1
timestamp 1698431365
transform 1 0 24192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__A1
timestamp 1698431365
transform 1 0 24528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__A1
timestamp 1698431365
transform 1 0 24864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2564__A1
timestamp 1698431365
transform -1 0 8624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2569__CLK
timestamp 1698431365
transform 1 0 7392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2570__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__CLK
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__CLK
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2574__CLK
timestamp 1698431365
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__CLK
timestamp 1698431365
transform 1 0 13104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__CLK
timestamp 1698431365
transform -1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__CLK
timestamp 1698431365
transform 1 0 12880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__CLK
timestamp 1698431365
transform 1 0 12432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__CLK
timestamp 1698431365
transform 1 0 20832 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2580__CLK
timestamp 1698431365
transform 1 0 22064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__CLK
timestamp 1698431365
transform 1 0 11760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__CLK
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__CLK
timestamp 1698431365
transform -1 0 15456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__CLK
timestamp 1698431365
transform 1 0 15232 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__CLK
timestamp 1698431365
transform 1 0 5712 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__CLK
timestamp 1698431365
transform -1 0 5152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2587__CLK
timestamp 1698431365
transform 1 0 47936 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2588__CLK
timestamp 1698431365
transform -1 0 28672 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__CLK
timestamp 1698431365
transform -1 0 14672 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__CLK
timestamp 1698431365
transform 1 0 12880 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2591__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__CLK
timestamp 1698431365
transform 1 0 8288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__CLK
timestamp 1698431365
transform -1 0 27664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__CLK
timestamp 1698431365
transform 1 0 13328 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__CLK
timestamp 1698431365
transform 1 0 18928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__CLK
timestamp 1698431365
transform 1 0 10976 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__CLK
timestamp 1698431365
transform 1 0 11424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2598__CLK
timestamp 1698431365
transform 1 0 9184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2599__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__CLK
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2601__CLK
timestamp 1698431365
transform 1 0 5824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2602__CLK
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2603__CLK
timestamp 1698431365
transform 1 0 5712 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2604__CLK
timestamp 1698431365
transform 1 0 5040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2605__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2606__CLK
timestamp 1698431365
transform 1 0 15232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__CLK
timestamp 1698431365
transform 1 0 20832 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__CLK
timestamp 1698431365
transform 1 0 26208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__CLK
timestamp 1698431365
transform 1 0 19264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__CLK
timestamp 1698431365
transform 1 0 16240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__CLK
timestamp 1698431365
transform 1 0 16800 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__CLK
timestamp 1698431365
transform 1 0 19488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2613__CLK
timestamp 1698431365
transform 1 0 27664 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__CLK
timestamp 1698431365
transform 1 0 31360 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__CLK
timestamp 1698431365
transform 1 0 32256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2616__CLK
timestamp 1698431365
transform 1 0 33824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__CLK
timestamp 1698431365
transform 1 0 34272 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__CLK
timestamp 1698431365
transform 1 0 34832 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2620__CLK
timestamp 1698431365
transform 1 0 42112 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__CLK
timestamp 1698431365
transform 1 0 45808 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2622__CLK
timestamp 1698431365
transform 1 0 30800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__CLK
timestamp 1698431365
transform 1 0 44464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__CLK
timestamp 1698431365
transform -1 0 48384 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__CLK
timestamp 1698431365
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__CLK
timestamp 1698431365
transform 1 0 49168 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__CLK
timestamp 1698431365
transform 1 0 49168 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2628__CLK
timestamp 1698431365
transform 1 0 51632 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__CLK
timestamp 1698431365
transform 1 0 48048 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__CLK
timestamp 1698431365
transform 1 0 52080 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__CLK
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__CLK
timestamp 1698431365
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__CLK
timestamp 1698431365
transform 1 0 43344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__CLK
timestamp 1698431365
transform 1 0 43008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__CLK
timestamp 1698431365
transform 1 0 43008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2636__CLK
timestamp 1698431365
transform 1 0 44912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__CLK
timestamp 1698431365
transform 1 0 42784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__CLK
timestamp 1698431365
transform -1 0 48720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__CLK
timestamp 1698431365
transform 1 0 48160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__CLK
timestamp 1698431365
transform -1 0 53536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__CLK
timestamp 1698431365
transform 1 0 45920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__CLK
timestamp 1698431365
transform -1 0 50848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2643__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__CLK
timestamp 1698431365
transform 1 0 57344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__CLK
timestamp 1698431365
transform 1 0 54432 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__CLK
timestamp 1698431365
transform 1 0 44912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__CLK
timestamp 1698431365
transform 1 0 54992 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__CLK
timestamp 1698431365
transform 1 0 54096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__CLK
timestamp 1698431365
transform 1 0 53648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2650__CLK
timestamp 1698431365
transform 1 0 50400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__CLK
timestamp 1698431365
transform 1 0 48160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__CLK
timestamp 1698431365
transform 1 0 48160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2653__CLK
timestamp 1698431365
transform 1 0 45136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2654__CLK
timestamp 1698431365
transform 1 0 41888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2655__CLK
timestamp 1698431365
transform 1 0 38528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2656__CLK
timestamp 1698431365
transform 1 0 38304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2657__CLK
timestamp 1698431365
transform 1 0 39424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2658__CLK
timestamp 1698431365
transform 1 0 35504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2659__CLK
timestamp 1698431365
transform 1 0 29568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__CLK
timestamp 1698431365
transform 1 0 29680 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__CLK
timestamp 1698431365
transform 1 0 35952 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__CLK
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__CLK
timestamp 1698431365
transform 1 0 48160 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2664__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2665__CLK
timestamp 1698431365
transform -1 0 35728 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2666__CLK
timestamp 1698431365
transform 1 0 19040 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2667__CLK
timestamp 1698431365
transform 1 0 19936 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2670__CLK
timestamp 1698431365
transform 1 0 32480 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__CLK
timestamp 1698431365
transform 1 0 32256 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__CLK
timestamp 1698431365
transform 1 0 34496 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__CLK
timestamp 1698431365
transform 1 0 34272 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2674__CLK
timestamp 1698431365
transform -1 0 32144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2675__CLK
timestamp 1698431365
transform 1 0 34720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__CLK
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2677__CLK
timestamp 1698431365
transform 1 0 37520 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__CLK
timestamp 1698431365
transform 1 0 34496 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2679__CLK
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__CLK
timestamp 1698431365
transform 1 0 34496 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__CLK
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__CLK
timestamp 1698431365
transform 1 0 34496 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__CLK
timestamp 1698431365
transform 1 0 7840 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__CLK
timestamp 1698431365
transform -1 0 11088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__CLK
timestamp 1698431365
transform 1 0 11872 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2686__CLK
timestamp 1698431365
transform 1 0 11312 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2687__CLK
timestamp 1698431365
transform 1 0 12320 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__CLK
timestamp 1698431365
transform 1 0 9856 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__CLK
timestamp 1698431365
transform 1 0 11872 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__CLK
timestamp 1698431365
transform 1 0 20944 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__CLK
timestamp 1698431365
transform 1 0 18704 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__CLK
timestamp 1698431365
transform 1 0 5040 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__CLK
timestamp 1698431365
transform 1 0 5040 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__CLK
timestamp 1698431365
transform 1 0 5040 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__CLK
timestamp 1698431365
transform 1 0 9296 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__CLK
timestamp 1698431365
transform 1 0 8736 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__CLK
timestamp 1698431365
transform 1 0 7840 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__CLK
timestamp 1698431365
transform 1 0 9408 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__CLK
timestamp 1698431365
transform 1 0 5040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__CLK
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__CLK
timestamp 1698431365
transform 1 0 8848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__CLK
timestamp 1698431365
transform -1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__CLK
timestamp 1698431365
transform 1 0 5712 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__CLK
timestamp 1698431365
transform 1 0 5040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__CLK
timestamp 1698431365
transform 1 0 5040 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2709__CLK
timestamp 1698431365
transform 1 0 29232 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__CLK
timestamp 1698431365
transform 1 0 26992 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__CLK
timestamp 1698431365
transform -1 0 24752 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__CLK
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__CLK
timestamp 1698431365
transform 1 0 14896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2714__CLK
timestamp 1698431365
transform 1 0 30016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2715__CLK
timestamp 1698431365
transform 1 0 22736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2716__CLK
timestamp 1698431365
transform 1 0 19600 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__CLK
timestamp 1698431365
transform 1 0 15568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2718__CLK
timestamp 1698431365
transform 1 0 15904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2719__CLK
timestamp 1698431365
transform 1 0 27440 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2720__CLK
timestamp 1698431365
transform 1 0 21392 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2721__CLK
timestamp 1698431365
transform -1 0 30576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2722__CLK
timestamp 1698431365
transform 1 0 28560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2723__CLK
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__CLK
timestamp 1698431365
transform 1 0 39088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2725__CLK
timestamp 1698431365
transform -1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__CLK
timestamp 1698431365
transform 1 0 23520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__CLK
timestamp 1698431365
transform -1 0 12992 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2728__CLK
timestamp 1698431365
transform 1 0 13440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2729__CLK
timestamp 1698431365
transform 1 0 32480 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2730__CLK
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__CLK
timestamp 1698431365
transform 1 0 20720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__CLK
timestamp 1698431365
transform -1 0 22736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__CLK
timestamp 1698431365
transform 1 0 34496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__CLK
timestamp 1698431365
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__CLK
timestamp 1698431365
transform 1 0 39648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__CLK
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2738__CLK
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2739__CLK
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2740__CLK
timestamp 1698431365
transform 1 0 28000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__CLK
timestamp 1698431365
transform 1 0 30800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2742__CLK
timestamp 1698431365
transform 1 0 37856 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__CLK
timestamp 1698431365
transform 1 0 23744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2744__CLK
timestamp 1698431365
transform 1 0 25312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__CLK
timestamp 1698431365
transform 1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2746__CLK
timestamp 1698431365
transform 1 0 26880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2747__CLK
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2748__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2749__CLK
timestamp 1698431365
transform 1 0 27776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2750__CLK
timestamp 1698431365
transform 1 0 27328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2751__CLK
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2752__CLK
timestamp 1698431365
transform 1 0 27888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2753__CLK
timestamp 1698431365
transform 1 0 30800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2754__CLK
timestamp 1698431365
transform 1 0 38864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2755__CLK
timestamp 1698431365
transform 1 0 6496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2756__CLK
timestamp 1698431365
transform 1 0 8512 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 28336 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 13216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 12544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 28000 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 8848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 9632 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 18032 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 20272 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 35168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 33936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 50288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 48832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 35504 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 34496 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 44576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 44912 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 21840 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 21280 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 15904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 15680 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 4704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output11_I
timestamp 1698431365
transform 1 0 29232 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30016 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_wb_clk_i asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1698431365
transform 1 0 23184 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1698431365
transform -1 0 28000 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1698431365
transform -1 0 8624 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1698431365
transform 1 0 6160 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1698431365
transform -1 0 18032 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1698431365
transform 1 0 15568 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1698431365
transform -1 0 38192 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1698431365
transform -1 0 37072 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1698431365
transform -1 0 50064 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1698431365
transform 1 0 32368 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1698431365
transform -1 0 33712 0 1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1698431365
transform -1 0 47712 0 -1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1698431365
transform -1 0 48048 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_158
timestamp 1698431365
transform 1 0 19040 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_166
timestamp 1698431365
transform 1 0 19936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_168
timestamp 1698431365
transform 1 0 20160 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_198
timestamp 1698431365
transform 1 0 23520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_202
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_123
timestamp 1698431365
transform 1 0 15120 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_155
timestamp 1698431365
transform 1 0 18704 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_163
timestamp 1698431365
transform 1 0 19600 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_167
timestamp 1698431365
transform 1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_212
timestamp 1698431365
transform 1 0 25088 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_216
timestamp 1698431365
transform 1 0 25536 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_224
timestamp 1698431365
transform 1 0 26432 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_230
timestamp 1698431365
transform 1 0 27104 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_238
timestamp 1698431365
transform 1 0 28000 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_242
timestamp 1698431365
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698431365
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_88
timestamp 1698431365
transform 1 0 11200 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_92
timestamp 1698431365
transform 1 0 11648 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_124
timestamp 1698431365
transform 1 0 15232 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_132
timestamp 1698431365
transform 1 0 16128 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_204
timestamp 1698431365
transform 1 0 24192 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_208
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_214
timestamp 1698431365
transform 1 0 25312 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_259
timestamp 1698431365
transform 1 0 30352 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_69
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_99
timestamp 1698431365
transform 1 0 12432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698431365
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_113
timestamp 1698431365
transform 1 0 14000 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_129
timestamp 1698431365
transform 1 0 15792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_131
timestamp 1698431365
transform 1 0 16016 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_134
timestamp 1698431365
transform 1 0 16352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_151
timestamp 1698431365
transform 1 0 18256 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_159
timestamp 1698431365
transform 1 0 19152 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_163
timestamp 1698431365
transform 1 0 19600 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_167
timestamp 1698431365
transform 1 0 20048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_185
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_191
timestamp 1698431365
transform 1 0 22736 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_199
timestamp 1698431365
transform 1 0 23632 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_203
timestamp 1698431365
transform 1 0 24080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_205
timestamp 1698431365
transform 1 0 24304 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_76
timestamp 1698431365
transform 1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_84
timestamp 1698431365
transform 1 0 10752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_100
timestamp 1698431365
transform 1 0 12544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_132
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_157
timestamp 1698431365
transform 1 0 18928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_159
timestamp 1698431365
transform 1 0 19152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_189
timestamp 1698431365
transform 1 0 22512 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_193
timestamp 1698431365
transform 1 0 22960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_197
timestamp 1698431365
transform 1 0 23408 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_205
timestamp 1698431365
transform 1 0 24304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_219
timestamp 1698431365
transform 1 0 25872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_221
timestamp 1698431365
transform 1 0 26096 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_226
timestamp 1698431365
transform 1 0 26656 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_230
timestamp 1698431365
transform 1 0 27104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_251
timestamp 1698431365
transform 1 0 29456 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_267
timestamp 1698431365
transform 1 0 31248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_275
timestamp 1698431365
transform 1 0 32144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698431365
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_85
timestamp 1698431365
transform 1 0 10864 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_89
timestamp 1698431365
transform 1 0 11312 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_92
timestamp 1698431365
transform 1 0 11648 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_100
timestamp 1698431365
transform 1 0 12544 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_123
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_165
timestamp 1698431365
transform 1 0 19824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_169
timestamp 1698431365
transform 1 0 20272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_204
timestamp 1698431365
transform 1 0 24192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_208
timestamp 1698431365
transform 1 0 24640 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_212
timestamp 1698431365
transform 1 0 25088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_220
timestamp 1698431365
transform 1 0 25984 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_228
timestamp 1698431365
transform 1 0 26880 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_234
timestamp 1698431365
transform 1 0 27552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_238
timestamp 1698431365
transform 1 0 28000 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_242
timestamp 1698431365
transform 1 0 28448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_257
timestamp 1698431365
transform 1 0 30128 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_289
timestamp 1698431365
transform 1 0 33712 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_305
timestamp 1698431365
transform 1 0 35504 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_313
timestamp 1698431365
transform 1 0 36400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_489
timestamp 1698431365
transform 1 0 56112 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_505
timestamp 1698431365
transform 1 0 57904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_36
timestamp 1698431365
transform 1 0 5376 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_78
timestamp 1698431365
transform 1 0 10080 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_94
timestamp 1698431365
transform 1 0 11872 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_110
timestamp 1698431365
transform 1 0 13664 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_126
timestamp 1698431365
transform 1 0 15456 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_134
timestamp 1698431365
transform 1 0 16352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_138
timestamp 1698431365
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_158
timestamp 1698431365
transform 1 0 19040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_162
timestamp 1698431365
transform 1 0 19488 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_166
timestamp 1698431365
transform 1 0 19936 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_168
timestamp 1698431365
transform 1 0 20160 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_231
timestamp 1698431365
transform 1 0 27216 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_233
timestamp 1698431365
transform 1 0 27440 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_263
timestamp 1698431365
transform 1 0 30800 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_51
timestamp 1698431365
transform 1 0 7056 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_59
timestamp 1698431365
transform 1 0 7952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_123
timestamp 1698431365
transform 1 0 15120 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_131
timestamp 1698431365
transform 1 0 16016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_135
timestamp 1698431365
transform 1 0 16464 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_143
timestamp 1698431365
transform 1 0 17360 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_236
timestamp 1698431365
transform 1 0 27776 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_243
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_286
timestamp 1698431365
transform 1 0 33376 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_302
timestamp 1698431365
transform 1 0 35168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_310
timestamp 1698431365
transform 1 0 36064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698431365
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_489
timestamp 1698431365
transform 1 0 56112 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_505
timestamp 1698431365
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_42
timestamp 1698431365
transform 1 0 6048 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_46
timestamp 1698431365
transform 1 0 6496 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_48
timestamp 1698431365
transform 1 0 6720 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_64
timestamp 1698431365
transform 1 0 8512 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_84
timestamp 1698431365
transform 1 0 10752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_88
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_172
timestamp 1698431365
transform 1 0 20608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_176
timestamp 1698431365
transform 1 0 21056 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_184
timestamp 1698431365
transform 1 0 21952 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_188
timestamp 1698431365
transform 1 0 22400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_196
timestamp 1698431365
transform 1 0 23296 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_233
timestamp 1698431365
transform 1 0 27440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_277
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698431365
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_10
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_14
timestamp 1698431365
transform 1 0 2912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_16
timestamp 1698431365
transform 1 0 3136 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_23
timestamp 1698431365
transform 1 0 3920 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_31
timestamp 1698431365
transform 1 0 4816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_49
timestamp 1698431365
transform 1 0 6832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_66
timestamp 1698431365
transform 1 0 8736 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_72
timestamp 1698431365
transform 1 0 9408 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_80
timestamp 1698431365
transform 1 0 10304 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_84
timestamp 1698431365
transform 1 0 10752 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_113
timestamp 1698431365
transform 1 0 14000 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_121
timestamp 1698431365
transform 1 0 14896 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_123
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_181
timestamp 1698431365
transform 1 0 21616 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_195
timestamp 1698431365
transform 1 0 23184 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_214
timestamp 1698431365
transform 1 0 25312 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_216
timestamp 1698431365
transform 1 0 25536 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_229
timestamp 1698431365
transform 1 0 26992 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_255
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_271
timestamp 1698431365
transform 1 0 31696 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_278
timestamp 1698431365
transform 1 0 32480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_297
timestamp 1698431365
transform 1 0 34608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_299
timestamp 1698431365
transform 1 0 34832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698431365
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_489
timestamp 1698431365
transform 1 0 56112 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_505
timestamp 1698431365
transform 1 0 57904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_6
timestamp 1698431365
transform 1 0 2016 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_36
timestamp 1698431365
transform 1 0 5376 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_40
timestamp 1698431365
transform 1 0 5824 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_101
timestamp 1698431365
transform 1 0 12656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_103
timestamp 1698431365
transform 1 0 12880 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_106
timestamp 1698431365
transform 1 0 13216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_125
timestamp 1698431365
transform 1 0 15344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_129
timestamp 1698431365
transform 1 0 15792 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_137
timestamp 1698431365
transform 1 0 16688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1698431365
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_158
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_162
timestamp 1698431365
transform 1 0 19488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_164
timestamp 1698431365
transform 1 0 19712 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_196
timestamp 1698431365
transform 1 0 23296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_200
timestamp 1698431365
transform 1 0 23744 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_216
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_230
timestamp 1698431365
transform 1 0 27104 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_238
timestamp 1698431365
transform 1 0 28000 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_249
timestamp 1698431365
transform 1 0 29232 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_265
timestamp 1698431365
transform 1 0 31024 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_273
timestamp 1698431365
transform 1 0 31920 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_340
timestamp 1698431365
transform 1 0 39424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_344
timestamp 1698431365
transform 1 0 39872 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_31
timestamp 1698431365
transform 1 0 4816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_58
timestamp 1698431365
transform 1 0 7840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_62
timestamp 1698431365
transform 1 0 8288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_122
timestamp 1698431365
transform 1 0 15008 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_138
timestamp 1698431365
transform 1 0 16800 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_146
timestamp 1698431365
transform 1 0 17696 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_153
timestamp 1698431365
transform 1 0 18480 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_155
timestamp 1698431365
transform 1 0 18704 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_191
timestamp 1698431365
transform 1 0 22736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_193
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_234
timestamp 1698431365
transform 1 0 27552 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_238
timestamp 1698431365
transform 1 0 28000 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_276
timestamp 1698431365
transform 1 0 32256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_280
timestamp 1698431365
transform 1 0 32704 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_296
timestamp 1698431365
transform 1 0 34496 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_310
timestamp 1698431365
transform 1 0 36064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698431365
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_489
timestamp 1698431365
transform 1 0 56112 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_505
timestamp 1698431365
transform 1 0 57904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_16
timestamp 1698431365
transform 1 0 3136 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_24
timestamp 1698431365
transform 1 0 4032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_28
timestamp 1698431365
transform 1 0 4480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_30
timestamp 1698431365
transform 1 0 4704 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_46
timestamp 1698431365
transform 1 0 6496 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_54
timestamp 1698431365
transform 1 0 7392 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_64
timestamp 1698431365
transform 1 0 8512 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_132
timestamp 1698431365
transform 1 0 16128 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_192
timestamp 1698431365
transform 1 0 22848 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_196
timestamp 1698431365
transform 1 0 23296 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698431365
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_238
timestamp 1698431365
transform 1 0 28000 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_242
timestamp 1698431365
transform 1 0 28448 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_244
timestamp 1698431365
transform 1 0 28672 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_253
timestamp 1698431365
transform 1 0 29680 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_269
timestamp 1698431365
transform 1 0 31472 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_297
timestamp 1698431365
transform 1 0 34608 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_301
timestamp 1698431365
transform 1 0 35056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_303
timestamp 1698431365
transform 1 0 35280 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_319
timestamp 1698431365
transform 1 0 37072 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_335
timestamp 1698431365
transform 1 0 38864 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_343
timestamp 1698431365
transform 1 0 39760 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698431365
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_31
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_39
timestamp 1698431365
transform 1 0 5712 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_42
timestamp 1698431365
transform 1 0 6048 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_46
timestamp 1698431365
transform 1 0 6496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_83
timestamp 1698431365
transform 1 0 10640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_100
timestamp 1698431365
transform 1 0 12544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_121
timestamp 1698431365
transform 1 0 14896 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_129
timestamp 1698431365
transform 1 0 15792 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_167
timestamp 1698431365
transform 1 0 20048 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_231
timestamp 1698431365
transform 1 0 27216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_294
timestamp 1698431365
transform 1 0 34272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_298
timestamp 1698431365
transform 1 0 34720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_489
timestamp 1698431365
transform 1 0 56112 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_505
timestamp 1698431365
transform 1 0 57904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_4
timestamp 1698431365
transform 1 0 1792 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_55
timestamp 1698431365
transform 1 0 7504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_59
timestamp 1698431365
transform 1 0 7952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_61
timestamp 1698431365
transform 1 0 8176 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_98
timestamp 1698431365
transform 1 0 12320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_102
timestamp 1698431365
transform 1 0 12768 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_106
timestamp 1698431365
transform 1 0 13216 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_112
timestamp 1698431365
transform 1 0 13888 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_118
timestamp 1698431365
transform 1 0 14560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_122
timestamp 1698431365
transform 1 0 15008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_124
timestamp 1698431365
transform 1 0 15232 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_127
timestamp 1698431365
transform 1 0 15568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_148
timestamp 1698431365
transform 1 0 17920 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_164
timestamp 1698431365
transform 1 0 19712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_195
timestamp 1698431365
transform 1 0 23184 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_199
timestamp 1698431365
transform 1 0 23632 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_234
timestamp 1698431365
transform 1 0 27552 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_250
timestamp 1698431365
transform 1 0 29344 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_258
timestamp 1698431365
transform 1 0 30240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_260
timestamp 1698431365
transform 1 0 30464 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_298
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_335
timestamp 1698431365
transform 1 0 38864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_339
timestamp 1698431365
transform 1 0 39312 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_347
timestamp 1698431365
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698431365
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_18
timestamp 1698431365
transform 1 0 3360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_26
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_91
timestamp 1698431365
transform 1 0 11536 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_95
timestamp 1698431365
transform 1 0 11984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_116
timestamp 1698431365
transform 1 0 14336 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_135
timestamp 1698431365
transform 1 0 16464 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_142
timestamp 1698431365
transform 1 0 17248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_146
timestamp 1698431365
transform 1 0 17696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_156
timestamp 1698431365
transform 1 0 18816 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_236
timestamp 1698431365
transform 1 0 27776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_240
timestamp 1698431365
transform 1 0 28224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_272
timestamp 1698431365
transform 1 0 31808 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_288
timestamp 1698431365
transform 1 0 33600 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_296
timestamp 1698431365
transform 1 0 34496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_489
timestamp 1698431365
transform 1 0 56112 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_505
timestamp 1698431365
transform 1 0 57904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_34
timestamp 1698431365
transform 1 0 5152 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_46
timestamp 1698431365
transform 1 0 6496 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_48
timestamp 1698431365
transform 1 0 6720 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_53
timestamp 1698431365
transform 1 0 7280 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_55
timestamp 1698431365
transform 1 0 7504 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_62
timestamp 1698431365
transform 1 0 8288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_76
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_82
timestamp 1698431365
transform 1 0 10528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_84
timestamp 1698431365
transform 1 0 10752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_89
timestamp 1698431365
transform 1 0 11312 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_105
timestamp 1698431365
transform 1 0 13104 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_112
timestamp 1698431365
transform 1 0 13888 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_116
timestamp 1698431365
transform 1 0 14336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_118
timestamp 1698431365
transform 1 0 14560 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_127
timestamp 1698431365
transform 1 0 15568 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_171
timestamp 1698431365
transform 1 0 20496 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_175
timestamp 1698431365
transform 1 0 20944 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_248
timestamp 1698431365
transform 1 0 29120 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_250
timestamp 1698431365
transform 1 0 29344 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_301
timestamp 1698431365
transform 1 0 35056 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_333
timestamp 1698431365
transform 1 0 38640 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698431365
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_31
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_52
timestamp 1698431365
transform 1 0 7168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_60
timestamp 1698431365
transform 1 0 8064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_74
timestamp 1698431365
transform 1 0 9632 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_78
timestamp 1698431365
transform 1 0 10080 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_86
timestamp 1698431365
transform 1 0 10976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_109
timestamp 1698431365
transform 1 0 13552 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_118
timestamp 1698431365
transform 1 0 14560 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_132
timestamp 1698431365
transform 1 0 16128 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_139
timestamp 1698431365
transform 1 0 16912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_143
timestamp 1698431365
transform 1 0 17360 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_182
timestamp 1698431365
transform 1 0 21728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_198
timestamp 1698431365
transform 1 0 23520 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_217
timestamp 1698431365
transform 1 0 25648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_237
timestamp 1698431365
transform 1 0 27888 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_257
timestamp 1698431365
transform 1 0 30128 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_264
timestamp 1698431365
transform 1 0 30912 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_268
timestamp 1698431365
transform 1 0 31360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_321
timestamp 1698431365
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_489
timestamp 1698431365
transform 1 0 56112 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_505
timestamp 1698431365
transform 1 0 57904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_82
timestamp 1698431365
transform 1 0 10528 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_106
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_108
timestamp 1698431365
transform 1 0 13440 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_127
timestamp 1698431365
transform 1 0 15568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698431365
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_187
timestamp 1698431365
transform 1 0 22288 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_191
timestamp 1698431365
transform 1 0 22736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_193
timestamp 1698431365
transform 1 0 22960 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698431365
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_222
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_230
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_234
timestamp 1698431365
transform 1 0 27552 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_236
timestamp 1698431365
transform 1 0 27776 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_243
timestamp 1698431365
transform 1 0 28560 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_257
timestamp 1698431365
transform 1 0 30128 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_261
timestamp 1698431365
transform 1 0 30576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_265
timestamp 1698431365
transform 1 0 31024 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_273
timestamp 1698431365
transform 1 0 31920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698431365
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_286
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_294
timestamp 1698431365
transform 1 0 34272 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_333
timestamp 1698431365
transform 1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_337
timestamp 1698431365
transform 1 0 39088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_345
timestamp 1698431365
transform 1 0 39984 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698431365
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698431365
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_18
timestamp 1698431365
transform 1 0 3360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_41
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_45
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_47
timestamp 1698431365
transform 1 0 6608 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_71
timestamp 1698431365
transform 1 0 9296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_79
timestamp 1698431365
transform 1 0 10192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_81
timestamp 1698431365
transform 1 0 10416 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_92
timestamp 1698431365
transform 1 0 11648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_94
timestamp 1698431365
transform 1 0 11872 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_111
timestamp 1698431365
transform 1 0 13776 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_126
timestamp 1698431365
transform 1 0 15456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_138
timestamp 1698431365
transform 1 0 16800 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_154
timestamp 1698431365
transform 1 0 18592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_156
timestamp 1698431365
transform 1 0 18816 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_163
timestamp 1698431365
transform 1 0 19600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_167
timestamp 1698431365
transform 1 0 20048 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_179
timestamp 1698431365
transform 1 0 21392 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_192
timestamp 1698431365
transform 1 0 22848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_194
timestamp 1698431365
transform 1 0 23072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_203
timestamp 1698431365
transform 1 0 24080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_207
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_209
timestamp 1698431365
transform 1 0 24752 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_212
timestamp 1698431365
transform 1 0 25088 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_220
timestamp 1698431365
transform 1 0 25984 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_224
timestamp 1698431365
transform 1 0 26432 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_231
timestamp 1698431365
transform 1 0 27216 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_235
timestamp 1698431365
transform 1 0 27664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_237
timestamp 1698431365
transform 1 0 27888 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_240
timestamp 1698431365
transform 1 0 28224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_262
timestamp 1698431365
transform 1 0 30688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_264
timestamp 1698431365
transform 1 0 30912 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_294
timestamp 1698431365
transform 1 0 34272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_298
timestamp 1698431365
transform 1 0 34720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_321
timestamp 1698431365
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698431365
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_489
timestamp 1698431365
transform 1 0 56112 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_505
timestamp 1698431365
transform 1 0 57904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_15
timestamp 1698431365
transform 1 0 3024 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_46
timestamp 1698431365
transform 1 0 6496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_56
timestamp 1698431365
transform 1 0 7616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_58
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_61
timestamp 1698431365
transform 1 0 8176 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_91
timestamp 1698431365
transform 1 0 11536 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_99
timestamp 1698431365
transform 1 0 12432 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_103
timestamp 1698431365
transform 1 0 12880 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_123
timestamp 1698431365
transform 1 0 15120 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_172
timestamp 1698431365
transform 1 0 20608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_176
timestamp 1698431365
transform 1 0 21056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_189
timestamp 1698431365
transform 1 0 22512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_221
timestamp 1698431365
transform 1 0 26096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_269
timestamp 1698431365
transform 1 0 31472 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_290
timestamp 1698431365
transform 1 0 33824 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_292
timestamp 1698431365
transform 1 0 34048 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_324
timestamp 1698431365
transform 1 0 37632 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_328
timestamp 1698431365
transform 1 0 38080 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_334
timestamp 1698431365
transform 1 0 38752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_338
timestamp 1698431365
transform 1 0 39200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_358
timestamp 1698431365
transform 1 0 41440 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_374
timestamp 1698431365
transform 1 0 43232 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_382
timestamp 1698431365
transform 1 0 44128 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_386
timestamp 1698431365
transform 1 0 44576 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_416
timestamp 1698431365
transform 1 0 47936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_31
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_52
timestamp 1698431365
transform 1 0 7168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_54
timestamp 1698431365
transform 1 0 7392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_71
timestamp 1698431365
transform 1 0 9296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_83
timestamp 1698431365
transform 1 0 10640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_91
timestamp 1698431365
transform 1 0 11536 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_99
timestamp 1698431365
transform 1 0 12432 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_103
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_117
timestamp 1698431365
transform 1 0 14448 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_135
timestamp 1698431365
transform 1 0 16464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_166
timestamp 1698431365
transform 1 0 19936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_168
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_181
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_189
timestamp 1698431365
transform 1 0 22512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_205
timestamp 1698431365
transform 1 0 24304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_209
timestamp 1698431365
transform 1 0 24752 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_239
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_253
timestamp 1698431365
transform 1 0 29680 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_269
timestamp 1698431365
transform 1 0 31472 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_273
timestamp 1698431365
transform 1 0 31920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_275
timestamp 1698431365
transform 1 0 32144 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_291
timestamp 1698431365
transform 1 0 33936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_293
timestamp 1698431365
transform 1 0 34160 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_319
timestamp 1698431365
transform 1 0 37072 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_371
timestamp 1698431365
transform 1 0 42896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_375
timestamp 1698431365
transform 1 0 43344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_379
timestamp 1698431365
transform 1 0 43792 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_416
timestamp 1698431365
transform 1 0 47936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_420
timestamp 1698431365
transform 1 0 48384 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_452
timestamp 1698431365
transform 1 0 51968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_454
timestamp 1698431365
transform 1 0 52192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_489
timestamp 1698431365
transform 1 0 56112 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_505
timestamp 1698431365
transform 1 0 57904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_6
timestamp 1698431365
transform 1 0 2016 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_36
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_40
timestamp 1698431365
transform 1 0 5824 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_48
timestamp 1698431365
transform 1 0 6720 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_80
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_104
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_108
timestamp 1698431365
transform 1 0 13440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_120
timestamp 1698431365
transform 1 0 14784 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_128
timestamp 1698431365
transform 1 0 15680 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_135
timestamp 1698431365
transform 1 0 16464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_146
timestamp 1698431365
transform 1 0 17696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_163
timestamp 1698431365
transform 1 0 19600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_176
timestamp 1698431365
transform 1 0 21056 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_183
timestamp 1698431365
transform 1 0 21840 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_185
timestamp 1698431365
transform 1 0 22064 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_196
timestamp 1698431365
transform 1 0 23296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_198
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_227
timestamp 1698431365
transform 1 0 26768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_231
timestamp 1698431365
transform 1 0 27216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_233
timestamp 1698431365
transform 1 0 27440 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_240
timestamp 1698431365
transform 1 0 28224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_244
timestamp 1698431365
transform 1 0 28672 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_248
timestamp 1698431365
transform 1 0 29120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_256
timestamp 1698431365
transform 1 0 30016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_260
timestamp 1698431365
transform 1 0 30464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_262
timestamp 1698431365
transform 1 0 30688 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_265
timestamp 1698431365
transform 1 0 31024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_297
timestamp 1698431365
transform 1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_299
timestamp 1698431365
transform 1 0 34832 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_394
timestamp 1698431365
transform 1 0 45472 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_402
timestamp 1698431365
transform 1 0 46368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_404
timestamp 1698431365
transform 1 0 46592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_418
timestamp 1698431365
transform 1 0 48160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_438
timestamp 1698431365
transform 1 0 50400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_444
timestamp 1698431365
transform 1 0 51072 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_476
timestamp 1698431365
transform 1 0 54656 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_484
timestamp 1698431365
transform 1 0 55552 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_488
timestamp 1698431365
transform 1 0 56000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1698431365
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_10
timestamp 1698431365
transform 1 0 2464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_14
timestamp 1698431365
transform 1 0 2912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_22
timestamp 1698431365
transform 1 0 3808 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_30
timestamp 1698431365
transform 1 0 4704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_58
timestamp 1698431365
transform 1 0 7840 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_74
timestamp 1698431365
transform 1 0 9632 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_78
timestamp 1698431365
transform 1 0 10080 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_85
timestamp 1698431365
transform 1 0 10864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_87
timestamp 1698431365
transform 1 0 11088 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_103
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_126
timestamp 1698431365
transform 1 0 15456 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_139
timestamp 1698431365
transform 1 0 16912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_143
timestamp 1698431365
transform 1 0 17360 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_155
timestamp 1698431365
transform 1 0 18704 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_161
timestamp 1698431365
transform 1 0 19376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698431365
transform 1 0 25312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_220
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_222
timestamp 1698431365
transform 1 0 26208 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_238
timestamp 1698431365
transform 1 0 28000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_240
timestamp 1698431365
transform 1 0 28224 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_262
timestamp 1698431365
transform 1 0 30688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_264
timestamp 1698431365
transform 1 0 30912 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_300
timestamp 1698431365
transform 1 0 34944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_332
timestamp 1698431365
transform 1 0 38528 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_366
timestamp 1698431365
transform 1 0 42336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_380
timestamp 1698431365
transform 1 0 43904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_382
timestamp 1698431365
transform 1 0 44128 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_401
timestamp 1698431365
transform 1 0 46256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_429
timestamp 1698431365
transform 1 0 49392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_433
timestamp 1698431365
transform 1 0 49840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_437
timestamp 1698431365
transform 1 0 50288 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_440
timestamp 1698431365
transform 1 0 50624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_454
timestamp 1698431365
transform 1 0 52192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_461
timestamp 1698431365
transform 1 0 52976 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_493
timestamp 1698431365
transform 1 0 56560 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_32
timestamp 1698431365
transform 1 0 4928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_49
timestamp 1698431365
transform 1 0 6832 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_64
timestamp 1698431365
transform 1 0 8512 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_101
timestamp 1698431365
transform 1 0 12656 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_127
timestamp 1698431365
transform 1 0 15568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_131
timestamp 1698431365
transform 1 0 16016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_148
timestamp 1698431365
transform 1 0 17920 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_168
timestamp 1698431365
transform 1 0 20160 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_241
timestamp 1698431365
transform 1 0 28336 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_271
timestamp 1698431365
transform 1 0 31696 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_286
timestamp 1698431365
transform 1 0 33376 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_335
timestamp 1698431365
transform 1 0 38864 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_403
timestamp 1698431365
transform 1 0 46480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_407
timestamp 1698431365
transform 1 0 46928 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_469
timestamp 1698431365
transform 1 0 53872 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_485
timestamp 1698431365
transform 1 0 55664 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_489
timestamp 1698431365
transform 1 0 56112 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_49
timestamp 1698431365
transform 1 0 6832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_51
timestamp 1698431365
transform 1 0 7056 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_61
timestamp 1698431365
transform 1 0 8176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_65
timestamp 1698431365
transform 1 0 8624 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_69
timestamp 1698431365
transform 1 0 9072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_71
timestamp 1698431365
transform 1 0 9296 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_76
timestamp 1698431365
transform 1 0 9856 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_92
timestamp 1698431365
transform 1 0 11648 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_96
timestamp 1698431365
transform 1 0 12096 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_136
timestamp 1698431365
transform 1 0 16576 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_140
timestamp 1698431365
transform 1 0 17024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_142
timestamp 1698431365
transform 1 0 17248 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_225
timestamp 1698431365
transform 1 0 26544 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_233
timestamp 1698431365
transform 1 0 27440 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_239
timestamp 1698431365
transform 1 0 28112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_253
timestamp 1698431365
transform 1 0 29680 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_269
timestamp 1698431365
transform 1 0 31472 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_277
timestamp 1698431365
transform 1 0 32368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_281
timestamp 1698431365
transform 1 0 32816 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_383
timestamp 1698431365
transform 1 0 44240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_415
timestamp 1698431365
transform 1 0 47824 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_439
timestamp 1698431365
transform 1 0 50512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_452
timestamp 1698431365
transform 1 0 51968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_454
timestamp 1698431365
transform 1 0 52192 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_471
timestamp 1698431365
transform 1 0 54096 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_475
timestamp 1698431365
transform 1 0 54544 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_507
timestamp 1698431365
transform 1 0 58128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_10
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_23
timestamp 1698431365
transform 1 0 3920 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_39
timestamp 1698431365
transform 1 0 5712 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_84
timestamp 1698431365
transform 1 0 10752 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_88
timestamp 1698431365
transform 1 0 11200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_90
timestamp 1698431365
transform 1 0 11424 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_97
timestamp 1698431365
transform 1 0 12208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_101
timestamp 1698431365
transform 1 0 12656 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_107
timestamp 1698431365
transform 1 0 13328 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_115
timestamp 1698431365
transform 1 0 14224 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_119
timestamp 1698431365
transform 1 0 14672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_123
timestamp 1698431365
transform 1 0 15120 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_176
timestamp 1698431365
transform 1 0 21056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_204
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_259
timestamp 1698431365
transform 1 0 30352 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_275
timestamp 1698431365
transform 1 0 32144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_343
timestamp 1698431365
transform 1 0 39760 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_400
timestamp 1698431365
transform 1 0 46144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_402
timestamp 1698431365
transform 1 0 46368 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_419
timestamp 1698431365
transform 1 0 48272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_465
timestamp 1698431365
transform 1 0 53424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_469
timestamp 1698431365
transform 1 0 53872 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_473
timestamp 1698431365
transform 1 0 54320 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_489
timestamp 1698431365
transform 1 0 56112 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698431365
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_41
timestamp 1698431365
transform 1 0 5936 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_100
timestamp 1698431365
transform 1 0 12544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_122
timestamp 1698431365
transform 1 0 15008 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_162
timestamp 1698431365
transform 1 0 19488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_166
timestamp 1698431365
transform 1 0 19936 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_212
timestamp 1698431365
transform 1 0 25088 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_228
timestamp 1698431365
transform 1 0 26880 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_232
timestamp 1698431365
transform 1 0 27328 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_251
timestamp 1698431365
transform 1 0 29456 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_380
timestamp 1698431365
transform 1 0 43904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_428
timestamp 1698431365
transform 1 0 49280 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_470
timestamp 1698431365
transform 1 0 53984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_474
timestamp 1698431365
transform 1 0 54432 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_478
timestamp 1698431365
transform 1 0 54880 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_494
timestamp 1698431365
transform 1 0 56672 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_502
timestamp 1698431365
transform 1 0 57568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_506
timestamp 1698431365
transform 1 0 58016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_508
timestamp 1698431365
transform 1 0 58240 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_18
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_22
timestamp 1698431365
transform 1 0 3808 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_52
timestamp 1698431365
transform 1 0 7168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_56
timestamp 1698431365
transform 1 0 7616 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_64
timestamp 1698431365
transform 1 0 8512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_130
timestamp 1698431365
transform 1 0 15904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_134
timestamp 1698431365
transform 1 0 16352 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_144
timestamp 1698431365
transform 1 0 17472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_173
timestamp 1698431365
transform 1 0 20720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698431365
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_218
timestamp 1698431365
transform 1 0 25760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_226
timestamp 1698431365
transform 1 0 26656 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_242
timestamp 1698431365
transform 1 0 28448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_254
timestamp 1698431365
transform 1 0 29792 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_270
timestamp 1698431365
transform 1 0 31584 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_304
timestamp 1698431365
transform 1 0 35392 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_340
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_416
timestamp 1698431365
transform 1 0 47936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_450
timestamp 1698431365
transform 1 0 51744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_452
timestamp 1698431365
transform 1 0 51968 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_482
timestamp 1698431365
transform 1 0 55328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698431365
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_508
timestamp 1698431365
transform 1 0 58240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_18
timestamp 1698431365
transform 1 0 3360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_43
timestamp 1698431365
transform 1 0 6160 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_48
timestamp 1698431365
transform 1 0 6720 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_85
timestamp 1698431365
transform 1 0 10864 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_113
timestamp 1698431365
transform 1 0 14000 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_121
timestamp 1698431365
transform 1 0 14896 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698431365
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_193
timestamp 1698431365
transform 1 0 22960 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_195
timestamp 1698431365
transform 1 0 23184 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_227
timestamp 1698431365
transform 1 0 26768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_231
timestamp 1698431365
transform 1 0 27216 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698431365
transform 1 0 28112 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_251
timestamp 1698431365
transform 1 0 29456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_271
timestamp 1698431365
transform 1 0 31696 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_279
timestamp 1698431365
transform 1 0 32592 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_299
timestamp 1698431365
transform 1 0 34832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_303
timestamp 1698431365
transform 1 0 35280 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_313
timestamp 1698431365
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_328
timestamp 1698431365
transform 1 0 38080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_332
timestamp 1698431365
transform 1 0 38528 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_362
timestamp 1698431365
transform 1 0 41888 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_467
timestamp 1698431365
transform 1 0 53648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_469
timestamp 1698431365
transform 1 0 53872 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_499
timestamp 1698431365
transform 1 0 57232 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_507
timestamp 1698431365
transform 1 0 58128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_10
timestamp 1698431365
transform 1 0 2464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_14
timestamp 1698431365
transform 1 0 2912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_16
timestamp 1698431365
transform 1 0 3136 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_65
timestamp 1698431365
transform 1 0 8624 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_95
timestamp 1698431365
transform 1 0 11984 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_127
timestamp 1698431365
transform 1 0 15568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_135
timestamp 1698431365
transform 1 0 16464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_168
timestamp 1698431365
transform 1 0 20160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_195
timestamp 1698431365
transform 1 0 23184 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_199
timestamp 1698431365
transform 1 0 23632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_201
timestamp 1698431365
transform 1 0 23856 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_248
timestamp 1698431365
transform 1 0 29120 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_302
timestamp 1698431365
transform 1 0 35168 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_356
timestamp 1698431365
transform 1 0 41216 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_368
timestamp 1698431365
transform 1 0 42560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_399
timestamp 1698431365
transform 1 0 46032 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_418
timestamp 1698431365
transform 1 0 48160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_456
timestamp 1698431365
transform 1 0 52416 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_466
timestamp 1698431365
transform 1 0 53536 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_488
timestamp 1698431365
transform 1 0 56000 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_496
timestamp 1698431365
transform 1 0 56896 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_504
timestamp 1698431365
transform 1 0 57792 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_49
timestamp 1698431365
transform 1 0 6832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_65
timestamp 1698431365
transform 1 0 8624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_67
timestamp 1698431365
transform 1 0 8848 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_97
timestamp 1698431365
transform 1 0 12208 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_123
timestamp 1698431365
transform 1 0 15120 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_127
timestamp 1698431365
transform 1 0 15568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_160
timestamp 1698431365
transform 1 0 19264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_164
timestamp 1698431365
transform 1 0 19712 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_189
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_193
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_206
timestamp 1698431365
transform 1 0 24416 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_232
timestamp 1698431365
transform 1 0 27328 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_276
timestamp 1698431365
transform 1 0 32256 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_292
timestamp 1698431365
transform 1 0 34048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_294
timestamp 1698431365
transform 1 0 34272 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_305
timestamp 1698431365
transform 1 0 35504 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_309
timestamp 1698431365
transform 1 0 35952 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_313
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_335
timestamp 1698431365
transform 1 0 38864 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_339
timestamp 1698431365
transform 1 0 39312 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_341
timestamp 1698431365
transform 1 0 39536 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_356
timestamp 1698431365
transform 1 0 41216 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_364
timestamp 1698431365
transform 1 0 42112 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_366
timestamp 1698431365
transform 1 0 42336 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_373
timestamp 1698431365
transform 1 0 43120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_377
timestamp 1698431365
transform 1 0 43568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_379
timestamp 1698431365
transform 1 0 43792 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_382
timestamp 1698431365
transform 1 0 44128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_435
timestamp 1698431365
transform 1 0 50064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_439
timestamp 1698431365
transform 1 0 50512 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_441
timestamp 1698431365
transform 1 0 50736 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_502
timestamp 1698431365
transform 1 0 57568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_506
timestamp 1698431365
transform 1 0 58016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_508
timestamp 1698431365
transform 1 0 58240 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_18
timestamp 1698431365
transform 1 0 3360 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_26
timestamp 1698431365
transform 1 0 4256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_30
timestamp 1698431365
transform 1 0 4704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_32
timestamp 1698431365
transform 1 0 4928 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_62
timestamp 1698431365
transform 1 0 8288 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_76
timestamp 1698431365
transform 1 0 9856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_93
timestamp 1698431365
transform 1 0 11760 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_101
timestamp 1698431365
transform 1 0 12656 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_131
timestamp 1698431365
transform 1 0 16016 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_135
timestamp 1698431365
transform 1 0 16464 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_146
timestamp 1698431365
transform 1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_148
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_153
timestamp 1698431365
transform 1 0 18480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_155
timestamp 1698431365
transform 1 0 18704 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_164
timestamp 1698431365
transform 1 0 19712 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_172
timestamp 1698431365
transform 1 0 20608 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_205
timestamp 1698431365
transform 1 0 24304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_228
timestamp 1698431365
transform 1 0 26880 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_236
timestamp 1698431365
transform 1 0 27776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_240
timestamp 1698431365
transform 1 0 28224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_242
timestamp 1698431365
transform 1 0 28448 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_265
timestamp 1698431365
transform 1 0 31024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_269
timestamp 1698431365
transform 1 0 31472 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_271
timestamp 1698431365
transform 1 0 31696 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_306
timestamp 1698431365
transform 1 0 35616 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_338
timestamp 1698431365
transform 1 0 39200 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_358
timestamp 1698431365
transform 1 0 41440 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_374
timestamp 1698431365
transform 1 0 43232 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_380
timestamp 1698431365
transform 1 0 43904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_384
timestamp 1698431365
transform 1 0 44352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_409
timestamp 1698431365
transform 1 0 47152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698431365
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_445
timestamp 1698431365
transform 1 0 51184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_447
timestamp 1698431365
transform 1 0 51408 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_477
timestamp 1698431365
transform 1 0 54768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_481
timestamp 1698431365
transform 1 0 55216 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_489
timestamp 1698431365
transform 1 0 56112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_508
timestamp 1698431365
transform 1 0 58240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_69
timestamp 1698431365
transform 1 0 9072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_71
timestamp 1698431365
transform 1 0 9296 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_78
timestamp 1698431365
transform 1 0 10080 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_94
timestamp 1698431365
transform 1 0 11872 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_102
timestamp 1698431365
transform 1 0 12768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_136
timestamp 1698431365
transform 1 0 16576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_140
timestamp 1698431365
transform 1 0 17024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_142
timestamp 1698431365
transform 1 0 17248 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_156
timestamp 1698431365
transform 1 0 18816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_162
timestamp 1698431365
transform 1 0 19488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_166
timestamp 1698431365
transform 1 0 19936 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_168
timestamp 1698431365
transform 1 0 20160 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_183
timestamp 1698431365
transform 1 0 21840 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_235
timestamp 1698431365
transform 1 0 27664 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_249
timestamp 1698431365
transform 1 0 29232 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_312
timestamp 1698431365
transform 1 0 36288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_323
timestamp 1698431365
transform 1 0 37520 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_325
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_378
timestamp 1698431365
transform 1 0 43680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_382
timestamp 1698431365
transform 1 0 44128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_471
timestamp 1698431365
transform 1 0 54096 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_503
timestamp 1698431365
transform 1 0 57680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_507
timestamp 1698431365
transform 1 0 58128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_101
timestamp 1698431365
transform 1 0 12656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_117
timestamp 1698431365
transform 1 0 14448 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_125
timestamp 1698431365
transform 1 0 15344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_127
timestamp 1698431365
transform 1 0 15568 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_146
timestamp 1698431365
transform 1 0 17696 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_148
timestamp 1698431365
transform 1 0 17920 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_244
timestamp 1698431365
transform 1 0 28672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_246
timestamp 1698431365
transform 1 0 28896 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_286
timestamp 1698431365
transform 1 0 33376 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_345
timestamp 1698431365
transform 1 0 39984 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_360
timestamp 1698431365
transform 1 0 41664 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_369
timestamp 1698431365
transform 1 0 42672 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_390
timestamp 1698431365
transform 1 0 45024 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1698431365
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_430
timestamp 1698431365
transform 1 0 49504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_472
timestamp 1698431365
transform 1 0 54208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_476
timestamp 1698431365
transform 1 0 54656 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_484
timestamp 1698431365
transform 1 0 55552 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_488
timestamp 1698431365
transform 1 0 56000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_508
timestamp 1698431365
transform 1 0 58240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_113
timestamp 1698431365
transform 1 0 14000 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_117
timestamp 1698431365
transform 1 0 14448 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_121
timestamp 1698431365
transform 1 0 14896 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_123
timestamp 1698431365
transform 1 0 15120 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_220
timestamp 1698431365
transform 1 0 25984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_238
timestamp 1698431365
transform 1 0 28000 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_242
timestamp 1698431365
transform 1 0 28448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_251
timestamp 1698431365
transform 1 0 29456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_253
timestamp 1698431365
transform 1 0 29680 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_260
timestamp 1698431365
transform 1 0 30464 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_276
timestamp 1698431365
transform 1 0 32256 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_284
timestamp 1698431365
transform 1 0 33152 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_286
timestamp 1698431365
transform 1 0 33376 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_300
timestamp 1698431365
transform 1 0 34944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_304
timestamp 1698431365
transform 1 0 35392 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_308
timestamp 1698431365
transform 1 0 35840 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_328
timestamp 1698431365
transform 1 0 38080 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_332
timestamp 1698431365
transform 1 0 38528 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_337
timestamp 1698431365
transform 1 0 39088 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_345
timestamp 1698431365
transform 1 0 39984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_353
timestamp 1698431365
transform 1 0 40880 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_391
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_395
timestamp 1698431365
transform 1 0 45584 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_404
timestamp 1698431365
transform 1 0 46592 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_411
timestamp 1698431365
transform 1 0 47376 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_421
timestamp 1698431365
transform 1 0 48496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_444
timestamp 1698431365
transform 1 0 51072 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_465
timestamp 1698431365
transform 1 0 53424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_467
timestamp 1698431365
transform 1 0 53648 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_497
timestamp 1698431365
transform 1 0 57008 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_505
timestamp 1698431365
transform 1 0 57904 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_125
timestamp 1698431365
transform 1 0 15344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_129
timestamp 1698431365
transform 1 0 15792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_194
timestamp 1698431365
transform 1 0 23072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_208
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_214
timestamp 1698431365
transform 1 0 25312 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_254
timestamp 1698431365
transform 1 0 29792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_258
timestamp 1698431365
transform 1 0 30240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_265
timestamp 1698431365
transform 1 0 31024 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_273
timestamp 1698431365
transform 1 0 31920 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_290
timestamp 1698431365
transform 1 0 33824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_306
timestamp 1698431365
transform 1 0 35616 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_314
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_316
timestamp 1698431365
transform 1 0 36736 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_335
timestamp 1698431365
transform 1 0 38864 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_343
timestamp 1698431365
transform 1 0 39760 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_347
timestamp 1698431365
transform 1 0 40208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698431365
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_364
timestamp 1698431365
transform 1 0 42112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_368
timestamp 1698431365
transform 1 0 42560 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_379
timestamp 1698431365
transform 1 0 43792 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_404
timestamp 1698431365
transform 1 0 46592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_406
timestamp 1698431365
transform 1 0 46816 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_415
timestamp 1698431365
transform 1 0 47824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_417
timestamp 1698431365
transform 1 0 48048 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_444
timestamp 1698431365
transform 1 0 51072 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_489
timestamp 1698431365
transform 1 0 56112 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_496
timestamp 1698431365
transform 1 0 56896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_500
timestamp 1698431365
transform 1 0 57344 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_508
timestamp 1698431365
transform 1 0 58240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_136
timestamp 1698431365
transform 1 0 16576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_144
timestamp 1698431365
transform 1 0 17472 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_153
timestamp 1698431365
transform 1 0 18480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_159
timestamp 1698431365
transform 1 0 19152 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_165
timestamp 1698431365
transform 1 0 19824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_167
timestamp 1698431365
transform 1 0 20048 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_170
timestamp 1698431365
transform 1 0 20384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_189
timestamp 1698431365
transform 1 0 22512 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_238
timestamp 1698431365
transform 1 0 28000 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_242
timestamp 1698431365
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_292
timestamp 1698431365
transform 1 0 34048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_296
timestamp 1698431365
transform 1 0 34496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_298
timestamp 1698431365
transform 1 0 34720 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_308
timestamp 1698431365
transform 1 0 35840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_310
timestamp 1698431365
transform 1 0 36064 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_350
timestamp 1698431365
transform 1 0 40544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_370
timestamp 1698431365
transform 1 0 42784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_372
timestamp 1698431365
transform 1 0 43008 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_395
timestamp 1698431365
transform 1 0 45584 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_407
timestamp 1698431365
transform 1 0 46928 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_423
timestamp 1698431365
transform 1 0 48720 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_430
timestamp 1698431365
transform 1 0 49504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_432
timestamp 1698431365
transform 1 0 49728 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_439
timestamp 1698431365
transform 1 0 50512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_445
timestamp 1698431365
transform 1 0 51184 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_479
timestamp 1698431365
transform 1 0 54992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_104
timestamp 1698431365
transform 1 0 12992 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_108
timestamp 1698431365
transform 1 0 13440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_110
timestamp 1698431365
transform 1 0 13664 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_117
timestamp 1698431365
transform 1 0 14448 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_121
timestamp 1698431365
transform 1 0 14896 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_125
timestamp 1698431365
transform 1 0 15344 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_128
timestamp 1698431365
transform 1 0 15680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_132
timestamp 1698431365
transform 1 0 16128 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_150
timestamp 1698431365
transform 1 0 18144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_158
timestamp 1698431365
transform 1 0 19040 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_188
timestamp 1698431365
transform 1 0 22400 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_192
timestamp 1698431365
transform 1 0 22848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_200
timestamp 1698431365
transform 1 0 23744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_216
timestamp 1698431365
transform 1 0 25536 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_232
timestamp 1698431365
transform 1 0 27328 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_235
timestamp 1698431365
transform 1 0 27664 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_239
timestamp 1698431365
transform 1 0 28112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_241
timestamp 1698431365
transform 1 0 28336 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_271
timestamp 1698431365
transform 1 0 31696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_275
timestamp 1698431365
transform 1 0 32144 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_311
timestamp 1698431365
transform 1 0 36176 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_345
timestamp 1698431365
transform 1 0 39984 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_360
timestamp 1698431365
transform 1 0 41664 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_364
timestamp 1698431365
transform 1 0 42112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_366
timestamp 1698431365
transform 1 0 42336 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_396
timestamp 1698431365
transform 1 0 45696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_400
timestamp 1698431365
transform 1 0 46144 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_424
timestamp 1698431365
transform 1 0 48832 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_474
timestamp 1698431365
transform 1 0 54432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_504
timestamp 1698431365
transform 1 0 57792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_508
timestamp 1698431365
transform 1 0 58240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_113
timestamp 1698431365
transform 1 0 14000 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_160
timestamp 1698431365
transform 1 0 19264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_170
timestamp 1698431365
transform 1 0 20384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_172
timestamp 1698431365
transform 1 0 20608 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_192
timestamp 1698431365
transform 1 0 22848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_200
timestamp 1698431365
transform 1 0 23744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_204
timestamp 1698431365
transform 1 0 24192 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_212
timestamp 1698431365
transform 1 0 25088 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_216
timestamp 1698431365
transform 1 0 25536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_218
timestamp 1698431365
transform 1 0 25760 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_261
timestamp 1698431365
transform 1 0 30576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_263
timestamp 1698431365
transform 1 0 30800 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_270
timestamp 1698431365
transform 1 0 31584 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_286
timestamp 1698431365
transform 1 0 33376 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_305
timestamp 1698431365
transform 1 0 35504 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_313
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_334
timestamp 1698431365
transform 1 0 38752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_336
timestamp 1698431365
transform 1 0 38976 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_366
timestamp 1698431365
transform 1 0 42336 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_373
timestamp 1698431365
transform 1 0 43120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_402
timestamp 1698431365
transform 1 0 46368 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_406
timestamp 1698431365
transform 1 0 46816 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_410
timestamp 1698431365
transform 1 0 47264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_412
timestamp 1698431365
transform 1 0 47488 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_88
timestamp 1698431365
transform 1 0 11200 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_92
timestamp 1698431365
transform 1 0 11648 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_122
timestamp 1698431365
transform 1 0 15008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_124
timestamp 1698431365
transform 1 0 15232 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_190
timestamp 1698431365
transform 1 0 22624 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_226
timestamp 1698431365
transform 1 0 26656 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_230
timestamp 1698431365
transform 1 0 27104 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_233
timestamp 1698431365
transform 1 0 27440 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_249
timestamp 1698431365
transform 1 0 29232 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_253
timestamp 1698431365
transform 1 0 29680 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_262
timestamp 1698431365
transform 1 0 30688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_272
timestamp 1698431365
transform 1 0 31808 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_290
timestamp 1698431365
transform 1 0 33824 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_306
timestamp 1698431365
transform 1 0 35616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_310
timestamp 1698431365
transform 1 0 36064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_312
timestamp 1698431365
transform 1 0 36288 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_344
timestamp 1698431365
transform 1 0 39872 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_348
timestamp 1698431365
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_368
timestamp 1698431365
transform 1 0 42560 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_372
timestamp 1698431365
transform 1 0 43008 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_375
timestamp 1698431365
transform 1 0 43344 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_411
timestamp 1698431365
transform 1 0 47376 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_488
timestamp 1698431365
transform 1 0 56000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_498
timestamp 1698431365
transform 1 0 57120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_502
timestamp 1698431365
transform 1 0 57568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_506
timestamp 1698431365
transform 1 0 58016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_115
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_149
timestamp 1698431365
transform 1 0 18032 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_183
timestamp 1698431365
transform 1 0 21840 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_231
timestamp 1698431365
transform 1 0 27216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_235
timestamp 1698431365
transform 1 0 27664 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_239
timestamp 1698431365
transform 1 0 28112 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_255
timestamp 1698431365
transform 1 0 29904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_277
timestamp 1698431365
transform 1 0 32368 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_281
timestamp 1698431365
transform 1 0 32816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_283
timestamp 1698431365
transform 1 0 33040 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_292
timestamp 1698431365
transform 1 0 34048 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_300
timestamp 1698431365
transform 1 0 34944 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_304
timestamp 1698431365
transform 1 0 35392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_306
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_338
timestamp 1698431365
transform 1 0 39200 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_340
timestamp 1698431365
transform 1 0 39424 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_370
timestamp 1698431365
transform 1 0 42784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_374
timestamp 1698431365
transform 1 0 43232 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_382
timestamp 1698431365
transform 1 0 44128 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_405
timestamp 1698431365
transform 1 0 46704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_433
timestamp 1698431365
transform 1 0 49840 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_454
timestamp 1698431365
transform 1 0 52192 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_467
timestamp 1698431365
transform 1 0 53648 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_471
timestamp 1698431365
transform 1 0 54096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_495
timestamp 1698431365
transform 1 0 56784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_499
timestamp 1698431365
transform 1 0 57232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_503
timestamp 1698431365
transform 1 0 57680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_507
timestamp 1698431365
transform 1 0 58128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_18
timestamp 1698431365
transform 1 0 3360 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_22
timestamp 1698431365
transform 1 0 3808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_24
timestamp 1698431365
transform 1 0 4032 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_33
timestamp 1698431365
transform 1 0 5040 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_65
timestamp 1698431365
transform 1 0 8624 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_69
timestamp 1698431365
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_101
timestamp 1698431365
transform 1 0 12656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_105
timestamp 1698431365
transform 1 0 13104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_109
timestamp 1698431365
transform 1 0 13552 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_113
timestamp 1698431365
transform 1 0 14000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_115
timestamp 1698431365
transform 1 0 14224 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_156
timestamp 1698431365
transform 1 0 18816 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_187
timestamp 1698431365
transform 1 0 22288 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_189
timestamp 1698431365
transform 1 0 22512 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_220
timestamp 1698431365
transform 1 0 25984 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_261
timestamp 1698431365
transform 1 0 30576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_277
timestamp 1698431365
transform 1 0 32368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_338
timestamp 1698431365
transform 1 0 39200 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_356
timestamp 1698431365
transform 1 0 41216 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_364
timestamp 1698431365
transform 1 0 42112 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_368
timestamp 1698431365
transform 1 0 42560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_398
timestamp 1698431365
transform 1 0 45920 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_406
timestamp 1698431365
transform 1 0 46816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_410
timestamp 1698431365
transform 1 0 47264 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_488
timestamp 1698431365
transform 1 0 56000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1698431365
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_31
timestamp 1698431365
transform 1 0 4816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_70
timestamp 1698431365
transform 1 0 9184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_74
timestamp 1698431365
transform 1 0 9632 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_126
timestamp 1698431365
transform 1 0 15456 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_157
timestamp 1698431365
transform 1 0 18928 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_167
timestamp 1698431365
transform 1 0 20048 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_185
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_209
timestamp 1698431365
transform 1 0 24752 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_242
timestamp 1698431365
transform 1 0 28448 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_249
timestamp 1698431365
transform 1 0 29232 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_256
timestamp 1698431365
transform 1 0 30016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_272
timestamp 1698431365
transform 1 0 31808 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_280
timestamp 1698431365
transform 1 0 32704 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_284
timestamp 1698431365
transform 1 0 33152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_286
timestamp 1698431365
transform 1 0 33376 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_301
timestamp 1698431365
transform 1 0 35056 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_309
timestamp 1698431365
transform 1 0 35952 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698431365
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_380
timestamp 1698431365
transform 1 0 43904 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_398
timestamp 1698431365
transform 1 0 45920 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_402
timestamp 1698431365
transform 1 0 46368 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_406
timestamp 1698431365
transform 1 0 46816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_410
timestamp 1698431365
transform 1 0 47264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_453
timestamp 1698431365
transform 1 0 52080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_465
timestamp 1698431365
transform 1 0 53424 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_497
timestamp 1698431365
transform 1 0 57008 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_505
timestamp 1698431365
transform 1 0 57904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_10
timestamp 1698431365
transform 1 0 2464 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_59
timestamp 1698431365
transform 1 0 7952 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_67
timestamp 1698431365
transform 1 0 8848 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_88
timestamp 1698431365
transform 1 0 11200 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_108
timestamp 1698431365
transform 1 0 13440 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_116
timestamp 1698431365
transform 1 0 14336 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_118
timestamp 1698431365
transform 1 0 14560 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_196
timestamp 1698431365
transform 1 0 23296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_204
timestamp 1698431365
transform 1 0 24192 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_208
timestamp 1698431365
transform 1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_218
timestamp 1698431365
transform 1 0 25760 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_224
timestamp 1698431365
transform 1 0 26432 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_238
timestamp 1698431365
transform 1 0 28000 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_246
timestamp 1698431365
transform 1 0 28896 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_250
timestamp 1698431365
transform 1 0 29344 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_266
timestamp 1698431365
transform 1 0 31136 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_287
timestamp 1698431365
transform 1 0 33488 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_303
timestamp 1698431365
transform 1 0 35280 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_311
timestamp 1698431365
transform 1 0 36176 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_315
timestamp 1698431365
transform 1 0 36624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_323
timestamp 1698431365
transform 1 0 37520 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_334
timestamp 1698431365
transform 1 0 38752 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_360
timestamp 1698431365
transform 1 0 41664 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_374
timestamp 1698431365
transform 1 0 43232 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_376
timestamp 1698431365
transform 1 0 43456 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_388
timestamp 1698431365
transform 1 0 44800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_390
timestamp 1698431365
transform 1 0 45024 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_399
timestamp 1698431365
transform 1 0 46032 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_440
timestamp 1698431365
transform 1 0 50624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_442
timestamp 1698431365
transform 1 0 50848 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_472
timestamp 1698431365
transform 1 0 54208 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_488
timestamp 1698431365
transform 1 0 56000 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_508
timestamp 1698431365
transform 1 0 58240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_31
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_44
timestamp 1698431365
transform 1 0 6272 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_57
timestamp 1698431365
transform 1 0 7728 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_61
timestamp 1698431365
transform 1 0 8176 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_93
timestamp 1698431365
transform 1 0 11760 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_113
timestamp 1698431365
transform 1 0 14000 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_128
timestamp 1698431365
transform 1 0 15680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_134
timestamp 1698431365
transform 1 0 16352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_145
timestamp 1698431365
transform 1 0 17584 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_151
timestamp 1698431365
transform 1 0 18256 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_169
timestamp 1698431365
transform 1 0 20272 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_191
timestamp 1698431365
transform 1 0 22736 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_195
timestamp 1698431365
transform 1 0 23184 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_198
timestamp 1698431365
transform 1 0 23520 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_206
timestamp 1698431365
transform 1 0 24416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_210
timestamp 1698431365
transform 1 0 24864 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_217
timestamp 1698431365
transform 1 0 25648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_221
timestamp 1698431365
transform 1 0 26096 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_231
timestamp 1698431365
transform 1 0 27216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_263
timestamp 1698431365
transform 1 0 30800 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_296
timestamp 1698431365
transform 1 0 34496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_300
timestamp 1698431365
transform 1 0 34944 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_308
timestamp 1698431365
transform 1 0 35840 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_312
timestamp 1698431365
transform 1 0 36288 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_346
timestamp 1698431365
transform 1 0 40096 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_350
timestamp 1698431365
transform 1 0 40544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_352
timestamp 1698431365
transform 1 0 40768 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_378
timestamp 1698431365
transform 1 0 43680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_409
timestamp 1698431365
transform 1 0 47152 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_413
timestamp 1698431365
transform 1 0 47600 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_427
timestamp 1698431365
transform 1 0 49168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_454
timestamp 1698431365
transform 1 0 52192 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_486
timestamp 1698431365
transform 1 0 55776 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_502
timestamp 1698431365
transform 1 0 57568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_506
timestamp 1698431365
transform 1 0 58016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_508
timestamp 1698431365
transform 1 0 58240 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_18
timestamp 1698431365
transform 1 0 3360 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_34
timestamp 1698431365
transform 1 0 5152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_65
timestamp 1698431365
transform 1 0 8624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_69
timestamp 1698431365
transform 1 0 9072 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_88
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_103
timestamp 1698431365
transform 1 0 12880 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_116
timestamp 1698431365
transform 1 0 14336 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_134
timestamp 1698431365
transform 1 0 16352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_138
timestamp 1698431365
transform 1 0 16800 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_146
timestamp 1698431365
transform 1 0 17696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_150
timestamp 1698431365
transform 1 0 18144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_154
timestamp 1698431365
transform 1 0 18592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_158
timestamp 1698431365
transform 1 0 19040 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_169
timestamp 1698431365
transform 1 0 20272 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_173
timestamp 1698431365
transform 1 0 20720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_192
timestamp 1698431365
transform 1 0 22848 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_200
timestamp 1698431365
transform 1 0 23744 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_207
timestamp 1698431365
transform 1 0 24528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_229
timestamp 1698431365
transform 1 0 26992 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_251
timestamp 1698431365
transform 1 0 29456 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_259
timestamp 1698431365
transform 1 0 30352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_261
timestamp 1698431365
transform 1 0 30576 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_290
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_294
timestamp 1698431365
transform 1 0 34272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_327
timestamp 1698431365
transform 1 0 37968 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_343
timestamp 1698431365
transform 1 0 39760 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_411
timestamp 1698431365
transform 1 0 47376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_415
timestamp 1698431365
transform 1 0 47824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_419
timestamp 1698431365
transform 1 0 48272 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_432
timestamp 1698431365
transform 1 0 49728 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_436
timestamp 1698431365
transform 1 0 50176 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_458
timestamp 1698431365
transform 1 0 52640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_462
timestamp 1698431365
transform 1 0 53088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_466
timestamp 1698431365
transform 1 0 53536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_470
timestamp 1698431365
transform 1 0 53984 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698431365
transform 1 0 55776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_10
timestamp 1698431365
transform 1 0 2464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_12
timestamp 1698431365
transform 1 0 2688 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_27
timestamp 1698431365
transform 1 0 4368 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_39
timestamp 1698431365
transform 1 0 5712 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_54
timestamp 1698431365
transform 1 0 7392 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_89
timestamp 1698431365
transform 1 0 11312 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_109
timestamp 1698431365
transform 1 0 13552 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_126
timestamp 1698431365
transform 1 0 15456 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_181
timestamp 1698431365
transform 1 0 21616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_210
timestamp 1698431365
transform 1 0 24864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_235
timestamp 1698431365
transform 1 0 27664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_263
timestamp 1698431365
transform 1 0 30800 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_271
timestamp 1698431365
transform 1 0 31696 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_329
timestamp 1698431365
transform 1 0 38192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_336
timestamp 1698431365
transform 1 0 38976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_346
timestamp 1698431365
transform 1 0 40096 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_354
timestamp 1698431365
transform 1 0 40992 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_356
timestamp 1698431365
transform 1 0 41216 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_389
timestamp 1698431365
transform 1 0 44912 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_419
timestamp 1698431365
transform 1 0 48272 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_423
timestamp 1698431365
transform 1 0 48720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_427
timestamp 1698431365
transform 1 0 49168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_454
timestamp 1698431365
transform 1 0 52192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_462
timestamp 1698431365
transform 1 0 53088 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_466
timestamp 1698431365
transform 1 0 53536 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_498
timestamp 1698431365
transform 1 0 57120 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_506
timestamp 1698431365
transform 1 0 58016 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_508
timestamp 1698431365
transform 1 0 58240 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_65
timestamp 1698431365
transform 1 0 8624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_69
timestamp 1698431365
transform 1 0 9072 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_76
timestamp 1698431365
transform 1 0 9856 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_84
timestamp 1698431365
transform 1 0 10752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_93
timestamp 1698431365
transform 1 0 11760 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_110
timestamp 1698431365
transform 1 0 13664 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_112
timestamp 1698431365
transform 1 0 13888 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_121
timestamp 1698431365
transform 1 0 14896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_123
timestamp 1698431365
transform 1 0 15120 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_159
timestamp 1698431365
transform 1 0 19152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_176
timestamp 1698431365
transform 1 0 21056 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_195
timestamp 1698431365
transform 1 0 23184 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_199
timestamp 1698431365
transform 1 0 23632 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_208
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_231
timestamp 1698431365
transform 1 0 27216 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_233
timestamp 1698431365
transform 1 0 27440 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_243
timestamp 1698431365
transform 1 0 28560 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_257
timestamp 1698431365
transform 1 0 30128 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_261
timestamp 1698431365
transform 1 0 30576 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_278
timestamp 1698431365
transform 1 0 32480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_288
timestamp 1698431365
transform 1 0 33600 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_294
timestamp 1698431365
transform 1 0 34272 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_356
timestamp 1698431365
transform 1 0 41216 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_358
timestamp 1698431365
transform 1 0 41440 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_407
timestamp 1698431365
transform 1 0 46928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_411
timestamp 1698431365
transform 1 0 47376 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698431365
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_474
timestamp 1698431365
transform 1 0 54432 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_18
timestamp 1698431365
transform 1 0 3360 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_27
timestamp 1698431365
transform 1 0 4368 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_33
timestamp 1698431365
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_41
timestamp 1698431365
transform 1 0 5936 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_57
timestamp 1698431365
transform 1 0 7728 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_88
timestamp 1698431365
transform 1 0 11200 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_103
timestamp 1698431365
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_116
timestamp 1698431365
transform 1 0 14336 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_120
timestamp 1698431365
transform 1 0 14784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_124
timestamp 1698431365
transform 1 0 15232 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_130
timestamp 1698431365
transform 1 0 15904 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_141
timestamp 1698431365
transform 1 0 17136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_143
timestamp 1698431365
transform 1 0 17360 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_162
timestamp 1698431365
transform 1 0 19488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_170
timestamp 1698431365
transform 1 0 20384 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_185
timestamp 1698431365
transform 1 0 22064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_187
timestamp 1698431365
transform 1 0 22288 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_208
timestamp 1698431365
transform 1 0 24640 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_221
timestamp 1698431365
transform 1 0 26096 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_229
timestamp 1698431365
transform 1 0 26992 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_231
timestamp 1698431365
transform 1 0 27216 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_239
timestamp 1698431365
transform 1 0 28112 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_243
timestamp 1698431365
transform 1 0 28560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_255
timestamp 1698431365
transform 1 0 29904 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_257
timestamp 1698431365
transform 1 0 30128 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_263
timestamp 1698431365
transform 1 0 30800 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_271
timestamp 1698431365
transform 1 0 31696 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_275
timestamp 1698431365
transform 1 0 32144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_277
timestamp 1698431365
transform 1 0 32368 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_280
timestamp 1698431365
transform 1 0 32704 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_288
timestamp 1698431365
transform 1 0 33600 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_290
timestamp 1698431365
transform 1 0 33824 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_323
timestamp 1698431365
transform 1 0 37520 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_339
timestamp 1698431365
transform 1 0 39312 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_343
timestamp 1698431365
transform 1 0 39760 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_345
timestamp 1698431365
transform 1 0 39984 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_356
timestamp 1698431365
transform 1 0 41216 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_360
timestamp 1698431365
transform 1 0 41664 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_377
timestamp 1698431365
transform 1 0 43568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_397
timestamp 1698431365
transform 1 0 45808 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_401
timestamp 1698431365
transform 1 0 46256 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_409
timestamp 1698431365
transform 1 0 47152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_416
timestamp 1698431365
transform 1 0 47936 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_430
timestamp 1698431365
transform 1 0 49504 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_454
timestamp 1698431365
transform 1 0 52192 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_462
timestamp 1698431365
transform 1 0 53088 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_494
timestamp 1698431365
transform 1 0 56672 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_502
timestamp 1698431365
transform 1 0 57568 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_506
timestamp 1698431365
transform 1 0 58016 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_508
timestamp 1698431365
transform 1 0 58240 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_74
timestamp 1698431365
transform 1 0 9632 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_90
timestamp 1698431365
transform 1 0 11424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_118
timestamp 1698431365
transform 1 0 14560 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_125
timestamp 1698431365
transform 1 0 15344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_127
timestamp 1698431365
transform 1 0 15568 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_144
timestamp 1698431365
transform 1 0 17472 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_152
timestamp 1698431365
transform 1 0 18368 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_190
timestamp 1698431365
transform 1 0 22624 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_208
timestamp 1698431365
transform 1 0 24640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_244
timestamp 1698431365
transform 1 0 28672 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_248
timestamp 1698431365
transform 1 0 29120 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_274
timestamp 1698431365
transform 1 0 32032 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_278
timestamp 1698431365
transform 1 0 32480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_288
timestamp 1698431365
transform 1 0 33600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_294
timestamp 1698431365
transform 1 0 34272 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_327
timestamp 1698431365
transform 1 0 37968 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_331
timestamp 1698431365
transform 1 0 38416 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_333
timestamp 1698431365
transform 1 0 38640 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_367
timestamp 1698431365
transform 1 0 42448 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_383
timestamp 1698431365
transform 1 0 44240 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_405
timestamp 1698431365
transform 1 0 46704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_409
timestamp 1698431365
transform 1 0 47152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_413
timestamp 1698431365
transform 1 0 47600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_417
timestamp 1698431365
transform 1 0 48048 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_456
timestamp 1698431365
transform 1 0 52416 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_488
timestamp 1698431365
transform 1 0 56000 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_32
timestamp 1698431365
transform 1 0 4928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_58
timestamp 1698431365
transform 1 0 7840 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_88
timestamp 1698431365
transform 1 0 11200 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_92
timestamp 1698431365
transform 1 0 11648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_96
timestamp 1698431365
transform 1 0 12096 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_103
timestamp 1698431365
transform 1 0 12880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_129
timestamp 1698431365
transform 1 0 15792 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_213
timestamp 1698431365
transform 1 0 25200 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_239
timestamp 1698431365
transform 1 0 28112 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_274
timestamp 1698431365
transform 1 0 32032 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_281
timestamp 1698431365
transform 1 0 32816 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_292
timestamp 1698431365
transform 1 0 34048 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_300
timestamp 1698431365
transform 1 0 34944 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_308
timestamp 1698431365
transform 1 0 35840 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_312
timestamp 1698431365
transform 1 0 36288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_321
timestamp 1698431365
transform 1 0 37296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_325
timestamp 1698431365
transform 1 0 37744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_335
timestamp 1698431365
transform 1 0 38864 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_372
timestamp 1698431365
transform 1 0 43008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_380
timestamp 1698431365
transform 1 0 43904 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1698431365
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_416
timestamp 1698431365
transform 1 0 47936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_420
timestamp 1698431365
transform 1 0 48384 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_452
timestamp 1698431365
transform 1 0 51968 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_454
timestamp 1698431365
transform 1 0 52192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_489
timestamp 1698431365
transform 1 0 56112 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_505
timestamp 1698431365
transform 1 0 57904 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_76
timestamp 1698431365
transform 1 0 9856 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_91
timestamp 1698431365
transform 1 0 11536 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_100
timestamp 1698431365
transform 1 0 12544 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_108
timestamp 1698431365
transform 1 0 13440 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_110
timestamp 1698431365
transform 1 0 13664 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_122
timestamp 1698431365
transform 1 0 15008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_126
timestamp 1698431365
transform 1 0 15456 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_128
timestamp 1698431365
transform 1 0 15680 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_131
timestamp 1698431365
transform 1 0 16016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_133
timestamp 1698431365
transform 1 0 16240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_151
timestamp 1698431365
transform 1 0 18256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_208
timestamp 1698431365
transform 1 0 24640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_246
timestamp 1698431365
transform 1 0 28896 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_257
timestamp 1698431365
transform 1 0 30128 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_278
timestamp 1698431365
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_323
timestamp 1698431365
transform 1 0 37520 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_325
timestamp 1698431365
transform 1 0 37744 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_332
timestamp 1698431365
transform 1 0 38528 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_336
timestamp 1698431365
transform 1 0 38976 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_387
timestamp 1698431365
transform 1 0 44688 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_391
timestamp 1698431365
transform 1 0 45136 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_407
timestamp 1698431365
transform 1 0 46928 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_415
timestamp 1698431365
transform 1 0 47824 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698431365
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_426
timestamp 1698431365
transform 1 0 49056 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_458
timestamp 1698431365
transform 1 0 52640 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698431365
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_31
timestamp 1698431365
transform 1 0 4816 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_59
timestamp 1698431365
transform 1 0 7952 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_67
timestamp 1698431365
transform 1 0 8848 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_71
timestamp 1698431365
transform 1 0 9296 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_73
timestamp 1698431365
transform 1 0 9520 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_80
timestamp 1698431365
transform 1 0 10304 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_84
timestamp 1698431365
transform 1 0 10752 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_86
timestamp 1698431365
transform 1 0 10976 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_96
timestamp 1698431365
transform 1 0 12096 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_98
timestamp 1698431365
transform 1 0 12320 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_124
timestamp 1698431365
transform 1 0 15232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_126
timestamp 1698431365
transform 1 0 15456 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_132
timestamp 1698431365
transform 1 0 16128 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_164
timestamp 1698431365
transform 1 0 19712 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_166
timestamp 1698431365
transform 1 0 19936 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_238
timestamp 1698431365
transform 1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_242
timestamp 1698431365
transform 1 0 28448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_244
timestamp 1698431365
transform 1 0 28672 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_262
timestamp 1698431365
transform 1 0 30688 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_272
timestamp 1698431365
transform 1 0 31808 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_276
timestamp 1698431365
transform 1 0 32256 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_303
timestamp 1698431365
transform 1 0 35280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_307
timestamp 1698431365
transform 1 0 35728 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_325
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_370
timestamp 1698431365
transform 1 0 42784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_374
timestamp 1698431365
transform 1 0 43232 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_382
timestamp 1698431365
transform 1 0 44128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_384
timestamp 1698431365
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_389
timestamp 1698431365
transform 1 0 44912 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_398
timestamp 1698431365
transform 1 0 45920 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_428
timestamp 1698431365
transform 1 0 49280 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_444
timestamp 1698431365
transform 1 0 51072 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_452
timestamp 1698431365
transform 1 0 51968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_454
timestamp 1698431365
transform 1 0 52192 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_489
timestamp 1698431365
transform 1 0 56112 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_505
timestamp 1698431365
transform 1 0 57904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_4
timestamp 1698431365
transform 1 0 1792 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_30
timestamp 1698431365
transform 1 0 4704 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_38
timestamp 1698431365
transform 1 0 5600 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_42
timestamp 1698431365
transform 1 0 6048 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_49
timestamp 1698431365
transform 1 0 6832 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_65
timestamp 1698431365
transform 1 0 8624 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_69
timestamp 1698431365
transform 1 0 9072 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_74
timestamp 1698431365
transform 1 0 9632 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_83
timestamp 1698431365
transform 1 0 10640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_97
timestamp 1698431365
transform 1 0 12208 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_99
timestamp 1698431365
transform 1 0 12432 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_137
timestamp 1698431365
transform 1 0 16688 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_139
timestamp 1698431365
transform 1 0 16912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_150
timestamp 1698431365
transform 1 0 18144 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_169
timestamp 1698431365
transform 1 0 20272 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_179
timestamp 1698431365
transform 1 0 21392 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_181
timestamp 1698431365
transform 1 0 21616 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_208
timestamp 1698431365
transform 1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_237
timestamp 1698431365
transform 1 0 27888 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_277
timestamp 1698431365
transform 1 0 32368 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_279
timestamp 1698431365
transform 1 0 32592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_290
timestamp 1698431365
transform 1 0 33824 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_294
timestamp 1698431365
transform 1 0 34272 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_298
timestamp 1698431365
transform 1 0 34720 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_302
timestamp 1698431365
transform 1 0 35168 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_304
timestamp 1698431365
transform 1 0 35392 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_336
timestamp 1698431365
transform 1 0 38976 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_344
timestamp 1698431365
transform 1 0 39872 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_358
timestamp 1698431365
transform 1 0 41440 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_374
timestamp 1698431365
transform 1 0 43232 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_382
timestamp 1698431365
transform 1 0 44128 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_399
timestamp 1698431365
transform 1 0 46032 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_401
timestamp 1698431365
transform 1 0 46256 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_442
timestamp 1698431365
transform 1 0 50848 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_446
timestamp 1698431365
transform 1 0 51296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_448
timestamp 1698431365
transform 1 0 51520 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_453
timestamp 1698431365
transform 1 0 52080 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_485
timestamp 1698431365
transform 1 0 55664 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_489
timestamp 1698431365
transform 1 0 56112 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1698431365
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_31
timestamp 1698431365
transform 1 0 4816 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_59
timestamp 1698431365
transform 1 0 7952 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_95
timestamp 1698431365
transform 1 0 11984 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_109
timestamp 1698431365
transform 1 0 13552 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_147
timestamp 1698431365
transform 1 0 17808 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_157
timestamp 1698431365
transform 1 0 18928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_161
timestamp 1698431365
transform 1 0 19376 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_181
timestamp 1698431365
transform 1 0 21616 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_183
timestamp 1698431365
transform 1 0 21840 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_192
timestamp 1698431365
transform 1 0 22848 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_200
timestamp 1698431365
transform 1 0 23744 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_216
timestamp 1698431365
transform 1 0 25536 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_223
timestamp 1698431365
transform 1 0 26320 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_227
timestamp 1698431365
transform 1 0 26768 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_231
timestamp 1698431365
transform 1 0 27216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_233
timestamp 1698431365
transform 1 0 27440 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_242
timestamp 1698431365
transform 1 0 28448 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_244
timestamp 1698431365
transform 1 0 28672 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_252
timestamp 1698431365
transform 1 0 29568 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_260
timestamp 1698431365
transform 1 0 30464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_262
timestamp 1698431365
transform 1 0 30688 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_303
timestamp 1698431365
transform 1 0 35280 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_307
timestamp 1698431365
transform 1 0 35728 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_349
timestamp 1698431365
transform 1 0 40432 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_353
timestamp 1698431365
transform 1 0 40880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_355
timestamp 1698431365
transform 1 0 41104 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_428
timestamp 1698431365
transform 1 0 49280 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_444
timestamp 1698431365
transform 1 0 51072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_448
timestamp 1698431365
transform 1 0 51520 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_452
timestamp 1698431365
transform 1 0 51968 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_454
timestamp 1698431365
transform 1 0 52192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_489
timestamp 1698431365
transform 1 0 56112 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_505
timestamp 1698431365
transform 1 0 57904 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_10
timestamp 1698431365
transform 1 0 2464 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_17
timestamp 1698431365
transform 1 0 3248 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_25
timestamp 1698431365
transform 1 0 4144 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_66
timestamp 1698431365
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_150
timestamp 1698431365
transform 1 0 18144 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_173
timestamp 1698431365
transform 1 0 20720 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_177
timestamp 1698431365
transform 1 0 21168 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_185
timestamp 1698431365
transform 1 0 22064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_200
timestamp 1698431365
transform 1 0 23744 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_228
timestamp 1698431365
transform 1 0 26880 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_254
timestamp 1698431365
transform 1 0 29792 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_277
timestamp 1698431365
transform 1 0 32368 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698431365
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_284
timestamp 1698431365
transform 1 0 33152 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_314
timestamp 1698431365
transform 1 0 36512 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_330
timestamp 1698431365
transform 1 0 38304 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_334
timestamp 1698431365
transform 1 0 38752 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_336
timestamp 1698431365
transform 1 0 38976 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_347
timestamp 1698431365
transform 1 0 40208 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_349
timestamp 1698431365
transform 1 0 40432 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_384
timestamp 1698431365
transform 1 0 44352 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_387
timestamp 1698431365
transform 1 0 44688 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_395
timestamp 1698431365
transform 1 0 45584 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_426
timestamp 1698431365
transform 1 0 49056 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_437
timestamp 1698431365
transform 1 0 50288 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_467
timestamp 1698431365
transform 1 0 53648 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_483
timestamp 1698431365
transform 1 0 55440 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_487
timestamp 1698431365
transform 1 0 55888 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_489
timestamp 1698431365
transform 1 0 56112 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698431365
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_55
timestamp 1698431365
transform 1 0 7504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_57
timestamp 1698431365
transform 1 0 7728 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_60
timestamp 1698431365
transform 1 0 8064 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_76
timestamp 1698431365
transform 1 0 9856 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_84
timestamp 1698431365
transform 1 0 10752 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_88
timestamp 1698431365
transform 1 0 11200 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_91
timestamp 1698431365
transform 1 0 11536 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_99
timestamp 1698431365
transform 1 0 12432 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_174
timestamp 1698431365
transform 1 0 20832 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_185
timestamp 1698431365
transform 1 0 22064 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_187
timestamp 1698431365
transform 1 0 22288 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_203
timestamp 1698431365
transform 1 0 24080 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_207
timestamp 1698431365
transform 1 0 24528 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_215
timestamp 1698431365
transform 1 0 25424 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_218
timestamp 1698431365
transform 1 0 25760 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_294
timestamp 1698431365
transform 1 0 34272 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_298
timestamp 1698431365
transform 1 0 34720 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_306
timestamp 1698431365
transform 1 0 35616 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_312
timestamp 1698431365
transform 1 0 36288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_314
timestamp 1698431365
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_333
timestamp 1698431365
transform 1 0 38640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_366
timestamp 1698431365
transform 1 0 42336 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_368
timestamp 1698431365
transform 1 0 42560 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_384
timestamp 1698431365
transform 1 0 44352 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_416
timestamp 1698431365
transform 1 0 47936 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_420
timestamp 1698431365
transform 1 0 48384 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_424
timestamp 1698431365
transform 1 0 48832 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_445
timestamp 1698431365
transform 1 0 51184 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_453
timestamp 1698431365
transform 1 0 52080 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_489
timestamp 1698431365
transform 1 0 56112 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_505
timestamp 1698431365
transform 1 0 57904 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_31
timestamp 1698431365
transform 1 0 4816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_35
timestamp 1698431365
transform 1 0 5264 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_56
timestamp 1698431365
transform 1 0 7616 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_64
timestamp 1698431365
transform 1 0 8512 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_68
timestamp 1698431365
transform 1 0 8960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_80
timestamp 1698431365
transform 1 0 10304 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_82
timestamp 1698431365
transform 1 0 10528 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_91
timestamp 1698431365
transform 1 0 11536 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_157
timestamp 1698431365
transform 1 0 18928 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_178
timestamp 1698431365
transform 1 0 21280 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_186
timestamp 1698431365
transform 1 0 22176 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_190
timestamp 1698431365
transform 1 0 22624 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_209
timestamp 1698431365
transform 1 0 24752 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_230
timestamp 1698431365
transform 1 0 27104 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_274
timestamp 1698431365
transform 1 0 32032 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_278
timestamp 1698431365
transform 1 0 32480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_286
timestamp 1698431365
transform 1 0 33376 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_302
timestamp 1698431365
transform 1 0 35168 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_329
timestamp 1698431365
transform 1 0 38192 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_331
timestamp 1698431365
transform 1 0 38416 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_348
timestamp 1698431365
transform 1 0 40320 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_370
timestamp 1698431365
transform 1 0 42784 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_382
timestamp 1698431365
transform 1 0 44128 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_414
timestamp 1698431365
transform 1 0 47712 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_418
timestamp 1698431365
transform 1 0 48160 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_455
timestamp 1698431365
transform 1 0 52304 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_487
timestamp 1698431365
transform 1 0 55888 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_489
timestamp 1698431365
transform 1 0 56112 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_508
timestamp 1698431365
transform 1 0 58240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_57
timestamp 1698431365
transform 1 0 7728 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_96
timestamp 1698431365
transform 1 0 12096 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_100
timestamp 1698431365
transform 1 0 12544 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_139
timestamp 1698431365
transform 1 0 16912 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_162
timestamp 1698431365
transform 1 0 19488 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_172
timestamp 1698431365
transform 1 0 20608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_174
timestamp 1698431365
transform 1 0 20832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_231
timestamp 1698431365
transform 1 0 27216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_276
timestamp 1698431365
transform 1 0 32256 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_280
timestamp 1698431365
transform 1 0 32704 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_284
timestamp 1698431365
transform 1 0 33152 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_361
timestamp 1698431365
transform 1 0 41776 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_363
timestamp 1698431365
transform 1 0 42000 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_382
timestamp 1698431365
transform 1 0 44128 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698431365
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_425
timestamp 1698431365
transform 1 0 48944 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_447
timestamp 1698431365
transform 1 0 51408 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_451
timestamp 1698431365
transform 1 0 51856 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_486
timestamp 1698431365
transform 1 0 55776 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_502
timestamp 1698431365
transform 1 0 57568 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_506
timestamp 1698431365
transform 1 0 58016 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_508
timestamp 1698431365
transform 1 0 58240 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_18
timestamp 1698431365
transform 1 0 3360 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_34
timestamp 1698431365
transform 1 0 5152 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_64
timestamp 1698431365
transform 1 0 8512 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_68
timestamp 1698431365
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_76
timestamp 1698431365
transform 1 0 9856 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_91
timestamp 1698431365
transform 1 0 11536 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_95
timestamp 1698431365
transform 1 0 11984 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_103
timestamp 1698431365
transform 1 0 12880 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_113
timestamp 1698431365
transform 1 0 14000 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_121
timestamp 1698431365
transform 1 0 14896 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_139
timestamp 1698431365
transform 1 0 16912 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_163
timestamp 1698431365
transform 1 0 19600 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_173
timestamp 1698431365
transform 1 0 20720 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_209
timestamp 1698431365
transform 1 0 24752 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_276
timestamp 1698431365
transform 1 0 32256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_286
timestamp 1698431365
transform 1 0 33376 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_288
timestamp 1698431365
transform 1 0 33600 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_323
timestamp 1698431365
transform 1 0 37520 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_325
timestamp 1698431365
transform 1 0 37744 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_349
timestamp 1698431365
transform 1 0 40432 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_382
timestamp 1698431365
transform 1 0 44128 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_386
timestamp 1698431365
transform 1 0 44576 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_472
timestamp 1698431365
transform 1 0 54208 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_488
timestamp 1698431365
transform 1 0 56000 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698431365
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_31
timestamp 1698431365
transform 1 0 4816 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_74
timestamp 1698431365
transform 1 0 9632 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_78
timestamp 1698431365
transform 1 0 10080 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_93
timestamp 1698431365
transform 1 0 11760 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_123
timestamp 1698431365
transform 1 0 15120 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_153
timestamp 1698431365
transform 1 0 18480 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_161
timestamp 1698431365
transform 1 0 19376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_172
timestamp 1698431365
transform 1 0 20608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_174
timestamp 1698431365
transform 1 0 20832 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_185
timestamp 1698431365
transform 1 0 22064 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_189
timestamp 1698431365
transform 1 0 22512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_198
timestamp 1698431365
transform 1 0 23520 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_200
timestamp 1698431365
transform 1 0 23744 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_210
timestamp 1698431365
transform 1 0 24864 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_241
timestamp 1698431365
transform 1 0 28336 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_255
timestamp 1698431365
transform 1 0 29904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_288
timestamp 1698431365
transform 1 0 33600 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_292
timestamp 1698431365
transform 1 0 34048 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_294
timestamp 1698431365
transform 1 0 34272 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_301
timestamp 1698431365
transform 1 0 35056 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_311
timestamp 1698431365
transform 1 0 36176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_321
timestamp 1698431365
transform 1 0 37296 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_323
timestamp 1698431365
transform 1 0 37520 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_349
timestamp 1698431365
transform 1 0 40432 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_380
timestamp 1698431365
transform 1 0 43904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_384
timestamp 1698431365
transform 1 0 44352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_391
timestamp 1698431365
transform 1 0 45136 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_393
timestamp 1698431365
transform 1 0 45360 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_420
timestamp 1698431365
transform 1 0 48384 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_447
timestamp 1698431365
transform 1 0 51408 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_489
timestamp 1698431365
transform 1 0 56112 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_505
timestamp 1698431365
transform 1 0 57904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_10
timestamp 1698431365
transform 1 0 2464 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_35
timestamp 1698431365
transform 1 0 5264 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_39
timestamp 1698431365
transform 1 0 5712 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_58
timestamp 1698431365
transform 1 0 7840 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_84
timestamp 1698431365
transform 1 0 10752 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_88
timestamp 1698431365
transform 1 0 11200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_120
timestamp 1698431365
transform 1 0 14784 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_128
timestamp 1698431365
transform 1 0 15680 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_132
timestamp 1698431365
transform 1 0 16128 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_138
timestamp 1698431365
transform 1 0 16800 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_189
timestamp 1698431365
transform 1 0 22512 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_218
timestamp 1698431365
transform 1 0 25760 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_222
timestamp 1698431365
transform 1 0 26208 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_230
timestamp 1698431365
transform 1 0 27104 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_234
timestamp 1698431365
transform 1 0 27552 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_236
timestamp 1698431365
transform 1 0 27776 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_266
timestamp 1698431365
transform 1 0 31136 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_270
timestamp 1698431365
transform 1 0 31584 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_317
timestamp 1698431365
transform 1 0 36848 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_319
timestamp 1698431365
transform 1 0 37072 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_349
timestamp 1698431365
transform 1 0 40432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_357
timestamp 1698431365
transform 1 0 41328 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_375
timestamp 1698431365
transform 1 0 43344 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_391
timestamp 1698431365
transform 1 0 45136 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_406
timestamp 1698431365
transform 1 0 46816 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_414
timestamp 1698431365
transform 1 0 47712 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_418
timestamp 1698431365
transform 1 0 48160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_440
timestamp 1698431365
transform 1 0 50624 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_472
timestamp 1698431365
transform 1 0 54208 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_488
timestamp 1698431365
transform 1 0 56000 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_508
timestamp 1698431365
transform 1 0 58240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_31
timestamp 1698431365
transform 1 0 4816 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_45
timestamp 1698431365
transform 1 0 6384 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_113
timestamp 1698431365
transform 1 0 14000 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_129
timestamp 1698431365
transform 1 0 15792 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_137
timestamp 1698431365
transform 1 0 16688 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_149
timestamp 1698431365
transform 1 0 18032 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_170
timestamp 1698431365
transform 1 0 20384 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_174
timestamp 1698431365
transform 1 0 20832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_181
timestamp 1698431365
transform 1 0 21616 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_185
timestamp 1698431365
transform 1 0 22064 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_187
timestamp 1698431365
transform 1 0 22288 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_214
timestamp 1698431365
transform 1 0 25312 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_218
timestamp 1698431365
transform 1 0 25760 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_226
timestamp 1698431365
transform 1 0 26656 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_228
timestamp 1698431365
transform 1 0 26880 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_233
timestamp 1698431365
transform 1 0 27440 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_241
timestamp 1698431365
transform 1 0 28336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_251
timestamp 1698431365
transform 1 0 29456 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_255
timestamp 1698431365
transform 1 0 29904 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_257
timestamp 1698431365
transform 1 0 30128 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_264
timestamp 1698431365
transform 1 0 30912 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_294
timestamp 1698431365
transform 1 0 34272 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_313
timestamp 1698431365
transform 1 0 36400 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_325
timestamp 1698431365
transform 1 0 37744 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_329
timestamp 1698431365
transform 1 0 38192 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_350
timestamp 1698431365
transform 1 0 40544 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_366
timestamp 1698431365
transform 1 0 42336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_382
timestamp 1698431365
transform 1 0 44128 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_384
timestamp 1698431365
transform 1 0 44352 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_416
timestamp 1698431365
transform 1 0 47936 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_418
timestamp 1698431365
transform 1 0 48160 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_448
timestamp 1698431365
transform 1 0 51520 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_452
timestamp 1698431365
transform 1 0 51968 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_454
timestamp 1698431365
transform 1 0 52192 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_489
timestamp 1698431365
transform 1 0 56112 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_505
timestamp 1698431365
transform 1 0 57904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_6
timestamp 1698431365
transform 1 0 2016 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_34
timestamp 1698431365
transform 1 0 5152 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_38
timestamp 1698431365
transform 1 0 5600 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_59
timestamp 1698431365
transform 1 0 7952 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_67
timestamp 1698431365
transform 1 0 8848 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_69
timestamp 1698431365
transform 1 0 9072 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_78
timestamp 1698431365
transform 1 0 10080 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_127
timestamp 1698431365
transform 1 0 15568 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_129
timestamp 1698431365
transform 1 0 15792 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_132
timestamp 1698431365
transform 1 0 16128 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_160
timestamp 1698431365
transform 1 0 19264 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_191
timestamp 1698431365
transform 1 0 22736 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_196
timestamp 1698431365
transform 1 0 23296 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_214
timestamp 1698431365
transform 1 0 25312 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_219
timestamp 1698431365
transform 1 0 25872 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_233
timestamp 1698431365
transform 1 0 27440 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_251
timestamp 1698431365
transform 1 0 29456 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_257
timestamp 1698431365
transform 1 0 30128 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_269
timestamp 1698431365
transform 1 0 31472 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_273
timestamp 1698431365
transform 1 0 31920 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_275
timestamp 1698431365
transform 1 0 32144 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_278
timestamp 1698431365
transform 1 0 32480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_286
timestamp 1698431365
transform 1 0 33376 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_296
timestamp 1698431365
transform 1 0 34496 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_298
timestamp 1698431365
transform 1 0 34720 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_330
timestamp 1698431365
transform 1 0 38304 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_334
timestamp 1698431365
transform 1 0 38752 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_336
timestamp 1698431365
transform 1 0 38976 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_341
timestamp 1698431365
transform 1 0 39536 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_345
timestamp 1698431365
transform 1 0 39984 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_347
timestamp 1698431365
transform 1 0 40208 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_362
timestamp 1698431365
transform 1 0 41888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_395
timestamp 1698431365
transform 1 0 45584 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_399
timestamp 1698431365
transform 1 0 46032 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_415
timestamp 1698431365
transform 1 0 47824 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_419
timestamp 1698431365
transform 1 0 48272 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698431365
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_31
timestamp 1698431365
transform 1 0 4816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_39
timestamp 1698431365
transform 1 0 5712 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_69
timestamp 1698431365
transform 1 0 9072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_73
timestamp 1698431365
transform 1 0 9520 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_123
timestamp 1698431365
transform 1 0 15120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_125
timestamp 1698431365
transform 1 0 15344 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_164
timestamp 1698431365
transform 1 0 19712 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_168
timestamp 1698431365
transform 1 0 20160 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_173
timestamp 1698431365
transform 1 0 20720 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_185
timestamp 1698431365
transform 1 0 22064 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_215
timestamp 1698431365
transform 1 0 25424 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_313
timestamp 1698431365
transform 1 0 36400 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_335
timestamp 1698431365
transform 1 0 38864 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_337
timestamp 1698431365
transform 1 0 39088 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_371
timestamp 1698431365
transform 1 0 42896 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_383
timestamp 1698431365
transform 1 0 44240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_451
timestamp 1698431365
transform 1 0 51856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_489
timestamp 1698431365
transform 1 0 56112 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_505
timestamp 1698431365
transform 1 0 57904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_18
timestamp 1698431365
transform 1 0 3360 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_26
timestamp 1698431365
transform 1 0 4256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_46
timestamp 1698431365
transform 1 0 6496 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_48
timestamp 1698431365
transform 1 0 6720 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_57
timestamp 1698431365
transform 1 0 7728 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_59
timestamp 1698431365
transform 1 0 7952 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_81
timestamp 1698431365
transform 1 0 10416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_93
timestamp 1698431365
transform 1 0 11760 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_101
timestamp 1698431365
transform 1 0 12656 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_159
timestamp 1698431365
transform 1 0 19152 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_176
timestamp 1698431365
transform 1 0 21056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_190
timestamp 1698431365
transform 1 0 22624 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_235
timestamp 1698431365
transform 1 0 27664 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_237
timestamp 1698431365
transform 1 0 27888 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_240
timestamp 1698431365
transform 1 0 28224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_242
timestamp 1698431365
transform 1 0 28448 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_257
timestamp 1698431365
transform 1 0 30128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_271
timestamp 1698431365
transform 1 0 31696 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_284
timestamp 1698431365
transform 1 0 33152 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_298
timestamp 1698431365
transform 1 0 34720 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_318
timestamp 1698431365
transform 1 0 36960 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_332
timestamp 1698431365
transform 1 0 38528 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_396
timestamp 1698431365
transform 1 0 45696 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_405
timestamp 1698431365
transform 1 0 46704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_407
timestamp 1698431365
transform 1 0 46928 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_418
timestamp 1698431365
transform 1 0 48160 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_420
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_429
timestamp 1698431365
transform 1 0 49392 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_441
timestamp 1698431365
transform 1 0 50736 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_444
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_453
timestamp 1698431365
transform 1 0 52080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_465
timestamp 1698431365
transform 1 0 53424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_473
timestamp 1698431365
transform 1 0 54320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_475
timestamp 1698431365
transform 1 0 54544 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_490
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_506
timestamp 1698431365
transform 1 0 58016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1698431365
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 19152 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 20384 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform 1 0 15232 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 15904 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output7 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22624 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output8
timestamp 1698431365
transform -1 0 24864 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output9
timestamp 1698431365
transform -1 0 24192 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output10
timestamp 1698431365
transform -1 0 27440 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output11
timestamp 1698431365
transform -1 0 29008 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output12 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28560 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output13
timestamp 1698431365
transform -1 0 31696 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output14
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output15
timestamp 1698431365
transform 1 0 33600 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output16
timestamp 1698431365
transform 1 0 35840 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output17
timestamp 1698431365
transform 1 0 37408 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output18
timestamp 1698431365
transform -1 0 38416 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output19
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output20
timestamp 1698431365
transform -1 0 42784 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_153
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_154
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_155
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_159
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_160
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_161
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_162
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_164
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_165
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_166
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_167
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_168
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_169
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_171
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_172
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_173
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_174
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_175
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_176
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_178
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_179
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_180
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_181
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_182
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_183
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_185
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_186
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_187
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_188
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_189
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_190
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_192
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_193
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_194
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_195
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_196
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_197
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_199
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_200
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_201
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_202
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_203
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_204
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_206
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_207
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_208
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_209
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_210
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_211
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_213
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_214
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_215
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_216
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_217
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_218
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_220
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_221
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_222
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_223
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_224
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_225
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_227
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_228
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_229
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_230
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_231
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_232
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_234
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_235
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_236
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_237
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_238
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_239
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_241
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_242
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_243
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_244
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_245
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_246
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_248
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_249
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_250
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_251
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_252
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_253
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_258
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_259
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_260
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_267
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_276
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_283
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_284
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_285
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_290
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_291
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_292
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_293
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_294
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_295
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_297
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_298
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_299
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_300
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_301
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_302
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_304
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_305
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_306
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_307
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_308
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_309
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_311
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_312
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_313
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_314
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_315
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_316
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_318
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_319
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_320
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_321
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_322
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_323
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_325
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_326
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_327
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_328
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_329
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_330
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_332
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_333
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_334
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_335
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_336
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_337
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_339
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_340
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_341
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_342
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_343
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_344
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_346
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_347
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_348
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_349
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_350
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_351
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_353
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_354
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_355
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_356
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_357
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_358
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_360
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_361
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_362
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_363
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_364
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_367
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_368
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_369
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_374
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_375
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_392
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_393
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_398
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_399
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_403
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_404
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_405
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_409
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_410
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_416
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_428
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_433
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_434
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_448
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_449
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_453
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_454
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_455
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_456
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_458
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_459
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_460
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_461
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_462
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_463
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_465
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_466
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_467
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_468
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_469
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_470
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_472
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_473
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_474
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_475
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_476
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_477
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_479
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_480
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_481
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_482
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_483
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_484
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_486
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_487
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_488
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_489
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_490
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_491
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_493
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_494
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_495
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_496
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_497
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_498
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_500
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_501
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_502
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_503
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_504
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_505
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_507
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_508
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_509
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_510
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_511
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_512
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_514
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_515
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_516
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_517
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_518
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_519
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_521
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_522
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_523
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_524
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_525
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_526
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_528
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_529
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_530
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_531
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_532
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_533
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_535
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_536
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_537
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_538
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_539
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_540
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_542
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_543
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_544
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_545
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_546
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_547
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_549
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_550
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_551
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_552
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_553
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_554
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_556
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_557
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_558
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_559
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_560
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_561
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_563
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_564
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_565
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_566
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_567
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_568
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_570
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_571
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_572
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_573
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_574
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_575
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_577
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_578
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_579
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_580
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_581
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_582
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_584
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_585
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_586
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_587
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_588
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_589
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_591
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_592
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_593
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_594
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_595
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_596
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_598
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_599
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_600
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_601
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_602
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_603
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_605
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_606
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_607
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_608
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_609
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_610
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_612
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_613
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_614
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_615
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_616
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_617
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_625
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_21 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22064 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_22
timestamp 1698431365
transform -1 0 23296 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_23
timestamp 1698431365
transform -1 0 25312 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_24
timestamp 1698431365
transform -1 0 25872 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_25
timestamp 1698431365
transform -1 0 27440 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_26
timestamp 1698431365
transform -1 0 29456 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_27
timestamp 1698431365
transform -1 0 30128 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_28
timestamp 1698431365
transform -1 0 31472 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_29
timestamp 1698431365
transform -1 0 32704 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_30
timestamp 1698431365
transform -1 0 35616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_31
timestamp 1698431365
transform -1 0 36400 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_32
timestamp 1698431365
transform -1 0 39424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_33
timestamp 1698431365
transform -1 0 38864 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_34
timestamp 1698431365
transform -1 0 39536 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_35
timestamp 1698431365
transform -1 0 6496 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_36
timestamp 1698431365
transform -1 0 7728 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_37
timestamp 1698431365
transform -1 0 8960 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_38
timestamp 1698431365
transform -1 0 10416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_39
timestamp 1698431365
transform -1 0 11760 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_40
timestamp 1698431365
transform -1 0 13440 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_41
timestamp 1698431365
transform -1 0 14336 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_42
timestamp 1698431365
transform 1 0 14784 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_43
timestamp 1698431365
transform 1 0 16128 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_44
timestamp 1698431365
transform 1 0 16912 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_45
timestamp 1698431365
transform -1 0 19712 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_46
timestamp 1698431365
transform -1 0 21056 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_47
timestamp 1698431365
transform -1 0 41888 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_48
timestamp 1698431365
transform -1 0 44352 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_49
timestamp 1698431365
transform -1 0 44240 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_50
timestamp 1698431365
transform -1 0 45696 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_51
timestamp 1698431365
transform -1 0 46704 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_52
timestamp 1698431365
transform -1 0 48160 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_53
timestamp 1698431365
transform -1 0 49392 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_54
timestamp 1698431365
transform -1 0 50736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_55
timestamp 1698431365
transform -1 0 52080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_56
timestamp 1698431365
transform -1 0 53424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_57
timestamp 1698431365
transform -1 0 55328 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_58
timestamp 1698431365
transform -1 0 56224 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_59 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_60
timestamp 1698431365
transform -1 0 7280 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_61
timestamp 1698431365
transform -1 0 8512 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_62
timestamp 1698431365
transform -1 0 9968 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_63
timestamp 1698431365
transform -1 0 11312 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_64
timestamp 1698431365
transform -1 0 12656 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_65
timestamp 1698431365
transform -1 0 13888 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_66
timestamp 1698431365
transform 1 0 14336 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_67
timestamp 1698431365
transform 1 0 15680 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_68
timestamp 1698431365
transform -1 0 19712 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_69
timestamp 1698431365
transform 1 0 18032 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_70
timestamp 1698431365
transform -1 0 20720 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_71
timestamp 1698431365
transform -1 0 43232 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_72
timestamp 1698431365
transform -1 0 43904 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_73
timestamp 1698431365
transform -1 0 44800 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_74
timestamp 1698431365
transform -1 0 45248 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_75
timestamp 1698431365
transform -1 0 46256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_76
timestamp 1698431365
transform -1 0 47712 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_77
timestamp 1698431365
transform -1 0 48944 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_78
timestamp 1698431365
transform -1 0 50288 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_79
timestamp 1698431365
transform -1 0 51632 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_80
timestamp 1698431365
transform -1 0 52976 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_81
timestamp 1698431365
transform -1 0 54320 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_82
timestamp 1698431365
transform -1 0 55776 0 -1 56448
box -86 -86 534 870
<< labels >>
flabel metal2 s 4928 59200 5040 60000 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 18368 59200 18480 60000 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 19712 59200 19824 60000 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 21056 59200 21168 60000 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 22400 59200 22512 60000 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 23744 59200 23856 60000 0 FreeSans 448 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 25088 59200 25200 60000 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 26432 59200 26544 60000 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 27776 59200 27888 60000 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 29120 59200 29232 60000 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 30464 59200 30576 60000 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 6272 59200 6384 60000 0 FreeSans 448 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 31808 59200 31920 60000 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 33152 59200 33264 60000 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 34496 59200 34608 60000 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 35840 59200 35952 60000 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 37184 59200 37296 60000 0 FreeSans 448 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 38528 59200 38640 60000 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 39872 59200 39984 60000 0 FreeSans 448 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 41216 59200 41328 60000 0 FreeSans 448 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 42560 59200 42672 60000 0 FreeSans 448 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 43904 59200 44016 60000 0 FreeSans 448 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 7616 59200 7728 60000 0 FreeSans 448 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 45248 59200 45360 60000 0 FreeSans 448 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 46592 59200 46704 60000 0 FreeSans 448 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 47936 59200 48048 60000 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 49280 59200 49392 60000 0 FreeSans 448 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 50624 59200 50736 60000 0 FreeSans 448 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 51968 59200 52080 60000 0 FreeSans 448 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 53312 59200 53424 60000 0 FreeSans 448 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 54656 59200 54768 60000 0 FreeSans 448 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 8960 59200 9072 60000 0 FreeSans 448 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 10304 59200 10416 60000 0 FreeSans 448 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 11648 59200 11760 60000 0 FreeSans 448 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 12992 59200 13104 60000 0 FreeSans 448 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 14336 59200 14448 60000 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 15680 59200 15792 60000 0 FreeSans 448 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 17024 59200 17136 60000 0 FreeSans 448 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 5376 59200 5488 60000 0 FreeSans 448 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 18816 59200 18928 60000 0 FreeSans 448 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 20160 59200 20272 60000 0 FreeSans 448 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 21504 59200 21616 60000 0 FreeSans 448 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 22848 59200 22960 60000 0 FreeSans 448 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 24192 59200 24304 60000 0 FreeSans 448 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 25536 59200 25648 60000 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 26880 59200 26992 60000 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 28224 59200 28336 60000 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 29568 59200 29680 60000 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 30912 59200 31024 60000 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 6720 59200 6832 60000 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 32256 59200 32368 60000 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 33600 59200 33712 60000 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 34944 59200 35056 60000 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 36288 59200 36400 60000 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 37632 59200 37744 60000 0 FreeSans 448 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 38976 59200 39088 60000 0 FreeSans 448 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 40320 59200 40432 60000 0 FreeSans 448 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 41664 59200 41776 60000 0 FreeSans 448 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 43008 59200 43120 60000 0 FreeSans 448 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 44352 59200 44464 60000 0 FreeSans 448 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 8064 59200 8176 60000 0 FreeSans 448 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 45696 59200 45808 60000 0 FreeSans 448 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 47040 59200 47152 60000 0 FreeSans 448 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 48384 59200 48496 60000 0 FreeSans 448 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 49728 59200 49840 60000 0 FreeSans 448 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 51072 59200 51184 60000 0 FreeSans 448 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 52416 59200 52528 60000 0 FreeSans 448 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 53760 59200 53872 60000 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 55104 59200 55216 60000 0 FreeSans 448 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 9408 59200 9520 60000 0 FreeSans 448 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 10752 59200 10864 60000 0 FreeSans 448 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 12096 59200 12208 60000 0 FreeSans 448 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 13440 59200 13552 60000 0 FreeSans 448 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 14784 59200 14896 60000 0 FreeSans 448 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 16128 59200 16240 60000 0 FreeSans 448 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 17472 59200 17584 60000 0 FreeSans 448 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 5824 59200 5936 60000 0 FreeSans 448 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 19264 59200 19376 60000 0 FreeSans 448 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 20608 59200 20720 60000 0 FreeSans 448 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 21952 59200 22064 60000 0 FreeSans 448 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 23296 59200 23408 60000 0 FreeSans 448 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 24640 59200 24752 60000 0 FreeSans 448 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 25984 59200 26096 60000 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 27328 59200 27440 60000 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 28672 59200 28784 60000 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 30016 59200 30128 60000 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 31360 59200 31472 60000 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 7168 59200 7280 60000 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 32704 59200 32816 60000 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 34048 59200 34160 60000 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 35392 59200 35504 60000 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 36736 59200 36848 60000 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 38080 59200 38192 60000 0 FreeSans 448 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 39424 59200 39536 60000 0 FreeSans 448 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 40768 59200 40880 60000 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 42112 59200 42224 60000 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 43456 59200 43568 60000 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 44800 59200 44912 60000 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 8512 59200 8624 60000 0 FreeSans 448 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 46144 59200 46256 60000 0 FreeSans 448 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 47488 59200 47600 60000 0 FreeSans 448 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 48832 59200 48944 60000 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 50176 59200 50288 60000 0 FreeSans 448 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 51520 59200 51632 60000 0 FreeSans 448 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 52864 59200 52976 60000 0 FreeSans 448 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 54208 59200 54320 60000 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 55552 59200 55664 60000 0 FreeSans 448 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 9856 59200 9968 60000 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 11200 59200 11312 60000 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 12544 59200 12656 60000 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 13888 59200 14000 60000 0 FreeSans 448 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 15232 59200 15344 60000 0 FreeSans 448 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 16576 59200 16688 60000 0 FreeSans 448 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 17920 59200 18032 60000 0 FreeSans 448 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 114 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 114 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 115 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 115 nsew ground bidirectional
flabel metal2 s 4032 59200 4144 60000 0 FreeSans 448 90 0 0 wb_clk_i
port 116 nsew signal input
flabel metal2 s 4480 59200 4592 60000 0 FreeSans 448 90 0 0 wb_rst_i
port 117 nsew signal input
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 16072 22288 16072 22288 0 _0000_
rlabel metal2 22344 20328 22344 20328 0 _0001_
rlabel metal2 15848 28084 15848 28084 0 _0002_
rlabel metal2 16352 28616 16352 28616 0 _0003_
rlabel metal2 15624 21168 15624 21168 0 _0004_
rlabel metal2 27496 38360 27496 38360 0 _0005_
rlabel metal3 13104 35112 13104 35112 0 _0006_
rlabel metal2 10360 37072 10360 37072 0 _0007_
rlabel metal2 17528 34552 17528 34552 0 _0008_
rlabel metal2 9464 40040 9464 40040 0 _0009_
rlabel metal2 26264 36848 26264 36848 0 _0010_
rlabel metal3 13216 38696 13216 38696 0 _0011_
rlabel metal2 21448 34440 21448 34440 0 _0012_
rlabel metal3 42056 55160 42056 55160 0 _0013_
rlabel metal3 44156 54600 44156 54600 0 _0014_
rlabel metal3 5264 26936 5264 26936 0 _0015_
rlabel metal2 7112 25592 7112 25592 0 _0016_
rlabel metal2 3080 21896 3080 21896 0 _0017_
rlabel metal2 2520 20440 2520 20440 0 _0018_
rlabel metal2 12936 26628 12936 26628 0 _0019_
rlabel metal2 10192 25592 10192 25592 0 _0020_
rlabel metal2 14280 24416 14280 24416 0 _0021_
rlabel metal2 10360 22624 10360 22624 0 _0022_
rlabel metal2 9912 30464 9912 30464 0 _0023_
rlabel metal2 9800 28280 9800 28280 0 _0024_
rlabel metal2 17584 20216 17584 20216 0 _0025_
rlabel metal2 19544 18760 19544 18760 0 _0026_
rlabel metal2 12936 6216 12936 6216 0 _0027_
rlabel metal2 10192 6776 10192 6776 0 _0028_
rlabel metal2 16408 5600 16408 5600 0 _0029_
rlabel metal2 16408 7896 16408 7896 0 _0030_
rlabel metal2 2968 24136 2968 24136 0 _0031_
rlabel metal2 2688 23240 2688 23240 0 _0032_
rlabel metal2 45640 53368 45640 53368 0 _0033_
rlabel metal2 13272 10920 13272 10920 0 _0034_
rlabel metal2 9576 9464 9576 9464 0 _0035_
rlabel metal2 6888 12488 6888 12488 0 _0036_
rlabel metal2 6440 9352 6440 9352 0 _0037_
rlabel metal2 2464 14616 2464 14616 0 _0038_
rlabel metal2 3528 15624 3528 15624 0 _0039_
rlabel metal2 2408 17752 2408 17752 0 _0040_
rlabel metal2 3416 18760 3416 18760 0 _0041_
rlabel metal2 2576 13048 2576 13048 0 _0042_
rlabel metal2 3360 11256 3360 11256 0 _0043_
rlabel metal2 16408 11032 16408 11032 0 _0044_
rlabel metal2 18424 10136 18424 10136 0 _0045_
rlabel metal2 28672 29176 28672 29176 0 _0046_
rlabel metal2 20440 30632 20440 30632 0 _0047_
rlabel metal2 13720 29736 13720 29736 0 _0048_
rlabel metal2 14280 30408 14280 30408 0 _0049_
rlabel metal3 16856 28728 16856 28728 0 _0050_
rlabel metal3 27720 37128 27720 37128 0 _0051_
rlabel metal2 45248 46536 45248 46536 0 _0052_
rlabel metal2 45640 48664 45640 48664 0 _0053_
rlabel metal2 48328 46424 48328 46424 0 _0054_
rlabel metal2 50232 46032 50232 46032 0 _0055_
rlabel metal2 51016 47656 51016 47656 0 _0056_
rlabel metal3 51968 51464 51968 51464 0 _0057_
rlabel metal2 49000 53368 49000 53368 0 _0058_
rlabel metal3 52528 50456 52528 50456 0 _0059_
rlabel metal2 33936 34216 33936 34216 0 _0060_
rlabel metal2 37688 32984 37688 32984 0 _0061_
rlabel metal2 40040 35224 40040 35224 0 _0062_
rlabel metal2 40488 36624 40488 36624 0 _0063_
rlabel metal2 41832 46200 41832 46200 0 _0064_
rlabel metal2 42392 44688 42392 44688 0 _0065_
rlabel metal3 43624 37912 43624 37912 0 _0066_
rlabel metal2 46648 40208 46648 40208 0 _0067_
rlabel metal2 49224 42000 49224 42000 0 _0068_
rlabel metal2 54824 39984 54824 39984 0 _0069_
rlabel metal3 44520 34216 44520 34216 0 _0070_
rlabel metal3 52136 38696 52136 38696 0 _0071_
rlabel metal2 54936 33768 54936 33768 0 _0072_
rlabel metal3 56840 35000 56840 35000 0 _0073_
rlabel metal3 54040 31640 54040 31640 0 _0074_
rlabel metal2 41888 31864 41888 31864 0 _0075_
rlabel metal2 46984 29008 46984 29008 0 _0076_
rlabel metal3 54152 26936 54152 26936 0 _0077_
rlabel metal2 50792 25424 50792 25424 0 _0078_
rlabel metal2 51632 23016 51632 23016 0 _0079_
rlabel metal2 45584 20104 45584 20104 0 _0080_
rlabel metal2 45696 20888 45696 20888 0 _0081_
rlabel metal3 45136 26488 45136 26488 0 _0082_
rlabel metal2 40936 27776 40936 27776 0 _0083_
rlabel metal2 39704 21168 39704 21168 0 _0084_
rlabel metal2 38696 25872 38696 25872 0 _0085_
rlabel metal2 36960 21672 36960 21672 0 _0086_
rlabel metal2 36456 26628 36456 26628 0 _0087_
rlabel metal2 30744 25872 30744 25872 0 _0088_
rlabel metal2 30184 28168 30184 28168 0 _0089_
rlabel metal2 34384 31080 34384 31080 0 _0090_
rlabel metal2 37632 31080 37632 31080 0 _0091_
rlabel metal2 46536 43904 46536 43904 0 _0092_
rlabel metal2 34888 47824 34888 47824 0 _0093_
rlabel metal3 35000 38696 35000 38696 0 _0094_
rlabel metal2 20216 53312 20216 53312 0 _0095_
rlabel metal3 19880 54376 19880 54376 0 _0096_
rlabel metal2 29848 30632 29848 30632 0 _0097_
rlabel metal3 30520 28728 30520 28728 0 _0098_
rlabel metal2 29792 50456 29792 50456 0 _0099_
rlabel metal2 26824 49392 26824 49392 0 _0100_
rlabel metal2 28896 48440 28896 48440 0 _0101_
rlabel metal2 31752 34048 31752 34048 0 _0102_
rlabel metal2 29400 34272 29400 34272 0 _0103_
rlabel metal2 32256 39032 32256 39032 0 _0104_
rlabel metal2 33880 37408 33880 37408 0 _0105_
rlabel metal2 35112 45192 35112 45192 0 _0106_
rlabel metal3 35112 43624 35112 43624 0 _0107_
rlabel metal2 37800 39872 37800 39872 0 _0108_
rlabel metal2 35672 40712 35672 40712 0 _0109_
rlabel metal2 36568 42112 36568 42112 0 _0110_
rlabel metal2 32760 41328 32760 41328 0 _0111_
rlabel metal2 9016 41720 9016 41720 0 _0112_
rlabel metal2 8904 43064 8904 43064 0 _0113_
rlabel metal3 9520 43624 9520 43624 0 _0114_
rlabel metal2 9016 47768 9016 47768 0 _0115_
rlabel metal3 10416 50456 10416 50456 0 _0116_
rlabel metal2 10024 53088 10024 53088 0 _0117_
rlabel metal2 14392 53368 14392 53368 0 _0118_
rlabel metal2 13272 52920 13272 52920 0 _0119_
rlabel metal2 17640 48664 17640 48664 0 _0120_
rlabel metal2 16296 51800 16296 51800 0 _0121_
rlabel metal2 2856 53368 2856 53368 0 _0122_
rlabel metal2 2520 54936 2520 54936 0 _0123_
rlabel metal2 4536 51800 4536 51800 0 _0124_
rlabel metal2 7784 54768 7784 54768 0 _0125_
rlabel metal2 6552 51016 6552 51016 0 _0126_
rlabel metal2 2520 50176 2520 50176 0 _0127_
rlabel metal2 6888 48048 6888 48048 0 _0128_
rlabel metal2 6216 44744 6216 44744 0 _0129_
rlabel metal3 7392 38136 7392 38136 0 _0130_
rlabel metal2 2520 38472 2520 38472 0 _0131_
rlabel metal2 2520 40152 2520 40152 0 _0132_
rlabel metal2 6552 40768 6552 40768 0 _0133_
rlabel metal2 2968 41608 2968 41608 0 _0134_
rlabel metal2 3864 43792 3864 43792 0 _0135_
rlabel metal2 3864 46424 3864 46424 0 _0136_
rlabel metal2 3864 47824 3864 47824 0 _0137_
rlabel metal2 27160 28168 27160 28168 0 _0138_
rlabel metal2 24304 26488 24304 26488 0 _0139_
rlabel metal2 22008 29064 22008 29064 0 _0140_
rlabel metal2 16296 27552 16296 27552 0 _0141_
rlabel metal2 16072 26376 16072 26376 0 _0142_
rlabel metal2 28840 32872 28840 32872 0 _0143_
rlabel metal2 24584 33656 24584 33656 0 _0144_
rlabel metal2 21336 31416 21336 31416 0 _0145_
rlabel metal3 13384 31864 13384 31864 0 _0146_
rlabel metal2 14224 33432 14224 33432 0 _0147_
rlabel metal3 25088 50456 25088 50456 0 _0148_
rlabel metal2 23072 53816 23072 53816 0 _0149_
rlabel metal2 24696 54712 24696 54712 0 _0150_
rlabel metal2 27384 52472 27384 52472 0 _0151_
rlabel metal3 34832 17752 34832 17752 0 _0152_
rlabel metal3 36680 15400 36680 15400 0 _0153_
rlabel metal2 17976 13608 17976 13608 0 _0154_
rlabel metal2 22568 11648 22568 11648 0 _0155_
rlabel metal2 15176 14056 15176 14056 0 _0156_
rlabel metal2 10360 13272 10360 13272 0 _0157_
rlabel metal3 29960 12824 29960 12824 0 _0158_
rlabel metal2 31080 10304 31080 10304 0 _0159_
rlabel metal2 18312 16352 18312 16352 0 _0160_
rlabel metal2 20888 15148 20888 15148 0 _0161_
rlabel metal2 31752 17192 31752 17192 0 _0162_
rlabel metal3 32088 14392 32088 14392 0 _0163_
rlabel metal3 33208 12264 33208 12264 0 _0164_
rlabel metal2 38472 12488 38472 12488 0 _0165_
rlabel metal2 9016 15736 9016 15736 0 _0166_
rlabel metal2 8008 14168 8008 14168 0 _0167_
rlabel metal2 25816 21280 25816 21280 0 _0168_
rlabel metal2 29176 20328 29176 20328 0 _0169_
rlabel metal2 32032 21784 32032 21784 0 _0170_
rlabel metal3 35056 20104 35056 20104 0 _0171_
rlabel metal2 21224 4648 21224 4648 0 _0172_
rlabel metal2 21672 5040 21672 5040 0 _0173_
rlabel metal2 25368 7168 25368 7168 0 _0174_
rlabel metal2 28056 6216 28056 6216 0 _0175_
rlabel metal2 20440 6944 20440 6944 0 _0176_
rlabel metal2 22232 10304 22232 10304 0 _0177_
rlabel metal2 25480 8904 25480 8904 0 _0178_
rlabel metal2 28504 9352 28504 9352 0 _0179_
rlabel metal2 26376 23464 26376 23464 0 _0180_
rlabel metal3 30128 23240 30128 23240 0 _0181_
rlabel metal2 32032 19320 32032 19320 0 _0182_
rlabel metal3 36456 18424 36456 18424 0 _0183_
rlabel metal2 4648 27104 4648 27104 0 _0184_
rlabel metal2 6328 28896 6328 28896 0 _0185_
rlabel metal2 26936 51632 26936 51632 0 _0186_
rlabel metal2 28840 53312 28840 53312 0 _0187_
rlabel metal2 30352 53480 30352 53480 0 _0188_
rlabel metal3 31612 52024 31612 52024 0 _0189_
rlabel metal2 32200 53368 32200 53368 0 _0190_
rlabel metal2 33656 54152 33656 54152 0 _0191_
rlabel metal2 35896 53984 35896 53984 0 _0192_
rlabel metal2 46312 31472 46312 31472 0 _0193_
rlabel metal2 44688 43400 44688 43400 0 _0194_
rlabel metal2 45080 36232 45080 36232 0 _0195_
rlabel metal3 45192 38696 45192 38696 0 _0196_
rlabel metal2 41496 30520 41496 30520 0 _0197_
rlabel metal2 45192 36848 45192 36848 0 _0198_
rlabel metal2 45752 37128 45752 37128 0 _0199_
rlabel metal2 42504 30464 42504 30464 0 _0200_
rlabel metal2 51576 27160 51576 27160 0 _0201_
rlabel metal2 52024 27608 52024 27608 0 _0202_
rlabel metal2 42168 40824 42168 40824 0 _0203_
rlabel metal2 43064 39704 43064 39704 0 _0204_
rlabel metal3 43848 40264 43848 40264 0 _0205_
rlabel metal2 45640 39928 45640 39928 0 _0206_
rlabel metal2 46200 39592 46200 39592 0 _0207_
rlabel metal2 43624 21392 43624 21392 0 _0208_
rlabel metal2 51520 40376 51520 40376 0 _0209_
rlabel metal2 45752 39144 45752 39144 0 _0210_
rlabel metal2 51128 41160 51128 41160 0 _0211_
rlabel metal2 43400 41832 43400 41832 0 _0212_
rlabel metal2 45080 42224 45080 42224 0 _0213_
rlabel metal3 42952 41048 42952 41048 0 _0214_
rlabel metal2 43960 40936 43960 40936 0 _0215_
rlabel metal2 43512 41104 43512 41104 0 _0216_
rlabel metal2 51968 42616 51968 42616 0 _0217_
rlabel metal2 48552 39648 48552 39648 0 _0218_
rlabel metal3 48664 31528 48664 31528 0 _0219_
rlabel metal3 48664 38808 48664 38808 0 _0220_
rlabel metal2 48272 39032 48272 39032 0 _0221_
rlabel metal2 49000 40040 49000 40040 0 _0222_
rlabel metal2 50456 38752 50456 38752 0 _0223_
rlabel metal2 50008 39200 50008 39200 0 _0224_
rlabel metal2 46816 39032 46816 39032 0 _0225_
rlabel metal2 51296 42616 51296 42616 0 _0226_
rlabel metal2 51800 42224 51800 42224 0 _0227_
rlabel metal3 53312 42504 53312 42504 0 _0228_
rlabel metal3 52360 42728 52360 42728 0 _0229_
rlabel metal2 52360 42448 52360 42448 0 _0230_
rlabel metal2 50792 41440 50792 41440 0 _0231_
rlabel metal2 50568 40096 50568 40096 0 _0232_
rlabel metal2 51912 40544 51912 40544 0 _0233_
rlabel metal3 47040 35672 47040 35672 0 _0234_
rlabel metal2 48664 36456 48664 36456 0 _0235_
rlabel metal2 49952 41384 49952 41384 0 _0236_
rlabel metal2 52136 42616 52136 42616 0 _0237_
rlabel metal2 52024 41720 52024 41720 0 _0238_
rlabel metal2 53144 40096 53144 40096 0 _0239_
rlabel metal2 53032 36736 53032 36736 0 _0240_
rlabel metal2 50680 35168 50680 35168 0 _0241_
rlabel metal2 45080 35224 45080 35224 0 _0242_
rlabel metal2 39144 20944 39144 20944 0 _0243_
rlabel metal2 43792 33544 43792 33544 0 _0244_
rlabel metal2 43624 34104 43624 34104 0 _0245_
rlabel metal2 46760 22792 46760 22792 0 _0246_
rlabel metal2 51128 36400 51128 36400 0 _0247_
rlabel metal2 50680 36512 50680 36512 0 _0248_
rlabel metal2 50904 36344 50904 36344 0 _0249_
rlabel metal3 49000 36232 49000 36232 0 _0250_
rlabel metal2 52192 35672 52192 35672 0 _0251_
rlabel metal2 49000 34384 49000 34384 0 _0252_
rlabel metal2 47768 36344 47768 36344 0 _0253_
rlabel metal2 47992 35672 47992 35672 0 _0254_
rlabel metal2 48216 36064 48216 36064 0 _0255_
rlabel metal2 47768 35728 47768 35728 0 _0256_
rlabel metal2 48104 36008 48104 36008 0 _0257_
rlabel metal2 54824 33600 54824 33600 0 _0258_
rlabel metal2 53760 34888 53760 34888 0 _0259_
rlabel metal2 54432 24024 54432 24024 0 _0260_
rlabel metal2 52584 36176 52584 36176 0 _0261_
rlabel metal2 53144 36176 53144 36176 0 _0262_
rlabel metal2 55048 36736 55048 36736 0 _0263_
rlabel metal2 50120 36456 50120 36456 0 _0264_
rlabel metal2 51464 35728 51464 35728 0 _0265_
rlabel metal2 52248 37744 52248 37744 0 _0266_
rlabel metal2 54712 37184 54712 37184 0 _0267_
rlabel metal2 56616 36064 56616 36064 0 _0268_
rlabel metal2 55216 34104 55216 34104 0 _0269_
rlabel metal2 54264 33544 54264 33544 0 _0270_
rlabel metal2 54432 34664 54432 34664 0 _0271_
rlabel metal2 55160 36400 55160 36400 0 _0272_
rlabel metal2 57288 34440 57288 34440 0 _0273_
rlabel metal3 56952 34328 56952 34328 0 _0274_
rlabel metal2 40040 28168 40040 28168 0 _0275_
rlabel metal2 50904 21000 50904 21000 0 _0276_
rlabel metal2 53480 29344 53480 29344 0 _0277_
rlabel metal2 52920 29232 52920 29232 0 _0278_
rlabel metal2 49952 30856 49952 30856 0 _0279_
rlabel metal2 52024 31080 52024 31080 0 _0280_
rlabel metal2 53256 34048 53256 34048 0 _0281_
rlabel metal2 51016 34384 51016 34384 0 _0282_
rlabel metal2 50512 30184 50512 30184 0 _0283_
rlabel metal2 50904 32256 50904 32256 0 _0284_
rlabel metal2 50344 32704 50344 32704 0 _0285_
rlabel metal3 51352 31976 51352 31976 0 _0286_
rlabel metal2 50904 22624 50904 22624 0 _0287_
rlabel metal2 47152 23128 47152 23128 0 _0288_
rlabel metal2 49784 25760 49784 25760 0 _0289_
rlabel metal2 44744 31024 44744 31024 0 _0290_
rlabel metal2 49784 30464 49784 30464 0 _0291_
rlabel metal3 53592 30184 53592 30184 0 _0292_
rlabel metal2 52136 30520 52136 30520 0 _0293_
rlabel metal2 50064 29288 50064 29288 0 _0294_
rlabel metal2 44856 30296 44856 30296 0 _0295_
rlabel metal2 45192 30016 45192 30016 0 _0296_
rlabel metal2 43512 31864 43512 31864 0 _0297_
rlabel metal3 42560 32424 42560 32424 0 _0298_
rlabel metal2 45640 28784 45640 28784 0 _0299_
rlabel metal2 50568 29512 50568 29512 0 _0300_
rlabel metal2 51128 28896 51128 28896 0 _0301_
rlabel metal2 45640 30968 45640 30968 0 _0302_
rlabel metal2 46536 27720 46536 27720 0 _0303_
rlabel metal2 45304 29680 45304 29680 0 _0304_
rlabel metal2 50232 28672 50232 28672 0 _0305_
rlabel metal2 49000 29960 49000 29960 0 _0306_
rlabel metal2 52248 25312 52248 25312 0 _0307_
rlabel metal2 48832 26376 48832 26376 0 _0308_
rlabel metal2 50008 26992 50008 26992 0 _0309_
rlabel metal2 52920 26824 52920 26824 0 _0310_
rlabel metal3 52416 25480 52416 25480 0 _0311_
rlabel metal3 51128 26264 51128 26264 0 _0312_
rlabel metal3 50288 26152 50288 26152 0 _0313_
rlabel metal2 50456 25816 50456 25816 0 _0314_
rlabel metal2 51128 25984 51128 25984 0 _0315_
rlabel metal2 52752 22568 52752 22568 0 _0316_
rlabel metal2 50120 24584 50120 24584 0 _0317_
rlabel metal2 53368 24808 53368 24808 0 _0318_
rlabel metal2 53144 28728 53144 28728 0 _0319_
rlabel metal2 55832 26152 55832 26152 0 _0320_
rlabel metal3 51576 23240 51576 23240 0 _0321_
rlabel metal2 53032 23800 53032 23800 0 _0322_
rlabel metal3 52696 23800 52696 23800 0 _0323_
rlabel metal2 51464 23128 51464 23128 0 _0324_
rlabel metal3 45752 23912 45752 23912 0 _0325_
rlabel metal2 44296 22568 44296 22568 0 _0326_
rlabel metal3 47040 22456 47040 22456 0 _0327_
rlabel metal2 51464 25312 51464 25312 0 _0328_
rlabel metal2 47320 24752 47320 24752 0 _0329_
rlabel metal2 45976 23072 45976 23072 0 _0330_
rlabel metal2 45976 24248 45976 24248 0 _0331_
rlabel metal2 48776 24360 48776 24360 0 _0332_
rlabel metal2 48104 25088 48104 25088 0 _0333_
rlabel metal2 47544 22848 47544 22848 0 _0334_
rlabel metal2 43848 23968 43848 23968 0 _0335_
rlabel metal2 50680 24360 50680 24360 0 _0336_
rlabel metal3 47320 25200 47320 25200 0 _0337_
rlabel metal3 43792 26264 43792 26264 0 _0338_
rlabel metal2 45752 23632 45752 23632 0 _0339_
rlabel metal2 45864 22400 45864 22400 0 _0340_
rlabel metal3 46704 22344 46704 22344 0 _0341_
rlabel metal2 47768 25816 47768 25816 0 _0342_
rlabel metal2 47208 26376 47208 26376 0 _0343_
rlabel metal3 47208 26376 47208 26376 0 _0344_
rlabel metal3 44464 26376 44464 26376 0 _0345_
rlabel metal2 47656 21504 47656 21504 0 _0346_
rlabel metal2 45192 22456 45192 22456 0 _0347_
rlabel metal2 43288 24864 43288 24864 0 _0348_
rlabel metal3 46424 23240 46424 23240 0 _0349_
rlabel via2 42392 23912 42392 23912 0 _0350_
rlabel metal3 42112 25368 42112 25368 0 _0351_
rlabel metal2 44072 26600 44072 26600 0 _0352_
rlabel metal3 43456 26600 43456 26600 0 _0353_
rlabel metal2 42280 26992 42280 26992 0 _0354_
rlabel metal2 42392 27384 42392 27384 0 _0355_
rlabel metal2 41720 27832 41720 27832 0 _0356_
rlabel metal3 41720 21560 41720 21560 0 _0357_
rlabel metal2 42504 21728 42504 21728 0 _0358_
rlabel metal2 41048 25816 41048 25816 0 _0359_
rlabel metal3 43400 20888 43400 20888 0 _0360_
rlabel metal3 43792 21448 43792 21448 0 _0361_
rlabel metal2 41272 24920 41272 24920 0 _0362_
rlabel metal2 42616 23688 42616 23688 0 _0363_
rlabel metal3 41048 23800 41048 23800 0 _0364_
rlabel metal2 41888 25480 41888 25480 0 _0365_
rlabel metal2 39928 24752 39928 24752 0 _0366_
rlabel metal2 41944 25144 41944 25144 0 _0367_
rlabel metal2 44744 25088 44744 25088 0 _0368_
rlabel metal2 38584 23184 38584 23184 0 _0369_
rlabel metal2 38696 24080 38696 24080 0 _0370_
rlabel metal3 40152 24920 40152 24920 0 _0371_
rlabel metal2 37352 21616 37352 21616 0 _0372_
rlabel metal2 37128 22232 37128 22232 0 _0373_
rlabel metal2 40376 23632 40376 23632 0 _0374_
rlabel metal2 35616 21784 35616 21784 0 _0375_
rlabel metal3 36344 22344 36344 22344 0 _0376_
rlabel metal2 38472 24360 38472 24360 0 _0377_
rlabel metal2 35560 23632 35560 23632 0 _0378_
rlabel metal3 36680 23800 36680 23800 0 _0379_
rlabel metal2 35224 23800 35224 23800 0 _0380_
rlabel metal2 37240 24360 37240 24360 0 _0381_
rlabel metal2 37912 25200 37912 25200 0 _0382_
rlabel metal3 36456 26712 36456 26712 0 _0383_
rlabel metal2 27608 32088 27608 32088 0 _0384_
rlabel metal3 33096 26320 33096 26320 0 _0385_
rlabel metal2 34216 25872 34216 25872 0 _0386_
rlabel metal3 34328 26264 34328 26264 0 _0387_
rlabel metal2 34552 22904 34552 22904 0 _0388_
rlabel metal2 35112 24584 35112 24584 0 _0389_
rlabel metal2 23912 40656 23912 40656 0 _0390_
rlabel metal2 32984 28224 32984 28224 0 _0391_
rlabel metal2 33320 27664 33320 27664 0 _0392_
rlabel metal2 34048 25368 34048 25368 0 _0393_
rlabel metal2 35448 29736 35448 29736 0 _0394_
rlabel metal2 34216 27832 34216 27832 0 _0395_
rlabel metal2 34552 28000 34552 28000 0 _0396_
rlabel metal2 34552 28952 34552 28952 0 _0397_
rlabel metal3 34384 29288 34384 29288 0 _0398_
rlabel metal2 34888 30016 34888 30016 0 _0399_
rlabel metal2 32424 30632 32424 30632 0 _0400_
rlabel metal2 34944 28616 34944 28616 0 _0401_
rlabel metal3 36624 30408 36624 30408 0 _0402_
rlabel metal2 45808 43512 45808 43512 0 _0403_
rlabel metal2 19544 49112 19544 49112 0 _0404_
rlabel metal2 20552 48384 20552 48384 0 _0405_
rlabel metal2 34384 47544 34384 47544 0 _0406_
rlabel metal2 30184 32424 30184 32424 0 _0407_
rlabel metal2 24808 43792 24808 43792 0 _0408_
rlabel metal2 20328 53032 20328 53032 0 _0409_
rlabel metal2 24360 43008 24360 43008 0 _0410_
rlabel metal2 24024 44744 24024 44744 0 _0411_
rlabel metal2 18984 44912 18984 44912 0 _0412_
rlabel metal2 29288 29624 29288 29624 0 _0413_
rlabel metal2 29960 29288 29960 29288 0 _0414_
rlabel metal2 28448 50456 28448 50456 0 _0415_
rlabel metal2 23240 46480 23240 46480 0 _0416_
rlabel metal2 24304 48216 24304 48216 0 _0417_
rlabel metal2 26376 49000 26376 49000 0 _0418_
rlabel metal2 24136 46256 24136 46256 0 _0419_
rlabel metal3 15344 49560 15344 49560 0 _0420_
rlabel metal3 16520 51464 16520 51464 0 _0421_
rlabel metal2 17976 51128 17976 51128 0 _0422_
rlabel metal3 15624 45640 15624 45640 0 _0423_
rlabel metal2 24360 45528 24360 45528 0 _0424_
rlabel metal2 21112 45080 21112 45080 0 _0425_
rlabel metal2 21784 44632 21784 44632 0 _0426_
rlabel metal4 24584 45696 24584 45696 0 _0427_
rlabel metal2 28952 48048 28952 48048 0 _0428_
rlabel metal3 28504 48776 28504 48776 0 _0429_
rlabel metal2 28168 50120 28168 50120 0 _0430_
rlabel metal2 31472 46872 31472 46872 0 _0431_
rlabel metal2 28784 50456 28784 50456 0 _0432_
rlabel metal2 28280 49840 28280 49840 0 _0433_
rlabel metal2 23352 46704 23352 46704 0 _0434_
rlabel metal3 22288 47208 22288 47208 0 _0435_
rlabel metal2 25424 47208 25424 47208 0 _0436_
rlabel metal2 27384 48440 27384 48440 0 _0437_
rlabel metal2 26488 48216 26488 48216 0 _0438_
rlabel metal2 29064 48160 29064 48160 0 _0439_
rlabel metal3 30352 45864 30352 45864 0 _0440_
rlabel metal2 30856 46312 30856 46312 0 _0441_
rlabel metal3 23240 46760 23240 46760 0 _0442_
rlabel metal2 22904 42168 22904 42168 0 _0443_
rlabel metal3 22064 40376 22064 40376 0 _0444_
rlabel metal2 22792 41216 22792 41216 0 _0445_
rlabel metal2 22232 40824 22232 40824 0 _0446_
rlabel metal2 23352 41440 23352 41440 0 _0447_
rlabel metal3 34888 37800 34888 37800 0 _0448_
rlabel metal2 29288 45472 29288 45472 0 _0449_
rlabel metal2 29400 45024 29400 45024 0 _0450_
rlabel metal3 32648 46648 32648 46648 0 _0451_
rlabel metal2 33208 44128 33208 44128 0 _0452_
rlabel metal2 31304 44240 31304 44240 0 _0453_
rlabel metal3 27160 46424 27160 46424 0 _0454_
rlabel metal2 27608 47152 27608 47152 0 _0455_
rlabel metal2 27832 46704 27832 46704 0 _0456_
rlabel metal2 30632 41104 30632 41104 0 _0457_
rlabel metal2 30912 40264 30912 40264 0 _0458_
rlabel metal2 31472 35112 31472 35112 0 _0459_
rlabel metal2 26936 41552 26936 41552 0 _0460_
rlabel metal2 29400 40880 29400 40880 0 _0461_
rlabel metal2 25592 39760 25592 39760 0 _0462_
rlabel metal2 24024 39592 24024 39592 0 _0463_
rlabel metal3 25144 41944 25144 41944 0 _0464_
rlabel metal2 26152 42056 26152 42056 0 _0465_
rlabel metal2 26600 40880 26600 40880 0 _0466_
rlabel metal2 26376 41776 26376 41776 0 _0467_
rlabel metal2 27048 46648 27048 46648 0 _0468_
rlabel metal2 12600 44632 12600 44632 0 _0469_
rlabel metal2 14504 45528 14504 45528 0 _0470_
rlabel metal2 25256 42672 25256 42672 0 _0471_
rlabel metal2 25536 42728 25536 42728 0 _0472_
rlabel metal2 25480 42224 25480 42224 0 _0473_
rlabel metal3 18984 44296 18984 44296 0 _0474_
rlabel metal3 31808 45192 31808 45192 0 _0475_
rlabel metal2 26376 43736 26376 43736 0 _0476_
rlabel metal2 27608 43400 27608 43400 0 _0477_
rlabel metal2 29960 38472 29960 38472 0 _0478_
rlabel metal2 30408 35336 30408 35336 0 _0479_
rlabel metal2 16464 46648 16464 46648 0 _0480_
rlabel metal2 22456 47208 22456 47208 0 _0481_
rlabel metal2 28896 40600 28896 40600 0 _0482_
rlabel metal2 27496 40320 27496 40320 0 _0483_
rlabel metal2 29176 43120 29176 43120 0 _0484_
rlabel metal3 30520 38808 30520 38808 0 _0485_
rlabel metal3 25004 41720 25004 41720 0 _0486_
rlabel metal2 32928 40488 32928 40488 0 _0487_
rlabel metal2 32816 38808 32816 38808 0 _0488_
rlabel metal3 33432 42056 33432 42056 0 _0489_
rlabel metal3 29792 39592 29792 39592 0 _0490_
rlabel metal2 28056 39592 28056 39592 0 _0491_
rlabel metal2 24472 46984 24472 46984 0 _0492_
rlabel metal2 24136 47544 24136 47544 0 _0493_
rlabel metal2 24808 45752 24808 45752 0 _0494_
rlabel metal2 28392 45360 28392 45360 0 _0495_
rlabel metal2 26600 44184 26600 44184 0 _0496_
rlabel metal2 25480 44016 25480 44016 0 _0497_
rlabel metal2 27160 43232 27160 43232 0 _0498_
rlabel metal3 31136 40152 31136 40152 0 _0499_
rlabel metal2 34328 38024 34328 38024 0 _0500_
rlabel metal3 25200 41160 25200 41160 0 _0501_
rlabel via2 25928 42392 25928 42392 0 _0502_
rlabel metal2 29400 42504 29400 42504 0 _0503_
rlabel metal2 26264 45808 26264 45808 0 _0504_
rlabel metal2 29736 43232 29736 43232 0 _0505_
rlabel metal2 29568 42840 29568 42840 0 _0506_
rlabel metal2 34216 44408 34216 44408 0 _0507_
rlabel metal2 26488 45920 26488 45920 0 _0508_
rlabel metal3 31024 44184 31024 44184 0 _0509_
rlabel metal2 33432 44352 33432 44352 0 _0510_
rlabel metal2 33656 44464 33656 44464 0 _0511_
rlabel metal2 30744 43288 30744 43288 0 _0512_
rlabel metal2 31136 40488 31136 40488 0 _0513_
rlabel metal3 34048 40936 34048 40936 0 _0514_
rlabel metal3 36344 42168 36344 42168 0 _0515_
rlabel metal3 36792 41048 36792 41048 0 _0516_
rlabel metal2 27552 42168 27552 42168 0 _0517_
rlabel metal2 28280 44520 28280 44520 0 _0518_
rlabel metal2 28392 42000 28392 42000 0 _0519_
rlabel metal2 27888 41160 27888 41160 0 _0520_
rlabel metal3 32144 41048 32144 41048 0 _0521_
rlabel metal2 15960 44296 15960 44296 0 _0522_
rlabel metal2 35168 41160 35168 41160 0 _0523_
rlabel metal2 29960 42280 29960 42280 0 _0524_
rlabel metal2 24920 43848 24920 43848 0 _0525_
rlabel metal2 27832 43232 27832 43232 0 _0526_
rlabel metal2 34328 43120 34328 43120 0 _0527_
rlabel metal3 35952 42616 35952 42616 0 _0528_
rlabel metal2 30632 44464 30632 44464 0 _0529_
rlabel metal2 27496 45360 27496 45360 0 _0530_
rlabel metal2 30072 44744 30072 44744 0 _0531_
rlabel metal2 31528 43120 31528 43120 0 _0532_
rlabel metal2 32760 41720 32760 41720 0 _0533_
rlabel metal2 14728 40768 14728 40768 0 _0534_
rlabel metal3 18368 42952 18368 42952 0 _0535_
rlabel metal3 17528 43288 17528 43288 0 _0536_
rlabel metal2 17528 44464 17528 44464 0 _0537_
rlabel metal3 16268 44408 16268 44408 0 _0538_
rlabel metal2 13104 41944 13104 41944 0 _0539_
rlabel metal2 7448 49616 7448 49616 0 _0540_
rlabel metal2 5768 46424 5768 46424 0 _0541_
rlabel metal2 3080 52976 3080 52976 0 _0542_
rlabel metal2 6552 46872 6552 46872 0 _0543_
rlabel metal2 5768 39928 5768 39928 0 _0544_
rlabel metal2 4984 41384 4984 41384 0 _0545_
rlabel metal2 2072 44800 2072 44800 0 _0546_
rlabel metal3 6216 45864 6216 45864 0 _0547_
rlabel metal3 8512 45752 8512 45752 0 _0548_
rlabel metal3 10752 43512 10752 43512 0 _0549_
rlabel metal2 12824 43120 12824 43120 0 _0550_
rlabel metal2 12432 41944 12432 41944 0 _0551_
rlabel metal2 14280 43736 14280 43736 0 _0552_
rlabel metal2 13832 44352 13832 44352 0 _0553_
rlabel metal2 16744 42336 16744 42336 0 _0554_
rlabel metal2 22680 42336 22680 42336 0 _0555_
rlabel metal2 16856 42112 16856 42112 0 _0556_
rlabel metal2 13608 42840 13608 42840 0 _0557_
rlabel metal2 13832 43456 13832 43456 0 _0558_
rlabel metal2 10248 47320 10248 47320 0 _0559_
rlabel metal2 10696 43792 10696 43792 0 _0560_
rlabel metal2 16856 43960 16856 43960 0 _0561_
rlabel metal2 15736 43960 15736 43960 0 _0562_
rlabel metal2 15288 44800 15288 44800 0 _0563_
rlabel metal2 10696 48048 10696 48048 0 _0564_
rlabel metal2 9912 47544 9912 47544 0 _0565_
rlabel metal2 14616 42336 14616 42336 0 _0566_
rlabel metal2 13720 43260 13720 43260 0 _0567_
rlabel metal2 11592 50960 11592 50960 0 _0568_
rlabel metal2 11256 51296 11256 51296 0 _0569_
rlabel metal2 11368 52696 11368 52696 0 _0570_
rlabel metal2 13384 52696 13384 52696 0 _0571_
rlabel metal2 16352 41944 16352 41944 0 _0572_
rlabel metal2 16352 42168 16352 42168 0 _0573_
rlabel metal3 13664 52808 13664 52808 0 _0574_
rlabel metal2 13552 51352 13552 51352 0 _0575_
rlabel metal2 16072 51128 16072 51128 0 _0576_
rlabel metal2 18144 50008 18144 50008 0 _0577_
rlabel metal2 17304 45696 17304 45696 0 _0578_
rlabel metal2 16520 51240 16520 51240 0 _0579_
rlabel metal2 17752 48496 17752 48496 0 _0580_
rlabel metal2 14392 38136 14392 38136 0 _0581_
rlabel metal2 17304 47656 17304 47656 0 _0582_
rlabel metal2 15848 52080 15848 52080 0 _0583_
rlabel metal2 5992 43456 5992 43456 0 _0584_
rlabel metal2 2744 53088 2744 53088 0 _0585_
rlabel metal2 2800 54488 2800 54488 0 _0586_
rlabel metal2 6384 46760 6384 46760 0 _0587_
rlabel metal2 5096 52584 5096 52584 0 _0588_
rlabel metal2 4424 51520 4424 51520 0 _0589_
rlabel metal2 7280 54488 7280 54488 0 _0590_
rlabel metal3 6440 49784 6440 49784 0 _0591_
rlabel metal2 7168 50568 7168 50568 0 _0592_
rlabel metal2 6048 50008 6048 50008 0 _0593_
rlabel metal2 7224 50120 7224 50120 0 _0594_
rlabel metal3 7448 48216 7448 48216 0 _0595_
rlabel metal2 8456 48272 8456 48272 0 _0596_
rlabel metal2 6440 40768 6440 40768 0 _0597_
rlabel metal2 6552 44632 6552 44632 0 _0598_
rlabel metal2 6944 44296 6944 44296 0 _0599_
rlabel metal2 6328 39256 6328 39256 0 _0600_
rlabel metal2 6664 39536 6664 39536 0 _0601_
rlabel metal3 4424 44184 4424 44184 0 _0602_
rlabel metal2 7672 39088 7672 39088 0 _0603_
rlabel metal3 3416 38920 3416 38920 0 _0604_
rlabel metal2 3976 39032 3976 39032 0 _0605_
rlabel metal2 5320 41552 5320 41552 0 _0606_
rlabel metal2 4480 39368 4480 39368 0 _0607_
rlabel metal3 6608 41160 6608 41160 0 _0608_
rlabel metal3 4480 41832 4480 41832 0 _0609_
rlabel metal2 3192 41720 3192 41720 0 _0610_
rlabel metal2 3528 41160 3528 41160 0 _0611_
rlabel metal3 4760 43624 4760 43624 0 _0612_
rlabel metal2 3304 45640 3304 45640 0 _0613_
rlabel metal2 2520 44912 2520 44912 0 _0614_
rlabel metal2 2744 46480 2744 46480 0 _0615_
rlabel metal2 2632 46984 2632 46984 0 _0616_
rlabel metal2 26376 29904 26376 29904 0 _0617_
rlabel metal3 21784 28504 21784 28504 0 _0618_
rlabel metal2 24416 26376 24416 26376 0 _0619_
rlabel metal2 25480 28336 25480 28336 0 _0620_
rlabel metal2 24024 26572 24024 26572 0 _0621_
rlabel metal3 22624 35784 22624 35784 0 _0622_
rlabel metal2 21616 24248 21616 24248 0 _0623_
rlabel metal2 22736 25480 22736 25480 0 _0624_
rlabel metal2 22344 28224 22344 28224 0 _0625_
rlabel metal2 20328 27384 20328 27384 0 _0626_
rlabel metal2 19432 27384 19432 27384 0 _0627_
rlabel metal2 20440 26572 20440 26572 0 _0628_
rlabel metal2 19544 26544 19544 26544 0 _0629_
rlabel metal2 24472 34272 24472 34272 0 _0630_
rlabel metal2 23800 50848 23800 50848 0 _0631_
rlabel metal2 23128 51184 23128 51184 0 _0632_
rlabel metal2 23520 51464 23520 51464 0 _0633_
rlabel metal2 23576 50092 23576 50092 0 _0634_
rlabel metal2 19320 41720 19320 41720 0 _0635_
rlabel metal3 20776 41944 20776 41944 0 _0636_
rlabel metal2 21504 49000 21504 49000 0 _0637_
rlabel metal3 20104 49784 20104 49784 0 _0638_
rlabel metal2 21336 48944 21336 48944 0 _0639_
rlabel metal3 21504 50456 21504 50456 0 _0640_
rlabel metal2 22792 50680 22792 50680 0 _0641_
rlabel metal2 23016 42896 23016 42896 0 _0642_
rlabel metal2 23576 47656 23576 47656 0 _0643_
rlabel metal2 22960 48440 22960 48440 0 _0644_
rlabel metal3 23912 49784 23912 49784 0 _0645_
rlabel metal2 22568 48552 22568 48552 0 _0646_
rlabel metal2 24864 42056 24864 42056 0 _0647_
rlabel metal3 23408 48888 23408 48888 0 _0648_
rlabel metal2 24136 40880 24136 40880 0 _0649_
rlabel metal2 23688 45024 23688 45024 0 _0650_
rlabel metal2 22792 49448 22792 49448 0 _0651_
rlabel metal3 21392 49672 21392 49672 0 _0652_
rlabel metal2 23352 53592 23352 53592 0 _0653_
rlabel metal2 23800 53536 23800 53536 0 _0654_
rlabel metal2 23912 49392 23912 49392 0 _0655_
rlabel metal2 23800 49756 23800 49756 0 _0656_
rlabel metal2 19880 51296 19880 51296 0 _0657_
rlabel metal3 20944 51240 20944 51240 0 _0658_
rlabel metal2 21896 52248 21896 52248 0 _0659_
rlabel metal2 24192 52808 24192 52808 0 _0660_
rlabel metal2 24192 50008 24192 50008 0 _0661_
rlabel metal2 19992 50904 19992 50904 0 _0662_
rlabel metal2 22568 51856 22568 51856 0 _0663_
rlabel metal2 24472 52472 24472 52472 0 _0664_
rlabel metal2 29960 11872 29960 11872 0 _0665_
rlabel metal2 35504 15064 35504 15064 0 _0666_
rlabel metal2 33656 17752 33656 17752 0 _0667_
rlabel metal2 31360 10584 31360 10584 0 _0668_
rlabel metal2 35168 14728 35168 14728 0 _0669_
rlabel metal2 13888 12824 13888 12824 0 _0670_
rlabel metal2 19768 13328 19768 13328 0 _0671_
rlabel metal2 18312 13216 18312 13216 0 _0672_
rlabel metal3 11256 13832 11256 13832 0 _0673_
rlabel metal3 21448 11368 21448 11368 0 _0674_
rlabel metal3 13048 12824 13048 12824 0 _0675_
rlabel metal2 14672 13160 14672 13160 0 _0676_
rlabel metal2 11256 12152 11256 12152 0 _0677_
rlabel metal2 24584 20160 24584 20160 0 _0678_
rlabel metal2 30296 12488 30296 12488 0 _0679_
rlabel metal2 29624 12432 29624 12432 0 _0680_
rlabel metal2 30296 10528 30296 10528 0 _0681_
rlabel metal2 21784 23072 21784 23072 0 _0682_
rlabel metal2 21952 20104 21952 20104 0 _0683_
rlabel metal3 20776 16072 20776 16072 0 _0684_
rlabel metal2 18928 15960 18928 15960 0 _0685_
rlabel metal2 21448 14000 21448 14000 0 _0686_
rlabel metal3 26040 15960 26040 15960 0 _0687_
rlabel metal2 26264 15512 26264 15512 0 _0688_
rlabel metal2 30408 16912 30408 16912 0 _0689_
rlabel metal2 30632 14784 30632 14784 0 _0690_
rlabel metal2 26936 11704 26936 11704 0 _0691_
rlabel metal2 33208 11648 33208 11648 0 _0692_
rlabel metal2 35392 11592 35392 11592 0 _0693_
rlabel metal2 12320 14504 12320 14504 0 _0694_
rlabel metal3 9968 14728 9968 14728 0 _0695_
rlabel metal3 9072 13720 9072 13720 0 _0696_
rlabel metal2 33768 20664 33768 20664 0 _0697_
rlabel metal2 27944 19544 27944 19544 0 _0698_
rlabel metal2 26824 20888 26824 20888 0 _0699_
rlabel metal2 36120 19880 36120 19880 0 _0700_
rlabel metal2 29288 20104 29288 20104 0 _0701_
rlabel metal2 33768 21560 33768 21560 0 _0702_
rlabel metal2 32816 21560 32816 21560 0 _0703_
rlabel metal3 34888 20776 34888 20776 0 _0704_
rlabel metal2 20888 7336 20888 7336 0 _0705_
rlabel metal2 22232 5936 22232 5936 0 _0706_
rlabel metal2 20440 5376 20440 5376 0 _0707_
rlabel metal2 28280 9520 28280 9520 0 _0708_
rlabel metal2 21336 5376 21336 5376 0 _0709_
rlabel metal2 26712 9408 26712 9408 0 _0710_
rlabel metal2 25704 6776 25704 6776 0 _0711_
rlabel metal2 27832 6944 27832 6944 0 _0712_
rlabel metal2 23576 9016 23576 9016 0 _0713_
rlabel metal2 20664 7728 20664 7728 0 _0714_
rlabel metal2 22232 9464 22232 9464 0 _0715_
rlabel metal2 26824 9856 26824 9856 0 _0716_
rlabel metal2 25816 8512 25816 8512 0 _0717_
rlabel metal2 28056 10080 28056 10080 0 _0718_
rlabel metal2 27720 22288 27720 22288 0 _0719_
rlabel metal2 26600 23240 26600 23240 0 _0720_
rlabel metal2 29288 23240 29288 23240 0 _0721_
rlabel metal3 24976 19992 24976 19992 0 _0722_
rlabel metal2 25928 19936 25928 19936 0 _0723_
rlabel metal2 32424 20328 32424 20328 0 _0724_
rlabel metal2 35000 18704 35000 18704 0 _0725_
rlabel metal2 7616 23912 7616 23912 0 _0726_
rlabel metal2 4984 27328 4984 27328 0 _0727_
rlabel metal3 6888 28616 6888 28616 0 _0728_
rlabel metal2 42504 51520 42504 51520 0 _0729_
rlabel metal2 49112 47768 49112 47768 0 _0730_
rlabel metal2 47432 51744 47432 51744 0 _0731_
rlabel metal3 48440 49896 48440 49896 0 _0732_
rlabel metal2 43960 50428 43960 50428 0 _0733_
rlabel metal3 42280 52024 42280 52024 0 _0734_
rlabel metal2 47096 51576 47096 51576 0 _0735_
rlabel metal2 46480 51352 46480 51352 0 _0736_
rlabel metal3 46648 51520 46648 51520 0 _0737_
rlabel metal3 50176 50568 50176 50568 0 _0738_
rlabel metal2 48328 51352 48328 51352 0 _0739_
rlabel metal2 43288 50624 43288 50624 0 _0740_
rlabel metal2 43736 51800 43736 51800 0 _0741_
rlabel metal2 42112 51464 42112 51464 0 _0742_
rlabel metal2 38472 53088 38472 53088 0 _0743_
rlabel metal3 40544 48776 40544 48776 0 _0744_
rlabel metal2 45640 51240 45640 51240 0 _0745_
rlabel metal2 42952 49504 42952 49504 0 _0746_
rlabel metal2 39984 51128 39984 51128 0 _0747_
rlabel metal2 42280 52976 42280 52976 0 _0748_
rlabel metal2 42616 50960 42616 50960 0 _0749_
rlabel metal2 42504 50736 42504 50736 0 _0750_
rlabel metal2 37464 50568 37464 50568 0 _0751_
rlabel metal2 43848 51520 43848 51520 0 _0752_
rlabel metal2 42504 49952 42504 49952 0 _0753_
rlabel metal2 41104 52136 41104 52136 0 _0754_
rlabel metal2 41944 50848 41944 50848 0 _0755_
rlabel metal2 43624 50064 43624 50064 0 _0756_
rlabel metal3 42336 49784 42336 49784 0 _0757_
rlabel metal3 38360 50456 38360 50456 0 _0758_
rlabel metal2 39256 48664 39256 48664 0 _0759_
rlabel metal3 41048 50456 41048 50456 0 _0760_
rlabel metal2 37352 51128 37352 51128 0 _0761_
rlabel metal2 38136 53200 38136 53200 0 _0762_
rlabel metal3 36792 50456 36792 50456 0 _0763_
rlabel metal2 35616 51912 35616 51912 0 _0764_
rlabel metal3 38640 51576 38640 51576 0 _0765_
rlabel metal2 39256 52752 39256 52752 0 _0766_
rlabel metal2 40264 51576 40264 51576 0 _0767_
rlabel metal2 40264 52248 40264 52248 0 _0768_
rlabel metal2 37912 52472 37912 52472 0 _0769_
rlabel metal3 43764 51128 43764 51128 0 _0770_
rlabel metal3 38808 51128 38808 51128 0 _0771_
rlabel metal2 39256 51240 39256 51240 0 _0772_
rlabel metal2 38808 52136 38808 52136 0 _0773_
rlabel metal3 34888 53032 34888 53032 0 _0774_
rlabel metal2 37688 52248 37688 52248 0 _0775_
rlabel metal2 35840 52920 35840 52920 0 _0776_
rlabel metal2 34216 52584 34216 52584 0 _0777_
rlabel metal2 40208 53480 40208 53480 0 _0778_
rlabel metal2 35336 50568 35336 50568 0 _0779_
rlabel metal2 36456 50792 36456 50792 0 _0780_
rlabel metal2 34440 52248 34440 52248 0 _0781_
rlabel metal2 35560 52976 35560 52976 0 _0782_
rlabel metal2 37128 51184 37128 51184 0 _0783_
rlabel metal2 36736 51352 36736 51352 0 _0784_
rlabel metal2 36344 52304 36344 52304 0 _0785_
rlabel metal2 36792 53368 36792 53368 0 _0786_
rlabel metal2 21560 39312 21560 39312 0 _0787_
rlabel metal2 31976 36848 31976 36848 0 _0788_
rlabel metal3 32984 36456 32984 36456 0 _0789_
rlabel metal3 19656 40600 19656 40600 0 _0790_
rlabel metal3 19544 40152 19544 40152 0 _0791_
rlabel metal2 22120 41104 22120 41104 0 _0792_
rlabel metal2 12432 48216 12432 48216 0 _0793_
rlabel metal2 14616 46592 14616 46592 0 _0794_
rlabel metal2 18200 51688 18200 51688 0 _0795_
rlabel metal3 18872 50344 18872 50344 0 _0796_
rlabel metal2 15960 49112 15960 49112 0 _0797_
rlabel metal2 15064 45584 15064 45584 0 _0798_
rlabel metal2 15848 46424 15848 46424 0 _0799_
rlabel metal2 12880 45752 12880 45752 0 _0800_
rlabel metal2 15736 46592 15736 46592 0 _0801_
rlabel metal2 13832 47208 13832 47208 0 _0802_
rlabel metal2 19824 48440 19824 48440 0 _0803_
rlabel metal2 16408 49392 16408 49392 0 _0804_
rlabel metal2 13104 48776 13104 48776 0 _0805_
rlabel metal2 14504 41664 14504 41664 0 _0806_
rlabel metal2 19432 41608 19432 41608 0 _0807_
rlabel metal3 22176 45864 22176 45864 0 _0808_
rlabel metal3 21448 46648 21448 46648 0 _0809_
rlabel metal2 18480 55496 18480 55496 0 _0810_
rlabel metal2 18648 48496 18648 48496 0 _0811_
rlabel metal2 19040 48328 19040 48328 0 _0812_
rlabel metal2 17416 41272 17416 41272 0 _0813_
rlabel metal2 13272 40712 13272 40712 0 _0814_
rlabel metal2 20440 44520 20440 44520 0 _0815_
rlabel metal3 13160 50568 13160 50568 0 _0816_
rlabel metal2 15400 52080 15400 52080 0 _0817_
rlabel metal2 12264 47880 12264 47880 0 _0818_
rlabel metal2 13496 46760 13496 46760 0 _0819_
rlabel metal3 19768 49560 19768 49560 0 _0820_
rlabel metal3 12824 46536 12824 46536 0 _0821_
rlabel metal3 11312 45640 11312 45640 0 _0822_
rlabel metal3 13048 46648 13048 46648 0 _0823_
rlabel metal2 17416 45808 17416 45808 0 _0824_
rlabel metal3 31416 46760 31416 46760 0 _0825_
rlabel metal3 20720 46536 20720 46536 0 _0826_
rlabel metal2 16632 38976 16632 38976 0 _0827_
rlabel metal2 17640 36736 17640 36736 0 _0828_
rlabel metal2 17752 34440 17752 34440 0 _0829_
rlabel metal2 18872 32200 18872 32200 0 _0830_
rlabel metal2 16632 31472 16632 31472 0 _0831_
rlabel metal2 16184 31528 16184 31528 0 _0832_
rlabel metal2 16352 30856 16352 30856 0 _0833_
rlabel metal2 17416 31640 17416 31640 0 _0834_
rlabel metal2 25480 29792 25480 29792 0 _0835_
rlabel metal2 26376 32648 26376 32648 0 _0836_
rlabel metal2 26488 29736 26488 29736 0 _0837_
rlabel metal3 24864 30184 24864 30184 0 _0838_
rlabel metal2 24248 31248 24248 31248 0 _0839_
rlabel metal2 23576 30352 23576 30352 0 _0840_
rlabel metal2 23240 29456 23240 29456 0 _0841_
rlabel metal2 25256 30856 25256 30856 0 _0842_
rlabel metal2 18312 32088 18312 32088 0 _0843_
rlabel metal3 17640 31640 17640 31640 0 _0844_
rlabel metal2 18536 33040 18536 33040 0 _0845_
rlabel metal3 18536 30968 18536 30968 0 _0846_
rlabel metal2 19264 31192 19264 31192 0 _0847_
rlabel metal2 18704 35672 18704 35672 0 _0848_
rlabel metal3 20272 35896 20272 35896 0 _0849_
rlabel metal3 20664 18984 20664 18984 0 _0850_
rlabel metal2 27496 14224 27496 14224 0 _0851_
rlabel metal2 24248 15904 24248 15904 0 _0852_
rlabel metal3 25536 15288 25536 15288 0 _0853_
rlabel metal2 27664 15288 27664 15288 0 _0854_
rlabel metal2 16184 16856 16184 16856 0 _0855_
rlabel metal2 22568 17584 22568 17584 0 _0856_
rlabel metal2 28840 12992 28840 12992 0 _0857_
rlabel metal2 30016 10024 30016 10024 0 _0858_
rlabel metal2 29736 18480 29736 18480 0 _0859_
rlabel metal2 29512 17248 29512 17248 0 _0860_
rlabel metal2 23240 18872 23240 18872 0 _0861_
rlabel metal3 23688 12936 23688 12936 0 _0862_
rlabel metal2 26824 15344 26824 15344 0 _0863_
rlabel metal2 27384 15064 27384 15064 0 _0864_
rlabel metal2 24808 15680 24808 15680 0 _0865_
rlabel metal3 31752 13720 31752 13720 0 _0866_
rlabel metal2 29176 8036 29176 8036 0 _0867_
rlabel metal2 31752 11536 31752 11536 0 _0868_
rlabel metal2 28504 11816 28504 11816 0 _0869_
rlabel metal2 27440 13496 27440 13496 0 _0870_
rlabel metal2 16128 16296 16128 16296 0 _0871_
rlabel metal2 27272 14280 27272 14280 0 _0872_
rlabel metal2 25032 14896 25032 14896 0 _0873_
rlabel metal2 24584 16016 24584 16016 0 _0874_
rlabel metal2 24920 16296 24920 16296 0 _0875_
rlabel metal2 28504 14784 28504 14784 0 _0876_
rlabel metal3 28896 17640 28896 17640 0 _0877_
rlabel metal3 29008 17864 29008 17864 0 _0878_
rlabel metal2 28112 14728 28112 14728 0 _0879_
rlabel metal2 27608 14616 27608 14616 0 _0880_
rlabel metal2 23912 12320 23912 12320 0 _0881_
rlabel metal2 23016 11088 23016 11088 0 _0882_
rlabel metal2 23688 12712 23688 12712 0 _0883_
rlabel metal2 24024 12824 24024 12824 0 _0884_
rlabel metal2 24080 15512 24080 15512 0 _0885_
rlabel metal2 23968 16968 23968 16968 0 _0886_
rlabel metal3 24752 16184 24752 16184 0 _0887_
rlabel metal2 25424 17864 25424 17864 0 _0888_
rlabel metal2 12376 17584 12376 17584 0 _0889_
rlabel metal2 12824 9464 12824 9464 0 _0890_
rlabel metal2 8680 15064 8680 15064 0 _0891_
rlabel metal2 9800 18480 9800 18480 0 _0892_
rlabel metal2 10360 18536 10360 18536 0 _0893_
rlabel metal2 14504 12320 14504 12320 0 _0894_
rlabel metal2 10976 19992 10976 19992 0 _0895_
rlabel metal3 10696 19992 10696 19992 0 _0896_
rlabel metal2 11536 18424 11536 18424 0 _0897_
rlabel metal3 15540 21672 15540 21672 0 _0898_
rlabel metal2 14056 17920 14056 17920 0 _0899_
rlabel metal2 11704 10864 11704 10864 0 _0900_
rlabel metal2 7168 17080 7168 17080 0 _0901_
rlabel metal2 15736 22064 15736 22064 0 _0902_
rlabel metal3 9184 18200 9184 18200 0 _0903_
rlabel metal3 11312 17864 11312 17864 0 _0904_
rlabel metal2 15624 17808 15624 17808 0 _0905_
rlabel metal2 12824 17528 12824 17528 0 _0906_
rlabel metal3 15400 20160 15400 20160 0 _0907_
rlabel metal2 12320 9240 12320 9240 0 _0908_
rlabel metal2 9632 20776 9632 20776 0 _0909_
rlabel metal3 9632 21000 9632 21000 0 _0910_
rlabel metal3 11368 19432 11368 19432 0 _0911_
rlabel metal2 12936 19152 12936 19152 0 _0912_
rlabel metal2 13720 21112 13720 21112 0 _0913_
rlabel metal2 13496 21056 13496 21056 0 _0914_
rlabel metal2 7784 17976 7784 17976 0 _0915_
rlabel metal2 8120 22596 8120 22596 0 _0916_
rlabel metal2 8512 21560 8512 21560 0 _0917_
rlabel via2 8232 21560 8232 21560 0 _0918_
rlabel metal2 13944 21112 13944 21112 0 _0919_
rlabel metal3 13496 19768 13496 19768 0 _0920_
rlabel metal2 13832 20440 13832 20440 0 _0921_
rlabel metal2 16408 20384 16408 20384 0 _0922_
rlabel metal2 23576 22512 23576 22512 0 _0923_
rlabel metal2 24192 38136 24192 38136 0 _0924_
rlabel metal2 24696 17472 24696 17472 0 _0925_
rlabel metal2 26376 16632 26376 16632 0 _0926_
rlabel metal2 25984 16632 25984 16632 0 _0927_
rlabel metal2 26600 15960 26600 15960 0 _0928_
rlabel metal3 20104 15400 20104 15400 0 _0929_
rlabel metal2 26376 18592 26376 18592 0 _0930_
rlabel metal2 25256 18032 25256 18032 0 _0931_
rlabel metal2 26712 17136 26712 17136 0 _0932_
rlabel metal2 25704 16408 25704 16408 0 _0933_
rlabel metal3 27048 14280 27048 14280 0 _0934_
rlabel metal2 26376 9240 26376 9240 0 _0935_
rlabel metal2 27048 13328 27048 13328 0 _0936_
rlabel metal2 26656 14504 26656 14504 0 _0937_
rlabel metal3 26096 14280 26096 14280 0 _0938_
rlabel metal2 25816 16576 25816 16576 0 _0939_
rlabel metal3 28392 17528 28392 17528 0 _0940_
rlabel metal2 26040 19376 26040 19376 0 _0941_
rlabel metal2 25592 19152 25592 19152 0 _0942_
rlabel metal2 24472 18256 24472 18256 0 _0943_
rlabel metal2 23800 17136 23800 17136 0 _0944_
rlabel metal2 22792 8960 22792 8960 0 _0945_
rlabel metal2 19096 13440 19096 13440 0 _0946_
rlabel metal2 22344 13272 22344 13272 0 _0947_
rlabel metal2 22624 14504 22624 14504 0 _0948_
rlabel metal3 23240 15624 23240 15624 0 _0949_
rlabel metal2 24472 16800 24472 16800 0 _0950_
rlabel metal2 24808 17976 24808 17976 0 _0951_
rlabel metal2 11536 13944 11536 13944 0 _0952_
rlabel metal2 11032 18144 11032 18144 0 _0953_
rlabel metal2 10976 20776 10976 20776 0 _0954_
rlabel metal2 11368 20048 11368 20048 0 _0955_
rlabel metal3 11816 18424 11816 18424 0 _0956_
rlabel metal3 14056 18424 14056 18424 0 _0957_
rlabel metal2 14952 16520 14952 16520 0 _0958_
rlabel metal2 6384 17080 6384 17080 0 _0959_
rlabel metal2 8008 18592 8008 18592 0 _0960_
rlabel metal2 13944 18480 13944 18480 0 _0961_
rlabel metal2 14392 18704 14392 18704 0 _0962_
rlabel metal2 15400 18816 15400 18816 0 _0963_
rlabel metal4 14728 8036 14728 8036 0 _0964_
rlabel metal2 7672 21560 7672 21560 0 _0965_
rlabel metal2 7448 19936 7448 19936 0 _0966_
rlabel metal2 14392 20160 14392 20160 0 _0967_
rlabel metal2 14840 19656 14840 19656 0 _0968_
rlabel metal2 13832 21952 13832 21952 0 _0969_
rlabel metal2 6944 26824 6944 26824 0 _0970_
rlabel metal2 7392 21560 7392 21560 0 _0971_
rlabel metal2 14280 21672 14280 21672 0 _0972_
rlabel metal2 14672 19208 14672 19208 0 _0973_
rlabel metal2 15288 19656 15288 19656 0 _0974_
rlabel metal2 15960 20496 15960 20496 0 _0975_
rlabel metal2 22736 26488 22736 26488 0 _0976_
rlabel metal2 23800 37632 23800 37632 0 _0977_
rlabel metal3 19880 37968 19880 37968 0 _0978_
rlabel metal3 20720 37016 20720 37016 0 _0979_
rlabel metal2 13496 49700 13496 49700 0 _0980_
rlabel metal2 13832 49728 13832 49728 0 _0981_
rlabel metal2 14168 49336 14168 49336 0 _0982_
rlabel metal3 17472 47432 17472 47432 0 _0983_
rlabel metal2 22008 39508 22008 39508 0 _0984_
rlabel metal2 19096 36792 19096 36792 0 _0985_
rlabel metal2 16184 37520 16184 37520 0 _0986_
rlabel metal2 26264 35672 26264 35672 0 _0987_
rlabel metal2 30856 38724 30856 38724 0 _0988_
rlabel metal2 20216 32760 20216 32760 0 _0989_
rlabel metal2 21728 33320 21728 33320 0 _0990_
rlabel metal2 21336 42504 21336 42504 0 _0991_
rlabel metal2 26152 39368 26152 39368 0 _0992_
rlabel metal2 26152 40936 26152 40936 0 _0993_
rlabel metal2 22120 44856 22120 44856 0 _0994_
rlabel metal2 21560 44072 21560 44072 0 _0995_
rlabel metal2 19992 37800 19992 37800 0 _0996_
rlabel metal4 19544 37016 19544 37016 0 _0997_
rlabel metal2 16240 39368 16240 39368 0 _0998_
rlabel metal2 19656 40936 19656 40936 0 _0999_
rlabel metal3 20776 40264 20776 40264 0 _1000_
rlabel metal2 22344 47656 22344 47656 0 _1001_
rlabel metal2 15288 43904 15288 43904 0 _1002_
rlabel metal4 14280 40432 14280 40432 0 _1003_
rlabel metal2 15568 40600 15568 40600 0 _1004_
rlabel metal2 15960 39144 15960 39144 0 _1005_
rlabel metal3 26152 35784 26152 35784 0 _1006_
rlabel metal2 21280 30184 21280 30184 0 _1007_
rlabel metal2 24360 41216 24360 41216 0 _1008_
rlabel metal2 23744 41048 23744 41048 0 _1009_
rlabel metal2 19432 45696 19432 45696 0 _1010_
rlabel metal2 25928 40824 25928 40824 0 _1011_
rlabel metal2 17808 55496 17808 55496 0 _1012_
rlabel metal2 17864 54040 17864 54040 0 _1013_
rlabel metal2 16464 54600 16464 54600 0 _1014_
rlabel metal3 18424 54264 18424 54264 0 _1015_
rlabel metal2 17528 40992 17528 40992 0 _1016_
rlabel metal2 18032 41384 18032 41384 0 _1017_
rlabel metal2 19096 44296 19096 44296 0 _1018_
rlabel metal3 20832 43400 20832 43400 0 _1019_
rlabel metal3 26824 37408 26824 37408 0 _1020_
rlabel metal3 19600 40376 19600 40376 0 _1021_
rlabel metal2 26040 44968 26040 44968 0 _1022_
rlabel metal2 26376 44520 26376 44520 0 _1023_
rlabel metal2 15288 37968 15288 37968 0 _1024_
rlabel metal2 15176 39088 15176 39088 0 _1025_
rlabel metal2 15176 43456 15176 43456 0 _1026_
rlabel metal2 15456 41944 15456 41944 0 _1027_
rlabel metal2 15624 37576 15624 37576 0 _1028_
rlabel metal2 14616 37856 14616 37856 0 _1029_
rlabel metal2 14840 37352 14840 37352 0 _1030_
rlabel metal2 24360 49168 24360 49168 0 _1031_
rlabel metal2 20552 31864 20552 31864 0 _1032_
rlabel metal2 15736 36400 15736 36400 0 _1033_
rlabel metal2 17416 39200 17416 39200 0 _1034_
rlabel metal2 15960 36344 15960 36344 0 _1035_
rlabel metal3 15372 35560 15372 35560 0 _1036_
rlabel metal2 42952 54488 42952 54488 0 _1037_
rlabel metal2 34048 50456 34048 50456 0 _1038_
rlabel metal2 34664 51352 34664 51352 0 _1039_
rlabel metal2 36344 50960 36344 50960 0 _1040_
rlabel metal2 34888 51856 34888 51856 0 _1041_
rlabel metal2 34552 51856 34552 51856 0 _1042_
rlabel metal2 40824 51296 40824 51296 0 _1043_
rlabel metal2 39144 52696 39144 52696 0 _1044_
rlabel metal2 39480 53424 39480 53424 0 _1045_
rlabel metal2 38640 52248 38640 52248 0 _1046_
rlabel metal2 30744 53368 30744 53368 0 _1047_
rlabel metal3 28280 29400 28280 29400 0 _1048_
rlabel metal3 20720 39480 20720 39480 0 _1049_
rlabel metal3 21112 39368 21112 39368 0 _1050_
rlabel metal2 23016 39200 23016 39200 0 _1051_
rlabel metal2 21840 39032 21840 39032 0 _1052_
rlabel metal3 19544 38920 19544 38920 0 _1053_
rlabel metal2 19544 40320 19544 40320 0 _1054_
rlabel metal3 18872 38864 18872 38864 0 _1055_
rlabel metal2 20552 37184 20552 37184 0 _1056_
rlabel metal2 22120 26152 22120 26152 0 _1057_
rlabel metal2 25032 30576 25032 30576 0 _1058_
rlabel metal2 28112 25480 28112 25480 0 _1059_
rlabel metal2 16184 26096 16184 26096 0 _1060_
rlabel metal2 6552 24696 6552 24696 0 _1061_
rlabel metal2 24584 24192 24584 24192 0 _1062_
rlabel metal2 24472 25872 24472 25872 0 _1063_
rlabel metal2 23464 23688 23464 23688 0 _1064_
rlabel metal2 19208 23184 19208 23184 0 _1065_
rlabel metal2 23912 23016 23912 23016 0 _1066_
rlabel metal2 18872 25536 18872 25536 0 _1067_
rlabel metal2 23016 24472 23016 24472 0 _1068_
rlabel metal3 20832 23912 20832 23912 0 _1069_
rlabel metal2 18088 23464 18088 23464 0 _1070_
rlabel metal2 18760 24752 18760 24752 0 _1071_
rlabel metal2 18480 25368 18480 25368 0 _1072_
rlabel metal2 6048 24920 6048 24920 0 _1073_
rlabel metal2 30352 29512 30352 29512 0 _1074_
rlabel metal2 29624 26096 29624 26096 0 _1075_
rlabel metal2 29792 11480 29792 11480 0 _1076_
rlabel metal3 9520 26824 9520 26824 0 _1077_
rlabel metal2 7784 25200 7784 25200 0 _1078_
rlabel metal2 15176 17304 15176 17304 0 _1079_
rlabel metal2 16744 22960 16744 22960 0 _1080_
rlabel metal2 23016 21896 23016 21896 0 _1081_
rlabel metal2 23128 20888 23128 20888 0 _1082_
rlabel metal2 6216 19936 6216 19936 0 _1083_
rlabel metal3 4704 21000 4704 21000 0 _1084_
rlabel metal3 20384 22232 20384 22232 0 _1085_
rlabel metal3 17864 22120 17864 22120 0 _1086_
rlabel metal3 3976 19992 3976 19992 0 _1087_
rlabel metal2 19992 26208 19992 26208 0 _1088_
rlabel metal2 19880 24752 19880 24752 0 _1089_
rlabel metal2 18872 23576 18872 23576 0 _1090_
rlabel metal2 12936 24472 12936 24472 0 _1091_
rlabel metal2 24472 24640 24472 24640 0 _1092_
rlabel metal2 22456 23464 22456 23464 0 _1093_
rlabel metal2 23352 19544 23352 19544 0 _1094_
rlabel metal2 12488 24136 12488 24136 0 _1095_
rlabel metal2 13608 26292 13608 26292 0 _1096_
rlabel metal3 10248 26264 10248 26264 0 _1097_
rlabel metal2 26488 25424 26488 25424 0 _1098_
rlabel metal3 24584 23912 24584 23912 0 _1099_
rlabel metal2 15848 22904 15848 22904 0 _1100_
rlabel metal2 13608 22568 13608 22568 0 _1101_
rlabel metal2 13832 24108 13832 24108 0 _1102_
rlabel metal2 10808 22344 10808 22344 0 _1103_
rlabel metal2 16296 42448 16296 42448 0 _1104_
rlabel metal2 17976 42840 17976 42840 0 _1105_
rlabel metal2 18424 29736 18424 29736 0 _1106_
rlabel metal2 10360 29848 10360 29848 0 _1107_
rlabel metal2 10360 27832 10360 27832 0 _1108_
rlabel metal3 21000 20552 21000 20552 0 _1109_
rlabel metal3 20944 23016 20944 23016 0 _1110_
rlabel metal2 20328 22736 20328 22736 0 _1111_
rlabel metal2 20664 21056 20664 21056 0 _1112_
rlabel metal2 19208 20776 19208 20776 0 _1113_
rlabel metal2 17864 20720 17864 20720 0 _1114_
rlabel metal2 19208 19488 19208 19488 0 _1115_
rlabel metal2 13384 7924 13384 7924 0 _1116_
rlabel metal2 14056 7616 14056 7616 0 _1117_
rlabel metal2 13552 6664 13552 6664 0 _1118_
rlabel metal2 11480 7672 11480 7672 0 _1119_
rlabel metal2 10864 7448 10864 7448 0 _1120_
rlabel metal2 23800 15848 23800 15848 0 _1121_
rlabel metal2 18032 7560 18032 7560 0 _1122_
rlabel metal2 16800 5992 16800 5992 0 _1123_
rlabel metal3 17136 7448 17136 7448 0 _1124_
rlabel metal3 6944 23128 6944 23128 0 _1125_
rlabel metal3 4592 23352 4592 23352 0 _1126_
rlabel metal2 2856 23520 2856 23520 0 _1127_
rlabel metal2 50792 47320 50792 47320 0 _1128_
rlabel metal2 45864 52696 45864 52696 0 _1129_
rlabel metal2 23016 25816 23016 25816 0 _1130_
rlabel metal2 15176 15792 15176 15792 0 _1131_
rlabel metal2 17304 19376 17304 19376 0 _1132_
rlabel metal2 14280 12208 14280 12208 0 _1133_
rlabel metal2 13720 10696 13720 10696 0 _1134_
rlabel metal3 10192 9016 10192 9016 0 _1135_
rlabel metal2 6776 12040 6776 12040 0 _1136_
rlabel metal2 8120 12936 8120 12936 0 _1137_
rlabel metal2 7392 11592 7392 11592 0 _1138_
rlabel metal2 6104 13776 6104 13776 0 _1139_
rlabel metal2 6888 10080 6888 10080 0 _1140_
rlabel metal2 24584 20496 24584 20496 0 _1141_
rlabel metal2 7056 16072 7056 16072 0 _1142_
rlabel metal2 2184 15568 2184 15568 0 _1143_
rlabel metal3 5096 15512 5096 15512 0 _1144_
rlabel metal2 7112 18592 7112 18592 0 _1145_
rlabel metal2 2072 18144 2072 18144 0 _1146_
rlabel metal3 5040 18424 5040 18424 0 _1147_
rlabel metal2 18088 16968 18088 16968 0 _1148_
rlabel metal2 6216 13888 6216 13888 0 _1149_
rlabel metal3 4368 13160 4368 13160 0 _1150_
rlabel metal2 3752 12152 3752 12152 0 _1151_
rlabel metal2 20664 21784 20664 21784 0 _1152_
rlabel metal2 19488 18312 19488 18312 0 _1153_
rlabel metal2 19768 10640 19768 10640 0 _1154_
rlabel metal3 17136 10584 17136 10584 0 _1155_
rlabel metal2 19208 11032 19208 11032 0 _1156_
rlabel metal2 17976 39368 17976 39368 0 _1157_
rlabel metal2 17528 38668 17528 38668 0 _1158_
rlabel metal2 19880 40096 19880 40096 0 _1159_
rlabel metal3 18872 39704 18872 39704 0 _1160_
rlabel metal2 19264 32760 19264 32760 0 _1161_
rlabel metal2 27048 32480 27048 32480 0 _1162_
rlabel metal2 23240 34328 23240 34328 0 _1163_
rlabel metal3 24752 33096 24752 33096 0 _1164_
rlabel metal2 27496 32648 27496 32648 0 _1165_
rlabel metal2 52136 32928 52136 32928 0 _1166_
rlabel metal3 21896 31808 21896 31808 0 _1167_
rlabel metal2 17864 32368 17864 32368 0 _1168_
rlabel metal2 24192 32536 24192 32536 0 _1169_
rlabel metal2 23688 32312 23688 32312 0 _1170_
rlabel metal2 21672 30576 21672 30576 0 _1171_
rlabel metal2 16520 32032 16520 32032 0 _1172_
rlabel metal2 16968 33880 16968 33880 0 _1173_
rlabel metal3 17752 32592 17752 32592 0 _1174_
rlabel metal2 51352 49504 51352 49504 0 _1175_
rlabel metal2 45640 46704 45640 46704 0 _1176_
rlabel metal3 45920 46648 45920 46648 0 _1177_
rlabel metal2 45752 46088 45752 46088 0 _1178_
rlabel metal2 47096 48272 47096 48272 0 _1179_
rlabel metal2 48272 47544 48272 47544 0 _1180_
rlabel metal3 46816 48104 46816 48104 0 _1181_
rlabel metal2 47992 46704 47992 46704 0 _1182_
rlabel metal3 48496 46648 48496 46648 0 _1183_
rlabel metal3 46592 47432 46592 47432 0 _1184_
rlabel metal2 50456 46872 50456 46872 0 _1185_
rlabel metal2 49952 46648 49952 46648 0 _1186_
rlabel metal2 50568 47824 50568 47824 0 _1187_
rlabel metal3 49224 51464 49224 51464 0 _1188_
rlabel metal2 50456 48216 50456 48216 0 _1189_
rlabel metal2 49784 51632 49784 51632 0 _1190_
rlabel metal2 50120 51240 50120 51240 0 _1191_
rlabel metal2 50344 51632 50344 51632 0 _1192_
rlabel metal2 50904 52472 50904 52472 0 _1193_
rlabel metal2 49280 52808 49280 52808 0 _1194_
rlabel metal2 49784 50120 49784 50120 0 _1195_
rlabel metal2 49784 51016 49784 51016 0 _1196_
rlabel metal2 51184 49784 51184 49784 0 _1197_
rlabel metal2 34104 35280 34104 35280 0 _1198_
rlabel metal2 41384 44576 41384 44576 0 _1199_
rlabel metal2 34664 34888 34664 34888 0 _1200_
rlabel metal2 39368 33320 39368 33320 0 _1201_
rlabel metal2 38248 34384 38248 34384 0 _1202_
rlabel metal2 37352 32424 37352 32424 0 _1203_
rlabel metal2 36680 33936 36680 33936 0 _1204_
rlabel metal2 38024 38920 38024 38920 0 _1205_
rlabel metal2 36904 37856 36904 37856 0 _1206_
rlabel metal2 39200 35672 39200 35672 0 _1207_
rlabel metal3 37744 38920 37744 38920 0 _1208_
rlabel metal2 36456 37576 36456 37576 0 _1209_
rlabel metal2 38696 36456 38696 36456 0 _1210_
rlabel metal2 38584 37240 38584 37240 0 _1211_
rlabel metal2 38920 36736 38920 36736 0 _1212_
rlabel metal2 40376 37968 40376 37968 0 _1213_
rlabel metal3 39480 37240 39480 37240 0 _1214_
rlabel metal2 39256 37128 39256 37128 0 _1215_
rlabel metal2 41104 46760 41104 46760 0 _1216_
rlabel metal2 37688 37688 37688 37688 0 _1217_
rlabel metal2 37912 37352 37912 37352 0 _1218_
rlabel metal2 38024 37296 38024 37296 0 _1219_
rlabel metal3 39256 45080 39256 45080 0 _1220_
rlabel metal2 40040 43792 40040 43792 0 _1221_
rlabel metal2 40376 45304 40376 45304 0 _1222_
rlabel metal3 42112 44296 42112 44296 0 _1223_
rlabel metal2 39032 42784 39032 42784 0 _1224_
rlabel metal2 39704 43680 39704 43680 0 _1225_
rlabel metal3 39872 43624 39872 43624 0 _1226_
rlabel metal3 41440 44072 41440 44072 0 _1227_
rlabel metal2 42728 44240 42728 44240 0 _1228_
rlabel metal2 42392 39816 42392 39816 0 _1229_
rlabel metal2 44856 38080 44856 38080 0 _1230_
rlabel metal2 40600 31752 40600 31752 0 _1231_
rlabel metal2 50568 42896 50568 42896 0 _1232_
rlabel metal2 39928 41608 39928 41608 0 _1233_
rlabel metal3 40712 40936 40712 40936 0 _1234_
rlabel metal2 43288 39984 43288 39984 0 _1235_
rlabel metal2 40264 43904 40264 43904 0 _1236_
rlabel metal2 39984 42056 39984 42056 0 _1237_
rlabel metal2 40264 41720 40264 41720 0 _1238_
rlabel metal2 41160 31024 41160 31024 0 _1239_
rlabel metal2 41272 29288 41272 29288 0 _1240_
rlabel metal2 46536 29456 46536 29456 0 _1241_
rlabel metal2 52696 28168 52696 28168 0 _1242_
rlabel metal3 48944 23912 48944 23912 0 _1243_
rlabel metal2 48552 22176 48552 22176 0 _1244_
rlabel metal2 47992 28616 47992 28616 0 _1245_
rlabel metal2 53312 32088 53312 32088 0 _1246_
rlabel metal2 51128 31080 51128 31080 0 _1247_
rlabel metal2 46200 40264 46200 40264 0 _1248_
rlabel metal2 46984 35280 46984 35280 0 _1249_
rlabel metal2 50792 42616 50792 42616 0 _1250_
rlabel metal3 51016 34440 51016 34440 0 _1251_
rlabel metal2 51968 32536 51968 32536 0 _1252_
rlabel metal2 52248 32928 52248 32928 0 _1253_
rlabel metal2 53368 34104 53368 34104 0 _1254_
rlabel metal2 53256 35448 53256 35448 0 _1255_
rlabel metal2 47096 33264 47096 33264 0 _1256_
rlabel metal2 46872 31304 46872 31304 0 _1257_
rlabel metal2 53256 27216 53256 27216 0 _1258_
rlabel metal2 51016 28784 51016 28784 0 _1259_
rlabel metal2 46760 28840 46760 28840 0 _1260_
rlabel metal2 46368 28056 46368 28056 0 _1261_
rlabel metal2 46984 30016 46984 30016 0 _1262_
rlabel metal2 45752 30352 45752 30352 0 _1263_
rlabel metal2 41944 33152 41944 33152 0 _1264_
rlabel metal2 46088 33264 46088 33264 0 _1265_
rlabel metal2 45080 33488 45080 33488 0 _1266_
rlabel via2 50680 27496 50680 27496 0 _1267_
rlabel metal2 45752 32648 45752 32648 0 _1268_
rlabel metal2 45416 32928 45416 32928 0 _1269_
rlabel metal2 46424 31472 46424 31472 0 _1270_
rlabel metal2 37576 31920 37576 31920 0 _1271_
rlabel metal3 35784 29400 35784 29400 0 _1272_
rlabel metal2 39816 20776 39816 20776 0 _1273_
rlabel metal2 39088 25032 39088 25032 0 _1274_
rlabel metal2 39480 29120 39480 29120 0 _1275_
rlabel metal2 45416 30576 45416 30576 0 _1276_
rlabel metal2 51240 35336 51240 35336 0 _1277_
rlabel metal2 49560 22456 49560 22456 0 _1278_
rlabel metal3 41776 39480 41776 39480 0 _1279_
rlabel metal3 41832 42504 41832 42504 0 _1280_
rlabel metal2 40264 43008 40264 43008 0 _1281_
rlabel metal2 40600 43120 40600 43120 0 _1282_
rlabel metal2 41944 43008 41944 43008 0 _1283_
rlabel metal2 42840 40544 42840 40544 0 _1284_
rlabel metal2 43736 39200 43736 39200 0 _1285_
rlabel metal2 45416 37968 45416 37968 0 _1286_
rlabel metal2 13160 13440 13160 13440 0 clknet_0_wb_clk_i
rlabel metal3 5936 12152 5936 12152 0 clknet_4_0_0_wb_clk_i
rlabel metal2 52360 26992 52360 26992 0 clknet_4_10_0_wb_clk_i
rlabel metal3 52136 40376 52136 40376 0 clknet_4_11_0_wb_clk_i
rlabel metal2 31808 41160 31808 41160 0 clknet_4_12_0_wb_clk_i
rlabel metal2 27720 54992 27720 54992 0 clknet_4_13_0_wb_clk_i
rlabel metal2 50568 48328 50568 48328 0 clknet_4_14_0_wb_clk_i
rlabel metal2 45416 54096 45416 54096 0 clknet_4_15_0_wb_clk_i
rlabel metal2 1848 20468 1848 20468 0 clknet_4_1_0_wb_clk_i
rlabel metal2 27272 5544 27272 5544 0 clknet_4_2_0_wb_clk_i
rlabel metal3 17864 18424 17864 18424 0 clknet_4_3_0_wb_clk_i
rlabel metal2 2296 25200 2296 25200 0 clknet_4_4_0_wb_clk_i
rlabel metal2 1848 54488 1848 54488 0 clknet_4_5_0_wb_clk_i
rlabel metal2 16016 34328 16016 34328 0 clknet_4_6_0_wb_clk_i
rlabel metal3 17920 49000 17920 49000 0 clknet_4_7_0_wb_clk_i
rlabel metal2 32312 12936 32312 12936 0 clknet_4_8_0_wb_clk_i
rlabel metal2 35784 25424 35784 25424 0 clknet_4_9_0_wb_clk_i
rlabel metal2 18984 56392 18984 56392 0 io_in[10]
rlabel metal2 20216 56616 20216 56616 0 io_in[11]
rlabel metal2 40936 54656 40936 54656 0 io_in[26]
rlabel metal2 15512 56336 15512 56336 0 io_in[8]
rlabel metal2 16072 56448 16072 56448 0 io_in[9]
rlabel metal2 22008 57610 22008 57610 0 io_out[12]
rlabel metal2 23912 55048 23912 55048 0 io_out[13]
rlabel metal3 23968 56280 23968 56280 0 io_out[14]
rlabel metal2 26432 54712 26432 54712 0 io_out[15]
rlabel metal2 27720 57400 27720 57400 0 io_out[16]
rlabel metal2 29400 56280 29400 56280 0 io_out[17]
rlabel metal3 30408 56280 30408 56280 0 io_out[18]
rlabel metal2 31416 57778 31416 57778 0 io_out[19]
rlabel metal2 34216 56504 34216 56504 0 io_out[20]
rlabel metal2 36456 56448 36456 56448 0 io_out[21]
rlabel metal2 38024 56504 38024 56504 0 io_out[22]
rlabel metal2 37464 55412 37464 55412 0 io_out[23]
rlabel metal2 40376 56280 40376 56280 0 io_out[24]
rlabel metal2 42056 56448 42056 56448 0 io_out[25]
rlabel metal2 18312 54208 18312 54208 0 net1
rlabel metal2 27272 53480 27272 53480 0 net10
rlabel metal2 29288 52360 29288 52360 0 net11
rlabel metal2 28616 55412 28616 55412 0 net12
rlabel metal2 31192 54152 31192 54152 0 net13
rlabel metal2 32088 55412 32088 55412 0 net14
rlabel metal2 33432 53844 33432 53844 0 net15
rlabel metal3 35056 55832 35056 55832 0 net16
rlabel metal3 36680 56056 36680 56056 0 net17
rlabel metal2 38136 54824 38136 54824 0 net18
rlabel metal2 39368 55412 39368 55412 0 net19
rlabel metal3 19376 55384 19376 55384 0 net2
rlabel metal2 42504 55216 42504 55216 0 net20
rlabel metal2 21784 56168 21784 56168 0 net21
rlabel metal2 22960 54712 22960 54712 0 net22
rlabel metal2 25032 55104 25032 55104 0 net23
rlabel metal2 25592 56994 25592 56994 0 net24
rlabel metal2 27160 54516 27160 54516 0 net25
rlabel metal3 28728 54712 28728 54712 0 net26
rlabel metal2 29736 56392 29736 56392 0 net27
rlabel metal2 31192 55076 31192 55076 0 net28
rlabel metal2 32424 55300 32424 55300 0 net29
rlabel metal3 41608 53032 41608 53032 0 net3
rlabel metal3 34496 56280 34496 56280 0 net30
rlabel metal3 35560 55160 35560 55160 0 net31
rlabel metal3 37744 56280 37744 56280 0 net32
rlabel metal2 38584 55300 38584 55300 0 net33
rlabel metal2 39256 55076 39256 55076 0 net34
rlabel metal2 6216 57008 6216 57008 0 net35
rlabel metal2 7336 56280 7336 56280 0 net36
rlabel metal2 8624 56280 8624 56280 0 net37
rlabel metal2 10024 56280 10024 56280 0 net38
rlabel metal2 11368 56280 11368 56280 0 net39
rlabel metal3 16688 56168 16688 56168 0 net4
rlabel metal2 13160 56672 13160 56672 0 net40
rlabel metal2 14000 56280 14000 56280 0 net41
rlabel metal2 15288 57778 15288 57778 0 net42
rlabel metal2 16408 55496 16408 55496 0 net43
rlabel metal2 17192 56448 17192 56448 0 net44
rlabel metal2 19376 56280 19376 56280 0 net45
rlabel metal2 20720 56280 20720 56280 0 net46
rlabel metal2 41608 55076 41608 55076 0 net47
rlabel metal2 42168 57778 42168 57778 0 net48
rlabel metal2 43960 55272 43960 55272 0 net49
rlabel metal3 16576 55160 16576 55160 0 net5
rlabel metal2 45360 56280 45360 56280 0 net50
rlabel metal2 46312 56280 46312 56280 0 net51
rlabel metal2 47880 57008 47880 57008 0 net52
rlabel metal2 49000 56280 49000 56280 0 net53
rlabel metal2 50344 56280 50344 56280 0 net54
rlabel metal2 51688 56280 51688 56280 0 net55
rlabel metal2 53032 56280 53032 56280 0 net56
rlabel metal2 55048 56560 55048 56560 0 net57
rlabel metal2 55944 56784 55944 56784 0 net58
rlabel metal2 4984 56392 4984 56392 0 net59
rlabel metal3 9968 40600 9968 40600 0 net6
rlabel metal2 6888 55944 6888 55944 0 net60
rlabel metal2 8176 55944 8176 55944 0 net61
rlabel metal2 9576 55944 9576 55944 0 net62
rlabel metal2 10920 55944 10920 55944 0 net63
rlabel metal2 12264 55944 12264 55944 0 net64
rlabel metal2 13552 55944 13552 55944 0 net65
rlabel metal2 14728 55944 14728 55944 0 net66
rlabel metal2 16072 55496 16072 55496 0 net67
rlabel metal2 19432 55776 19432 55776 0 net68
rlabel metal3 18592 55832 18592 55832 0 net69
rlabel metal2 24584 51576 24584 51576 0 net7
rlabel metal2 20440 56448 20440 56448 0 net70
rlabel metal2 42952 56392 42952 56392 0 net71
rlabel metal2 43624 56504 43624 56504 0 net72
rlabel metal2 43064 57610 43064 57610 0 net73
rlabel metal2 44968 56280 44968 56280 0 net74
rlabel metal2 45864 55944 45864 55944 0 net75
rlabel metal2 47264 55944 47264 55944 0 net76
rlabel metal2 48552 55944 48552 55944 0 net77
rlabel metal2 49896 55944 49896 55944 0 net78
rlabel metal2 51240 55944 51240 55944 0 net79
rlabel metal3 24136 54488 24136 54488 0 net8
rlabel metal2 52584 55944 52584 55944 0 net80
rlabel metal2 53928 55944 53928 55944 0 net81
rlabel metal2 55384 56056 55384 56056 0 net82
rlabel metal2 24080 56056 24080 56056 0 net9
rlabel metal2 11200 41944 11200 41944 0 simon1.millis_counter\[0\]
rlabel metal2 13048 43176 13048 43176 0 simon1.millis_counter\[1\]
rlabel metal3 16632 48944 16632 48944 0 simon1.millis_counter\[2\]
rlabel metal2 15176 48664 15176 48664 0 simon1.millis_counter\[3\]
rlabel metal3 11592 50344 11592 50344 0 simon1.millis_counter\[4\]
rlabel metal2 12936 50428 12936 50428 0 simon1.millis_counter\[5\]
rlabel metal2 12936 53760 12936 53760 0 simon1.millis_counter\[6\]
rlabel metal2 16184 50064 16184 50064 0 simon1.millis_counter\[7\]
rlabel metal2 19992 49560 19992 49560 0 simon1.millis_counter\[8\]
rlabel metal2 19208 51632 19208 51632 0 simon1.millis_counter\[9\]
rlabel metal2 29568 30072 29568 30072 0 simon1.next_random\[0\]
rlabel metal3 29848 29512 29848 29512 0 simon1.next_random\[1\]
rlabel metal2 35112 33320 35112 33320 0 simon1.play1.freq\[0\]
rlabel metal2 31528 34216 31528 34216 0 simon1.play1.freq\[1\]
rlabel metal3 33768 39032 33768 39032 0 simon1.play1.freq\[2\]
rlabel metal2 36064 36456 36064 36456 0 simon1.play1.freq\[3\]
rlabel metal2 38360 45584 38360 45584 0 simon1.play1.freq\[4\]
rlabel metal2 39480 44184 39480 44184 0 simon1.play1.freq\[5\]
rlabel metal2 39928 39648 39928 39648 0 simon1.play1.freq\[6\]
rlabel metal2 38808 40656 38808 40656 0 simon1.play1.freq\[7\]
rlabel metal2 47432 42392 47432 42392 0 simon1.play1.freq\[8\]
rlabel metal3 53088 40936 53088 40936 0 simon1.play1.freq\[9\]
rlabel metal2 36008 33656 36008 33656 0 simon1.play1.tick_counter\[0\]
rlabel metal2 51352 35672 51352 35672 0 simon1.play1.tick_counter\[10\]
rlabel metal2 51744 38024 51744 38024 0 simon1.play1.tick_counter\[11\]
rlabel metal2 54712 32928 54712 32928 0 simon1.play1.tick_counter\[12\]
rlabel metal2 55272 34664 55272 34664 0 simon1.play1.tick_counter\[13\]
rlabel metal3 53480 30968 53480 30968 0 simon1.play1.tick_counter\[14\]
rlabel metal2 52696 31808 52696 31808 0 simon1.play1.tick_counter\[15\]
rlabel metal3 54152 29400 54152 29400 0 simon1.play1.tick_counter\[16\]
rlabel metal2 57064 27496 57064 27496 0 simon1.play1.tick_counter\[17\]
rlabel metal3 52360 27832 52360 27832 0 simon1.play1.tick_counter\[18\]
rlabel metal2 52024 25536 52024 25536 0 simon1.play1.tick_counter\[19\]
rlabel metal2 40376 33768 40376 33768 0 simon1.play1.tick_counter\[1\]
rlabel metal2 47656 24192 47656 24192 0 simon1.play1.tick_counter\[20\]
rlabel metal2 48888 22792 48888 22792 0 simon1.play1.tick_counter\[21\]
rlabel metal2 46536 25368 46536 25368 0 simon1.play1.tick_counter\[22\]
rlabel metal3 45304 25480 45304 25480 0 simon1.play1.tick_counter\[23\]
rlabel metal3 41496 20104 41496 20104 0 simon1.play1.tick_counter\[24\]
rlabel metal2 40600 25312 40600 25312 0 simon1.play1.tick_counter\[25\]
rlabel metal2 39312 21784 39312 21784 0 simon1.play1.tick_counter\[26\]
rlabel metal2 38752 28504 38752 28504 0 simon1.play1.tick_counter\[27\]
rlabel metal2 32928 25592 32928 25592 0 simon1.play1.tick_counter\[28\]
rlabel metal2 34216 27272 34216 27272 0 simon1.play1.tick_counter\[29\]
rlabel metal3 41608 35000 41608 35000 0 simon1.play1.tick_counter\[2\]
rlabel metal3 36792 30184 36792 30184 0 simon1.play1.tick_counter\[30\]
rlabel metal2 39816 31248 39816 31248 0 simon1.play1.tick_counter\[31\]
rlabel metal2 42616 36736 42616 36736 0 simon1.play1.tick_counter\[3\]
rlabel metal3 41664 43288 41664 43288 0 simon1.play1.tick_counter\[4\]
rlabel metal2 44408 42504 44408 42504 0 simon1.play1.tick_counter\[5\]
rlabel metal3 42560 38024 42560 38024 0 simon1.play1.tick_counter\[6\]
rlabel metal2 45192 40936 45192 40936 0 simon1.play1.tick_counter\[7\]
rlabel metal3 49504 42728 49504 42728 0 simon1.play1.tick_counter\[8\]
rlabel metal2 51352 40320 51352 40320 0 simon1.play1.tick_counter\[9\]
rlabel metal2 47768 52976 47768 52976 0 simon1.score1.active_digit
rlabel metal2 48888 50484 48888 50484 0 simon1.score1.ena
rlabel metal3 41608 46536 41608 46536 0 simon1.score1.inc
rlabel metal2 44296 48216 44296 48216 0 simon1.score1.ones\[0\]
rlabel metal2 47208 51408 47208 51408 0 simon1.score1.ones\[1\]
rlabel metal2 46760 51268 46760 51268 0 simon1.score1.ones\[2\]
rlabel metal2 52472 45136 52472 45136 0 simon1.score1.ones\[3\]
rlabel metal2 50904 48944 50904 48944 0 simon1.score1.tens\[0\]
rlabel metal3 45472 52136 45472 52136 0 simon1.score1.tens\[1\]
rlabel metal2 50120 53368 50120 53368 0 simon1.score1.tens\[2\]
rlabel metal2 52024 50624 52024 50624 0 simon1.score1.tens\[3\]
rlabel metal2 30408 37072 30408 37072 0 simon1.score_rst
rlabel metal2 11256 21056 11256 21056 0 simon1.seq\[0\]\[0\]
rlabel metal2 11200 21672 11200 21672 0 simon1.seq\[0\]\[1\]
rlabel metal2 16408 23744 16408 23744 0 simon1.seq\[10\]\[0\]
rlabel metal3 12152 22568 12152 22568 0 simon1.seq\[10\]\[1\]
rlabel metal2 14504 24248 14504 24248 0 simon1.seq\[11\]\[0\]
rlabel metal2 12376 25032 12376 25032 0 simon1.seq\[11\]\[1\]
rlabel metal2 6104 20440 6104 20440 0 simon1.seq\[12\]\[0\]
rlabel metal2 5432 20160 5432 20160 0 simon1.seq\[12\]\[1\]
rlabel metal2 7280 24808 7280 24808 0 simon1.seq\[13\]\[0\]
rlabel metal2 8904 24416 8904 24416 0 simon1.seq\[13\]\[1\]
rlabel metal3 16800 6552 16800 6552 0 simon1.seq\[14\]\[0\]
rlabel metal2 18536 8736 18536 8736 0 simon1.seq\[14\]\[1\]
rlabel metal2 15064 6496 15064 6496 0 simon1.seq\[15\]\[0\]
rlabel metal2 12264 7168 12264 7168 0 simon1.seq\[15\]\[1\]
rlabel metal2 19768 20720 19768 20720 0 simon1.seq\[16\]\[0\]
rlabel metal2 21672 18256 21672 18256 0 simon1.seq\[16\]\[1\]
rlabel metal2 25704 22512 25704 22512 0 simon1.seq\[17\]\[0\]
rlabel metal3 29064 22456 29064 22456 0 simon1.seq\[17\]\[1\]
rlabel metal2 33544 21168 33544 21168 0 simon1.seq\[18\]\[0\]
rlabel metal2 37464 19376 37464 19376 0 simon1.seq\[18\]\[1\]
rlabel metal2 33432 17360 33432 17360 0 simon1.seq\[19\]\[0\]
rlabel metal2 36008 14392 36008 14392 0 simon1.seq\[19\]\[1\]
rlabel metal2 11424 16184 11424 16184 0 simon1.seq\[1\]\[0\]
rlabel metal2 9800 14784 9800 14784 0 simon1.seq\[1\]\[1\]
rlabel metal2 18984 13440 18984 13440 0 simon1.seq\[20\]\[0\]
rlabel metal3 22344 13160 22344 13160 0 simon1.seq\[20\]\[1\]
rlabel metal2 18536 12152 18536 12152 0 simon1.seq\[21\]\[0\]
rlabel metal2 20328 10976 20328 10976 0 simon1.seq\[21\]\[1\]
rlabel metal2 22008 6440 22008 6440 0 simon1.seq\[22\]\[0\]
rlabel metal2 24976 5208 24976 5208 0 simon1.seq\[22\]\[1\]
rlabel via2 22344 8344 22344 8344 0 simon1.seq\[23\]\[0\]
rlabel metal2 24360 9520 24360 9520 0 simon1.seq\[23\]\[1\]
rlabel metal2 27160 20440 27160 20440 0 simon1.seq\[24\]\[0\]
rlabel metal2 29624 19656 29624 19656 0 simon1.seq\[24\]\[1\]
rlabel via2 27272 9912 27272 9912 0 simon1.seq\[25\]\[0\]
rlabel metal3 29400 9912 29400 9912 0 simon1.seq\[25\]\[1\]
rlabel metal2 29624 16352 29624 16352 0 simon1.seq\[26\]\[0\]
rlabel metal2 31080 14616 31080 14616 0 simon1.seq\[26\]\[1\]
rlabel metal2 20328 16520 20328 16520 0 simon1.seq\[27\]\[0\]
rlabel metal3 24808 15176 24808 15176 0 simon1.seq\[27\]\[1\]
rlabel metal2 29176 12656 29176 12656 0 simon1.seq\[28\]\[0\]
rlabel metal2 32088 10304 32088 10304 0 simon1.seq\[28\]\[1\]
rlabel metal2 27496 6832 27496 6832 0 simon1.seq\[29\]\[0\]
rlabel metal2 29288 6552 29288 6552 0 simon1.seq\[29\]\[1\]
rlabel metal2 13048 13384 13048 13384 0 simon1.seq\[2\]\[0\]
rlabel metal2 11592 12208 11592 12208 0 simon1.seq\[2\]\[1\]
rlabel metal2 34216 12544 34216 12544 0 simon1.seq\[30\]\[0\]
rlabel metal2 36344 12208 36344 12208 0 simon1.seq\[30\]\[1\]
rlabel metal2 34104 19040 34104 19040 0 simon1.seq\[31\]\[0\]
rlabel metal2 36120 13720 36120 13720 0 simon1.seq\[31\]\[1\]
rlabel metal3 5376 13048 5376 13048 0 simon1.seq\[3\]\[0\]
rlabel metal2 5432 13384 5432 13384 0 simon1.seq\[3\]\[1\]
rlabel metal3 6440 17864 6440 17864 0 simon1.seq\[4\]\[0\]
rlabel metal2 6328 18760 6328 18760 0 simon1.seq\[4\]\[1\]
rlabel metal2 4760 14616 4760 14616 0 simon1.seq\[5\]\[0\]
rlabel metal2 6440 16072 6440 16072 0 simon1.seq\[5\]\[1\]
rlabel metal2 7672 11760 7672 11760 0 simon1.seq\[6\]\[0\]
rlabel metal2 7448 9632 7448 9632 0 simon1.seq\[6\]\[1\]
rlabel metal2 14728 11312 14728 11312 0 simon1.seq\[7\]\[0\]
rlabel metal3 11648 9912 11648 9912 0 simon1.seq\[7\]\[1\]
rlabel metal2 5768 22736 5768 22736 0 simon1.seq\[8\]\[0\]
rlabel metal2 6104 22736 6104 22736 0 simon1.seq\[8\]\[1\]
rlabel metal3 6720 27720 6720 27720 0 simon1.seq\[9\]\[0\]
rlabel metal2 7560 28280 7560 28280 0 simon1.seq\[9\]\[1\]
rlabel metal3 24304 30968 24304 30968 0 simon1.seq_counter\[0\]
rlabel via2 24920 32536 24920 32536 0 simon1.seq_counter\[1\]
rlabel metal2 23128 31416 23128 31416 0 simon1.seq_counter\[2\]
rlabel metal2 16408 31808 16408 31808 0 simon1.seq_counter\[3\]
rlabel metal2 16408 33096 16408 33096 0 simon1.seq_counter\[4\]
rlabel metal2 25704 25032 25704 25032 0 simon1.seq_length\[0\]
rlabel via1 26600 27173 26600 27173 0 simon1.seq_length\[1\]
rlabel metal2 21560 26208 21560 26208 0 simon1.seq_length\[2\]
rlabel metal2 17976 24080 17976 24080 0 simon1.seq_length\[3\]
rlabel metal2 21448 25256 21448 25256 0 simon1.seq_length\[4\]
rlabel metal3 23128 38136 23128 38136 0 simon1.state\[0\]
rlabel metal3 15176 35672 15176 35672 0 simon1.state\[1\]
rlabel metal2 22232 39200 22232 39200 0 simon1.state\[2\]
rlabel metal2 18648 36848 18648 36848 0 simon1.state\[3\]
rlabel metal2 12376 39592 12376 39592 0 simon1.state\[4\]
rlabel metal3 20832 36456 20832 36456 0 simon1.state\[5\]
rlabel metal2 19432 38472 19432 38472 0 simon1.state\[6\]
rlabel metal2 19488 33992 19488 33992 0 simon1.state\[7\]
rlabel metal2 4648 53872 4648 53872 0 simon1.tick_counter\[0\]
rlabel metal2 5544 39648 5544 39648 0 simon1.tick_counter\[10\]
rlabel metal2 5544 41552 5544 41552 0 simon1.tick_counter\[11\]
rlabel metal2 4256 42840 4256 42840 0 simon1.tick_counter\[12\]
rlabel metal2 1960 44016 1960 44016 0 simon1.tick_counter\[13\]
rlabel metal2 2184 46704 2184 46704 0 simon1.tick_counter\[14\]
rlabel metal2 3080 45920 3080 45920 0 simon1.tick_counter\[15\]
rlabel metal2 3752 52416 3752 52416 0 simon1.tick_counter\[1\]
rlabel metal2 4760 52920 4760 52920 0 simon1.tick_counter\[2\]
rlabel metal2 7448 52864 7448 52864 0 simon1.tick_counter\[3\]
rlabel metal3 7056 52920 7056 52920 0 simon1.tick_counter\[4\]
rlabel metal2 5544 48552 5544 48552 0 simon1.tick_counter\[5\]
rlabel metal2 6104 48888 6104 48888 0 simon1.tick_counter\[6\]
rlabel metal2 7560 46536 7560 46536 0 simon1.tick_counter\[7\]
rlabel metal3 6496 38808 6496 38808 0 simon1.tick_counter\[8\]
rlabel metal2 2856 38920 2856 38920 0 simon1.tick_counter\[9\]
rlabel metal2 31976 50680 31976 50680 0 simon1.tone_sequence_counter\[0\]
rlabel metal2 30072 47880 30072 47880 0 simon1.tone_sequence_counter\[1\]
rlabel metal2 30856 48328 30856 48328 0 simon1.tone_sequence_counter\[2\]
rlabel metal2 24528 47432 24528 47432 0 simon1.user_input\[0\]
rlabel metal2 22736 47208 22736 47208 0 simon1.user_input\[1\]
rlabel metal2 9016 48104 9016 48104 0 wb_clk_i
rlabel metal2 4592 56280 4592 56280 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
