* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuD

* Black-box entry subcircuit for urish_simon_says abstract view
.subckt urish_simon_says io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vdd vss wb_clk_i wb_rst_i
.ends

* Black-box entry subcircuit for top_design_mux abstract view
.subckt top_design_mux diego_clk diego_ena diego_io_in[0] diego_io_in[10] diego_io_in[11]
+ diego_io_in[12] diego_io_in[13] diego_io_in[14] diego_io_in[15] diego_io_in[16]
+ diego_io_in[17] diego_io_in[18] diego_io_in[19] diego_io_in[1] diego_io_in[20] diego_io_in[21]
+ diego_io_in[22] diego_io_in[23] diego_io_in[24] diego_io_in[25] diego_io_in[26]
+ diego_io_in[27] diego_io_in[28] diego_io_in[29] diego_io_in[2] diego_io_in[30] diego_io_in[31]
+ diego_io_in[32] diego_io_in[33] diego_io_in[34] diego_io_in[35] diego_io_in[36]
+ diego_io_in[37] diego_io_in[3] diego_io_in[4] diego_io_in[5] diego_io_in[6] diego_io_in[7]
+ diego_io_in[8] diego_io_in[9] diego_io_oeb[0] diego_io_oeb[10] diego_io_oeb[11]
+ diego_io_oeb[12] diego_io_oeb[13] diego_io_oeb[14] diego_io_oeb[15] diego_io_oeb[16]
+ diego_io_oeb[17] diego_io_oeb[18] diego_io_oeb[19] diego_io_oeb[1] diego_io_oeb[20]
+ diego_io_oeb[21] diego_io_oeb[22] diego_io_oeb[23] diego_io_oeb[24] diego_io_oeb[25]
+ diego_io_oeb[26] diego_io_oeb[27] diego_io_oeb[28] diego_io_oeb[29] diego_io_oeb[2]
+ diego_io_oeb[30] diego_io_oeb[31] diego_io_oeb[3] diego_io_oeb[4] diego_io_oeb[5]
+ diego_io_oeb[6] diego_io_oeb[7] diego_io_oeb[8] diego_io_oeb[9] diego_io_out[0]
+ diego_io_out[10] diego_io_out[11] diego_io_out[12] diego_io_out[13] diego_io_out[14]
+ diego_io_out[15] diego_io_out[16] diego_io_out[17] diego_io_out[18] diego_io_out[19]
+ diego_io_out[1] diego_io_out[20] diego_io_out[21] diego_io_out[22] diego_io_out[23]
+ diego_io_out[24] diego_io_out[25] diego_io_out[26] diego_io_out[27] diego_io_out[28]
+ diego_io_out[29] diego_io_out[2] diego_io_out[30] diego_io_out[31] diego_io_out[3]
+ diego_io_out[4] diego_io_out[5] diego_io_out[6] diego_io_out[7] diego_io_out[8]
+ diego_io_out[9] diego_rst i_design_reset[0] i_design_reset[1] i_design_reset[2]
+ i_design_reset[3] i_design_reset[4] i_design_reset[5] i_design_reset[6] i_design_reset[7]
+ i_mux_auto_reset_enb i_mux_io5_reset_enb i_mux_sel[0] i_mux_sel[1] i_mux_sel[2]
+ i_mux_sel[3] i_mux_sys_reset_enb io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la_in[0] la_in[10] la_in[11] la_in[12] la_in[13] la_in[14] la_in[15]
+ la_in[1] la_in[2] la_in[3] la_in[4] la_in[5] la_in[6] la_in[7] la_in[8] la_in[9]
+ mux_conf_clk pawel_clk pawel_ena pawel_io_in[0] pawel_io_in[10] pawel_io_in[11]
+ pawel_io_in[12] pawel_io_in[13] pawel_io_in[14] pawel_io_in[15] pawel_io_in[16]
+ pawel_io_in[17] pawel_io_in[18] pawel_io_in[19] pawel_io_in[1] pawel_io_in[20] pawel_io_in[21]
+ pawel_io_in[22] pawel_io_in[23] pawel_io_in[24] pawel_io_in[25] pawel_io_in[26]
+ pawel_io_in[27] pawel_io_in[28] pawel_io_in[29] pawel_io_in[2] pawel_io_in[30] pawel_io_in[31]
+ pawel_io_in[32] pawel_io_in[33] pawel_io_in[34] pawel_io_in[35] pawel_io_in[36]
+ pawel_io_in[37] pawel_io_in[3] pawel_io_in[4] pawel_io_in[5] pawel_io_in[6] pawel_io_in[7]
+ pawel_io_in[8] pawel_io_in[9] pawel_io_oeb[0] pawel_io_oeb[10] pawel_io_oeb[11]
+ pawel_io_oeb[12] pawel_io_oeb[1] pawel_io_oeb[2] pawel_io_oeb[3] pawel_io_oeb[4]
+ pawel_io_oeb[5] pawel_io_oeb[6] pawel_io_oeb[7] pawel_io_oeb[8] pawel_io_oeb[9]
+ pawel_io_out[0] pawel_io_out[10] pawel_io_out[11] pawel_io_out[12] pawel_io_out[1]
+ pawel_io_out[2] pawel_io_out[3] pawel_io_out[4] pawel_io_out[5] pawel_io_out[6]
+ pawel_io_out[7] pawel_io_out[8] pawel_io_out[9] pawel_rst solos_clk solos_ena solos_gpio_ready
+ solos_io_in[0] solos_io_in[10] solos_io_in[11] solos_io_in[12] solos_io_in[13] solos_io_in[14]
+ solos_io_in[15] solos_io_in[16] solos_io_in[17] solos_io_in[18] solos_io_in[19]
+ solos_io_in[1] solos_io_in[20] solos_io_in[21] solos_io_in[22] solos_io_in[23] solos_io_in[24]
+ solos_io_in[25] solos_io_in[26] solos_io_in[27] solos_io_in[28] solos_io_in[29]
+ solos_io_in[2] solos_io_in[30] solos_io_in[31] solos_io_in[32] solos_io_in[33] solos_io_in[34]
+ solos_io_in[35] solos_io_in[36] solos_io_in[37] solos_io_in[3] solos_io_in[4] solos_io_in[5]
+ solos_io_in[6] solos_io_in[7] solos_io_in[8] solos_io_in[9] solos_io_out[0] solos_io_out[10]
+ solos_io_out[11] solos_io_out[12] solos_io_out[1] solos_io_out[2] solos_io_out[3]
+ solos_io_out[4] solos_io_out[5] solos_io_out[6] solos_io_out[7] solos_io_out[8]
+ solos_io_out[9] solos_rst trzf2_clk trzf2_ena trzf2_io_in[0] trzf2_io_in[10] trzf2_io_in[11]
+ trzf2_io_in[12] trzf2_io_in[13] trzf2_io_in[14] trzf2_io_in[15] trzf2_io_in[16]
+ trzf2_io_in[17] trzf2_io_in[18] trzf2_io_in[19] trzf2_io_in[1] trzf2_io_in[20] trzf2_io_in[21]
+ trzf2_io_in[22] trzf2_io_in[23] trzf2_io_in[24] trzf2_io_in[25] trzf2_io_in[26]
+ trzf2_io_in[27] trzf2_io_in[28] trzf2_io_in[29] trzf2_io_in[2] trzf2_io_in[30] trzf2_io_in[31]
+ trzf2_io_in[32] trzf2_io_in[33] trzf2_io_in[34] trzf2_io_in[35] trzf2_io_in[36]
+ trzf2_io_in[37] trzf2_io_in[3] trzf2_io_in[4] trzf2_io_in[5] trzf2_io_in[6] trzf2_io_in[7]
+ trzf2_io_in[8] trzf2_io_in[9] trzf2_la_in[0] trzf2_la_in[10] trzf2_la_in[11] trzf2_la_in[12]
+ trzf2_la_in[1] trzf2_la_in[2] trzf2_la_in[3] trzf2_la_in[4] trzf2_la_in[5] trzf2_la_in[6]
+ trzf2_la_in[7] trzf2_la_in[8] trzf2_la_in[9] trzf2_o_gpout[0] trzf2_o_gpout[1] trzf2_o_gpout[2]
+ trzf2_o_hsync trzf2_o_rgb[0] trzf2_o_rgb[1] trzf2_o_rgb[2] trzf2_o_rgb[3] trzf2_o_rgb[4]
+ trzf2_o_rgb[5] trzf2_o_tex_csb trzf2_o_tex_oeb0 trzf2_o_tex_out0 trzf2_o_tex_sclk
+ trzf2_o_vsync trzf2_rst trzf_clk trzf_ena trzf_io_in[0] trzf_io_in[10] trzf_io_in[11]
+ trzf_io_in[12] trzf_io_in[13] trzf_io_in[14] trzf_io_in[15] trzf_io_in[16] trzf_io_in[17]
+ trzf_io_in[18] trzf_io_in[19] trzf_io_in[1] trzf_io_in[20] trzf_io_in[21] trzf_io_in[22]
+ trzf_io_in[23] trzf_io_in[24] trzf_io_in[25] trzf_io_in[26] trzf_io_in[27] trzf_io_in[28]
+ trzf_io_in[29] trzf_io_in[2] trzf_io_in[30] trzf_io_in[31] trzf_io_in[32] trzf_io_in[33]
+ trzf_io_in[34] trzf_io_in[35] trzf_io_in[36] trzf_io_in[37] trzf_io_in[3] trzf_io_in[4]
+ trzf_io_in[5] trzf_io_in[6] trzf_io_in[7] trzf_io_in[8] trzf_io_in[9] trzf_la_in[0]
+ trzf_la_in[10] trzf_la_in[11] trzf_la_in[12] trzf_la_in[1] trzf_la_in[2] trzf_la_in[3]
+ trzf_la_in[4] trzf_la_in[5] trzf_la_in[6] trzf_la_in[7] trzf_la_in[8] trzf_la_in[9]
+ trzf_o_gpout[0] trzf_o_gpout[1] trzf_o_gpout[2] trzf_o_hsync trzf_o_rgb[0] trzf_o_rgb[1]
+ trzf_o_rgb[2] trzf_o_rgb[3] trzf_o_rgb[4] trzf_o_rgb[5] trzf_o_tex_csb trzf_o_tex_oeb0
+ trzf_o_tex_out0 trzf_o_tex_sclk trzf_o_vsync trzf_rst uri_clk uri_ena uri_io_in[0]
+ uri_io_in[10] uri_io_in[11] uri_io_in[12] uri_io_in[13] uri_io_in[14] uri_io_in[15]
+ uri_io_in[16] uri_io_in[17] uri_io_in[18] uri_io_in[19] uri_io_in[1] uri_io_in[20]
+ uri_io_in[21] uri_io_in[22] uri_io_in[23] uri_io_in[24] uri_io_in[25] uri_io_in[26]
+ uri_io_in[27] uri_io_in[28] uri_io_in[29] uri_io_in[2] uri_io_in[30] uri_io_in[31]
+ uri_io_in[32] uri_io_in[33] uri_io_in[34] uri_io_in[35] uri_io_in[36] uri_io_in[37]
+ uri_io_in[3] uri_io_in[4] uri_io_in[5] uri_io_in[6] uri_io_in[7] uri_io_in[8] uri_io_in[9]
+ uri_io_oeb[0] uri_io_oeb[10] uri_io_oeb[11] uri_io_oeb[12] uri_io_oeb[13] uri_io_oeb[14]
+ uri_io_oeb[15] uri_io_oeb[16] uri_io_oeb[17] uri_io_oeb[18] uri_io_oeb[1] uri_io_oeb[2]
+ uri_io_oeb[3] uri_io_oeb[4] uri_io_oeb[5] uri_io_oeb[6] uri_io_oeb[7] uri_io_oeb[8]
+ uri_io_oeb[9] uri_io_out[0] uri_io_out[10] uri_io_out[11] uri_io_out[12] uri_io_out[13]
+ uri_io_out[14] uri_io_out[15] uri_io_out[16] uri_io_out[17] uri_io_out[18] uri_io_out[1]
+ uri_io_out[2] uri_io_out[3] uri_io_out[4] uri_io_out[5] uri_io_out[6] uri_io_out[7]
+ uri_io_out[8] uri_io_out[9] uri_rst vdd vgasp_clk vgasp_io_in[0] vgasp_io_in[10]
+ vgasp_io_in[11] vgasp_io_in[12] vgasp_io_in[13] vgasp_io_in[14] vgasp_io_in[15]
+ vgasp_io_in[16] vgasp_io_in[17] vgasp_io_in[18] vgasp_io_in[19] vgasp_io_in[1] vgasp_io_in[20]
+ vgasp_io_in[21] vgasp_io_in[22] vgasp_io_in[23] vgasp_io_in[24] vgasp_io_in[25]
+ vgasp_io_in[26] vgasp_io_in[27] vgasp_io_in[28] vgasp_io_in[29] vgasp_io_in[2] vgasp_io_in[30]
+ vgasp_io_in[31] vgasp_io_in[32] vgasp_io_in[33] vgasp_io_in[34] vgasp_io_in[35]
+ vgasp_io_in[36] vgasp_io_in[37] vgasp_io_in[3] vgasp_io_in[4] vgasp_io_in[5] vgasp_io_in[6]
+ vgasp_io_in[7] vgasp_io_in[8] vgasp_io_in[9] vgasp_rst vgasp_uio_oe[0] vgasp_uio_oe[1]
+ vgasp_uio_oe[2] vgasp_uio_oe[3] vgasp_uio_oe[4] vgasp_uio_oe[5] vgasp_uio_oe[6]
+ vgasp_uio_oe[7] vgasp_uio_out[0] vgasp_uio_out[1] vgasp_uio_out[2] vgasp_uio_out[3]
+ vgasp_uio_out[4] vgasp_uio_out[5] vgasp_uio_out[6] vgasp_uio_out[7] vgasp_uo_out[0]
+ vgasp_uo_out[1] vgasp_uo_out[2] vgasp_uo_out[3] vgasp_uo_out[4] vgasp_uo_out[5]
+ vgasp_uo_out[6] vgasp_uo_out[7] vss wb_clk_i wb_rst_i
.ends

* Black-box entry subcircuit for top_raybox_zero_fsm abstract view
.subckt top_raybox_zero_fsm i_clk i_debug_map_overlay i_debug_trace_overlay i_debug_vec_overlay
+ i_gpout0_sel[0] i_gpout0_sel[1] i_gpout0_sel[2] i_gpout0_sel[3] i_gpout1_sel[0]
+ i_gpout1_sel[1] i_gpout1_sel[2] i_gpout1_sel[3] i_gpout2_sel[0] i_gpout2_sel[1]
+ i_gpout2_sel[2] i_gpout2_sel[3] i_mode[0] i_mode[1] i_mode[2] i_reg_csb i_reg_mosi
+ i_reg_outs_enb i_reg_sclk i_reset i_tex_in[0] i_tex_in[1] i_tex_in[2] i_tex_in[3]
+ i_vec_csb i_vec_mosi i_vec_sclk o_gpout[0] o_gpout[1] o_gpout[2] o_hsync o_rgb[0]
+ o_rgb[1] o_rgb[2] o_rgb[3] o_rgb[4] o_rgb[5] o_tex_csb o_tex_oeb0 o_tex_out0 o_tex_sclk
+ o_vsync vdd vss
.ends

* Black-box entry subcircuit for top_vga_spi_rom abstract view
.subckt top_vga_spi_rom clk rst ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5]
+ ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6]
+ uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6]
+ uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6]
+ uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] vdd vss
.ends

* Black-box entry subcircuit for wrapped_wb_hyperram abstract view
.subckt wrapped_wb_hyperram io_in[0] io_in[10] io_in[11] io_in[12] io_in[1] io_in[2]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6]
+ io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[1]
+ io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ rst_i vdd vss wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for user_proj_cpu abstract view
.subckt user_proj_cpu io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for top_solo_squash abstract view
.subckt top_solo_squash clk gpio_ready io_in[0] io_in[10] io_in[11] io_in[12] io_in[1]
+ io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] rst vdd vss
.ends

.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xurish_simon_says uri_io_in\[0\] uri_io_in\[10\] uri_io_in\[11\] uri_io_in\[12\] uri_io_in\[13\]
+ uri_io_in\[14\] uri_io_in\[15\] uri_io_in\[16\] uri_io_in\[17\] uri_io_in\[18\]
+ uri_io_in\[19\] uri_io_in\[1\] uri_io_in\[20\] uri_io_in\[21\] uri_io_in\[22\] uri_io_in\[23\]
+ uri_io_in\[24\] uri_io_in\[25\] uri_io_in\[26\] uri_io_in\[27\] uri_io_in\[28\]
+ uri_io_in\[29\] uri_io_in\[2\] uri_io_in\[30\] uri_io_in\[31\] uri_io_in\[32\] uri_io_in\[33\]
+ uri_io_in\[34\] uri_io_in\[35\] uri_io_in\[36\] uri_io_in\[37\] uri_io_in\[3\] uri_io_in\[4\]
+ uri_io_in\[5\] uri_io_in\[6\] uri_io_in\[7\] uri_io_in\[8\] uri_io_in\[9\] urish_simon_says/io_oeb[0]
+ uri_io_oeb\[10\] uri_io_oeb\[11\] uri_io_oeb\[12\] uri_io_oeb\[13\] uri_io_oeb\[14\]
+ uri_io_oeb\[15\] uri_io_oeb\[16\] uri_io_oeb\[17\] uri_io_oeb\[18\] uri_io_oeb\[19\]
+ urish_simon_says/io_oeb[1] uri_io_oeb\[20\] uri_io_oeb\[21\] uri_io_oeb\[22\] uri_io_oeb\[23\]
+ uri_io_oeb\[24\] uri_io_oeb\[25\] uri_io_oeb\[26\] urish_simon_says/io_oeb[27] urish_simon_says/io_oeb[28]
+ urish_simon_says/io_oeb[29] urish_simon_says/io_oeb[2] urish_simon_says/io_oeb[30]
+ urish_simon_says/io_oeb[31] urish_simon_says/io_oeb[32] urish_simon_says/io_oeb[33]
+ urish_simon_says/io_oeb[34] urish_simon_says/io_oeb[35] urish_simon_says/io_oeb[36]
+ urish_simon_says/io_oeb[37] urish_simon_says/io_oeb[3] urish_simon_says/io_oeb[4]
+ urish_simon_says/io_oeb[5] urish_simon_says/io_oeb[6] urish_simon_says/io_oeb[7]
+ uri_io_oeb\[8\] uri_io_oeb\[9\] urish_simon_says/io_out[0] uri_io_out\[10\] uri_io_out\[11\]
+ uri_io_out\[12\] uri_io_out\[13\] uri_io_out\[14\] uri_io_out\[15\] uri_io_out\[16\]
+ uri_io_out\[17\] uri_io_out\[18\] uri_io_out\[19\] urish_simon_says/io_out[1] uri_io_out\[20\]
+ uri_io_out\[21\] uri_io_out\[22\] uri_io_out\[23\] uri_io_out\[24\] uri_io_out\[25\]
+ uri_io_out\[26\] urish_simon_says/io_out[27] urish_simon_says/io_out[28] urish_simon_says/io_out[29]
+ urish_simon_says/io_out[2] urish_simon_says/io_out[30] urish_simon_says/io_out[31]
+ urish_simon_says/io_out[32] urish_simon_says/io_out[33] urish_simon_says/io_out[34]
+ urish_simon_says/io_out[35] urish_simon_says/io_out[36] urish_simon_says/io_out[37]
+ urish_simon_says/io_out[3] urish_simon_says/io_out[4] urish_simon_says/io_out[5]
+ urish_simon_says/io_out[6] urish_simon_says/io_out[7] uri_io_out\[8\] uri_io_out\[9\]
+ vdd vss uri_clk uri_rst urish_simon_says
Xtop_design_mux diego_clk top_design_mux/diego_ena top_design_mux/diego_io_in[0] diego_io_in_all38\[10\]
+ diego_io_in_all38\[11\] diego_io_in_all38\[12\] diego_io_in_all38\[13\] diego_io_in_all38\[14\]
+ diego_io_in_all38\[15\] diego_io_in_all38\[16\] diego_io_in_all38\[17\] diego_io_in_all38\[18\]
+ diego_io_in_all38\[19\] top_design_mux/diego_io_in[1] diego_io_in_all38\[20\] diego_io_in_all38\[21\]
+ diego_io_in_all38\[22\] diego_io_in_all38\[23\] diego_io_in_all38\[24\] diego_io_in_all38\[25\]
+ diego_io_in_all38\[26\] diego_io_in_all38\[27\] diego_io_in_all38\[28\] diego_io_in_all38\[29\]
+ top_design_mux/diego_io_in[2] diego_io_in_all38\[30\] diego_io_in_all38\[31\] diego_io_in_all38\[32\]
+ diego_io_in_all38\[33\] diego_io_in_all38\[34\] diego_io_in_all38\[35\] diego_io_in_all38\[36\]
+ diego_io_in_all38\[37\] top_design_mux/diego_io_in[3] top_design_mux/diego_io_in[4]
+ top_design_mux/diego_io_in[5] diego_io_in_all38\[6\] diego_io_in_all38\[7\] diego_io_in_all38\[8\]
+ diego_io_in_all38\[9\] diego_io_oeb\[0\] diego_io_oeb\[10\] diego_io_oeb\[11\] diego_io_oeb\[12\]
+ diego_io_oeb\[13\] diego_io_oeb\[14\] diego_io_oeb\[15\] diego_io_oeb\[16\] diego_io_oeb\[17\]
+ diego_io_oeb\[18\] diego_io_oeb\[19\] diego_io_oeb\[1\] diego_io_oeb\[20\] diego_io_oeb\[21\]
+ diego_io_oeb\[22\] diego_io_oeb\[23\] diego_io_oeb\[24\] diego_io_oeb\[25\] diego_io_oeb\[26\]
+ diego_io_oeb\[27\] diego_io_oeb\[28\] diego_io_oeb\[29\] diego_io_oeb\[2\] diego_io_oeb\[30\]
+ diego_io_oeb\[31\] diego_io_oeb\[3\] diego_io_oeb\[4\] diego_io_oeb\[5\] diego_io_oeb\[6\]
+ diego_io_oeb\[7\] diego_io_oeb\[8\] diego_io_oeb\[9\] diego_io_out\[0\] diego_io_out\[10\]
+ diego_io_out\[11\] diego_io_out\[12\] diego_io_out\[13\] diego_io_out\[14\] diego_io_out\[15\]
+ diego_io_out\[16\] diego_io_out\[17\] diego_io_out\[18\] diego_io_out\[19\] diego_io_out\[1\]
+ diego_io_out\[20\] diego_io_out\[21\] diego_io_out\[22\] diego_io_out\[23\] diego_io_out\[24\]
+ diego_io_out\[25\] diego_io_out\[26\] diego_io_out\[27\] diego_io_out\[28\] diego_io_out\[29\]
+ diego_io_out\[2\] diego_io_out\[30\] diego_io_out\[31\] diego_io_out\[3\] diego_io_out\[4\]
+ diego_io_out\[5\] diego_io_out\[6\] diego_io_out\[7\] diego_io_out\[8\] diego_io_out\[9\]
+ top_design_mux/diego_rst la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[54] la_data_in[48]
+ la_data_in[49] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] io_in[0]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ top_design_mux/io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] top_design_mux/io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] top_design_mux/io_out[2] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] top_design_mux/io_out[3]
+ top_design_mux/io_out[4] top_design_mux/io_out[5] top_design_mux/io_out[6] top_design_mux/io_out[7]
+ io_out[8] io_out[9] la_data_in[8] la_data_in[18] la_data_in[19] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[9] la_data_in[10] la_data_in[11] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[63]
+ top_design_mux/pawel_clk top_design_mux/pawel_ena top_design_mux/pawel_io_in[0]
+ top_design_mux/pawel_io_in[10] top_design_mux/pawel_io_in[11] top_design_mux/pawel_io_in[12]
+ top_design_mux/pawel_io_in[13] top_design_mux/pawel_io_in[14] top_design_mux/pawel_io_in[15]
+ top_design_mux/pawel_io_in[16] top_design_mux/pawel_io_in[17] top_design_mux/pawel_io_in[18]
+ top_design_mux/pawel_io_in[19] top_design_mux/pawel_io_in[1] top_design_mux/pawel_io_in[20]
+ top_design_mux/pawel_io_in[21] top_design_mux/pawel_io_in[22] top_design_mux/pawel_io_in[23]
+ top_design_mux/pawel_io_in[24] pawel_io_in_all38\[25\] pawel_io_in_all38\[26\] pawel_io_in_all38\[27\]
+ pawel_io_in_all38\[28\] pawel_io_in_all38\[29\] top_design_mux/pawel_io_in[2] pawel_io_in_all38\[30\]
+ pawel_io_in_all38\[31\] pawel_io_in_all38\[32\] pawel_io_in_all38\[33\] pawel_io_in_all38\[34\]
+ pawel_io_in_all38\[35\] pawel_io_in_all38\[36\] pawel_io_in_all38\[37\] top_design_mux/pawel_io_in[3]
+ top_design_mux/pawel_io_in[4] top_design_mux/pawel_io_in[5] top_design_mux/pawel_io_in[6]
+ top_design_mux/pawel_io_in[7] top_design_mux/pawel_io_in[8] top_design_mux/pawel_io_in[9]
+ pawel_io_oeb\[0\] pawel_io_oeb\[10\] pawel_io_oeb\[11\] pawel_io_oeb\[12\] pawel_io_oeb\[1\]
+ pawel_io_oeb\[2\] pawel_io_oeb\[3\] pawel_io_oeb\[4\] pawel_io_oeb\[5\] pawel_io_oeb\[6\]
+ pawel_io_oeb\[7\] pawel_io_oeb\[8\] pawel_io_oeb\[9\] pawel_io_out\[0\] pawel_io_out\[10\]
+ pawel_io_out\[11\] pawel_io_out\[12\] pawel_io_out\[1\] pawel_io_out\[2\] pawel_io_out\[3\]
+ pawel_io_out\[4\] pawel_io_out\[5\] pawel_io_out\[6\] pawel_io_out\[7\] pawel_io_out\[8\]
+ pawel_io_out\[9\] pawel_mux_rst solos_clk top_design_mux/solos_ena solos_gpio_ready
+ top_design_mux/solos_io_in[0] solos_io_in_all38\[10\] solos_io_in_all38\[11\] solos_io_in_all38\[12\]
+ solos_io_in_all38\[13\] solos_io_in_all38\[14\] solos_io_in_all38\[15\] solos_io_in_all38\[16\]
+ solos_io_in_all38\[17\] solos_io_in_all38\[18\] solos_io_in_all38\[19\] top_design_mux/solos_io_in[1]
+ solos_io_in_all38\[20\] top_design_mux/solos_io_in[21] top_design_mux/solos_io_in[22]
+ top_design_mux/solos_io_in[23] top_design_mux/solos_io_in[24] top_design_mux/solos_io_in[25]
+ top_design_mux/solos_io_in[26] top_design_mux/solos_io_in[27] top_design_mux/solos_io_in[28]
+ top_design_mux/solos_io_in[29] top_design_mux/solos_io_in[2] top_design_mux/solos_io_in[30]
+ top_design_mux/solos_io_in[31] top_design_mux/solos_io_in[32] top_design_mux/solos_io_in[33]
+ top_design_mux/solos_io_in[34] top_design_mux/solos_io_in[35] top_design_mux/solos_io_in[36]
+ top_design_mux/solos_io_in[37] top_design_mux/solos_io_in[3] top_design_mux/solos_io_in[4]
+ top_design_mux/solos_io_in[5] top_design_mux/solos_io_in[6] top_design_mux/solos_io_in[7]
+ solos_io_in_all38\[8\] solos_io_in_all38\[9\] solos_io_out\[0\] solos_io_out\[10\]
+ solos_io_out\[11\] solos_io_out\[12\] solos_io_out\[1\] solos_io_out\[2\] solos_io_out\[3\]
+ solos_io_out\[4\] solos_io_out\[5\] solos_io_out\[6\] solos_io_out\[7\] solos_io_out\[8\]
+ solos_io_out\[9\] solos_rst trzf2_clk top_design_mux/trzf2_ena top_design_mux/trzf2_io_in[0]
+ top_design_mux/trzf2_io_in[10] top_design_mux/trzf2_io_in[11] top_design_mux/trzf2_io_in[12]
+ top_design_mux/trzf2_io_in[13] top_design_mux/trzf2_io_in[14] top_design_mux/trzf2_io_in[15]
+ top_design_mux/trzf2_io_in[16] top_design_mux/trzf2_io_in[17] trzf2_io_in\[18\]
+ trzf2_io_in\[19\] top_design_mux/trzf2_io_in[1] trzf2_io_in\[20\] trzf2_io_in\[21\]
+ trzf2_io_in\[22\] trzf2_io_in\[23\] trzf2_io_in\[24\] trzf2_io_in\[25\] trzf2_io_in\[26\]
+ trzf2_io_in\[27\] trzf2_io_in\[28\] trzf2_io_in\[29\] top_design_mux/trzf2_io_in[2]
+ trzf2_io_in\[30\] trzf2_io_in\[31\] trzf2_io_in\[32\] trzf2_io_in\[33\] trzf2_io_in\[34\]
+ top_design_mux/trzf2_io_in[35] top_design_mux/trzf2_io_in[36] top_design_mux/trzf2_io_in[37]
+ top_design_mux/trzf2_io_in[3] top_design_mux/trzf2_io_in[4] top_design_mux/trzf2_io_in[5]
+ top_design_mux/trzf2_io_in[6] top_design_mux/trzf2_io_in[7] top_design_mux/trzf2_io_in[8]
+ top_design_mux/trzf2_io_in[9] top_design_mux/trzf2_la_in[0] trzf2_la_in\[10\] trzf2_la_in\[11\]
+ trzf2_la_in\[12\] trzf2_la_in\[1\] trzf2_la_in\[2\] trzf2_la_in\[3\] trzf2_la_in\[4\]
+ trzf2_la_in\[5\] trzf2_la_in\[6\] trzf2_la_in\[7\] trzf2_la_in\[8\] trzf2_la_in\[9\]
+ trzf2_o_gpout\[0\] trzf2_o_gpout\[1\] trzf2_o_gpout\[2\] trzf2_o_hsync trzf2_o_rgb\[0\]
+ trzf2_o_rgb\[1\] trzf2_o_rgb\[2\] trzf2_o_rgb\[3\] trzf2_o_rgb\[4\] trzf2_o_rgb\[5\]
+ trzf2_o_tex_csb trzf2_o_tex_oeb0 trzf2_o_tex_out0 trzf2_o_tex_sclk trzf2_o_vsync
+ trzf2_rst trzf_clk top_design_mux/trzf_ena top_design_mux/trzf_io_in[0] top_design_mux/trzf_io_in[10]
+ top_design_mux/trzf_io_in[11] top_design_mux/trzf_io_in[12] top_design_mux/trzf_io_in[13]
+ top_design_mux/trzf_io_in[14] top_design_mux/trzf_io_in[15] top_design_mux/trzf_io_in[16]
+ top_design_mux/trzf_io_in[17] trzf_io_in\[18\] trzf_io_in\[19\] top_design_mux/trzf_io_in[1]
+ trzf_io_in\[20\] trzf_io_in\[21\] trzf_io_in\[22\] trzf_io_in\[23\] trzf_io_in\[24\]
+ trzf_io_in\[25\] trzf_io_in\[26\] trzf_io_in\[27\] trzf_io_in\[28\] trzf_io_in\[29\]
+ top_design_mux/trzf_io_in[2] trzf_io_in\[30\] trzf_io_in\[31\] trzf_io_in\[32\]
+ trzf_io_in\[33\] trzf_io_in\[34\] top_design_mux/trzf_io_in[35] top_design_mux/trzf_io_in[36]
+ top_design_mux/trzf_io_in[37] top_design_mux/trzf_io_in[3] top_design_mux/trzf_io_in[4]
+ top_design_mux/trzf_io_in[5] top_design_mux/trzf_io_in[6] top_design_mux/trzf_io_in[7]
+ top_design_mux/trzf_io_in[8] top_design_mux/trzf_io_in[9] top_design_mux/trzf_la_in[0]
+ trzf_la_in\[10\] trzf_la_in\[11\] trzf_la_in\[12\] trzf_la_in\[1\] trzf_la_in\[2\]
+ trzf_la_in\[3\] trzf_la_in\[4\] trzf_la_in\[5\] trzf_la_in\[6\] trzf_la_in\[7\]
+ trzf_la_in\[8\] trzf_la_in\[9\] trzf_o_gpout\[0\] trzf_o_gpout\[1\] trzf_o_gpout\[2\]
+ trzf_o_hsync trzf_o_rgb\[0\] trzf_o_rgb\[1\] trzf_o_rgb\[2\] trzf_o_rgb\[3\] trzf_o_rgb\[4\]
+ trzf_o_rgb\[5\] trzf_o_tex_csb trzf_o_tex_oeb0 trzf_o_tex_out0 trzf_o_tex_sclk trzf_o_vsync
+ trzf_rst uri_clk top_design_mux/uri_ena uri_io_in\[0\] uri_io_in\[10\] uri_io_in\[11\]
+ uri_io_in\[12\] uri_io_in\[13\] uri_io_in\[14\] uri_io_in\[15\] uri_io_in\[16\]
+ uri_io_in\[17\] uri_io_in\[18\] uri_io_in\[19\] uri_io_in\[1\] uri_io_in\[20\] uri_io_in\[21\]
+ uri_io_in\[22\] uri_io_in\[23\] uri_io_in\[24\] uri_io_in\[25\] uri_io_in\[26\]
+ uri_io_in\[27\] uri_io_in\[28\] uri_io_in\[29\] uri_io_in\[2\] uri_io_in\[30\] uri_io_in\[31\]
+ uri_io_in\[32\] uri_io_in\[33\] uri_io_in\[34\] uri_io_in\[35\] uri_io_in\[36\]
+ uri_io_in\[37\] uri_io_in\[3\] uri_io_in\[4\] uri_io_in\[5\] uri_io_in\[6\] uri_io_in\[7\]
+ uri_io_in\[8\] uri_io_in\[9\] uri_io_oeb\[8\] uri_io_oeb\[18\] uri_io_oeb\[19\]
+ uri_io_oeb\[20\] uri_io_oeb\[21\] uri_io_oeb\[22\] uri_io_oeb\[23\] uri_io_oeb\[24\]
+ uri_io_oeb\[25\] uri_io_oeb\[26\] uri_io_oeb\[9\] uri_io_oeb\[10\] uri_io_oeb\[11\]
+ uri_io_oeb\[12\] uri_io_oeb\[13\] uri_io_oeb\[14\] uri_io_oeb\[15\] uri_io_oeb\[16\]
+ uri_io_oeb\[17\] uri_io_out\[8\] uri_io_out\[18\] uri_io_out\[19\] uri_io_out\[20\]
+ uri_io_out\[21\] uri_io_out\[22\] uri_io_out\[23\] uri_io_out\[24\] uri_io_out\[25\]
+ uri_io_out\[26\] uri_io_out\[9\] uri_io_out\[10\] uri_io_out\[11\] uri_io_out\[12\]
+ uri_io_out\[13\] uri_io_out\[14\] uri_io_out\[15\] uri_io_out\[16\] uri_io_out\[17\]
+ uri_rst vdd vgasp_clk top_design_mux/vgasp_io_in[0] top_design_mux/vgasp_io_in[10]
+ top_design_mux/vgasp_io_in[11] top_design_mux/vgasp_io_in[12] top_design_mux/vgasp_io_in[13]
+ top_design_mux/vgasp_io_in[14] top_design_mux/vgasp_io_in[15] top_design_mux/vgasp_io_in[16]
+ top_design_mux/vgasp_io_in[17] vgasp_io_in\[18\] vgasp_io_in\[19\] top_design_mux/vgasp_io_in[1]
+ vgasp_io_in\[20\] vgasp_io_in\[21\] vgasp_io_in\[22\] vgasp_io_in\[23\] vgasp_io_in\[24\]
+ vgasp_io_in\[25\] vgasp_io_in\[26\] vgasp_io_in\[27\] vgasp_io_in\[28\] vgasp_io_in\[29\]
+ top_design_mux/vgasp_io_in[2] vgasp_io_in\[30\] vgasp_io_in\[31\] vgasp_io_in\[32\]
+ top_design_mux/vgasp_io_in[33] top_design_mux/vgasp_io_in[34] top_design_mux/vgasp_io_in[35]
+ top_design_mux/vgasp_io_in[36] vgasp_io_in\[37\] top_design_mux/vgasp_io_in[3] top_design_mux/vgasp_io_in[4]
+ top_design_mux/vgasp_io_in[5] top_design_mux/vgasp_io_in[6] top_design_mux/vgasp_io_in[7]
+ top_design_mux/vgasp_io_in[8] top_design_mux/vgasp_io_in[9] vgasp_rst vgasp_uio_oe\[0\]
+ vgasp_uio_oe\[1\] vgasp_uio_oe\[2\] vgasp_uio_oe\[3\] vgasp_uio_oe\[4\] vgasp_uio_oe\[5\]
+ vgasp_uio_oe\[6\] vgasp_uio_oe\[7\] vgasp_uio_out\[0\] vgasp_uio_out\[1\] vgasp_uio_out\[2\]
+ vgasp_uio_out\[3\] vgasp_uio_out\[4\] vgasp_uio_out\[5\] vgasp_uio_out\[6\] vgasp_uio_out\[7\]
+ vgasp_uo_out\[0\] vgasp_uo_out\[1\] vgasp_uo_out\[2\] vgasp_uo_out\[3\] vgasp_uo_out\[4\]
+ vgasp_uo_out\[5\] vgasp_uo_out\[6\] vgasp_uo_out\[7\] vss wb_clk_i wb_rst_i top_design_mux
Xtop_raybox_zero_fsm trzf_clk trzf_io_in\[29\] trzf_io_in\[30\] trzf_io_in\[28\] trzf_la_in\[1\]
+ trzf_la_in\[2\] trzf_la_in\[3\] trzf_la_in\[4\] trzf_la_in\[5\] trzf_la_in\[6\]
+ trzf_la_in\[7\] trzf_la_in\[8\] trzf_la_in\[9\] trzf_la_in\[10\] trzf_la_in\[11\]
+ trzf_la_in\[12\] trzf_io_in\[32\] trzf_io_in\[33\] trzf_io_in\[34\] trzf_io_in\[25\]
+ trzf_io_in\[27\] trzf_io_in\[31\] trzf_io_in\[26\] trzf_rst trzf_io_in\[18\] trzf_io_in\[19\]
+ trzf_io_in\[20\] trzf_io_in\[21\] trzf_io_in\[22\] trzf_io_in\[24\] trzf_io_in\[23\]
+ trzf_o_gpout\[0\] trzf_o_gpout\[1\] trzf_o_gpout\[2\] trzf_o_hsync trzf_o_rgb\[0\]
+ trzf_o_rgb\[1\] trzf_o_rgb\[2\] trzf_o_rgb\[3\] trzf_o_rgb\[4\] trzf_o_rgb\[5\]
+ trzf_o_tex_csb trzf_o_tex_oeb0 trzf_o_tex_out0 trzf_o_tex_sclk trzf_o_vsync vdd
+ vss top_raybox_zero_fsm
Xtop_raybox_zero_fsm2 trzf2_clk trzf2_io_in\[29\] trzf2_io_in\[30\] trzf2_io_in\[28\]
+ trzf2_la_in\[1\] trzf2_la_in\[2\] trzf2_la_in\[3\] trzf2_la_in\[4\] trzf2_la_in\[5\]
+ trzf2_la_in\[6\] trzf2_la_in\[7\] trzf2_la_in\[8\] trzf2_la_in\[9\] trzf2_la_in\[10\]
+ trzf2_la_in\[11\] trzf2_la_in\[12\] trzf2_io_in\[32\] trzf2_io_in\[33\] trzf2_io_in\[34\]
+ trzf2_io_in\[25\] trzf2_io_in\[27\] trzf2_io_in\[31\] trzf2_io_in\[26\] trzf2_rst
+ trzf2_io_in\[18\] trzf2_io_in\[19\] trzf2_io_in\[20\] trzf2_io_in\[21\] trzf2_io_in\[22\]
+ trzf2_io_in\[24\] trzf2_io_in\[23\] trzf2_o_gpout\[0\] trzf2_o_gpout\[1\] trzf2_o_gpout\[2\]
+ trzf2_o_hsync trzf2_o_rgb\[0\] trzf2_o_rgb\[1\] trzf2_o_rgb\[2\] trzf2_o_rgb\[3\]
+ trzf2_o_rgb\[4\] trzf2_o_rgb\[5\] trzf2_o_tex_csb trzf2_o_tex_oeb0 trzf2_o_tex_out0
+ trzf2_o_tex_sclk trzf2_o_vsync vdd vss top_raybox_zero_fsm
Xtop_vga_spi_rom vgasp_clk vgasp_rst vgasp_io_in\[22\] vgasp_io_in\[23\] vgasp_io_in\[24\]
+ vgasp_io_in\[28\] vgasp_io_in\[29\] vgasp_io_in\[25\] vgasp_io_in\[26\] vgasp_io_in\[27\]
+ vgasp_io_in\[32\] vgasp_io_in\[18\] vgasp_io_in\[19\] vgasp_io_in\[30\] vgasp_io_in\[31\]
+ vgasp_io_in\[37\] vgasp_io_in\[20\] vgasp_io_in\[21\] vgasp_uio_oe\[0\] vgasp_uio_oe\[1\]
+ vgasp_uio_oe\[2\] vgasp_uio_oe\[3\] vgasp_uio_oe\[4\] vgasp_uio_oe\[5\] vgasp_uio_oe\[6\]
+ vgasp_uio_oe\[7\] vgasp_uio_out\[0\] vgasp_uio_out\[1\] vgasp_uio_out\[2\] vgasp_uio_out\[3\]
+ vgasp_uio_out\[4\] vgasp_uio_out\[5\] vgasp_uio_out\[6\] vgasp_uio_out\[7\] vgasp_uo_out\[0\]
+ vgasp_uo_out\[1\] vgasp_uo_out\[2\] vgasp_uo_out\[3\] vgasp_uo_out\[4\] vgasp_uo_out\[5\]
+ vgasp_uo_out\[6\] vgasp_uo_out\[7\] vdd vss top_vga_spi_rom
Xwrapped_wb_hyperram pawel_io_in_all38\[25\] pawel_io_in_all38\[35\] pawel_io_in_all38\[36\]
+ pawel_io_in_all38\[37\] pawel_io_in_all38\[26\] pawel_io_in_all38\[27\] pawel_io_in_all38\[28\]
+ pawel_io_in_all38\[29\] pawel_io_in_all38\[30\] pawel_io_in_all38\[31\] pawel_io_in_all38\[32\]
+ pawel_io_in_all38\[33\] pawel_io_in_all38\[34\] pawel_io_oeb\[0\] pawel_io_oeb\[10\]
+ pawel_io_oeb\[11\] pawel_io_oeb\[12\] pawel_io_oeb\[1\] pawel_io_oeb\[2\] pawel_io_oeb\[3\]
+ pawel_io_oeb\[4\] pawel_io_oeb\[5\] pawel_io_oeb\[6\] pawel_io_oeb\[7\] pawel_io_oeb\[8\]
+ pawel_io_oeb\[9\] pawel_io_out\[0\] pawel_io_out\[10\] pawel_io_out\[11\] pawel_io_out\[12\]
+ pawel_io_out\[1\] pawel_io_out\[2\] pawel_io_out\[3\] pawel_io_out\[4\] pawel_io_out\[5\]
+ pawel_io_out\[6\] pawel_io_out\[7\] pawel_io_out\[8\] pawel_io_out\[9\] pawel_mux_rst
+ vdd vss wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i wrapped_wb_hyperram
Xuser_proj_cpu diego_io_in_all38\[6\] diego_io_in_all38\[16\] diego_io_in_all38\[17\]
+ diego_io_in_all38\[18\] diego_io_in_all38\[19\] diego_io_in_all38\[20\] diego_io_in_all38\[21\]
+ diego_io_in_all38\[22\] diego_io_in_all38\[23\] diego_io_in_all38\[24\] diego_io_in_all38\[25\]
+ diego_io_in_all38\[7\] diego_io_in_all38\[26\] diego_io_in_all38\[27\] diego_io_in_all38\[28\]
+ diego_io_in_all38\[29\] diego_io_in_all38\[30\] diego_io_in_all38\[31\] diego_io_in_all38\[32\]
+ diego_io_in_all38\[33\] diego_io_in_all38\[34\] diego_io_in_all38\[35\] diego_io_in_all38\[8\]
+ diego_io_in_all38\[36\] diego_io_in_all38\[37\] diego_io_in_all38\[9\] diego_io_in_all38\[10\]
+ diego_io_in_all38\[11\] diego_io_in_all38\[12\] diego_io_in_all38\[13\] diego_io_in_all38\[14\]
+ diego_io_in_all38\[15\] diego_io_oeb\[0\] diego_io_oeb\[10\] diego_io_oeb\[11\]
+ diego_io_oeb\[12\] diego_io_oeb\[13\] diego_io_oeb\[14\] diego_io_oeb\[15\] diego_io_oeb\[16\]
+ diego_io_oeb\[17\] diego_io_oeb\[18\] diego_io_oeb\[19\] diego_io_oeb\[1\] diego_io_oeb\[20\]
+ diego_io_oeb\[21\] diego_io_oeb\[22\] diego_io_oeb\[23\] diego_io_oeb\[24\] diego_io_oeb\[25\]
+ diego_io_oeb\[26\] diego_io_oeb\[27\] diego_io_oeb\[28\] diego_io_oeb\[29\] diego_io_oeb\[2\]
+ diego_io_oeb\[30\] diego_io_oeb\[31\] diego_io_oeb\[3\] diego_io_oeb\[4\] diego_io_oeb\[5\]
+ diego_io_oeb\[6\] diego_io_oeb\[7\] diego_io_oeb\[8\] diego_io_oeb\[9\] diego_io_out\[0\]
+ diego_io_out\[10\] diego_io_out\[11\] diego_io_out\[12\] diego_io_out\[13\] diego_io_out\[14\]
+ diego_io_out\[15\] diego_io_out\[16\] diego_io_out\[17\] diego_io_out\[18\] diego_io_out\[19\]
+ diego_io_out\[1\] diego_io_out\[20\] diego_io_out\[21\] diego_io_out\[22\] diego_io_out\[23\]
+ diego_io_out\[24\] diego_io_out\[25\] diego_io_out\[26\] diego_io_out\[27\] diego_io_out\[28\]
+ diego_io_out\[29\] diego_io_out\[2\] diego_io_out\[30\] diego_io_out\[31\] diego_io_out\[3\]
+ diego_io_out\[4\] diego_io_out\[5\] diego_io_out\[6\] diego_io_out\[7\] diego_io_out\[8\]
+ diego_io_out\[9\] vdd vss diego_clk user_proj_cpu
Xtop_solo_squash solos_clk solos_gpio_ready solos_io_in_all38\[8\] solos_io_in_all38\[18\]
+ solos_io_in_all38\[19\] solos_io_in_all38\[20\] solos_io_in_all38\[9\] solos_io_in_all38\[10\]
+ solos_io_in_all38\[11\] solos_io_in_all38\[12\] solos_io_in_all38\[13\] solos_io_in_all38\[14\]
+ solos_io_in_all38\[15\] solos_io_in_all38\[16\] solos_io_in_all38\[17\] solos_io_out\[0\]
+ solos_io_out\[10\] solos_io_out\[11\] solos_io_out\[12\] solos_io_out\[1\] solos_io_out\[2\]
+ solos_io_out\[3\] solos_io_out\[4\] solos_io_out\[5\] solos_io_out\[6\] solos_io_out\[7\]
+ solos_io_out\[8\] solos_io_out\[9\] solos_rst vdd vss top_solo_squash
.ends

