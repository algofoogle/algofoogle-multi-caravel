module asic_hat_logo(
`ifdef USE_POWER_PINS
	inout vdd,
	inout vss
`endif
);
endmodule
